module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 ;
  assign n256 = x240 ^ x61 ^ 1'b0 ;
  assign n257 = x103 & n256 ;
  assign n258 = x112 & x132 ;
  assign n259 = n258 ^ x153 ^ 1'b0 ;
  assign n260 = x25 & x235 ;
  assign n261 = ~x13 & n260 ;
  assign n262 = x42 ^ x9 ^ 1'b0 ;
  assign n263 = x128 & n262 ;
  assign n264 = ( x8 & x52 ) | ( x8 & ~x108 ) | ( x52 & ~x108 ) ;
  assign n265 = x125 & n264 ;
  assign n266 = n265 ^ x253 ^ 1'b0 ;
  assign n267 = ( ~x30 & x196 ) | ( ~x30 & x218 ) | ( x196 & x218 ) ;
  assign n268 = n267 ^ x108 ^ x45 ;
  assign n269 = ( ~x151 & x223 ) | ( ~x151 & x249 ) | ( x223 & x249 ) ;
  assign n270 = x171 ^ x102 ^ x31 ;
  assign n271 = ( x10 & x49 ) | ( x10 & ~x179 ) | ( x49 & ~x179 ) ;
  assign n272 = x61 & n271 ;
  assign n273 = n272 ^ x114 ^ 1'b0 ;
  assign n278 = ( ~x31 & x140 ) | ( ~x31 & x147 ) | ( x140 & x147 ) ;
  assign n274 = x232 ^ x169 ^ x41 ;
  assign n275 = n274 ^ x225 ^ x202 ;
  assign n276 = x113 & n275 ;
  assign n277 = n276 ^ x104 ^ 1'b0 ;
  assign n279 = n278 ^ n277 ^ x144 ;
  assign n282 = ( x53 & ~x54 ) | ( x53 & x65 ) | ( ~x54 & x65 ) ;
  assign n280 = ( x28 & ~x95 ) | ( x28 & x234 ) | ( ~x95 & x234 ) ;
  assign n281 = x238 & n280 ;
  assign n283 = n282 ^ n281 ^ 1'b0 ;
  assign n284 = n283 ^ n271 ^ x146 ;
  assign n285 = x109 & x192 ;
  assign n286 = n285 ^ n274 ^ 1'b0 ;
  assign n287 = ( x100 & ~x126 ) | ( x100 & x215 ) | ( ~x126 & x215 ) ;
  assign n288 = ( x108 & x195 ) | ( x108 & ~x219 ) | ( x195 & ~x219 ) ;
  assign n289 = ( x58 & ~x188 ) | ( x58 & n288 ) | ( ~x188 & n288 ) ;
  assign n290 = n289 ^ x176 ^ x3 ;
  assign n291 = x254 ^ x73 ^ x45 ;
  assign n292 = x55 & ~n291 ;
  assign n293 = n292 ^ x75 ^ 1'b0 ;
  assign n294 = x113 & x157 ;
  assign n295 = n294 ^ x82 ^ 1'b0 ;
  assign n299 = x225 ^ x212 ^ x76 ;
  assign n296 = x167 & ~n263 ;
  assign n297 = x105 & n296 ;
  assign n298 = n297 ^ x188 ^ 1'b0 ;
  assign n300 = n299 ^ n298 ^ x162 ;
  assign n301 = ( x26 & x236 ) | ( x26 & n300 ) | ( x236 & n300 ) ;
  assign n302 = x129 ^ x47 ^ x29 ;
  assign n303 = x89 & x97 ;
  assign n304 = n302 & n303 ;
  assign n305 = x128 ^ x123 ^ 1'b0 ;
  assign n306 = x247 & n305 ;
  assign n307 = x30 & n306 ;
  assign n308 = n307 ^ x145 ^ 1'b0 ;
  assign n309 = x4 & x170 ;
  assign n310 = n309 ^ x144 ^ 1'b0 ;
  assign n311 = n310 ^ x163 ^ x94 ;
  assign n312 = ( x34 & ~x65 ) | ( x34 & x160 ) | ( ~x65 & x160 ) ;
  assign n313 = n312 ^ n291 ^ n268 ;
  assign n314 = n313 ^ x182 ^ 1'b0 ;
  assign n315 = n311 & ~n314 ;
  assign n318 = ( x9 & x11 ) | ( x9 & ~x76 ) | ( x11 & ~x76 ) ;
  assign n316 = x221 ^ x105 ^ 1'b0 ;
  assign n317 = x145 & n316 ;
  assign n319 = n318 ^ n317 ^ 1'b0 ;
  assign n320 = x78 & n319 ;
  assign n321 = ( x17 & x153 ) | ( x17 & ~x241 ) | ( x153 & ~x241 ) ;
  assign n322 = x28 & n321 ;
  assign n323 = n322 ^ x177 ^ 1'b0 ;
  assign n324 = ( ~x14 & x32 ) | ( ~x14 & x126 ) | ( x32 & x126 ) ;
  assign n325 = x222 ^ x207 ^ x107 ;
  assign n326 = ( x66 & ~x120 ) | ( x66 & x239 ) | ( ~x120 & x239 ) ;
  assign n327 = ( ~x77 & x101 ) | ( ~x77 & n326 ) | ( x101 & n326 ) ;
  assign n328 = ( x65 & n325 ) | ( x65 & n327 ) | ( n325 & n327 ) ;
  assign n329 = x226 & n293 ;
  assign n330 = ( x4 & ~x92 ) | ( x4 & x135 ) | ( ~x92 & x135 ) ;
  assign n331 = ( x161 & ~x185 ) | ( x161 & n330 ) | ( ~x185 & n330 ) ;
  assign n332 = ( x210 & ~x230 ) | ( x210 & n257 ) | ( ~x230 & n257 ) ;
  assign n340 = ( x33 & x136 ) | ( x33 & ~x179 ) | ( x136 & ~x179 ) ;
  assign n335 = x251 ^ x140 ^ 1'b0 ;
  assign n336 = x57 & n335 ;
  assign n337 = ( ~x106 & x144 ) | ( ~x106 & x177 ) | ( x144 & x177 ) ;
  assign n338 = n337 ^ x100 ^ 1'b0 ;
  assign n339 = n336 & n338 ;
  assign n341 = n340 ^ n339 ^ n337 ;
  assign n333 = x230 ^ x122 ^ x31 ;
  assign n334 = ( x12 & ~x40 ) | ( x12 & n333 ) | ( ~x40 & n333 ) ;
  assign n342 = n341 ^ n334 ^ x37 ;
  assign n343 = ~x235 & x243 ;
  assign n348 = ( ~x95 & x187 ) | ( ~x95 & x252 ) | ( x187 & x252 ) ;
  assign n349 = n348 ^ x155 ^ x104 ;
  assign n346 = ( x42 & x89 ) | ( x42 & ~x223 ) | ( x89 & ~x223 ) ;
  assign n345 = x209 ^ x168 ^ x120 ;
  assign n347 = n346 ^ n345 ^ x203 ;
  assign n344 = x211 & ~n291 ;
  assign n350 = n349 ^ n347 ^ n344 ;
  assign n351 = x249 ^ x152 ^ 1'b0 ;
  assign n352 = x146 & ~n351 ;
  assign n353 = x164 ^ x92 ^ 1'b0 ;
  assign n354 = x35 & x210 ;
  assign n355 = ~x148 & n354 ;
  assign n356 = ( x187 & n353 ) | ( x187 & n355 ) | ( n353 & n355 ) ;
  assign n357 = n304 ^ n283 ^ x97 ;
  assign n358 = ( ~x132 & n278 ) | ( ~x132 & n318 ) | ( n278 & n318 ) ;
  assign n359 = ( ~x178 & n277 ) | ( ~x178 & n358 ) | ( n277 & n358 ) ;
  assign n360 = n359 ^ x252 ^ x145 ;
  assign n361 = x229 ^ x122 ^ x75 ;
  assign n362 = n318 & ~n361 ;
  assign n363 = n362 ^ n326 ^ 1'b0 ;
  assign n364 = x178 & ~x247 ;
  assign n365 = ( x57 & n270 ) | ( x57 & n364 ) | ( n270 & n364 ) ;
  assign n367 = ( ~x0 & x132 ) | ( ~x0 & x135 ) | ( x132 & x135 ) ;
  assign n368 = n367 ^ x241 ^ x34 ;
  assign n366 = n321 ^ x161 ^ x35 ;
  assign n369 = n368 ^ n366 ^ n357 ;
  assign n370 = x68 & x112 ;
  assign n371 = n323 ^ x183 ^ 1'b0 ;
  assign n372 = ( x233 & ~n370 ) | ( x233 & n371 ) | ( ~n370 & n371 ) ;
  assign n373 = n372 ^ x129 ^ x127 ;
  assign n374 = ( x163 & ~n278 ) | ( x163 & n311 ) | ( ~n278 & n311 ) ;
  assign n375 = ~x10 & n374 ;
  assign n376 = n375 ^ x118 ^ 1'b0 ;
  assign n377 = n331 ^ n306 ^ 1'b0 ;
  assign n378 = x93 & n377 ;
  assign n379 = n311 ^ x247 ^ x190 ;
  assign n380 = x244 ^ x183 ^ x66 ;
  assign n381 = ( x155 & ~n379 ) | ( x155 & n380 ) | ( ~n379 & n380 ) ;
  assign n388 = x115 & x142 ;
  assign n389 = n388 ^ x104 ^ 1'b0 ;
  assign n390 = ( x2 & n275 ) | ( x2 & n389 ) | ( n275 & n389 ) ;
  assign n382 = n318 ^ x228 ^ x148 ;
  assign n384 = ( x151 & ~x178 ) | ( x151 & x198 ) | ( ~x178 & x198 ) ;
  assign n383 = ( x71 & x169 ) | ( x71 & ~x182 ) | ( x169 & ~x182 ) ;
  assign n385 = n384 ^ n383 ^ x79 ;
  assign n386 = n382 | n385 ;
  assign n387 = x102 | n386 ;
  assign n391 = n390 ^ n387 ^ n315 ;
  assign n395 = ( ~x197 & x221 ) | ( ~x197 & n349 ) | ( x221 & n349 ) ;
  assign n392 = x70 & x146 ;
  assign n393 = n392 ^ x17 ^ 1'b0 ;
  assign n394 = n393 ^ n264 ^ x141 ;
  assign n396 = n395 ^ n394 ^ x10 ;
  assign n397 = x45 ^ x8 ^ 1'b0 ;
  assign n398 = ( x104 & x142 ) | ( x104 & n290 ) | ( x142 & n290 ) ;
  assign n399 = ( ~x205 & x206 ) | ( ~x205 & x232 ) | ( x206 & x232 ) ;
  assign n400 = n399 ^ n373 ^ x92 ;
  assign n401 = ( x30 & ~x54 ) | ( x30 & x145 ) | ( ~x54 & x145 ) ;
  assign n402 = x250 ^ x90 ^ x49 ;
  assign n403 = n402 ^ n296 ^ 1'b0 ;
  assign n404 = n401 & ~n403 ;
  assign n405 = x135 ^ x64 ^ x56 ;
  assign n406 = ( x140 & ~x147 ) | ( x140 & x237 ) | ( ~x147 & x237 ) ;
  assign n407 = ( ~x81 & x116 ) | ( ~x81 & x121 ) | ( x116 & x121 ) ;
  assign n408 = ( x158 & ~n320 ) | ( x158 & n407 ) | ( ~n320 & n407 ) ;
  assign n409 = ( n405 & ~n406 ) | ( n405 & n408 ) | ( ~n406 & n408 ) ;
  assign n412 = x88 ^ x34 ^ x25 ;
  assign n413 = x107 ^ x14 ^ 1'b0 ;
  assign n414 = ~n412 & n413 ;
  assign n410 = ( ~x127 & x138 ) | ( ~x127 & n280 ) | ( x138 & n280 ) ;
  assign n411 = n263 & n410 ;
  assign n415 = n414 ^ n411 ^ 1'b0 ;
  assign n416 = ( x145 & x154 ) | ( x145 & ~x187 ) | ( x154 & ~x187 ) ;
  assign n417 = x32 & x131 ;
  assign n418 = ~n278 & n417 ;
  assign n419 = ( x163 & n416 ) | ( x163 & n418 ) | ( n416 & n418 ) ;
  assign n420 = ( x41 & x45 ) | ( x41 & ~x236 ) | ( x45 & ~x236 ) ;
  assign n421 = ( x52 & x149 ) | ( x52 & ~n420 ) | ( x149 & ~n420 ) ;
  assign n422 = n346 ^ n313 ^ x96 ;
  assign n423 = n421 & n422 ;
  assign n424 = ( x223 & n408 ) | ( x223 & ~n423 ) | ( n408 & ~n423 ) ;
  assign n425 = ( x71 & ~x99 ) | ( x71 & x135 ) | ( ~x99 & x135 ) ;
  assign n426 = n425 ^ x24 ^ 1'b0 ;
  assign n427 = x188 & n426 ;
  assign n428 = n326 ^ x163 ^ 1'b0 ;
  assign n429 = x9 & n428 ;
  assign n430 = ( n393 & n427 ) | ( n393 & ~n429 ) | ( n427 & ~n429 ) ;
  assign n431 = x233 ^ x111 ^ x19 ;
  assign n432 = n312 ^ x192 ^ 1'b0 ;
  assign n433 = x145 & n432 ;
  assign n434 = n433 ^ n311 ^ x139 ;
  assign n435 = x192 ^ x157 ^ 1'b0 ;
  assign n436 = x43 & n435 ;
  assign n437 = x227 ^ x18 ^ 1'b0 ;
  assign n438 = n436 & n437 ;
  assign n439 = n308 ^ x134 ^ 1'b0 ;
  assign n440 = n438 & ~n439 ;
  assign n441 = ~x131 & n336 ;
  assign n442 = x235 ^ x206 ^ x68 ;
  assign n443 = n321 & ~n442 ;
  assign n444 = ~x127 & n443 ;
  assign n445 = n298 ^ x139 ^ 1'b0 ;
  assign n446 = n444 | n445 ;
  assign n447 = ( x100 & x111 ) | ( x100 & ~x168 ) | ( x111 & ~x168 ) ;
  assign n448 = x31 & ~n261 ;
  assign n449 = ~x17 & n448 ;
  assign n450 = n447 | n449 ;
  assign n451 = x235 & n450 ;
  assign n452 = n446 & n451 ;
  assign n453 = n444 ^ x93 ^ 1'b0 ;
  assign n454 = x13 & x106 ;
  assign n455 = n454 ^ x126 ^ 1'b0 ;
  assign n456 = ( x45 & x108 ) | ( x45 & n310 ) | ( x108 & n310 ) ;
  assign n457 = n456 ^ x15 ^ 1'b0 ;
  assign n458 = n356 & n457 ;
  assign n459 = x165 ^ x101 ^ x7 ;
  assign n460 = ( x7 & x120 ) | ( x7 & n459 ) | ( x120 & n459 ) ;
  assign n461 = x69 ^ x20 ^ 1'b0 ;
  assign n462 = n447 ^ n306 ^ x215 ;
  assign n463 = x12 & n462 ;
  assign n464 = x81 & x199 ;
  assign n465 = n464 ^ x121 ^ 1'b0 ;
  assign n466 = ( x79 & x198 ) | ( x79 & ~x202 ) | ( x198 & ~x202 ) ;
  assign n469 = n275 ^ x227 ^ x105 ;
  assign n470 = n469 ^ x196 ^ x115 ;
  assign n468 = ( x41 & x58 ) | ( x41 & ~x170 ) | ( x58 & ~x170 ) ;
  assign n471 = n470 ^ n468 ^ x246 ;
  assign n467 = n288 ^ x14 ^ 1'b0 ;
  assign n472 = n471 ^ n467 ^ 1'b0 ;
  assign n473 = n466 & ~n472 ;
  assign n474 = ( x132 & n465 ) | ( x132 & ~n473 ) | ( n465 & ~n473 ) ;
  assign n477 = x8 & x215 ;
  assign n478 = n477 ^ x249 ^ 1'b0 ;
  assign n475 = ( ~x126 & x169 ) | ( ~x126 & x236 ) | ( x169 & x236 ) ;
  assign n476 = ~n320 & n475 ;
  assign n479 = n478 ^ n476 ^ 1'b0 ;
  assign n480 = x71 & n479 ;
  assign n481 = x196 ^ x17 ^ 1'b0 ;
  assign n482 = ( n357 & n433 ) | ( n357 & ~n481 ) | ( n433 & ~n481 ) ;
  assign n483 = x7 & n339 ;
  assign n484 = ~x229 & n483 ;
  assign n485 = n277 ^ x214 ^ x89 ;
  assign n486 = n484 & n485 ;
  assign n488 = ( x110 & x156 ) | ( x110 & ~x220 ) | ( x156 & ~x220 ) ;
  assign n487 = n449 ^ n423 ^ n329 ;
  assign n489 = n488 ^ n487 ^ x92 ;
  assign n490 = ( x86 & x219 ) | ( x86 & ~n489 ) | ( x219 & ~n489 ) ;
  assign n491 = ( x49 & ~x104 ) | ( x49 & n320 ) | ( ~x104 & n320 ) ;
  assign n492 = ( ~x107 & n320 ) | ( ~x107 & n491 ) | ( n320 & n491 ) ;
  assign n493 = x35 & ~n442 ;
  assign n494 = n493 ^ x207 ^ 1'b0 ;
  assign n495 = ( ~x240 & n367 ) | ( ~x240 & n494 ) | ( n367 & n494 ) ;
  assign n496 = x158 ^ x98 ^ x75 ;
  assign n497 = ( ~x52 & x62 ) | ( ~x52 & n442 ) | ( x62 & n442 ) ;
  assign n498 = ( x122 & n496 ) | ( x122 & ~n497 ) | ( n496 & ~n497 ) ;
  assign n499 = n498 ^ x141 ^ 1'b0 ;
  assign n500 = n499 ^ n414 ^ n278 ;
  assign n501 = ( ~x114 & n387 ) | ( ~x114 & n433 ) | ( n387 & n433 ) ;
  assign n502 = ( x212 & n500 ) | ( x212 & ~n501 ) | ( n500 & ~n501 ) ;
  assign n503 = ( x15 & x36 ) | ( x15 & n291 ) | ( x36 & n291 ) ;
  assign n504 = n465 ^ x226 ^ x59 ;
  assign n505 = n340 ^ x223 ^ x170 ;
  assign n506 = n383 ^ x199 ^ 1'b0 ;
  assign n507 = x12 & n506 ;
  assign n508 = ( n504 & n505 ) | ( n504 & n507 ) | ( n505 & n507 ) ;
  assign n509 = ( ~n424 & n503 ) | ( ~n424 & n508 ) | ( n503 & n508 ) ;
  assign n510 = n509 ^ x143 ^ 1'b0 ;
  assign n511 = n502 & n510 ;
  assign n512 = x156 & x245 ;
  assign n513 = ~x31 & n512 ;
  assign n522 = ( x157 & ~x175 ) | ( x157 & n286 ) | ( ~x175 & n286 ) ;
  assign n523 = x79 & n327 ;
  assign n524 = ( n259 & n269 ) | ( n259 & ~n523 ) | ( n269 & ~n523 ) ;
  assign n525 = ( ~n290 & n522 ) | ( ~n290 & n524 ) | ( n522 & n524 ) ;
  assign n516 = n346 ^ x131 ^ x11 ;
  assign n514 = x105 & n312 ;
  assign n515 = n514 ^ n390 ^ 1'b0 ;
  assign n517 = n516 ^ n515 ^ n301 ;
  assign n518 = n415 ^ n374 ^ 1'b0 ;
  assign n519 = n517 | n518 ;
  assign n520 = ~x157 & n499 ;
  assign n521 = n519 | n520 ;
  assign n526 = n525 ^ n521 ^ 1'b0 ;
  assign n527 = n513 & n526 ;
  assign n529 = x147 ^ x64 ^ 1'b0 ;
  assign n530 = ( ~x102 & x209 ) | ( ~x102 & n529 ) | ( x209 & n529 ) ;
  assign n528 = ~x179 & n279 ;
  assign n531 = n530 ^ n528 ^ n358 ;
  assign n532 = ( ~x98 & x235 ) | ( ~x98 & n530 ) | ( x235 & n530 ) ;
  assign n533 = x43 & n532 ;
  assign n534 = n533 ^ n516 ^ 1'b0 ;
  assign n535 = n534 ^ x202 ^ 1'b0 ;
  assign n537 = n356 ^ x164 ^ 1'b0 ;
  assign n536 = n367 ^ x233 ^ 1'b0 ;
  assign n538 = n537 ^ n536 ^ n441 ;
  assign n539 = x183 ^ x84 ^ x7 ;
  assign n540 = n539 ^ n344 ^ x81 ;
  assign n541 = x195 ^ x9 ^ 1'b0 ;
  assign n542 = ( ~x15 & x69 ) | ( ~x15 & x105 ) | ( x69 & x105 ) ;
  assign n543 = x31 & n542 ;
  assign n544 = n543 ^ n534 ^ 1'b0 ;
  assign n545 = ( n298 & n449 ) | ( n298 & ~n544 ) | ( n449 & ~n544 ) ;
  assign n546 = ( n327 & n394 ) | ( n327 & n545 ) | ( n394 & n545 ) ;
  assign n547 = x171 & n410 ;
  assign n548 = ( x68 & ~x143 ) | ( x68 & x225 ) | ( ~x143 & x225 ) ;
  assign n549 = n548 ^ n458 ^ x62 ;
  assign n550 = n270 ^ n261 ^ x14 ;
  assign n551 = x142 ^ x96 ^ 1'b0 ;
  assign n552 = x12 & n551 ;
  assign n553 = ( ~x111 & n315 ) | ( ~x111 & n364 ) | ( n315 & n364 ) ;
  assign n554 = n513 | n553 ;
  assign n555 = n552 | n554 ;
  assign n556 = ( x7 & ~x47 ) | ( x7 & x184 ) | ( ~x47 & x184 ) ;
  assign n557 = n336 ^ n277 ^ x179 ;
  assign n558 = ( x162 & x204 ) | ( x162 & ~n557 ) | ( x204 & ~n557 ) ;
  assign n559 = ( ~n321 & n556 ) | ( ~n321 & n558 ) | ( n556 & n558 ) ;
  assign n560 = ( x111 & ~x167 ) | ( x111 & n482 ) | ( ~x167 & n482 ) ;
  assign n561 = n492 ^ n409 ^ 1'b0 ;
  assign n562 = n485 ^ x197 ^ x141 ;
  assign n563 = ( x133 & ~n277 ) | ( x133 & n562 ) | ( ~n277 & n562 ) ;
  assign n564 = x140 & x174 ;
  assign n565 = n564 ^ x67 ^ 1'b0 ;
  assign n566 = ( x85 & ~n353 ) | ( x85 & n565 ) | ( ~n353 & n565 ) ;
  assign n567 = n374 ^ n267 ^ 1'b0 ;
  assign n568 = x188 & n567 ;
  assign n569 = ~n261 & n568 ;
  assign n570 = n566 & n569 ;
  assign n571 = ( ~x90 & x121 ) | ( ~x90 & x154 ) | ( x121 & x154 ) ;
  assign n572 = ( x46 & x147 ) | ( x46 & ~n571 ) | ( x147 & ~n571 ) ;
  assign n573 = n572 ^ n387 ^ x72 ;
  assign n574 = n429 | n573 ;
  assign n582 = ( x138 & ~x201 ) | ( x138 & x222 ) | ( ~x201 & x222 ) ;
  assign n579 = x198 ^ x71 ^ x14 ;
  assign n580 = ( x28 & x189 ) | ( x28 & n579 ) | ( x189 & n579 ) ;
  assign n581 = ( n382 & n390 ) | ( n382 & ~n580 ) | ( n390 & ~n580 ) ;
  assign n577 = n438 ^ x90 ^ 1'b0 ;
  assign n578 = x233 & n577 ;
  assign n583 = n582 ^ n581 ^ n578 ;
  assign n575 = n282 ^ x39 ^ x8 ;
  assign n576 = ( x127 & n519 ) | ( x127 & n575 ) | ( n519 & n575 ) ;
  assign n584 = n583 ^ n576 ^ 1'b0 ;
  assign n585 = n346 & ~n584 ;
  assign n586 = ( x187 & n321 ) | ( x187 & n365 ) | ( n321 & n365 ) ;
  assign n593 = ( ~x172 & x208 ) | ( ~x172 & n383 ) | ( x208 & n383 ) ;
  assign n587 = ( ~x182 & x212 ) | ( ~x182 & n385 ) | ( x212 & n385 ) ;
  assign n588 = x95 & x186 ;
  assign n589 = n588 ^ x118 ^ 1'b0 ;
  assign n590 = x89 & ~n589 ;
  assign n591 = n590 ^ x56 ^ 1'b0 ;
  assign n592 = ( x155 & ~n587 ) | ( x155 & n591 ) | ( ~n587 & n591 ) ;
  assign n594 = n593 ^ n592 ^ n391 ;
  assign n595 = n594 ^ n578 ^ n358 ;
  assign n596 = n586 & ~n595 ;
  assign n597 = n596 ^ n519 ^ 1'b0 ;
  assign n598 = ( ~x14 & x125 ) | ( ~x14 & n496 ) | ( x125 & n496 ) ;
  assign n599 = ( x82 & ~x132 ) | ( x82 & n598 ) | ( ~x132 & n598 ) ;
  assign n600 = n599 ^ n466 ^ x90 ;
  assign n601 = x65 & x159 ;
  assign n602 = ~x187 & n601 ;
  assign n603 = n289 ^ x223 ^ x128 ;
  assign n604 = ( n600 & n602 ) | ( n600 & n603 ) | ( n602 & n603 ) ;
  assign n605 = ( x39 & ~x69 ) | ( x39 & x115 ) | ( ~x69 & x115 ) ;
  assign n606 = x126 ^ x116 ^ x108 ;
  assign n607 = ( x30 & x112 ) | ( x30 & n606 ) | ( x112 & n606 ) ;
  assign n608 = x142 & ~n607 ;
  assign n609 = x151 & ~n608 ;
  assign n610 = n609 ^ x32 ^ 1'b0 ;
  assign n611 = n508 & ~n610 ;
  assign n612 = n611 ^ x85 ^ 1'b0 ;
  assign n613 = x94 & x146 ;
  assign n614 = ~x53 & n613 ;
  assign n615 = ( ~x117 & x133 ) | ( ~x117 & x146 ) | ( x133 & x146 ) ;
  assign n616 = n615 ^ x234 ^ x178 ;
  assign n617 = ( ~n497 & n525 ) | ( ~n497 & n616 ) | ( n525 & n616 ) ;
  assign n618 = ~n614 & n617 ;
  assign n619 = n618 ^ x133 ^ 1'b0 ;
  assign n620 = ( x46 & ~n488 ) | ( x46 & n619 ) | ( ~n488 & n619 ) ;
  assign n621 = x251 ^ x206 ^ x14 ;
  assign n630 = n615 ^ n583 ^ n497 ;
  assign n632 = ( n363 & n526 ) | ( n363 & ~n630 ) | ( n526 & ~n630 ) ;
  assign n622 = ( x106 & x212 ) | ( x106 & ~n498 ) | ( x212 & ~n498 ) ;
  assign n625 = x56 & x216 ;
  assign n626 = ~x97 & n625 ;
  assign n627 = n334 & ~n626 ;
  assign n623 = x6 & ~n366 ;
  assign n624 = ~x207 & n623 ;
  assign n628 = n627 ^ n624 ^ x67 ;
  assign n629 = n622 & ~n628 ;
  assign n631 = n630 ^ n629 ^ 1'b0 ;
  assign n633 = n632 ^ n631 ^ n530 ;
  assign n634 = n535 ^ x185 ^ x164 ;
  assign n635 = n553 ^ x214 ^ x6 ;
  assign n636 = ( n404 & ~n456 ) | ( n404 & n465 ) | ( ~n456 & n465 ) ;
  assign n637 = ( n277 & n635 ) | ( n277 & n636 ) | ( n635 & n636 ) ;
  assign n638 = n302 | n637 ;
  assign n639 = n638 ^ n259 ^ 1'b0 ;
  assign n640 = n478 ^ x250 ^ x2 ;
  assign n641 = n640 ^ x43 ^ 1'b0 ;
  assign n642 = ( ~x7 & x216 ) | ( ~x7 & n641 ) | ( x216 & n641 ) ;
  assign n643 = ( n492 & n639 ) | ( n492 & ~n642 ) | ( n639 & ~n642 ) ;
  assign n646 = x180 ^ x79 ^ 1'b0 ;
  assign n647 = x147 & n646 ;
  assign n644 = ( ~x22 & x121 ) | ( ~x22 & x152 ) | ( x121 & x152 ) ;
  assign n645 = n644 ^ n579 ^ n383 ;
  assign n648 = n647 ^ n645 ^ 1'b0 ;
  assign n650 = ( x51 & ~x89 ) | ( x51 & n326 ) | ( ~x89 & n326 ) ;
  assign n651 = n650 ^ x238 ^ 1'b0 ;
  assign n652 = x24 & n651 ;
  assign n649 = n321 ^ x149 ^ x65 ;
  assign n653 = n652 ^ n649 ^ x7 ;
  assign n655 = n268 ^ x221 ^ x157 ;
  assign n656 = n655 ^ x174 ^ x143 ;
  assign n657 = n326 & ~n656 ;
  assign n654 = x111 & x218 ;
  assign n658 = n657 ^ n654 ^ 1'b0 ;
  assign n659 = n570 ^ n301 ^ x15 ;
  assign n660 = n531 & n659 ;
  assign n661 = n660 ^ n442 ^ 1'b0 ;
  assign n662 = x226 & ~n447 ;
  assign n668 = n320 ^ x152 ^ x143 ;
  assign n665 = ( ~x85 & x98 ) | ( ~x85 & x204 ) | ( x98 & x204 ) ;
  assign n663 = n344 & n356 ;
  assign n664 = n663 ^ n283 ^ 1'b0 ;
  assign n666 = n665 ^ n664 ^ n394 ;
  assign n667 = x98 & n666 ;
  assign n669 = n668 ^ n667 ^ 1'b0 ;
  assign n670 = n410 ^ x196 ^ x134 ;
  assign n671 = x21 & x235 ;
  assign n672 = ~n574 & n671 ;
  assign n673 = x170 ^ x93 ^ x39 ;
  assign n674 = ( x47 & ~x67 ) | ( x47 & n673 ) | ( ~x67 & n673 ) ;
  assign n675 = x62 & x122 ;
  assign n676 = n675 ^ x245 ^ 1'b0 ;
  assign n677 = ( x132 & ~n674 ) | ( x132 & n676 ) | ( ~n674 & n676 ) ;
  assign n678 = ( x21 & x192 ) | ( x21 & ~x245 ) | ( x192 & ~x245 ) ;
  assign n679 = x138 & ~n261 ;
  assign n680 = ~x120 & n679 ;
  assign n681 = ( n391 & n678 ) | ( n391 & ~n680 ) | ( n678 & ~n680 ) ;
  assign n684 = x146 ^ x123 ^ x91 ;
  assign n685 = x135 ^ x51 ^ 1'b0 ;
  assign n686 = x98 & n685 ;
  assign n687 = ( x168 & n684 ) | ( x168 & n686 ) | ( n684 & n686 ) ;
  assign n688 = ( x99 & n268 ) | ( x99 & ~n687 ) | ( n268 & ~n687 ) ;
  assign n689 = ( n401 & ~n404 ) | ( n401 & n688 ) | ( ~n404 & n688 ) ;
  assign n682 = ( x168 & n397 ) | ( x168 & n500 ) | ( n397 & n500 ) ;
  assign n683 = n682 ^ n361 ^ x37 ;
  assign n690 = n689 ^ n683 ^ n399 ;
  assign n691 = ( x37 & x69 ) | ( x37 & ~x126 ) | ( x69 & ~x126 ) ;
  assign n692 = ( ~n373 & n559 ) | ( ~n373 & n691 ) | ( n559 & n691 ) ;
  assign n693 = x161 & n575 ;
  assign n694 = n693 ^ n306 ^ x202 ;
  assign n696 = n532 ^ n313 ^ x181 ;
  assign n695 = x230 & n324 ;
  assign n697 = n696 ^ n695 ^ 1'b0 ;
  assign n698 = n697 ^ n447 ^ x93 ;
  assign n700 = n291 ^ n257 ^ x101 ;
  assign n701 = n700 ^ n652 ^ 1'b0 ;
  assign n702 = x220 & n701 ;
  assign n699 = n522 ^ n450 ^ x97 ;
  assign n703 = n702 ^ n699 ^ 1'b0 ;
  assign n704 = n698 & ~n703 ;
  assign n705 = x146 & ~n290 ;
  assign n706 = n705 ^ x91 ^ 1'b0 ;
  assign n707 = ( n421 & n496 ) | ( n421 & ~n706 ) | ( n496 & ~n706 ) ;
  assign n708 = ( x182 & n560 ) | ( x182 & n707 ) | ( n560 & n707 ) ;
  assign n709 = n326 & ~n497 ;
  assign n710 = n709 ^ n603 ^ 1'b0 ;
  assign n730 = x50 & x136 ;
  assign n731 = n730 ^ x198 ^ 1'b0 ;
  assign n732 = n731 ^ n575 ^ n371 ;
  assign n711 = x221 ^ x202 ^ 1'b0 ;
  assign n712 = x149 & n711 ;
  assign n713 = ~x86 & n712 ;
  assign n714 = x161 & x219 ;
  assign n715 = n713 & n714 ;
  assign n716 = n366 ^ n365 ^ x190 ;
  assign n717 = n716 ^ n306 ^ x65 ;
  assign n720 = ( x2 & x158 ) | ( x2 & ~x217 ) | ( x158 & ~x217 ) ;
  assign n721 = n720 ^ x227 ^ x68 ;
  assign n718 = x188 ^ x24 ^ 1'b0 ;
  assign n719 = x198 & n718 ;
  assign n722 = n721 ^ n719 ^ x25 ;
  assign n723 = ( x58 & x97 ) | ( x58 & ~n722 ) | ( x97 & ~n722 ) ;
  assign n724 = ( ~n269 & n717 ) | ( ~n269 & n723 ) | ( n717 & n723 ) ;
  assign n725 = ( x120 & n525 ) | ( x120 & ~n724 ) | ( n525 & ~n724 ) ;
  assign n726 = x232 ^ x50 ^ 1'b0 ;
  assign n727 = n726 ^ n481 ^ n289 ;
  assign n728 = n727 ^ n605 ^ x216 ;
  assign n729 = ( n715 & n725 ) | ( n715 & ~n728 ) | ( n725 & ~n728 ) ;
  assign n733 = n732 ^ n729 ^ n458 ;
  assign n734 = n733 ^ n344 ^ 1'b0 ;
  assign n735 = n710 & n734 ;
  assign n741 = x141 & ~n268 ;
  assign n742 = n602 & n741 ;
  assign n743 = x216 & ~n742 ;
  assign n744 = n743 ^ n382 ^ 1'b0 ;
  assign n736 = ( n293 & n327 ) | ( n293 & ~n330 ) | ( n327 & ~n330 ) ;
  assign n737 = n674 | n736 ;
  assign n738 = n737 ^ x214 ^ 1'b0 ;
  assign n739 = n738 ^ n583 ^ 1'b0 ;
  assign n740 = n739 ^ x237 ^ x218 ;
  assign n745 = n744 ^ n740 ^ x152 ;
  assign n746 = n673 ^ n478 ^ 1'b0 ;
  assign n747 = ~n598 & n746 ;
  assign n748 = n747 ^ n284 ^ x221 ;
  assign n749 = n402 ^ x122 ^ x54 ;
  assign n750 = ~n475 & n749 ;
  assign n751 = x169 | n750 ;
  assign n753 = x218 ^ x35 ^ 1'b0 ;
  assign n754 = x37 & n753 ;
  assign n755 = n754 ^ n277 ^ n268 ;
  assign n752 = ( x127 & ~x194 ) | ( x127 & n431 ) | ( ~x194 & n431 ) ;
  assign n756 = n755 ^ n752 ^ x135 ;
  assign n757 = n756 ^ n379 ^ x89 ;
  assign n758 = n282 ^ n263 ^ x50 ;
  assign n759 = n758 ^ x210 ^ x149 ;
  assign n762 = ( x171 & ~x208 ) | ( x171 & n310 ) | ( ~x208 & n310 ) ;
  assign n760 = n758 ^ n552 ^ n357 ;
  assign n761 = n664 & n760 ;
  assign n763 = n762 ^ n761 ^ 1'b0 ;
  assign n764 = ~n759 & n763 ;
  assign n765 = n645 ^ n581 ^ x59 ;
  assign n766 = ( x158 & ~n346 ) | ( x158 & n765 ) | ( ~n346 & n765 ) ;
  assign n767 = n348 & n600 ;
  assign n768 = n767 ^ x76 ^ 1'b0 ;
  assign n769 = x200 & ~n768 ;
  assign n770 = ~n766 & n769 ;
  assign n771 = ( x25 & x64 ) | ( x25 & ~x137 ) | ( x64 & ~x137 ) ;
  assign n772 = n771 ^ n347 ^ x154 ;
  assign n773 = n355 & ~n772 ;
  assign n774 = n486 ^ n395 ^ x92 ;
  assign n775 = n522 ^ n501 ^ x131 ;
  assign n776 = n775 ^ n744 ^ 1'b0 ;
  assign n777 = n774 | n776 ;
  assign n778 = ( x116 & ~x197 ) | ( x116 & n298 ) | ( ~x197 & n298 ) ;
  assign n779 = n647 ^ n301 ^ n261 ;
  assign n780 = ~n341 & n779 ;
  assign n781 = ~x13 & n780 ;
  assign n782 = n778 | n781 ;
  assign n783 = n607 | n782 ;
  assign n784 = ~x117 & x252 ;
  assign n785 = n652 ^ x158 ^ x118 ;
  assign n786 = ( n270 & ~n310 ) | ( n270 & n785 ) | ( ~n310 & n785 ) ;
  assign n787 = n656 ^ n503 ^ x62 ;
  assign n788 = n465 ^ n433 ^ n414 ;
  assign n789 = ( x144 & n313 ) | ( x144 & n788 ) | ( n313 & n788 ) ;
  assign n790 = ( n275 & ~n787 ) | ( n275 & n789 ) | ( ~n787 & n789 ) ;
  assign n791 = ( ~n310 & n471 ) | ( ~n310 & n656 ) | ( n471 & n656 ) ;
  assign n793 = ( x58 & x92 ) | ( x58 & ~n327 ) | ( x92 & ~n327 ) ;
  assign n794 = n793 ^ x161 ^ x101 ;
  assign n795 = n794 ^ n293 ^ n290 ;
  assign n796 = ( n400 & ~n556 ) | ( n400 & n795 ) | ( ~n556 & n795 ) ;
  assign n797 = n796 ^ n614 ^ x166 ;
  assign n792 = n726 & ~n773 ;
  assign n798 = n797 ^ n792 ^ 1'b0 ;
  assign n801 = ( x36 & x40 ) | ( x36 & ~n436 ) | ( x40 & ~n436 ) ;
  assign n799 = ( ~x38 & x189 ) | ( ~x38 & n376 ) | ( x189 & n376 ) ;
  assign n800 = n799 ^ n318 ^ 1'b0 ;
  assign n802 = n801 ^ n800 ^ 1'b0 ;
  assign n803 = ( x243 & ~x248 ) | ( x243 & n592 ) | ( ~x248 & n592 ) ;
  assign n804 = n656 ^ x74 ^ 1'b0 ;
  assign n805 = x102 & ~n804 ;
  assign n806 = n805 ^ x117 ^ 1'b0 ;
  assign n807 = n321 & n806 ;
  assign n808 = ( ~x11 & x111 ) | ( ~x11 & x222 ) | ( x111 & x222 ) ;
  assign n809 = n808 ^ n720 ^ n488 ;
  assign n810 = x179 & ~n809 ;
  assign n811 = n800 & n810 ;
  assign n812 = ( x59 & n427 ) | ( x59 & n794 ) | ( n427 & n794 ) ;
  assign n813 = n438 ^ x77 ^ x26 ;
  assign n814 = ( n650 & n779 ) | ( n650 & n813 ) | ( n779 & n813 ) ;
  assign n815 = n812 & n814 ;
  assign n816 = n644 ^ n536 ^ 1'b0 ;
  assign n817 = n815 & ~n816 ;
  assign n818 = n817 ^ n658 ^ n467 ;
  assign n819 = ( n499 & n560 ) | ( n499 & n768 ) | ( n560 & n768 ) ;
  assign n820 = ( x54 & ~x221 ) | ( x54 & n819 ) | ( ~x221 & n819 ) ;
  assign n821 = n357 ^ n278 ^ 1'b0 ;
  assign n822 = ( n310 & n640 ) | ( n310 & ~n690 ) | ( n640 & ~n690 ) ;
  assign n826 = n697 ^ x126 ^ 1'b0 ;
  assign n827 = n449 | n826 ;
  assign n824 = x137 & x252 ;
  assign n825 = ~x243 & n824 ;
  assign n823 = n684 ^ x135 ^ x80 ;
  assign n828 = n827 ^ n825 ^ n823 ;
  assign n829 = ( n634 & ~n759 ) | ( n634 & n828 ) | ( ~n759 & n828 ) ;
  assign n830 = n353 | n469 ;
  assign n831 = ( ~x7 & x208 ) | ( ~x7 & n626 ) | ( x208 & n626 ) ;
  assign n832 = n532 & ~n831 ;
  assign n833 = ~n353 & n832 ;
  assign n834 = ( x74 & n401 ) | ( x74 & n833 ) | ( n401 & n833 ) ;
  assign n835 = n657 ^ x227 ^ x92 ;
  assign n836 = ( x27 & ~n834 ) | ( x27 & n835 ) | ( ~n834 & n835 ) ;
  assign n837 = ( n284 & n830 ) | ( n284 & n836 ) | ( n830 & n836 ) ;
  assign n838 = n837 ^ n752 ^ n732 ;
  assign n846 = n313 ^ x179 ^ x38 ;
  assign n844 = n348 ^ x238 ^ 1'b0 ;
  assign n845 = x92 & n844 ;
  assign n847 = n846 ^ n845 ^ x223 ;
  assign n842 = n429 ^ n382 ^ x72 ;
  assign n843 = x231 & n842 ;
  assign n848 = n847 ^ n843 ^ x88 ;
  assign n849 = n848 ^ n465 ^ x197 ;
  assign n839 = n333 | n341 ;
  assign n840 = n839 ^ x61 ^ 1'b0 ;
  assign n841 = n840 ^ n678 ^ n370 ;
  assign n850 = n849 ^ n841 ^ x248 ;
  assign n851 = n673 ^ n339 ^ 1'b0 ;
  assign n852 = x18 & ~n851 ;
  assign n853 = ( x69 & n270 ) | ( x69 & n852 ) | ( n270 & n852 ) ;
  assign n854 = n665 ^ n356 ^ n352 ;
  assign n855 = n854 ^ x165 ^ 1'b0 ;
  assign n856 = n853 & n855 ;
  assign n857 = x27 & ~n856 ;
  assign n858 = n607 ^ x225 ^ x136 ;
  assign n859 = n401 ^ x56 ^ 1'b0 ;
  assign n860 = ( n466 & ~n711 ) | ( n466 & n859 ) | ( ~n711 & n859 ) ;
  assign n861 = x222 ^ x68 ^ 1'b0 ;
  assign n862 = n861 ^ n586 ^ 1'b0 ;
  assign n863 = n860 & n862 ;
  assign n864 = ( n857 & ~n858 ) | ( n857 & n863 ) | ( ~n858 & n863 ) ;
  assign n865 = ( x83 & x254 ) | ( x83 & ~n864 ) | ( x254 & ~n864 ) ;
  assign n866 = x101 | n689 ;
  assign n867 = n725 ^ n592 ^ 1'b0 ;
  assign n868 = n866 & n867 ;
  assign n869 = ( ~n326 & n535 ) | ( ~n326 & n868 ) | ( n535 & n868 ) ;
  assign n870 = n423 ^ n328 ^ 1'b0 ;
  assign n875 = x8 & n562 ;
  assign n872 = n571 ^ n264 ^ x200 ;
  assign n871 = n412 ^ n259 ^ 1'b0 ;
  assign n873 = n872 ^ n871 ^ x177 ;
  assign n874 = ( n586 & n628 ) | ( n586 & n873 ) | ( n628 & n873 ) ;
  assign n876 = n875 ^ n874 ^ n259 ;
  assign n877 = n469 | n771 ;
  assign n879 = x222 & n264 ;
  assign n880 = n879 ^ n720 ^ 1'b0 ;
  assign n881 = ( x136 & ~x227 ) | ( x136 & n880 ) | ( ~x227 & n880 ) ;
  assign n878 = x52 & n278 ;
  assign n882 = n881 ^ n878 ^ 1'b0 ;
  assign n883 = ( n834 & n877 ) | ( n834 & ~n882 ) | ( n877 & ~n882 ) ;
  assign n884 = x186 & n883 ;
  assign n885 = n884 ^ n722 ^ 1'b0 ;
  assign n886 = x132 & ~n885 ;
  assign n887 = n637 ^ n519 ^ n427 ;
  assign n888 = n628 ^ n520 ^ 1'b0 ;
  assign n889 = n542 & n888 ;
  assign n890 = n889 ^ n749 ^ n515 ;
  assign n891 = n517 ^ n345 ^ x155 ;
  assign n892 = n891 ^ n470 ^ 1'b0 ;
  assign n893 = x189 & ~n602 ;
  assign n894 = n893 ^ n383 ^ 1'b0 ;
  assign n895 = x115 & ~n894 ;
  assign n896 = n677 | n895 ;
  assign n897 = n751 ^ n565 ^ x78 ;
  assign n904 = n656 ^ n344 ^ x48 ;
  assign n899 = ~x236 & n466 ;
  assign n900 = n637 | n899 ;
  assign n901 = n446 & ~n900 ;
  assign n902 = n901 ^ n304 ^ x158 ;
  assign n898 = x82 & n279 ;
  assign n903 = n902 ^ n898 ^ n301 ;
  assign n905 = n904 ^ n903 ^ n845 ;
  assign n907 = n615 ^ n504 ^ n438 ;
  assign n908 = ( x193 & ~n542 ) | ( x193 & n907 ) | ( ~n542 & n907 ) ;
  assign n906 = n504 ^ n434 ^ n271 ;
  assign n909 = n908 ^ n906 ^ 1'b0 ;
  assign n910 = x252 ^ x226 ^ x95 ;
  assign n911 = n910 ^ n284 ^ x127 ;
  assign n912 = n911 ^ x139 ^ 1'b0 ;
  assign n913 = n912 ^ n783 ^ n591 ;
  assign n914 = x62 & n446 ;
  assign n915 = ( x57 & ~n488 ) | ( x57 & n914 ) | ( ~n488 & n914 ) ;
  assign n916 = n915 ^ n574 ^ n261 ;
  assign n918 = n532 ^ x44 ^ 1'b0 ;
  assign n917 = n783 ^ n329 ^ x97 ;
  assign n919 = n918 ^ n917 ^ n456 ;
  assign n920 = ( n744 & n770 ) | ( n744 & n919 ) | ( n770 & n919 ) ;
  assign n921 = ( x151 & n459 ) | ( x151 & ~n604 ) | ( n459 & ~n604 ) ;
  assign n922 = ( ~x99 & n542 ) | ( ~x99 & n912 ) | ( n542 & n912 ) ;
  assign n923 = n922 ^ n572 ^ 1'b0 ;
  assign n924 = n801 & n923 ;
  assign n925 = ~x127 & n924 ;
  assign n927 = n361 ^ x210 ^ x179 ;
  assign n928 = n927 ^ n391 ^ x150 ;
  assign n926 = x117 & ~n850 ;
  assign n929 = n928 ^ n926 ^ 1'b0 ;
  assign n930 = ~x147 & x234 ;
  assign n931 = ( x72 & n369 ) | ( x72 & ~n756 ) | ( n369 & ~n756 ) ;
  assign n932 = n931 ^ n901 ^ 1'b0 ;
  assign n933 = ( n301 & n488 ) | ( n301 & n755 ) | ( n488 & n755 ) ;
  assign n934 = n750 ^ n503 ^ 1'b0 ;
  assign n935 = ( x190 & n933 ) | ( x190 & n934 ) | ( n933 & n934 ) ;
  assign n936 = n935 ^ n328 ^ 1'b0 ;
  assign n938 = x190 & n760 ;
  assign n937 = n420 & n687 ;
  assign n939 = n938 ^ n937 ^ 1'b0 ;
  assign n940 = x184 & n475 ;
  assign n941 = ~x59 & n940 ;
  assign n942 = ~n797 & n941 ;
  assign n943 = x197 & ~n364 ;
  assign n944 = n943 ^ n269 ^ 1'b0 ;
  assign n945 = n870 & ~n944 ;
  assign n954 = x84 & ~n487 ;
  assign n955 = n954 ^ x89 ^ 1'b0 ;
  assign n953 = n412 ^ x241 ^ x90 ;
  assign n948 = n289 ^ x151 ^ x129 ;
  assign n949 = n302 | n948 ;
  assign n950 = n949 ^ x113 ^ 1'b0 ;
  assign n951 = ( n341 & n459 ) | ( n341 & n950 ) | ( n459 & n950 ) ;
  assign n947 = n578 ^ n496 ^ x88 ;
  assign n952 = n951 ^ n947 ^ n274 ;
  assign n956 = n955 ^ n953 ^ n952 ;
  assign n957 = n655 & ~n956 ;
  assign n958 = n334 & n957 ;
  assign n946 = ~n495 & n840 ;
  assign n959 = n958 ^ n946 ^ 1'b0 ;
  assign n960 = n326 & ~n539 ;
  assign n961 = ~x93 & n960 ;
  assign n962 = ( ~x67 & n312 ) | ( ~x67 & n961 ) | ( n312 & n961 ) ;
  assign n963 = ( n553 & n575 ) | ( n553 & ~n962 ) | ( n575 & ~n962 ) ;
  assign n965 = x118 & ~n517 ;
  assign n966 = n371 & n965 ;
  assign n964 = x61 & n423 ;
  assign n967 = n966 ^ n964 ^ 1'b0 ;
  assign n968 = n967 ^ n649 ^ 1'b0 ;
  assign n969 = x163 | n944 ;
  assign n970 = n969 ^ n827 ^ n694 ;
  assign n972 = x196 & ~n444 ;
  assign n973 = n972 ^ x202 ^ 1'b0 ;
  assign n971 = ( n325 & n425 ) | ( n325 & n677 ) | ( n425 & n677 ) ;
  assign n974 = n973 ^ n971 ^ x254 ;
  assign n977 = ( x74 & ~x105 ) | ( x74 & n813 ) | ( ~x105 & n813 ) ;
  assign n978 = n548 | n977 ;
  assign n975 = x83 ^ x16 ^ 1'b0 ;
  assign n976 = x162 & ~n975 ;
  assign n979 = n978 ^ n976 ^ 1'b0 ;
  assign n1003 = n393 ^ x242 ^ x189 ;
  assign n1004 = n1003 ^ x31 ^ 1'b0 ;
  assign n1005 = ~n575 & n1004 ;
  assign n1000 = n614 ^ x160 ^ x40 ;
  assign n1001 = n494 ^ n470 ^ x250 ;
  assign n1002 = ( x57 & n1000 ) | ( x57 & ~n1001 ) | ( n1000 & ~n1001 ) ;
  assign n1006 = n1005 ^ n1002 ^ n349 ;
  assign n998 = n278 ^ x235 ^ 1'b0 ;
  assign n999 = ~n576 & n998 ;
  assign n981 = n537 ^ n444 ^ n360 ;
  assign n980 = x45 & x152 ;
  assign n982 = n981 ^ n980 ^ 1'b0 ;
  assign n983 = n982 ^ n353 ^ x69 ;
  assign n984 = ( x192 & n382 ) | ( x192 & ~n793 ) | ( n382 & ~n793 ) ;
  assign n985 = x160 & ~n984 ;
  assign n986 = n342 & n985 ;
  assign n987 = n986 ^ n684 ^ n603 ;
  assign n988 = ( ~x47 & n795 ) | ( ~x47 & n987 ) | ( n795 & n987 ) ;
  assign n993 = ( n527 & n559 ) | ( n527 & n948 ) | ( n559 & n948 ) ;
  assign n989 = ~x141 & x239 ;
  assign n990 = n989 ^ n349 ^ 1'b0 ;
  assign n991 = ~n452 & n990 ;
  assign n992 = ( n332 & n473 ) | ( n332 & ~n991 ) | ( n473 & ~n991 ) ;
  assign n994 = n993 ^ n992 ^ 1'b0 ;
  assign n995 = ( ~x206 & n988 ) | ( ~x206 & n994 ) | ( n988 & n994 ) ;
  assign n996 = ~n349 & n995 ;
  assign n997 = ~n983 & n996 ;
  assign n1007 = n1006 ^ n999 ^ n997 ;
  assign n1008 = x133 & n1006 ;
  assign n1009 = ~n287 & n1008 ;
  assign n1010 = x165 ^ x68 ^ 1'b0 ;
  assign n1011 = x119 & n1010 ;
  assign n1012 = n1011 ^ n805 ^ n375 ;
  assign n1013 = n657 ^ n471 ^ 1'b0 ;
  assign n1014 = n1012 & ~n1013 ;
  assign n1016 = ( x180 & n302 ) | ( x180 & n412 ) | ( n302 & n412 ) ;
  assign n1015 = n984 ^ x182 ^ 1'b0 ;
  assign n1017 = n1016 ^ n1015 ^ n645 ;
  assign n1018 = n1017 ^ x211 ^ x20 ;
  assign n1019 = ( x9 & ~n321 ) | ( x9 & n614 ) | ( ~n321 & n614 ) ;
  assign n1020 = n1019 ^ n312 ^ x9 ;
  assign n1021 = n500 & n1020 ;
  assign n1022 = n626 & n1021 ;
  assign n1023 = ( x110 & x222 ) | ( x110 & n313 ) | ( x222 & n313 ) ;
  assign n1024 = ( x53 & n795 ) | ( x53 & ~n1023 ) | ( n795 & ~n1023 ) ;
  assign n1025 = x49 & ~n1024 ;
  assign n1026 = ( ~n331 & n882 ) | ( ~n331 & n1025 ) | ( n882 & n1025 ) ;
  assign n1027 = n948 ^ n755 ^ x155 ;
  assign n1028 = n1027 ^ n801 ^ 1'b0 ;
  assign n1029 = n1028 ^ n345 ^ x115 ;
  assign n1030 = n418 ^ x71 ^ 1'b0 ;
  assign n1031 = n286 & ~n1030 ;
  assign n1032 = n678 & ~n1031 ;
  assign n1033 = n578 ^ x187 ^ x3 ;
  assign n1034 = n724 ^ x246 ^ 1'b0 ;
  assign n1035 = n1002 ^ x227 ^ x150 ;
  assign n1036 = n282 & ~n1035 ;
  assign n1037 = ~n532 & n1036 ;
  assign n1038 = n1037 ^ n492 ^ n431 ;
  assign n1039 = n1038 ^ n341 ^ x245 ;
  assign n1040 = x223 ^ x74 ^ 1'b0 ;
  assign n1041 = n582 ^ n571 ^ x186 ;
  assign n1042 = ( ~x156 & x248 ) | ( ~x156 & n1041 ) | ( x248 & n1041 ) ;
  assign n1043 = x227 ^ x25 ^ 1'b0 ;
  assign n1044 = ~n1042 & n1043 ;
  assign n1045 = n1040 & n1044 ;
  assign n1046 = n901 & n1045 ;
  assign n1047 = n1046 ^ n1007 ^ n820 ;
  assign n1051 = x62 & n438 ;
  assign n1052 = ~x9 & n1051 ;
  assign n1053 = n1052 ^ x210 ^ 1'b0 ;
  assign n1054 = n894 | n1053 ;
  assign n1050 = n907 ^ n640 ^ x199 ;
  assign n1055 = n1054 ^ n1050 ^ n393 ;
  assign n1056 = ( x108 & ~n756 ) | ( x108 & n1055 ) | ( ~n756 & n1055 ) ;
  assign n1048 = n433 ^ n273 ^ x26 ;
  assign n1049 = x204 & n1048 ;
  assign n1057 = n1056 ^ n1049 ^ 1'b0 ;
  assign n1060 = n989 ^ x9 ^ 1'b0 ;
  assign n1061 = x161 ^ x63 ^ x46 ;
  assign n1062 = ( x54 & n320 ) | ( x54 & n1061 ) | ( n320 & n1061 ) ;
  assign n1063 = ( ~n257 & n1060 ) | ( ~n257 & n1062 ) | ( n1060 & n1062 ) ;
  assign n1064 = ( x218 & ~n507 ) | ( x218 & n877 ) | ( ~n507 & n877 ) ;
  assign n1065 = n1064 ^ n334 ^ 1'b0 ;
  assign n1066 = n1063 | n1065 ;
  assign n1058 = n371 ^ x144 ^ x91 ;
  assign n1059 = x88 & n1058 ;
  assign n1067 = n1066 ^ n1059 ^ 1'b0 ;
  assign n1068 = ( x9 & ~x166 ) | ( x9 & n264 ) | ( ~x166 & n264 ) ;
  assign n1069 = ~n831 & n1068 ;
  assign n1070 = n1069 ^ n459 ^ 1'b0 ;
  assign n1071 = ~x143 & n1070 ;
  assign n1072 = ( ~x106 & x146 ) | ( ~x106 & n665 ) | ( x146 & n665 ) ;
  assign n1073 = ~x146 & n1072 ;
  assign n1074 = ~x16 & n1073 ;
  assign n1075 = x135 & n328 ;
  assign n1076 = n1074 & n1075 ;
  assign n1077 = n831 ^ n424 ^ x232 ;
  assign n1078 = ( x223 & n385 ) | ( x223 & n1077 ) | ( n385 & n1077 ) ;
  assign n1079 = ( ~x34 & n433 ) | ( ~x34 & n1061 ) | ( n433 & n1061 ) ;
  assign n1080 = n1079 ^ n672 ^ x197 ;
  assign n1081 = ~n858 & n903 ;
  assign n1082 = n1081 ^ n597 ^ 1'b0 ;
  assign n1083 = x13 & ~n372 ;
  assign n1084 = ~n407 & n1083 ;
  assign n1085 = n1084 ^ n406 ^ x67 ;
  assign n1086 = n859 & ~n1085 ;
  assign n1087 = n1086 ^ n485 ^ 1'b0 ;
  assign n1088 = n1082 | n1087 ;
  assign n1089 = n337 ^ x116 ^ 1'b0 ;
  assign n1090 = ~n345 & n1089 ;
  assign n1091 = n1090 ^ x151 ^ 1'b0 ;
  assign n1092 = n278 ^ x129 ^ 1'b0 ;
  assign n1093 = n1091 & n1092 ;
  assign n1094 = x29 & x164 ;
  assign n1095 = ~n1093 & n1094 ;
  assign n1099 = ( x5 & ~x138 ) | ( x5 & n268 ) | ( ~x138 & n268 ) ;
  assign n1100 = ( ~x6 & x44 ) | ( ~x6 & n1099 ) | ( x44 & n1099 ) ;
  assign n1097 = x24 & n594 ;
  assign n1096 = n1037 ^ n1019 ^ 1'b0 ;
  assign n1098 = n1097 ^ n1096 ^ n639 ;
  assign n1101 = n1100 ^ n1098 ^ n523 ;
  assign n1102 = ( x91 & x183 ) | ( x91 & ~n1101 ) | ( x183 & ~n1101 ) ;
  assign n1103 = n885 ^ x253 ^ 1'b0 ;
  assign n1104 = n895 & ~n1103 ;
  assign n1105 = n630 & n1104 ;
  assign n1106 = n1038 & n1105 ;
  assign n1107 = ( x94 & x101 ) | ( x94 & n579 ) | ( x101 & n579 ) ;
  assign n1108 = n1107 ^ n1052 ^ n486 ;
  assign n1109 = x201 & n1108 ;
  assign n1113 = ( x196 & n389 ) | ( x196 & ~n604 ) | ( n389 & ~n604 ) ;
  assign n1111 = n358 ^ x224 ^ x24 ;
  assign n1112 = n1111 ^ n887 ^ n843 ;
  assign n1110 = ( n415 & n643 ) | ( n415 & n969 ) | ( n643 & n969 ) ;
  assign n1114 = n1113 ^ n1112 ^ n1110 ;
  assign n1115 = n572 ^ x193 ^ 1'b0 ;
  assign n1116 = n1115 ^ n371 ^ n304 ;
  assign n1117 = ( x92 & n298 ) | ( x92 & n1011 ) | ( n298 & n1011 ) ;
  assign n1118 = ( ~x252 & n414 ) | ( ~x252 & n1117 ) | ( n414 & n1117 ) ;
  assign n1123 = x187 ^ x68 ^ x61 ;
  assign n1124 = n1123 ^ n650 ^ n298 ;
  assign n1119 = ( ~x216 & n833 ) | ( ~x216 & n854 ) | ( n833 & n854 ) ;
  assign n1120 = ( n740 & n794 ) | ( n740 & ~n1119 ) | ( n794 & ~n1119 ) ;
  assign n1121 = n425 | n1120 ;
  assign n1122 = n540 & ~n1121 ;
  assign n1125 = n1124 ^ n1122 ^ n817 ;
  assign n1126 = ( n1116 & ~n1118 ) | ( n1116 & n1125 ) | ( ~n1118 & n1125 ) ;
  assign n1127 = n1095 ^ n931 ^ 1'b0 ;
  assign n1128 = x108 ^ x70 ^ 1'b0 ;
  assign n1129 = x197 & n1128 ;
  assign n1130 = n494 | n678 ;
  assign n1131 = ( n581 & ~n1129 ) | ( n581 & n1130 ) | ( ~n1129 & n1130 ) ;
  assign n1132 = n955 ^ n494 ^ x242 ;
  assign n1133 = ( x97 & ~n1131 ) | ( x97 & n1132 ) | ( ~n1131 & n1132 ) ;
  assign n1134 = n978 & ~n1133 ;
  assign n1135 = x104 & ~x227 ;
  assign n1136 = n535 & ~n1016 ;
  assign n1137 = n811 ^ n279 ^ 1'b0 ;
  assign n1141 = ( x9 & n344 ) | ( x9 & n716 ) | ( n344 & n716 ) ;
  assign n1138 = n400 ^ n320 ^ 1'b0 ;
  assign n1139 = x103 & ~n1138 ;
  assign n1140 = ( n327 & n355 ) | ( n327 & n1139 ) | ( n355 & n1139 ) ;
  assign n1142 = n1141 ^ n1140 ^ n961 ;
  assign n1143 = ( x175 & n1137 ) | ( x175 & ~n1142 ) | ( n1137 & ~n1142 ) ;
  assign n1144 = ~x4 & n444 ;
  assign n1145 = n1139 ^ x186 ^ 1'b0 ;
  assign n1146 = n321 & n1145 ;
  assign n1147 = ( ~n462 & n1144 ) | ( ~n462 & n1146 ) | ( n1144 & n1146 ) ;
  assign n1148 = n903 & n1147 ;
  assign n1149 = n1148 ^ n1117 ^ 1'b0 ;
  assign n1150 = x142 & ~n680 ;
  assign n1151 = n1150 ^ n449 ^ 1'b0 ;
  assign n1152 = ( ~n390 & n997 ) | ( ~n390 & n1151 ) | ( n997 & n1151 ) ;
  assign n1153 = n383 & ~n1016 ;
  assign n1154 = x245 ^ x156 ^ x28 ;
  assign n1155 = n1154 ^ n1130 ^ 1'b0 ;
  assign n1156 = ( ~x179 & n1153 ) | ( ~x179 & n1155 ) | ( n1153 & n1155 ) ;
  assign n1157 = x227 | n1156 ;
  assign n1158 = x130 | n1157 ;
  assign n1159 = n1158 ^ n647 ^ 1'b0 ;
  assign n1160 = x18 & x32 ;
  assign n1161 = n1160 ^ x233 ^ 1'b0 ;
  assign n1162 = x158 ^ x52 ^ 1'b0 ;
  assign n1163 = n1162 ^ n795 ^ 1'b0 ;
  assign n1164 = ~n1161 & n1163 ;
  assign n1167 = ( x38 & x239 ) | ( x38 & n1019 ) | ( x239 & n1019 ) ;
  assign n1168 = n1167 ^ x232 ^ x186 ;
  assign n1165 = n399 ^ x85 ^ 1'b0 ;
  assign n1166 = n353 & n1165 ;
  assign n1169 = n1168 ^ n1166 ^ 1'b0 ;
  assign n1174 = x65 & n784 ;
  assign n1175 = ~n640 & n1174 ;
  assign n1176 = n394 ^ n321 ^ 1'b0 ;
  assign n1177 = ~n1175 & n1176 ;
  assign n1171 = n891 ^ n599 ^ 1'b0 ;
  assign n1172 = ~n364 & n1171 ;
  assign n1170 = n944 ^ n731 ^ x118 ;
  assign n1173 = n1172 ^ n1170 ^ x107 ;
  assign n1178 = n1177 ^ n1173 ^ 1'b0 ;
  assign n1179 = n1169 & ~n1178 ;
  assign n1180 = ( x34 & n919 ) | ( x34 & ~n1107 ) | ( n919 & ~n1107 ) ;
  assign n1181 = ( ~x130 & x171 ) | ( ~x130 & n320 ) | ( x171 & n320 ) ;
  assign n1182 = n1181 ^ x127 ^ 1'b0 ;
  assign n1183 = ( ~x147 & n333 ) | ( ~x147 & n1117 ) | ( n333 & n1117 ) ;
  assign n1184 = n425 ^ x134 ^ x3 ;
  assign n1185 = ( x6 & x170 ) | ( x6 & ~n571 ) | ( x170 & ~n571 ) ;
  assign n1186 = ( n283 & ~n1184 ) | ( n283 & n1185 ) | ( ~n1184 & n1185 ) ;
  assign n1187 = ~n777 & n1186 ;
  assign n1188 = n1183 & n1187 ;
  assign n1189 = ( x38 & ~x122 ) | ( x38 & n408 ) | ( ~x122 & n408 ) ;
  assign n1190 = n401 & n1189 ;
  assign n1191 = n1190 ^ n659 ^ 1'b0 ;
  assign n1192 = ( x198 & ~n1188 ) | ( x198 & n1191 ) | ( ~n1188 & n1191 ) ;
  assign n1193 = ~n684 & n1192 ;
  assign n1194 = n930 & n1193 ;
  assign n1195 = ( x45 & n600 ) | ( x45 & ~n738 ) | ( n600 & ~n738 ) ;
  assign n1196 = n856 | n1042 ;
  assign n1197 = ( ~n315 & n1023 ) | ( ~n315 & n1196 ) | ( n1023 & n1196 ) ;
  assign n1198 = n1195 & n1197 ;
  assign n1199 = x8 & ~n329 ;
  assign n1200 = n1199 ^ n313 ^ 1'b0 ;
  assign n1201 = ( n756 & ~n896 ) | ( n756 & n1200 ) | ( ~n896 & n1200 ) ;
  assign n1202 = x147 ^ x126 ^ x52 ;
  assign n1203 = x217 & ~n1202 ;
  assign n1204 = n469 & n1203 ;
  assign n1205 = ( x3 & ~x110 ) | ( x3 & n348 ) | ( ~x110 & n348 ) ;
  assign n1206 = n1205 ^ n684 ^ x78 ;
  assign n1207 = n872 ^ x227 ^ 1'b0 ;
  assign n1208 = n1207 ^ n1096 ^ n975 ;
  assign n1209 = ( x247 & n365 ) | ( x247 & ~n505 ) | ( n365 & ~n505 ) ;
  assign n1210 = n827 ^ n298 ^ x202 ;
  assign n1211 = n868 ^ n582 ^ x10 ;
  assign n1212 = n1211 ^ n991 ^ n321 ;
  assign n1213 = n1212 ^ n628 ^ n414 ;
  assign n1214 = ( n1209 & n1210 ) | ( n1209 & ~n1213 ) | ( n1210 & ~n1213 ) ;
  assign n1215 = ( x73 & ~n542 ) | ( x73 & n1011 ) | ( ~n542 & n1011 ) ;
  assign n1216 = n1215 ^ n612 ^ 1'b0 ;
  assign n1217 = n656 | n1216 ;
  assign n1218 = n1168 ^ n829 ^ x78 ;
  assign n1219 = ( n529 & ~n1217 ) | ( n529 & n1218 ) | ( ~n1217 & n1218 ) ;
  assign n1226 = ( x43 & x114 ) | ( x43 & n302 ) | ( x114 & n302 ) ;
  assign n1224 = n1019 ^ n474 ^ x227 ;
  assign n1221 = n598 ^ n378 ^ 1'b0 ;
  assign n1222 = ( x250 & ~n263 ) | ( x250 & n1221 ) | ( ~n263 & n1221 ) ;
  assign n1223 = n1222 ^ x162 ^ 1'b0 ;
  assign n1225 = n1224 ^ n1223 ^ n1188 ;
  assign n1220 = x160 & ~n920 ;
  assign n1227 = n1226 ^ n1225 ^ n1220 ;
  assign n1229 = ~n515 & n768 ;
  assign n1228 = x0 & n390 ;
  assign n1230 = n1229 ^ n1228 ^ 1'b0 ;
  assign n1231 = n1014 ^ n410 ^ n401 ;
  assign n1232 = n830 ^ n324 ^ 1'b0 ;
  assign n1233 = ~n1231 & n1232 ;
  assign n1239 = n405 | n1015 ;
  assign n1240 = n270 & ~n1239 ;
  assign n1236 = ( x26 & ~n299 ) | ( x26 & n825 ) | ( ~n299 & n825 ) ;
  assign n1234 = ~n478 & n705 ;
  assign n1235 = ~x131 & n1234 ;
  assign n1237 = n1236 ^ n1235 ^ n647 ;
  assign n1238 = ( ~x38 & n803 ) | ( ~x38 & n1237 ) | ( n803 & n1237 ) ;
  assign n1241 = n1240 ^ n1238 ^ n1232 ;
  assign n1242 = n261 ^ x119 ^ x27 ;
  assign n1243 = n835 & ~n1202 ;
  assign n1244 = ( n615 & n1242 ) | ( n615 & ~n1243 ) | ( n1242 & ~n1243 ) ;
  assign n1245 = n1244 ^ n640 ^ n619 ;
  assign n1246 = x138 ^ x116 ^ x107 ;
  assign n1247 = ( n560 & n1112 ) | ( n560 & n1246 ) | ( n1112 & n1246 ) ;
  assign n1249 = n1161 ^ x242 ^ 1'b0 ;
  assign n1250 = x8 & ~n1249 ;
  assign n1248 = ( ~x16 & x45 ) | ( ~x16 & x47 ) | ( x45 & x47 ) ;
  assign n1251 = n1250 ^ n1248 ^ n423 ;
  assign n1252 = ( x32 & n379 ) | ( x32 & ~n891 ) | ( n379 & ~n891 ) ;
  assign n1253 = x118 & ~n488 ;
  assign n1254 = ~n1252 & n1253 ;
  assign n1255 = n1251 | n1254 ;
  assign n1256 = n1255 ^ x201 ^ 1'b0 ;
  assign n1257 = n591 ^ n312 ^ x106 ;
  assign n1260 = n808 ^ n412 ^ n298 ;
  assign n1258 = n641 ^ n631 ^ x246 ;
  assign n1259 = n429 & ~n1258 ;
  assign n1261 = n1260 ^ n1259 ^ 1'b0 ;
  assign n1262 = n1261 ^ n332 ^ n280 ;
  assign n1263 = n1257 & ~n1262 ;
  assign n1264 = n1263 ^ x190 ^ 1'b0 ;
  assign n1265 = ( x120 & n857 ) | ( x120 & n1003 ) | ( n857 & n1003 ) ;
  assign n1267 = n891 ^ n691 ^ x112 ;
  assign n1266 = ( ~n421 & n594 ) | ( ~n421 & n883 ) | ( n594 & n883 ) ;
  assign n1268 = n1267 ^ n1266 ^ n404 ;
  assign n1269 = x124 ^ x96 ^ x71 ;
  assign n1270 = n1269 ^ x176 ^ 1'b0 ;
  assign n1271 = n1064 & ~n1270 ;
  assign n1272 = n1271 ^ n822 ^ 1'b0 ;
  assign n1275 = ~n295 & n597 ;
  assign n1276 = ~n1243 & n1275 ;
  assign n1273 = n556 ^ n542 ^ x156 ;
  assign n1274 = ( n803 & n966 ) | ( n803 & ~n1273 ) | ( n966 & ~n1273 ) ;
  assign n1277 = n1276 ^ n1274 ^ 1'b0 ;
  assign n1278 = n594 & ~n1277 ;
  assign n1279 = n1278 ^ n375 ^ x47 ;
  assign n1280 = n691 ^ x172 ^ x146 ;
  assign n1281 = n1280 ^ n1090 ^ 1'b0 ;
  assign n1282 = x80 & ~n1281 ;
  assign n1283 = ( ~x102 & n488 ) | ( ~x102 & n1282 ) | ( n488 & n1282 ) ;
  assign n1284 = ( x44 & ~x131 ) | ( x44 & n1283 ) | ( ~x131 & n1283 ) ;
  assign n1285 = n758 ^ n598 ^ x43 ;
  assign n1286 = n1285 ^ n1044 ^ 1'b0 ;
  assign n1287 = n391 | n1286 ;
  assign n1288 = x45 | n1287 ;
  assign n1289 = n346 & n1288 ;
  assign n1290 = n1284 & n1289 ;
  assign n1291 = n1172 ^ n1108 ^ n708 ;
  assign n1296 = ( n516 & ~n763 ) | ( n516 & n993 ) | ( ~n763 & n993 ) ;
  assign n1295 = n969 ^ x146 ^ 1'b0 ;
  assign n1292 = ( n484 & n576 ) | ( n484 & ~n881 ) | ( n576 & ~n881 ) ;
  assign n1293 = ( n691 & ~n882 ) | ( n691 & n1292 ) | ( ~n882 & n1292 ) ;
  assign n1294 = ( ~x49 & n594 ) | ( ~x49 & n1293 ) | ( n594 & n1293 ) ;
  assign n1297 = n1296 ^ n1295 ^ n1294 ;
  assign n1314 = x208 & ~n270 ;
  assign n1315 = ~n320 & n1314 ;
  assign n1310 = n1260 ^ n910 ^ n547 ;
  assign n1311 = n749 & ~n1310 ;
  assign n1312 = n1311 ^ n414 ^ 1'b0 ;
  assign n1306 = n754 ^ x200 ^ x142 ;
  assign n1307 = ( ~n608 & n772 ) | ( ~n608 & n1306 ) | ( n772 & n1306 ) ;
  assign n1308 = ( x45 & n327 ) | ( x45 & n1307 ) | ( n327 & n1307 ) ;
  assign n1309 = ( ~x248 & n1141 ) | ( ~x248 & n1308 ) | ( n1141 & n1308 ) ;
  assign n1313 = n1312 ^ n1309 ^ n845 ;
  assign n1301 = n369 ^ x37 ^ 1'b0 ;
  assign n1302 = n1301 ^ x252 ^ 1'b0 ;
  assign n1303 = n696 ^ n541 ^ 1'b0 ;
  assign n1304 = n1302 & n1303 ;
  assign n1298 = ( ~x46 & x212 ) | ( ~x46 & n687 ) | ( x212 & n687 ) ;
  assign n1299 = x50 & ~n632 ;
  assign n1300 = n1298 & n1299 ;
  assign n1305 = n1304 ^ n1300 ^ 1'b0 ;
  assign n1316 = n1315 ^ n1313 ^ n1305 ;
  assign n1317 = n860 ^ n552 ^ x203 ;
  assign n1318 = n1317 ^ x109 ^ 1'b0 ;
  assign n1319 = n1186 & ~n1318 ;
  assign n1320 = n1319 ^ n326 ^ x34 ;
  assign n1321 = ( n275 & n365 ) | ( n275 & ~n1320 ) | ( n365 & ~n1320 ) ;
  assign n1322 = n1254 ^ n604 ^ x14 ;
  assign n1323 = n1236 ^ n1003 ^ 1'b0 ;
  assign n1335 = x120 & x121 ;
  assign n1336 = n1335 ^ x80 ^ 1'b0 ;
  assign n1337 = n1336 ^ x157 ^ 1'b0 ;
  assign n1331 = x162 ^ x145 ^ x126 ;
  assign n1332 = x67 & n450 ;
  assign n1333 = n1332 ^ n573 ^ 1'b0 ;
  assign n1334 = n1331 | n1333 ;
  assign n1338 = n1337 ^ n1334 ^ n1060 ;
  assign n1326 = ( x46 & x151 ) | ( x46 & ~x210 ) | ( x151 & ~x210 ) ;
  assign n1327 = n715 ^ n710 ^ x127 ;
  assign n1328 = n1326 & n1327 ;
  assign n1329 = ~n950 & n1328 ;
  assign n1330 = n1329 ^ n617 ^ x87 ;
  assign n1324 = n1261 ^ n1096 ^ x235 ;
  assign n1325 = n1324 ^ n1099 ^ n438 ;
  assign n1339 = n1338 ^ n1330 ^ n1325 ;
  assign n1350 = ( ~x181 & n350 ) | ( ~x181 & n981 ) | ( n350 & n981 ) ;
  assign n1351 = ( ~x23 & n330 ) | ( ~x23 & n1350 ) | ( n330 & n1350 ) ;
  assign n1340 = n295 ^ x203 ^ x68 ;
  assign n1341 = n1189 ^ n507 ^ n396 ;
  assign n1342 = n759 & ~n1341 ;
  assign n1343 = ~n1340 & n1342 ;
  assign n1344 = n863 ^ n785 ^ n687 ;
  assign n1345 = n864 ^ n368 ^ 1'b0 ;
  assign n1346 = n1344 & n1345 ;
  assign n1347 = n1346 ^ n446 ^ x160 ;
  assign n1348 = n587 | n1347 ;
  assign n1349 = n1343 & ~n1348 ;
  assign n1352 = n1351 ^ n1349 ^ x231 ;
  assign n1356 = ( n805 & ~n896 ) | ( n805 & n1350 ) | ( ~n896 & n1350 ) ;
  assign n1353 = x218 & n532 ;
  assign n1354 = n376 & n1353 ;
  assign n1355 = n1354 ^ x113 ^ 1'b0 ;
  assign n1357 = n1356 ^ n1355 ^ x155 ;
  assign n1358 = ( x206 & ~n794 ) | ( x206 & n973 ) | ( ~n794 & n973 ) ;
  assign n1359 = ( x101 & ~n913 ) | ( x101 & n1358 ) | ( ~n913 & n1358 ) ;
  assign n1361 = x191 | n977 ;
  assign n1360 = n955 ^ n691 ^ x163 ;
  assign n1362 = n1361 ^ n1360 ^ n570 ;
  assign n1365 = ( x55 & ~x106 ) | ( x55 & x236 ) | ( ~x106 & x236 ) ;
  assign n1366 = ( n300 & ~n390 ) | ( n300 & n1365 ) | ( ~n390 & n1365 ) ;
  assign n1363 = x56 ^ x55 ^ 1'b0 ;
  assign n1364 = n944 & ~n1363 ;
  assign n1367 = n1366 ^ n1364 ^ 1'b0 ;
  assign n1368 = n910 ^ x170 ^ x140 ;
  assign n1369 = n341 | n1368 ;
  assign n1373 = n1100 ^ n652 ^ n332 ;
  assign n1374 = n367 & n1373 ;
  assign n1375 = ~n344 & n1374 ;
  assign n1370 = x2 & ~n1218 ;
  assign n1371 = n973 & n1370 ;
  assign n1372 = n1371 ^ n1012 ^ 1'b0 ;
  assign n1376 = n1375 ^ n1372 ^ n580 ;
  assign n1377 = n1006 ^ n339 ^ 1'b0 ;
  assign n1378 = ~n1029 & n1377 ;
  assign n1379 = n1378 ^ n655 ^ 1'b0 ;
  assign n1380 = ( x219 & ~n398 ) | ( x219 & n485 ) | ( ~n398 & n485 ) ;
  assign n1381 = n1380 ^ n1260 ^ n511 ;
  assign n1382 = x190 ^ x103 ^ 1'b0 ;
  assign n1383 = ( x253 & n1381 ) | ( x253 & ~n1382 ) | ( n1381 & ~n1382 ) ;
  assign n1384 = x125 & ~n520 ;
  assign n1385 = n1384 ^ n1002 ^ n414 ;
  assign n1386 = n895 & ~n1385 ;
  assign n1387 = n1386 ^ n453 ^ 1'b0 ;
  assign n1388 = ~n1349 & n1387 ;
  assign n1389 = ~n1383 & n1388 ;
  assign n1390 = n1308 ^ n747 ^ x209 ;
  assign n1391 = ( x47 & ~x217 ) | ( x47 & n1285 ) | ( ~x217 & n1285 ) ;
  assign n1392 = n579 ^ n269 ^ x176 ;
  assign n1393 = n647 & n1392 ;
  assign n1394 = n1393 ^ n1344 ^ 1'b0 ;
  assign n1395 = n1391 | n1394 ;
  assign n1396 = n910 | n1202 ;
  assign n1397 = n1396 ^ n301 ^ 1'b0 ;
  assign n1398 = n951 ^ x148 ^ 1'b0 ;
  assign n1399 = ( x239 & n1397 ) | ( x239 & n1398 ) | ( n1397 & n1398 ) ;
  assign n1400 = ( n818 & n1395 ) | ( n818 & n1399 ) | ( n1395 & n1399 ) ;
  assign n1401 = n1400 ^ n1242 ^ 1'b0 ;
  assign n1402 = ( n430 & ~n599 ) | ( n430 & n602 ) | ( ~n599 & n602 ) ;
  assign n1403 = n1402 ^ n858 ^ n503 ;
  assign n1404 = n1403 ^ n488 ^ 1'b0 ;
  assign n1405 = n602 & n635 ;
  assign n1406 = ( ~n325 & n1299 ) | ( ~n325 & n1405 ) | ( n1299 & n1405 ) ;
  assign n1407 = n1406 ^ n744 ^ n667 ;
  assign n1408 = ~n829 & n1407 ;
  assign n1409 = n1408 ^ n1326 ^ n681 ;
  assign n1411 = x205 ^ x107 ^ 1'b0 ;
  assign n1412 = x70 & n1411 ;
  assign n1414 = ( x91 & ~x220 ) | ( x91 & n1280 ) | ( ~x220 & n1280 ) ;
  assign n1413 = x141 & x249 ;
  assign n1415 = n1414 ^ n1413 ^ 1'b0 ;
  assign n1416 = n1412 & ~n1415 ;
  assign n1417 = ( n904 & n987 ) | ( n904 & ~n1416 ) | ( n987 & ~n1416 ) ;
  assign n1410 = n911 ^ x219 ^ 1'b0 ;
  assign n1418 = n1417 ^ n1410 ^ n1362 ;
  assign n1423 = n1002 ^ x242 ^ x236 ;
  assign n1422 = n1023 ^ n935 ^ 1'b0 ;
  assign n1419 = x1 & n628 ;
  assign n1420 = ( n522 & n1077 ) | ( n522 & n1419 ) | ( n1077 & n1419 ) ;
  assign n1421 = n1420 ^ n287 ^ x48 ;
  assign n1424 = n1423 ^ n1422 ^ n1421 ;
  assign n1425 = x251 & ~n471 ;
  assign n1426 = n645 ^ n358 ^ x123 ;
  assign n1427 = n1426 ^ n1146 ^ 1'b0 ;
  assign n1428 = x145 & ~n1427 ;
  assign n1429 = ( x81 & ~n387 ) | ( x81 & n700 ) | ( ~n387 & n700 ) ;
  assign n1430 = n1022 ^ x188 ^ 1'b0 ;
  assign n1431 = n626 | n1430 ;
  assign n1432 = n1429 & ~n1431 ;
  assign n1433 = n1432 ^ n971 ^ 1'b0 ;
  assign n1434 = ( ~n462 & n1223 ) | ( ~n462 & n1265 ) | ( n1223 & n1265 ) ;
  assign n1435 = n1108 ^ n707 ^ x4 ;
  assign n1436 = n1189 ^ n866 ^ x82 ;
  assign n1437 = ( ~x32 & n973 ) | ( ~x32 & n1302 ) | ( n973 & n1302 ) ;
  assign n1438 = n1437 ^ n1162 ^ x3 ;
  assign n1439 = ( n808 & n1436 ) | ( n808 & n1438 ) | ( n1436 & n1438 ) ;
  assign n1440 = ( ~n1195 & n1435 ) | ( ~n1195 & n1439 ) | ( n1435 & n1439 ) ;
  assign n1441 = n491 ^ n286 ^ 1'b0 ;
  assign n1442 = x14 & n1441 ;
  assign n1448 = n831 ^ x215 ^ 1'b0 ;
  assign n1449 = n1448 ^ n666 ^ n527 ;
  assign n1451 = x1 | n1108 ;
  assign n1450 = n430 & n988 ;
  assign n1452 = n1451 ^ n1450 ^ n754 ;
  assign n1453 = ( ~x116 & n1449 ) | ( ~x116 & n1452 ) | ( n1449 & n1452 ) ;
  assign n1454 = ( x10 & ~x128 ) | ( x10 & n1453 ) | ( ~x128 & n1453 ) ;
  assign n1447 = n419 & n1003 ;
  assign n1443 = ~n418 & n645 ;
  assign n1444 = ~n481 & n1443 ;
  assign n1445 = n1087 | n1444 ;
  assign n1446 = n1445 ^ n1063 ^ 1'b0 ;
  assign n1455 = n1454 ^ n1447 ^ n1446 ;
  assign n1456 = n1412 ^ n552 ^ x192 ;
  assign n1457 = x105 ^ x87 ^ x31 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = n1458 ^ x42 ^ 1'b0 ;
  assign n1460 = n858 ^ n732 ^ 1'b0 ;
  assign n1461 = n1460 ^ n1347 ^ n418 ;
  assign n1462 = n1459 & ~n1461 ;
  assign n1463 = n1462 ^ n1354 ^ 1'b0 ;
  assign n1464 = n1361 ^ n842 ^ n691 ;
  assign n1465 = n436 | n1464 ;
  assign n1468 = x31 & n582 ;
  assign n1469 = ~x230 & n1468 ;
  assign n1470 = n1469 ^ n488 ^ 1'b0 ;
  assign n1471 = x55 & ~n1470 ;
  assign n1466 = n517 ^ n458 ^ x113 ;
  assign n1467 = ( n343 & n562 ) | ( n343 & n1466 ) | ( n562 & n1466 ) ;
  assign n1472 = n1471 ^ n1467 ^ n566 ;
  assign n1473 = x99 & ~n1067 ;
  assign n1474 = x79 & n1473 ;
  assign n1475 = n781 ^ n369 ^ 1'b0 ;
  assign n1476 = ~n941 & n1475 ;
  assign n1477 = ( ~x250 & n296 ) | ( ~x250 & n1242 ) | ( n296 & n1242 ) ;
  assign n1478 = x245 & n1477 ;
  assign n1479 = n1478 ^ n573 ^ 1'b0 ;
  assign n1480 = ( x244 & n579 ) | ( x244 & n1479 ) | ( n579 & n1479 ) ;
  assign n1481 = n1218 ^ n1192 ^ n934 ;
  assign n1482 = n1481 ^ n1413 ^ 1'b0 ;
  assign n1483 = n1131 ^ x212 ^ 1'b0 ;
  assign n1484 = n997 | n1483 ;
  assign n1485 = ( x82 & n267 ) | ( x82 & ~n529 ) | ( n267 & ~n529 ) ;
  assign n1486 = n1485 ^ x139 ^ 1'b0 ;
  assign n1487 = n1484 & ~n1486 ;
  assign n1488 = n835 ^ n416 ^ x73 ;
  assign n1490 = ( ~x69 & x97 ) | ( ~x69 & n1147 ) | ( x97 & n1147 ) ;
  assign n1489 = x211 & n416 ;
  assign n1491 = n1490 ^ n1489 ^ 1'b0 ;
  assign n1492 = ( ~x245 & n1488 ) | ( ~x245 & n1491 ) | ( n1488 & n1491 ) ;
  assign n1497 = n270 & n548 ;
  assign n1493 = n667 & ~n1491 ;
  assign n1494 = n732 & ~n1493 ;
  assign n1495 = n1494 ^ n798 ^ 1'b0 ;
  assign n1496 = n1495 ^ n871 ^ n647 ;
  assign n1498 = n1497 ^ n1496 ^ n669 ;
  assign n1499 = x206 ^ x179 ^ x9 ;
  assign n1500 = ( n344 & ~n993 ) | ( n344 & n1499 ) | ( ~n993 & n1499 ) ;
  assign n1501 = x186 & n1130 ;
  assign n1502 = n1501 ^ n420 ^ 1'b0 ;
  assign n1503 = ( ~x175 & n394 ) | ( ~x175 & n842 ) | ( n394 & n842 ) ;
  assign n1504 = n808 ^ n363 ^ 1'b0 ;
  assign n1505 = n716 & n904 ;
  assign n1506 = n374 & ~n1505 ;
  assign n1507 = n1506 ^ n725 ^ 1'b0 ;
  assign n1508 = ( n659 & ~n1504 ) | ( n659 & n1507 ) | ( ~n1504 & n1507 ) ;
  assign n1509 = ( n599 & ~n853 ) | ( n599 & n1508 ) | ( ~n853 & n1508 ) ;
  assign n1510 = n1503 & n1509 ;
  assign n1511 = ( ~n1500 & n1502 ) | ( ~n1500 & n1510 ) | ( n1502 & n1510 ) ;
  assign n1512 = x81 & n1107 ;
  assign n1513 = ~x71 & n1512 ;
  assign n1514 = n1513 ^ n1217 ^ 1'b0 ;
  assign n1515 = n565 ^ x223 ^ x156 ;
  assign n1516 = n1515 ^ n984 ^ n875 ;
  assign n1517 = n1516 ^ n829 ^ x94 ;
  assign n1518 = n1471 ^ n740 ^ n487 ;
  assign n1519 = ( ~n562 & n1236 ) | ( ~n562 & n1518 ) | ( n1236 & n1518 ) ;
  assign n1527 = ( ~x74 & n524 ) | ( ~x74 & n1392 ) | ( n524 & n1392 ) ;
  assign n1521 = x223 ^ x199 ^ x0 ;
  assign n1522 = n418 ^ x164 ^ 1'b0 ;
  assign n1523 = n589 | n1522 ;
  assign n1524 = ( n1449 & ~n1521 ) | ( n1449 & n1523 ) | ( ~n1521 & n1523 ) ;
  assign n1520 = n1485 ^ n876 ^ n444 ;
  assign n1525 = n1524 ^ n1520 ^ 1'b0 ;
  assign n1526 = x1 & ~n1525 ;
  assign n1528 = n1527 ^ n1526 ^ n765 ;
  assign n1529 = n1528 ^ n1331 ^ x40 ;
  assign n1543 = x34 & n1477 ;
  assign n1544 = n1543 ^ n726 ^ 1'b0 ;
  assign n1545 = x201 & n306 ;
  assign n1546 = n1544 & n1545 ;
  assign n1547 = n1546 ^ n710 ^ 1'b0 ;
  assign n1548 = n726 & ~n1547 ;
  assign n1549 = n1129 & n1548 ;
  assign n1540 = x141 & n1297 ;
  assign n1541 = n1540 ^ n331 ^ 1'b0 ;
  assign n1542 = n1541 ^ n1410 ^ x224 ;
  assign n1530 = ( x63 & n597 ) | ( x63 & ~n969 ) | ( n597 & ~n969 ) ;
  assign n1534 = n796 ^ n553 ^ x195 ;
  assign n1531 = n441 ^ x48 ^ 1'b0 ;
  assign n1532 = n1504 | n1531 ;
  assign n1533 = n647 & ~n1532 ;
  assign n1535 = n1534 ^ n1533 ^ 1'b0 ;
  assign n1536 = ( x60 & n431 ) | ( x60 & ~n1285 ) | ( n431 & ~n1285 ) ;
  assign n1537 = n1536 ^ n941 ^ x160 ;
  assign n1538 = n1537 ^ n508 ^ 1'b0 ;
  assign n1539 = ( n1530 & n1535 ) | ( n1530 & ~n1538 ) | ( n1535 & ~n1538 ) ;
  assign n1550 = n1549 ^ n1542 ^ n1539 ;
  assign n1552 = n1315 ^ n541 ^ x216 ;
  assign n1553 = ( n614 & n1144 ) | ( n614 & n1552 ) | ( n1144 & n1552 ) ;
  assign n1551 = x42 & ~n901 ;
  assign n1554 = n1553 ^ n1551 ^ 1'b0 ;
  assign n1555 = ( x74 & ~n687 ) | ( x74 & n1554 ) | ( ~n687 & n1554 ) ;
  assign n1556 = ( n368 & ~n1266 ) | ( n368 & n1555 ) | ( ~n1266 & n1555 ) ;
  assign n1557 = x199 & n1139 ;
  assign n1558 = ~n1350 & n1557 ;
  assign n1559 = n1558 ^ n825 ^ x232 ;
  assign n1560 = n482 & n1559 ;
  assign n1569 = n545 ^ n358 ^ 1'b0 ;
  assign n1570 = n1569 ^ n883 ^ n333 ;
  assign n1561 = n1072 ^ n300 ^ x56 ;
  assign n1562 = ( ~x118 & n843 ) | ( ~x118 & n1091 ) | ( n843 & n1091 ) ;
  assign n1563 = n1561 & ~n1562 ;
  assign n1564 = n1563 ^ x42 ^ 1'b0 ;
  assign n1565 = n1564 ^ n1381 ^ n616 ;
  assign n1566 = n908 | n1200 ;
  assign n1567 = n1565 & ~n1566 ;
  assign n1568 = n1567 ^ x202 ^ 1'b0 ;
  assign n1571 = n1570 ^ n1568 ^ n346 ;
  assign n1572 = ( n873 & ~n1134 ) | ( n873 & n1217 ) | ( ~n1134 & n1217 ) ;
  assign n1573 = ( x16 & x182 ) | ( x16 & n716 ) | ( x182 & n716 ) ;
  assign n1574 = ( n396 & n1020 ) | ( n396 & ~n1573 ) | ( n1020 & ~n1573 ) ;
  assign n1575 = n1574 ^ n1265 ^ x132 ;
  assign n1576 = n1197 ^ n750 ^ n719 ;
  assign n1577 = n1576 ^ n548 ^ 1'b0 ;
  assign n1578 = n749 ^ x128 ^ 1'b0 ;
  assign n1579 = ( ~n529 & n1488 ) | ( ~n529 & n1578 ) | ( n1488 & n1578 ) ;
  assign n1580 = n1579 ^ n1197 ^ 1'b0 ;
  assign n1581 = n987 & ~n1580 ;
  assign n1584 = n854 & ~n1269 ;
  assign n1585 = n455 & n1584 ;
  assign n1586 = n1585 ^ n366 ^ x39 ;
  assign n1583 = n911 ^ x164 ^ 1'b0 ;
  assign n1587 = n1586 ^ n1583 ^ 1'b0 ;
  assign n1582 = n927 ^ x245 ^ x64 ;
  assign n1588 = n1587 ^ n1582 ^ 1'b0 ;
  assign n1589 = ( n366 & n1274 ) | ( n366 & ~n1346 ) | ( n1274 & ~n1346 ) ;
  assign n1590 = n916 ^ n547 ^ 1'b0 ;
  assign n1591 = n1267 ^ n953 ^ n868 ;
  assign n1592 = ( n829 & ~n1419 ) | ( n829 & n1591 ) | ( ~n1419 & n1591 ) ;
  assign n1593 = ( n1589 & ~n1590 ) | ( n1589 & n1592 ) | ( ~n1590 & n1592 ) ;
  assign n1594 = n1593 ^ n1552 ^ n901 ;
  assign n1595 = n886 ^ n607 ^ n605 ;
  assign n1596 = ( n368 & n603 ) | ( n368 & ~n908 ) | ( n603 & ~n908 ) ;
  assign n1597 = n1027 | n1596 ;
  assign n1598 = n1597 ^ n485 ^ 1'b0 ;
  assign n1599 = ( x48 & n273 ) | ( x48 & n1116 ) | ( n273 & n1116 ) ;
  assign n1600 = ( x130 & ~n368 ) | ( x130 & n573 ) | ( ~n368 & n573 ) ;
  assign n1601 = ( n643 & n835 ) | ( n643 & n1600 ) | ( n835 & n1600 ) ;
  assign n1602 = ( ~n997 & n1599 ) | ( ~n997 & n1601 ) | ( n1599 & n1601 ) ;
  assign n1603 = n608 ^ n311 ^ x47 ;
  assign n1604 = x235 & n1603 ;
  assign n1605 = n1285 | n1604 ;
  assign n1606 = x88 | n956 ;
  assign n1607 = ( n528 & n659 ) | ( n528 & n1606 ) | ( n659 & n1606 ) ;
  assign n1608 = x33 & n1607 ;
  assign n1609 = n1608 ^ n1237 ^ 1'b0 ;
  assign n1610 = ( ~n977 & n1211 ) | ( ~n977 & n1609 ) | ( n1211 & n1609 ) ;
  assign n1611 = ( x84 & n1184 ) | ( x84 & n1602 ) | ( n1184 & n1602 ) ;
  assign n1615 = n833 ^ n576 ^ 1'b0 ;
  assign n1616 = ~n641 & n1615 ;
  assign n1617 = n1616 ^ n1188 ^ 1'b0 ;
  assign n1618 = n903 & ~n1617 ;
  assign n1612 = n296 ^ x182 ^ 1'b0 ;
  assign n1613 = n1351 ^ n934 ^ 1'b0 ;
  assign n1614 = n1612 & ~n1613 ;
  assign n1619 = n1618 ^ n1614 ^ n1471 ;
  assign n1620 = n825 ^ n581 ^ n414 ;
  assign n1621 = x154 & ~n825 ;
  assign n1622 = n1620 & n1621 ;
  assign n1623 = n1405 ^ n441 ^ 1'b0 ;
  assign n1624 = ~n1622 & n1623 ;
  assign n1625 = n1619 & n1624 ;
  assign n1629 = ( x183 & x211 ) | ( x183 & n538 ) | ( x211 & n538 ) ;
  assign n1626 = n326 ^ x215 ^ x21 ;
  assign n1627 = n1626 ^ n1226 ^ n828 ;
  assign n1628 = n1627 ^ n1207 ^ 1'b0 ;
  assign n1630 = n1629 ^ n1628 ^ 1'b0 ;
  assign n1631 = n1143 | n1630 ;
  assign n1632 = n786 ^ x153 ^ x52 ;
  assign n1633 = ( x70 & ~n412 ) | ( x70 & n606 ) | ( ~n412 & n606 ) ;
  assign n1634 = x167 & ~n317 ;
  assign n1635 = ( ~n834 & n1633 ) | ( ~n834 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1636 = ( ~n983 & n1020 ) | ( ~n983 & n1635 ) | ( n1020 & n1635 ) ;
  assign n1637 = ( n1444 & n1632 ) | ( n1444 & ~n1636 ) | ( n1632 & ~n1636 ) ;
  assign n1638 = n1637 ^ n1484 ^ 1'b0 ;
  assign n1649 = ~x14 & x192 ;
  assign n1647 = n1116 ^ x242 ^ 1'b0 ;
  assign n1648 = n747 & ~n1647 ;
  assign n1650 = n1649 ^ n1648 ^ 1'b0 ;
  assign n1639 = n315 ^ n267 ^ x98 ;
  assign n1640 = n1070 ^ x230 ^ 1'b0 ;
  assign n1641 = ~n1639 & n1640 ;
  assign n1642 = n1641 ^ n773 ^ x135 ;
  assign n1643 = ~x185 & n1642 ;
  assign n1644 = n1620 ^ n1378 ^ 1'b0 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1646 = ~n978 & n1645 ;
  assign n1651 = n1650 ^ n1646 ^ n312 ;
  assign n1658 = n1111 ^ n953 ^ n887 ;
  assign n1657 = ( n405 & ~n665 ) | ( n405 & n1212 ) | ( ~n665 & n1212 ) ;
  assign n1652 = n350 ^ x240 ^ x204 ;
  assign n1653 = ( n636 & n1211 ) | ( n636 & ~n1652 ) | ( n1211 & ~n1652 ) ;
  assign n1654 = n895 & ~n1502 ;
  assign n1655 = n1654 ^ n1058 ^ 1'b0 ;
  assign n1656 = ( x225 & n1653 ) | ( x225 & n1655 ) | ( n1653 & n1655 ) ;
  assign n1659 = n1658 ^ n1657 ^ n1656 ;
  assign n1662 = n339 & n499 ;
  assign n1663 = ~n296 & n1662 ;
  assign n1660 = n1268 ^ x87 ^ 1'b0 ;
  assign n1661 = x121 & ~n1660 ;
  assign n1664 = n1663 ^ n1661 ^ 1'b0 ;
  assign n1665 = ( x205 & ~n760 ) | ( x205 & n768 ) | ( ~n760 & n768 ) ;
  assign n1666 = n1665 ^ x121 ^ x6 ;
  assign n1667 = n1477 ^ n1273 ^ 1'b0 ;
  assign n1668 = n1252 & ~n1667 ;
  assign n1669 = x227 & n1668 ;
  assign n1670 = n1015 & n1669 ;
  assign n1671 = n1670 ^ x121 ^ 1'b0 ;
  assign n1672 = n1666 & ~n1671 ;
  assign n1673 = n1041 ^ n524 ^ 1'b0 ;
  assign n1679 = ( n744 & n766 ) | ( n744 & n1015 ) | ( n766 & n1015 ) ;
  assign n1674 = ( n356 & n470 ) | ( n356 & n515 ) | ( n470 & n515 ) ;
  assign n1675 = n989 ^ n349 ^ n327 ;
  assign n1676 = ( n542 & ~n901 ) | ( n542 & n1675 ) | ( ~n901 & n1675 ) ;
  assign n1677 = ( x201 & ~n1674 ) | ( x201 & n1676 ) | ( ~n1674 & n1676 ) ;
  assign n1678 = ( x140 & ~n548 ) | ( x140 & n1677 ) | ( ~n548 & n1677 ) ;
  assign n1680 = n1679 ^ n1678 ^ 1'b0 ;
  assign n1681 = ( n269 & n794 ) | ( n269 & n1426 ) | ( n794 & n1426 ) ;
  assign n1682 = ( x50 & ~n397 ) | ( x50 & n955 ) | ( ~n397 & n955 ) ;
  assign n1683 = n1682 ^ n1011 ^ x88 ;
  assign n1684 = n296 & n450 ;
  assign n1685 = ~n927 & n1684 ;
  assign n1686 = n414 ^ n382 ^ n293 ;
  assign n1687 = n1117 ^ n373 ^ 1'b0 ;
  assign n1688 = x19 & n1687 ;
  assign n1689 = n490 | n1544 ;
  assign n1690 = ( ~n622 & n1688 ) | ( ~n622 & n1689 ) | ( n1688 & n1689 ) ;
  assign n1691 = ( n814 & n1686 ) | ( n814 & ~n1690 ) | ( n1686 & ~n1690 ) ;
  assign n1692 = n1691 ^ n349 ^ 1'b0 ;
  assign n1693 = n497 & ~n1692 ;
  assign n1694 = ( x143 & n1685 ) | ( x143 & n1693 ) | ( n1685 & n1693 ) ;
  assign n1695 = ( n409 & n1683 ) | ( n409 & ~n1694 ) | ( n1683 & ~n1694 ) ;
  assign n1696 = n589 ^ n396 ^ 1'b0 ;
  assign n1697 = x185 & ~n1696 ;
  assign n1698 = n1313 ^ x216 ^ 1'b0 ;
  assign n1699 = n1697 & ~n1698 ;
  assign n1700 = n1699 ^ n458 ^ 1'b0 ;
  assign n1701 = n785 ^ n336 ^ x96 ;
  assign n1702 = n1701 ^ n397 ^ x120 ;
  assign n1703 = n1702 ^ x225 ^ 1'b0 ;
  assign n1704 = x63 & n1703 ;
  assign n1705 = n1704 ^ n414 ^ 1'b0 ;
  assign n1706 = ~n1084 & n1705 ;
  assign n1707 = n507 ^ n436 ^ x217 ;
  assign n1708 = ( n420 & ~n1541 ) | ( n420 & n1707 ) | ( ~n1541 & n1707 ) ;
  assign n1709 = n1310 ^ n1154 ^ x25 ;
  assign n1710 = n1709 ^ n958 ^ n840 ;
  assign n1711 = n1710 ^ n720 ^ n503 ;
  assign n1712 = n1692 ^ n1093 ^ 1'b0 ;
  assign n1713 = n1712 ^ n1390 ^ n930 ;
  assign n1714 = n837 ^ x173 ^ x59 ;
  assign n1715 = n740 ^ n593 ^ 1'b0 ;
  assign n1716 = n1714 | n1715 ;
  assign n1717 = n1227 ^ n995 ^ 1'b0 ;
  assign n1718 = n476 ^ x25 ^ 1'b0 ;
  assign n1719 = n1718 ^ n866 ^ n595 ;
  assign n1720 = ( x163 & ~n320 ) | ( x163 & n1719 ) | ( ~n320 & n1719 ) ;
  assign n1721 = n436 & n947 ;
  assign n1722 = ~n1515 & n1721 ;
  assign n1723 = n1722 ^ x35 ^ 1'b0 ;
  assign n1724 = n1027 | n1723 ;
  assign n1725 = n778 ^ n380 ^ x200 ;
  assign n1726 = ( n694 & ~n1054 ) | ( n694 & n1725 ) | ( ~n1054 & n1725 ) ;
  assign n1727 = n1165 ^ n773 ^ n698 ;
  assign n1728 = n1456 ^ x168 ^ x38 ;
  assign n1729 = n1728 ^ n1485 ^ n778 ;
  assign n1730 = ( n299 & n315 ) | ( n299 & ~n1729 ) | ( n315 & ~n1729 ) ;
  assign n1731 = n263 & n423 ;
  assign n1732 = n1730 & n1731 ;
  assign n1733 = ( ~n1535 & n1727 ) | ( ~n1535 & n1732 ) | ( n1727 & n1732 ) ;
  assign n1734 = n1527 ^ x225 ^ 1'b0 ;
  assign n1735 = n1734 ^ n1144 ^ 1'b0 ;
  assign n1736 = ( n1726 & n1733 ) | ( n1726 & ~n1735 ) | ( n1733 & ~n1735 ) ;
  assign n1737 = ( ~n1720 & n1724 ) | ( ~n1720 & n1736 ) | ( n1724 & n1736 ) ;
  assign n1738 = n1599 ^ n1412 ^ x60 ;
  assign n1739 = n1691 ^ x2 ^ 1'b0 ;
  assign n1740 = n1739 ^ n1691 ^ n897 ;
  assign n1741 = ( n642 & n1738 ) | ( n642 & ~n1740 ) | ( n1738 & ~n1740 ) ;
  assign n1742 = n1116 | n1527 ;
  assign n1743 = n1742 ^ n1017 ^ 1'b0 ;
  assign n1744 = n1273 ^ n1033 ^ 1'b0 ;
  assign n1745 = n925 & n1744 ;
  assign n1746 = n586 & ~n1745 ;
  assign n1747 = n899 | n1258 ;
  assign n1748 = ( n395 & n1169 ) | ( n395 & n1747 ) | ( n1169 & n1747 ) ;
  assign n1749 = x2 & ~n520 ;
  assign n1750 = n891 & n1749 ;
  assign n1751 = n1750 ^ n727 ^ n326 ;
  assign n1752 = ( ~n1260 & n1623 ) | ( ~n1260 & n1751 ) | ( n1623 & n1751 ) ;
  assign n1753 = n814 ^ n766 ^ n469 ;
  assign n1754 = n622 ^ x90 ^ 1'b0 ;
  assign n1755 = n1754 ^ n882 ^ n264 ;
  assign n1756 = n1107 ^ n664 ^ n497 ;
  assign n1757 = n447 ^ x29 ^ 1'b0 ;
  assign n1758 = n1757 ^ n1221 ^ n634 ;
  assign n1759 = ( x36 & x64 ) | ( x36 & n478 ) | ( x64 & n478 ) ;
  assign n1760 = ( x74 & ~n1282 ) | ( x74 & n1759 ) | ( ~n1282 & n1759 ) ;
  assign n1761 = ( ~n1756 & n1758 ) | ( ~n1756 & n1760 ) | ( n1758 & n1760 ) ;
  assign n1762 = n1761 ^ n1616 ^ n842 ;
  assign n1763 = ( ~n351 & n1196 ) | ( ~n351 & n1762 ) | ( n1196 & n1762 ) ;
  assign n1764 = n1755 & n1763 ;
  assign n1765 = x189 & ~n1041 ;
  assign n1766 = ~n895 & n1765 ;
  assign n1767 = x166 & ~n1766 ;
  assign n1768 = n1767 ^ x178 ^ 1'b0 ;
  assign n1769 = n1768 ^ n607 ^ x64 ;
  assign n1770 = ( n561 & n798 ) | ( n561 & n1769 ) | ( n798 & n1769 ) ;
  assign n1771 = ( n866 & n1206 ) | ( n866 & ~n1770 ) | ( n1206 & ~n1770 ) ;
  assign n1772 = n1771 ^ n935 ^ 1'b0 ;
  assign n1773 = x95 & n1772 ;
  assign n1774 = ( x87 & n636 ) | ( x87 & ~n1355 ) | ( n636 & ~n1355 ) ;
  assign n1775 = n1636 ^ n931 ^ n566 ;
  assign n1776 = ( n828 & n1774 ) | ( n828 & ~n1775 ) | ( n1774 & ~n1775 ) ;
  assign n1777 = n1431 ^ n1227 ^ x172 ;
  assign n1778 = ( n289 & ~n525 ) | ( n289 & n969 ) | ( ~n525 & n969 ) ;
  assign n1779 = n1675 ^ n1382 ^ 1'b0 ;
  assign n1780 = n1778 & ~n1779 ;
  assign n1782 = x43 & ~n459 ;
  assign n1783 = n762 & n1782 ;
  assign n1781 = ~n274 & n578 ;
  assign n1784 = n1783 ^ n1781 ^ 1'b0 ;
  assign n1785 = n1784 ^ n580 ^ 1'b0 ;
  assign n1786 = n1202 | n1513 ;
  assign n1787 = n1785 | n1786 ;
  assign n1788 = n1787 ^ n1392 ^ 1'b0 ;
  assign n1789 = ~x131 & n1788 ;
  assign n1790 = ( x137 & ~n1244 ) | ( x137 & n1555 ) | ( ~n1244 & n1555 ) ;
  assign n1791 = x158 | n982 ;
  assign n1792 = n1791 ^ n308 ^ 1'b0 ;
  assign n1793 = n918 & n1792 ;
  assign n1795 = n430 ^ x143 ^ x108 ;
  assign n1796 = n1795 ^ n442 ^ 1'b0 ;
  assign n1794 = n617 ^ n568 ^ n478 ;
  assign n1797 = n1796 ^ n1794 ^ n1298 ;
  assign n1798 = ~n1405 & n1797 ;
  assign n1799 = n517 & n1798 ;
  assign n1800 = n1793 & ~n1799 ;
  assign n1801 = n1800 ^ n438 ^ 1'b0 ;
  assign n1802 = n414 & n1801 ;
  assign n1803 = n1553 & n1802 ;
  assign n1804 = x111 & n1371 ;
  assign n1806 = ( x247 & ~n710 ) | ( x247 & n1435 ) | ( ~n710 & n1435 ) ;
  assign n1805 = n1724 ^ n515 ^ 1'b0 ;
  assign n1807 = n1806 ^ n1805 ^ n1710 ;
  assign n1808 = ( n656 & ~n720 ) | ( n656 & n1002 ) | ( ~n720 & n1002 ) ;
  assign n1809 = ( ~x245 & n959 ) | ( ~x245 & n1808 ) | ( n959 & n1808 ) ;
  assign n1810 = n1809 ^ x200 ^ 1'b0 ;
  assign n1811 = n1502 | n1810 ;
  assign n1812 = n1248 ^ x96 ^ 1'b0 ;
  assign n1813 = ~n434 & n1812 ;
  assign n1814 = ( ~x166 & x231 ) | ( ~x166 & n394 ) | ( x231 & n394 ) ;
  assign n1816 = n530 ^ x46 ^ x25 ;
  assign n1815 = n546 & n1040 ;
  assign n1817 = n1816 ^ n1815 ^ 1'b0 ;
  assign n1818 = n1817 ^ x143 ^ 1'b0 ;
  assign n1819 = ( n886 & ~n1814 ) | ( n886 & n1818 ) | ( ~n1814 & n1818 ) ;
  assign n1820 = ( ~n607 & n1813 ) | ( ~n607 & n1819 ) | ( n1813 & n1819 ) ;
  assign n1821 = n416 & ~n591 ;
  assign n1822 = n1192 ^ n890 ^ x187 ;
  assign n1823 = ( n913 & n1821 ) | ( n913 & n1822 ) | ( n1821 & n1822 ) ;
  assign n1825 = n1172 & n1304 ;
  assign n1826 = ~n1261 & n1825 ;
  assign n1824 = n594 ^ x45 ^ 1'b0 ;
  assign n1827 = n1826 ^ n1824 ^ x40 ;
  assign n1828 = n583 ^ n345 ^ 1'b0 ;
  assign n1829 = n664 & n1828 ;
  assign n1830 = n1709 & n1829 ;
  assign n1831 = n269 & n870 ;
  assign n1832 = n825 & n1831 ;
  assign n1833 = n992 & n1832 ;
  assign n1834 = n1664 ^ n970 ^ 1'b0 ;
  assign n1835 = n871 & ~n1834 ;
  assign n1836 = ~x173 & n1381 ;
  assign n1837 = n1181 & n1836 ;
  assign n1838 = n755 & n1837 ;
  assign n1839 = n1838 ^ n1729 ^ n1251 ;
  assign n1840 = n1839 ^ n1777 ^ 1'b0 ;
  assign n1841 = n370 ^ x180 ^ 1'b0 ;
  assign n1842 = ~n602 & n1841 ;
  assign n1843 = n1842 ^ x240 ^ 1'b0 ;
  assign n1844 = ( ~x250 & n414 ) | ( ~x250 & n1843 ) | ( n414 & n1843 ) ;
  assign n1845 = n1716 ^ n779 ^ n429 ;
  assign n1846 = ( n1391 & n1787 ) | ( n1391 & n1845 ) | ( n1787 & n1845 ) ;
  assign n1859 = x103 ^ x64 ^ 1'b0 ;
  assign n1860 = x16 & n1859 ;
  assign n1861 = n975 ^ x44 ^ 1'b0 ;
  assign n1862 = n1860 & ~n1861 ;
  assign n1847 = x233 & n1682 ;
  assign n1848 = ~n503 & n1847 ;
  assign n1853 = ( ~x47 & n323 ) | ( ~x47 & n571 ) | ( n323 & n571 ) ;
  assign n1854 = n1853 ^ n1207 ^ 1'b0 ;
  assign n1855 = n1377 & ~n1854 ;
  assign n1851 = n473 ^ n333 ^ x170 ;
  assign n1852 = n1515 & ~n1851 ;
  assign n1849 = n664 & ~n1345 ;
  assign n1850 = n1849 ^ n344 ^ 1'b0 ;
  assign n1856 = n1855 ^ n1852 ^ n1850 ;
  assign n1857 = x78 & n1856 ;
  assign n1858 = n1848 & n1857 ;
  assign n1863 = n1862 ^ n1858 ^ n927 ;
  assign n1865 = x208 ^ x187 ^ 1'b0 ;
  assign n1866 = n1865 ^ n1284 ^ 1'b0 ;
  assign n1864 = ~n649 & n1397 ;
  assign n1867 = n1866 ^ n1864 ^ 1'b0 ;
  assign n1880 = n565 ^ n529 ^ x18 ;
  assign n1868 = ( ~x2 & n453 ) | ( ~x2 & n1044 ) | ( n453 & n1044 ) ;
  assign n1869 = n355 ^ x73 ^ x34 ;
  assign n1870 = n1282 & ~n1869 ;
  assign n1871 = ( n517 & ~n1868 ) | ( n517 & n1870 ) | ( ~n1868 & n1870 ) ;
  assign n1872 = x99 & ~n1871 ;
  assign n1873 = ~n1406 & n1872 ;
  assign n1874 = n1582 ^ x212 ^ 1'b0 ;
  assign n1875 = n798 | n1874 ;
  assign n1876 = n1875 ^ n1583 ^ n1344 ;
  assign n1877 = n1876 ^ n788 ^ 1'b0 ;
  assign n1878 = n1873 | n1877 ;
  assign n1879 = n1878 ^ n1352 ^ 1'b0 ;
  assign n1881 = n1880 ^ n1879 ^ 1'b0 ;
  assign n1882 = n1867 & n1881 ;
  assign n1883 = n269 ^ x222 ^ 1'b0 ;
  assign n1884 = ( x16 & x23 ) | ( x16 & ~x192 ) | ( x23 & ~x192 ) ;
  assign n1885 = n1814 ^ x73 ^ 1'b0 ;
  assign n1886 = n1884 & n1885 ;
  assign n1887 = ~n1883 & n1886 ;
  assign n1888 = x35 & n1312 ;
  assign n1889 = n1888 ^ n856 ^ 1'b0 ;
  assign n1890 = ~n1887 & n1889 ;
  assign n1891 = n1890 ^ n1002 ^ n731 ;
  assign n1892 = ( ~n389 & n829 ) | ( ~n389 & n1891 ) | ( n829 & n1891 ) ;
  assign n1893 = ( n325 & n716 ) | ( n325 & ~n794 ) | ( n716 & ~n794 ) ;
  assign n1894 = ( x224 & ~n440 ) | ( x224 & n1893 ) | ( ~n440 & n1893 ) ;
  assign n1895 = n731 | n1448 ;
  assign n1896 = n1895 ^ n799 ^ 1'b0 ;
  assign n1897 = n1896 ^ n766 ^ x114 ;
  assign n1898 = n1897 ^ n1292 ^ n755 ;
  assign n1899 = n469 | n887 ;
  assign n1900 = ( ~n591 & n1898 ) | ( ~n591 & n1899 ) | ( n1898 & n1899 ) ;
  assign n1901 = ( n902 & ~n908 ) | ( n902 & n966 ) | ( ~n908 & n966 ) ;
  assign n1902 = n928 ^ n578 ^ n277 ;
  assign n1903 = ( x116 & n1901 ) | ( x116 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = ( ~n1062 & n1116 ) | ( ~n1062 & n1903 ) | ( n1116 & n1903 ) ;
  assign n1905 = ( n1894 & n1900 ) | ( n1894 & ~n1904 ) | ( n1900 & ~n1904 ) ;
  assign n1906 = n1756 ^ n831 ^ n674 ;
  assign n1907 = n1906 ^ n1399 ^ n376 ;
  assign n1908 = n458 & ~n1907 ;
  assign n1909 = ~n931 & n1908 ;
  assign n1910 = n1909 ^ n1759 ^ n270 ;
  assign n1911 = n1503 ^ x80 ^ 1'b0 ;
  assign n1912 = n291 | n872 ;
  assign n1913 = n1912 ^ x39 ^ 1'b0 ;
  assign n1914 = ( ~n360 & n365 ) | ( ~n360 & n1913 ) | ( n365 & n1913 ) ;
  assign n1915 = ( n728 & n1124 ) | ( n728 & n1914 ) | ( n1124 & n1914 ) ;
  assign n1916 = n516 ^ n355 ^ x175 ;
  assign n1917 = n1916 ^ n1754 ^ n1285 ;
  assign n1918 = ( ~x113 & n729 ) | ( ~x113 & n1917 ) | ( n729 & n1917 ) ;
  assign n1926 = n1129 ^ n526 ^ x201 ;
  assign n1927 = ( x64 & n598 ) | ( x64 & n1926 ) | ( n598 & n1926 ) ;
  assign n1924 = n899 ^ n645 ^ n503 ;
  assign n1925 = ( n334 & ~n1759 ) | ( n334 & n1924 ) | ( ~n1759 & n1924 ) ;
  assign n1928 = n1927 ^ n1925 ^ n1168 ;
  assign n1923 = x164 & ~n1591 ;
  assign n1929 = n1928 ^ n1923 ^ 1'b0 ;
  assign n1919 = x178 & ~n756 ;
  assign n1920 = n1919 ^ x108 ^ 1'b0 ;
  assign n1921 = x207 & n1920 ;
  assign n1922 = n1071 & ~n1921 ;
  assign n1930 = n1929 ^ n1922 ^ 1'b0 ;
  assign n1931 = ( ~n1508 & n1918 ) | ( ~n1508 & n1930 ) | ( n1918 & n1930 ) ;
  assign n1932 = n1915 | n1931 ;
  assign n1933 = x163 & ~n1932 ;
  assign n1934 = ( n853 & n1911 ) | ( n853 & n1933 ) | ( n1911 & n1933 ) ;
  assign n1935 = ~n656 & n894 ;
  assign n1936 = ( x103 & n375 ) | ( x103 & n396 ) | ( n375 & n396 ) ;
  assign n1937 = n1735 ^ n271 ^ 1'b0 ;
  assign n1938 = n1936 & ~n1937 ;
  assign n1949 = n1144 ^ x156 ^ 1'b0 ;
  assign n1939 = ( n523 & n550 ) | ( n523 & n827 ) | ( n550 & n827 ) ;
  assign n1940 = n1939 ^ n568 ^ 1'b0 ;
  assign n1941 = n977 | n1940 ;
  assign n1942 = n1941 ^ n269 ^ 1'b0 ;
  assign n1945 = n1558 ^ n1460 ^ n516 ;
  assign n1943 = n842 ^ x126 ^ 1'b0 ;
  assign n1944 = n1943 ^ n882 ^ 1'b0 ;
  assign n1946 = n1945 ^ n1944 ^ n722 ;
  assign n1947 = n1942 & ~n1946 ;
  assign n1948 = ( n379 & ~n1134 ) | ( n379 & n1947 ) | ( ~n1134 & n1947 ) ;
  assign n1950 = n1949 ^ n1948 ^ 1'b0 ;
  assign n1951 = n797 ^ x128 ^ 1'b0 ;
  assign n1952 = ~n383 & n607 ;
  assign n1953 = n1604 & ~n1952 ;
  assign n1954 = ( x87 & n1951 ) | ( x87 & n1953 ) | ( n1951 & n1953 ) ;
  assign n1955 = x61 & ~n799 ;
  assign n1956 = n1955 ^ n1487 ^ 1'b0 ;
  assign n1957 = x104 & n1336 ;
  assign n1958 = x16 | n802 ;
  assign n1962 = n1197 ^ n1001 ^ n438 ;
  assign n1959 = n1652 ^ n1385 ^ x240 ;
  assign n1960 = ( n366 & n794 ) | ( n366 & n1959 ) | ( n794 & n1959 ) ;
  assign n1961 = ~n1838 & n1960 ;
  assign n1963 = n1962 ^ n1961 ^ x216 ;
  assign n1964 = x201 & ~n1963 ;
  assign n1965 = ~n1958 & n1964 ;
  assign n1970 = n1054 ^ n535 ^ n526 ;
  assign n1971 = n1970 ^ n1901 ^ n1248 ;
  assign n1972 = n1971 ^ n868 ^ 1'b0 ;
  assign n1969 = n670 | n1054 ;
  assign n1973 = n1972 ^ n1969 ^ 1'b0 ;
  assign n1967 = n1309 ^ n1279 ^ n444 ;
  assign n1966 = n549 ^ n460 ^ x89 ;
  assign n1968 = n1967 ^ n1966 ^ n529 ;
  assign n1974 = n1973 ^ n1968 ^ n594 ;
  assign n1975 = n1965 | n1974 ;
  assign n1976 = n1975 ^ n1503 ^ 1'b0 ;
  assign n1977 = ( ~n798 & n1957 ) | ( ~n798 & n1976 ) | ( n1957 & n1976 ) ;
  assign n1995 = ( n659 & n717 ) | ( n659 & n1041 ) | ( n717 & n1041 ) ;
  assign n1978 = ~n785 & n1729 ;
  assign n1979 = ~x199 & n1978 ;
  assign n1980 = n1087 ^ n562 ^ n407 ;
  assign n1981 = ( n661 & n945 ) | ( n661 & n1237 ) | ( n945 & n1237 ) ;
  assign n1982 = n1096 & ~n1219 ;
  assign n1983 = ( n1980 & n1981 ) | ( n1980 & ~n1982 ) | ( n1981 & ~n1982 ) ;
  assign n1985 = n757 ^ n542 ^ 1'b0 ;
  assign n1986 = n1985 ^ n300 ^ 1'b0 ;
  assign n1987 = ~n929 & n1986 ;
  assign n1988 = n1674 ^ n982 ^ x233 ;
  assign n1989 = n1988 ^ n1256 ^ 1'b0 ;
  assign n1990 = n1987 & n1989 ;
  assign n1984 = n955 | n1926 ;
  assign n1991 = n1990 ^ n1984 ^ 1'b0 ;
  assign n1992 = ( ~n1185 & n1983 ) | ( ~n1185 & n1991 ) | ( n1983 & n1991 ) ;
  assign n1993 = n1992 ^ n1025 ^ 1'b0 ;
  assign n1994 = n1979 | n1993 ;
  assign n1996 = n1995 ^ n1994 ^ n606 ;
  assign n1997 = ( n476 & ~n948 ) | ( n476 & n1496 ) | ( ~n948 & n1496 ) ;
  assign n1998 = ( x163 & x198 ) | ( x163 & n1997 ) | ( x198 & n1997 ) ;
  assign n1999 = ~x197 & n1213 ;
  assign n2000 = n501 & ~n1870 ;
  assign n2001 = ~n931 & n2000 ;
  assign n2002 = n355 | n1144 ;
  assign n2003 = n2002 ^ n961 ^ x235 ;
  assign n2004 = ( n538 & n1186 ) | ( n538 & n2003 ) | ( n1186 & n2003 ) ;
  assign n2005 = ( n1349 & n2001 ) | ( n1349 & ~n2004 ) | ( n2001 & ~n2004 ) ;
  assign n2006 = n1720 ^ n885 ^ x7 ;
  assign n2007 = n2006 ^ n1307 ^ n495 ;
  assign n2008 = n2007 ^ n1629 ^ x90 ;
  assign n2009 = x238 & ~n605 ;
  assign n2011 = n812 ^ n423 ^ 1'b0 ;
  assign n2012 = n2011 ^ n1573 ^ x75 ;
  assign n2010 = n698 ^ n482 ^ n441 ;
  assign n2013 = n2012 ^ n2010 ^ 1'b0 ;
  assign n2014 = n836 | n2013 ;
  assign n2015 = n2014 ^ n2010 ^ n620 ;
  assign n2018 = n1403 ^ n1337 ^ x67 ;
  assign n2016 = ( n1142 & ~n1181 ) | ( n1142 & n1634 ) | ( ~n1181 & n1634 ) ;
  assign n2017 = n2016 ^ n1945 ^ n1155 ;
  assign n2019 = n2018 ^ n2017 ^ 1'b0 ;
  assign n2020 = n1931 ^ n643 ^ n460 ;
  assign n2021 = n1221 ^ n799 ^ x138 ;
  assign n2022 = n2021 ^ n1119 ^ n466 ;
  assign n2023 = n2022 ^ n1344 ^ 1'b0 ;
  assign n2024 = x13 & ~n2023 ;
  assign n2025 = ( ~n574 & n864 ) | ( ~n574 & n1997 ) | ( n864 & n1997 ) ;
  assign n2026 = n752 & n771 ;
  assign n2027 = n1903 & n2026 ;
  assign n2028 = ( n849 & ~n1118 ) | ( n849 & n1734 ) | ( ~n1118 & n1734 ) ;
  assign n2029 = ( x94 & ~n424 ) | ( x94 & n994 ) | ( ~n424 & n994 ) ;
  assign n2030 = n605 ^ x188 ^ 1'b0 ;
  assign n2031 = n2029 & n2030 ;
  assign n2032 = n1261 ^ n828 ^ n781 ;
  assign n2033 = ( ~n536 & n565 ) | ( ~n536 & n1622 ) | ( n565 & n1622 ) ;
  assign n2034 = ( ~n662 & n1336 ) | ( ~n662 & n2033 ) | ( n1336 & n2033 ) ;
  assign n2035 = ~n2032 & n2034 ;
  assign n2036 = n720 ^ n467 ^ 1'b0 ;
  assign n2037 = ~n1061 & n2036 ;
  assign n2038 = n2037 ^ n846 ^ 1'b0 ;
  assign n2039 = n2038 ^ n1778 ^ n1033 ;
  assign n2040 = ( x65 & ~n1032 ) | ( x65 & n2039 ) | ( ~n1032 & n2039 ) ;
  assign n2041 = n2040 ^ n995 ^ n919 ;
  assign n2042 = ( n593 & n2035 ) | ( n593 & ~n2041 ) | ( n2035 & ~n2041 ) ;
  assign n2043 = ( ~n790 & n1435 ) | ( ~n790 & n1777 ) | ( n1435 & n1777 ) ;
  assign n2044 = n376 & ~n2043 ;
  assign n2045 = n355 ^ x123 ^ x43 ;
  assign n2046 = n1123 | n2045 ;
  assign n2047 = n756 | n1637 ;
  assign n2064 = ~x254 & n1337 ;
  assign n2065 = n1345 ^ n1040 ^ 1'b0 ;
  assign n2066 = n2064 | n2065 ;
  assign n2067 = n2066 ^ n700 ^ 1'b0 ;
  assign n2049 = n717 ^ n707 ^ 1'b0 ;
  assign n2050 = n719 & ~n2049 ;
  assign n2058 = n1573 ^ x236 ^ x219 ;
  assign n2055 = n1209 ^ n277 ^ x245 ;
  assign n2056 = n912 & n2055 ;
  assign n2057 = ~x10 & n2056 ;
  assign n2059 = n2058 ^ n2057 ^ n442 ;
  assign n2060 = n2059 ^ n1310 ^ n604 ;
  assign n2052 = n591 ^ n548 ^ x200 ;
  assign n2051 = ( x68 & ~n1515 ) | ( x68 & n1725 ) | ( ~n1515 & n1725 ) ;
  assign n2053 = n2052 ^ n2051 ^ n587 ;
  assign n2054 = ( n1262 & ~n1273 ) | ( n1262 & n2053 ) | ( ~n1273 & n2053 ) ;
  assign n2061 = n2060 ^ n2054 ^ 1'b0 ;
  assign n2062 = n2050 & n2061 ;
  assign n2063 = n534 & n2062 ;
  assign n2068 = n2067 ^ n2063 ^ 1'b0 ;
  assign n2048 = ~n799 & n1112 ;
  assign n2069 = n2068 ^ n2048 ^ 1'b0 ;
  assign n2070 = ( ~x227 & n1172 ) | ( ~x227 & n1306 ) | ( n1172 & n1306 ) ;
  assign n2071 = n1205 ^ n1084 ^ x249 ;
  assign n2072 = ~n1853 & n2071 ;
  assign n2073 = ( n1714 & n1972 ) | ( n1714 & n2072 ) | ( n1972 & n2072 ) ;
  assign n2074 = x70 | n2073 ;
  assign n2075 = n1233 ^ x122 ^ 1'b0 ;
  assign n2076 = n1980 | n2075 ;
  assign n2077 = ( n1424 & n1843 ) | ( n1424 & ~n2076 ) | ( n1843 & ~n2076 ) ;
  assign n2078 = ( x136 & ~n1988 ) | ( x136 & n2077 ) | ( ~n1988 & n2077 ) ;
  assign n2080 = n390 ^ x239 ^ x134 ;
  assign n2081 = ( ~x191 & n853 ) | ( ~x191 & n2080 ) | ( n853 & n2080 ) ;
  assign n2079 = n620 & n723 ;
  assign n2082 = n2081 ^ n2079 ^ n1282 ;
  assign n2083 = n1518 ^ n693 ^ n357 ;
  assign n2084 = n396 ^ x104 ^ 1'b0 ;
  assign n2085 = ( ~n318 & n455 ) | ( ~n318 & n2084 ) | ( n455 & n2084 ) ;
  assign n2086 = n1677 & ~n2085 ;
  assign n2087 = n2086 ^ n1757 ^ 1'b0 ;
  assign n2088 = ( n736 & ~n1688 ) | ( n736 & n2087 ) | ( ~n1688 & n2087 ) ;
  assign n2089 = ( n778 & n1308 ) | ( n778 & ~n1916 ) | ( n1308 & ~n1916 ) ;
  assign n2090 = n1727 & ~n2089 ;
  assign n2091 = n2090 ^ n889 ^ x15 ;
  assign n2092 = n733 ^ n470 ^ x141 ;
  assign n2093 = x26 & ~n463 ;
  assign n2094 = n2093 ^ x86 ^ 1'b0 ;
  assign n2095 = ~n631 & n1350 ;
  assign n2096 = n2094 & n2095 ;
  assign n2097 = ( ~n1906 & n1970 ) | ( ~n1906 & n2096 ) | ( n1970 & n2096 ) ;
  assign n2098 = ( x95 & n1218 ) | ( x95 & n2097 ) | ( n1218 & n2097 ) ;
  assign n2099 = n2092 & ~n2098 ;
  assign n2100 = n702 & n1988 ;
  assign n2104 = n1024 ^ x180 ^ 1'b0 ;
  assign n2102 = x46 & n572 ;
  assign n2103 = n2102 ^ n2052 ^ 1'b0 ;
  assign n2105 = n2104 ^ n2103 ^ 1'b0 ;
  assign n2106 = ( ~x13 & n1077 ) | ( ~x13 & n2105 ) | ( n1077 & n2105 ) ;
  assign n2101 = n1023 ^ n799 ^ n348 ;
  assign n2107 = n2106 ^ n2101 ^ 1'b0 ;
  assign n2108 = n1006 ^ x236 ^ x81 ;
  assign n2109 = n2108 ^ n1860 ^ x136 ;
  assign n2110 = n2109 ^ n1763 ^ n993 ;
  assign n2111 = n2110 ^ n2055 ^ 1'b0 ;
  assign n2112 = x173 & ~n684 ;
  assign n2113 = ~n279 & n2112 ;
  assign n2114 = n2113 ^ n1929 ^ n1312 ;
  assign n2115 = ( ~n1970 & n1971 ) | ( ~n1970 & n2114 ) | ( n1971 & n2114 ) ;
  assign n2116 = n2115 ^ n835 ^ x233 ;
  assign n2117 = n300 | n412 ;
  assign n2118 = n1835 | n2117 ;
  assign n2122 = ( x40 & n1123 ) | ( x40 & ~n1523 ) | ( n1123 & ~n1523 ) ;
  assign n2119 = ~n412 & n640 ;
  assign n2120 = n2119 ^ n857 ^ 1'b0 ;
  assign n2121 = ~n1532 & n2120 ;
  assign n2123 = n2122 ^ n2121 ^ 1'b0 ;
  assign n2124 = n863 ^ x105 ^ 1'b0 ;
  assign n2125 = ( ~x125 & n823 ) | ( ~x125 & n2124 ) | ( n823 & n2124 ) ;
  assign n2126 = ( n1179 & n2123 ) | ( n1179 & n2125 ) | ( n2123 & n2125 ) ;
  assign n2138 = n489 & n657 ;
  assign n2139 = n2138 ^ n1795 ^ 1'b0 ;
  assign n2127 = ( x84 & n475 ) | ( x84 & n1221 ) | ( n475 & n1221 ) ;
  assign n2128 = ( ~x14 & n447 ) | ( ~x14 & n2127 ) | ( n447 & n2127 ) ;
  assign n2129 = ( x163 & ~n1884 ) | ( x163 & n2128 ) | ( ~n1884 & n2128 ) ;
  assign n2131 = x212 & ~n290 ;
  assign n2132 = n2131 ^ x28 ^ 1'b0 ;
  assign n2133 = ( x68 & ~x194 ) | ( x68 & n2132 ) | ( ~x194 & n2132 ) ;
  assign n2134 = n1184 ^ n1117 ^ x50 ;
  assign n2135 = ( n339 & n2133 ) | ( n339 & n2134 ) | ( n2133 & n2134 ) ;
  assign n2130 = ( n1162 & ~n1379 ) | ( n1162 & n1568 ) | ( ~n1379 & n1568 ) ;
  assign n2136 = n2135 ^ n2130 ^ 1'b0 ;
  assign n2137 = ~n2129 & n2136 ;
  assign n2140 = n2139 ^ n2137 ^ 1'b0 ;
  assign n2141 = ( n805 & ~n1495 ) | ( n805 & n1961 ) | ( ~n1495 & n1961 ) ;
  assign n2142 = ( ~n2126 & n2140 ) | ( ~n2126 & n2141 ) | ( n2140 & n2141 ) ;
  assign n2148 = ( ~x149 & n481 ) | ( ~x149 & n705 ) | ( n481 & n705 ) ;
  assign n2149 = n951 ^ x6 ^ 1'b0 ;
  assign n2150 = n1284 | n2149 ;
  assign n2151 = ( n624 & n2148 ) | ( n624 & n2150 ) | ( n2148 & n2150 ) ;
  assign n2152 = n2151 ^ n559 ^ 1'b0 ;
  assign n2153 = ~n1338 & n2152 ;
  assign n2154 = n2153 ^ n1354 ^ 1'b0 ;
  assign n2155 = n2154 ^ n548 ^ 1'b0 ;
  assign n2156 = ~n1619 & n2155 ;
  assign n2147 = n1629 ^ n1394 ^ n1127 ;
  assign n2143 = n948 ^ n425 ^ x139 ;
  assign n2144 = ~n885 & n2143 ;
  assign n2145 = n2144 ^ n698 ^ n630 ;
  assign n2146 = ( n655 & ~n2010 ) | ( n655 & n2145 ) | ( ~n2010 & n2145 ) ;
  assign n2157 = n2156 ^ n2147 ^ n2146 ;
  assign n2158 = ( x143 & n1330 ) | ( x143 & ~n2078 ) | ( n1330 & ~n2078 ) ;
  assign n2159 = n1869 ^ n925 ^ 1'b0 ;
  assign n2160 = n1865 & n2159 ;
  assign n2161 = ( x241 & n932 ) | ( x241 & ~n2160 ) | ( n932 & ~n2160 ) ;
  assign n2173 = ( ~n469 & n999 ) | ( ~n469 & n1386 ) | ( n999 & n1386 ) ;
  assign n2162 = ( x167 & ~n257 ) | ( x167 & n539 ) | ( ~n257 & n539 ) ;
  assign n2163 = ( ~x136 & n1019 ) | ( ~x136 & n1130 ) | ( n1019 & n1130 ) ;
  assign n2164 = n2162 | n2163 ;
  assign n2170 = n429 & n1129 ;
  assign n2165 = ~n505 & n548 ;
  assign n2166 = ~x222 & n2165 ;
  assign n2167 = n394 ^ x78 ^ 1'b0 ;
  assign n2168 = ~n2166 & n2167 ;
  assign n2169 = ( n400 & n863 ) | ( n400 & ~n2168 ) | ( n863 & ~n2168 ) ;
  assign n2171 = n2170 ^ n2169 ^ 1'b0 ;
  assign n2172 = ~n2164 & n2171 ;
  assign n2174 = n2173 ^ n2172 ^ 1'b0 ;
  assign n2175 = ( n817 & n2161 ) | ( n817 & ~n2174 ) | ( n2161 & ~n2174 ) ;
  assign n2176 = ( n597 & ~n798 ) | ( n597 & n2175 ) | ( ~n798 & n2175 ) ;
  assign n2185 = n1380 ^ n652 ^ x227 ;
  assign n2186 = n2185 ^ n330 ^ x166 ;
  assign n2183 = n360 ^ x230 ^ x219 ;
  assign n2182 = ( x110 & n2032 ) | ( x110 & n2033 ) | ( n2032 & n2033 ) ;
  assign n2184 = n2183 ^ n2182 ^ x175 ;
  assign n2178 = ( x46 & ~x116 ) | ( x46 & n330 ) | ( ~x116 & n330 ) ;
  assign n2179 = n2178 ^ n1883 ^ n1766 ;
  assign n2180 = n2179 ^ n1310 ^ n909 ;
  assign n2177 = n1822 ^ n515 ^ 1'b0 ;
  assign n2181 = n2180 ^ n2177 ^ n458 ;
  assign n2187 = n2186 ^ n2184 ^ n2181 ;
  assign n2188 = n2015 ^ x221 ^ x20 ;
  assign n2193 = n1347 ^ n763 ^ n520 ;
  assign n2189 = ( n602 & ~n853 ) | ( n602 & n2120 ) | ( ~n853 & n2120 ) ;
  assign n2190 = n2189 ^ n1499 ^ n617 ;
  assign n2191 = n332 & ~n2190 ;
  assign n2192 = n524 & n2191 ;
  assign n2194 = n2193 ^ n2192 ^ n1326 ;
  assign n2195 = ( x211 & x241 ) | ( x211 & ~n1151 ) | ( x241 & ~n1151 ) ;
  assign n2196 = x196 ^ x70 ^ 1'b0 ;
  assign n2197 = n817 & n2196 ;
  assign n2198 = ( n342 & ~n2195 ) | ( n342 & n2197 ) | ( ~n2195 & n2197 ) ;
  assign n2199 = ( ~x180 & n1795 ) | ( ~x180 & n1860 ) | ( n1795 & n1860 ) ;
  assign n2200 = ( n351 & n616 ) | ( n351 & n726 ) | ( n616 & n726 ) ;
  assign n2201 = n2200 ^ x145 ^ 1'b0 ;
  assign n2202 = n399 & n2201 ;
  assign n2203 = ( x163 & ~n2199 ) | ( x163 & n2202 ) | ( ~n2199 & n2202 ) ;
  assign n2204 = n978 & n2203 ;
  assign n2205 = n2198 & n2204 ;
  assign n2206 = ( n525 & n1900 ) | ( n525 & n2205 ) | ( n1900 & n2205 ) ;
  assign n2207 = x209 & n357 ;
  assign n2208 = n570 & n2207 ;
  assign n2209 = n1564 ^ n361 ^ 1'b0 ;
  assign n2210 = n2209 ^ n1076 ^ n723 ;
  assign n2211 = n1635 | n2210 ;
  assign n2212 = x62 | n2211 ;
  assign n2213 = n2133 ^ n535 ^ 1'b0 ;
  assign n2215 = x5 & x86 ;
  assign n2216 = n941 & n2215 ;
  assign n2217 = ( ~n434 & n1041 ) | ( ~n434 & n2216 ) | ( n1041 & n2216 ) ;
  assign n2218 = ( n431 & n870 ) | ( n431 & ~n2217 ) | ( n870 & ~n2217 ) ;
  assign n2214 = ( x174 & n610 ) | ( x174 & n635 ) | ( n610 & n635 ) ;
  assign n2219 = n2218 ^ n2214 ^ 1'b0 ;
  assign n2220 = n2213 & n2219 ;
  assign n2221 = ( n715 & n2212 ) | ( n715 & n2220 ) | ( n2212 & n2220 ) ;
  assign n2222 = n1905 ^ n1276 ^ n500 ;
  assign n2224 = n1186 ^ n1100 ^ n822 ;
  assign n2223 = n1850 ^ n1597 ^ n1569 ;
  assign n2225 = n2224 ^ n2223 ^ 1'b0 ;
  assign n2226 = ~n987 & n2225 ;
  assign n2227 = n1880 ^ n290 ^ x208 ;
  assign n2228 = n2227 ^ n1410 ^ 1'b0 ;
  assign n2229 = n2228 ^ x27 ^ 1'b0 ;
  assign n2230 = x221 & n2229 ;
  assign n2231 = ( n505 & n1274 ) | ( n505 & ~n1718 ) | ( n1274 & ~n1718 ) ;
  assign n2232 = n1521 ^ n615 ^ n390 ;
  assign n2233 = ( x240 & ~n696 ) | ( x240 & n2232 ) | ( ~n696 & n2232 ) ;
  assign n2234 = n1581 ^ x116 ^ x85 ;
  assign n2235 = n1552 ^ n967 ^ n406 ;
  assign n2236 = n973 ^ n634 ^ 1'b0 ;
  assign n2237 = x112 & ~n2236 ;
  assign n2238 = n340 & n2237 ;
  assign n2239 = ~x166 & n2238 ;
  assign n2240 = ~n2235 & n2239 ;
  assign n2241 = ( n261 & n1392 ) | ( n261 & n2240 ) | ( n1392 & n2240 ) ;
  assign n2243 = x28 & ~n1412 ;
  assign n2242 = n1224 ^ n681 ^ n460 ;
  assign n2244 = n2243 ^ n2242 ^ n412 ;
  assign n2245 = n1616 ^ n894 ^ 1'b0 ;
  assign n2246 = ~n619 & n1862 ;
  assign n2247 = n2246 ^ n1848 ^ 1'b0 ;
  assign n2248 = n1361 ^ n1084 ^ n414 ;
  assign n2249 = n2248 ^ n1725 ^ 1'b0 ;
  assign n2250 = n1056 & ~n2249 ;
  assign n2251 = ( n2245 & n2247 ) | ( n2245 & n2250 ) | ( n2247 & n2250 ) ;
  assign n2252 = ( ~n1435 & n1609 ) | ( ~n1435 & n2005 ) | ( n1609 & n2005 ) ;
  assign n2254 = n1240 ^ n861 ^ x32 ;
  assign n2253 = n889 & n1365 ;
  assign n2255 = n2254 ^ n2253 ^ 1'b0 ;
  assign n2256 = ( n587 & n673 ) | ( n587 & ~n2255 ) | ( n673 & ~n2255 ) ;
  assign n2257 = n2256 ^ x75 ^ 1'b0 ;
  assign n2258 = n2257 ^ n1313 ^ n1133 ;
  assign n2263 = ( x156 & n1507 ) | ( x156 & ~n1633 ) | ( n1507 & ~n1633 ) ;
  assign n2264 = ( n310 & n1044 ) | ( n310 & n2263 ) | ( n1044 & n2263 ) ;
  assign n2261 = n943 & ~n1313 ;
  assign n2262 = n2261 ^ n865 ^ 1'b0 ;
  assign n2259 = ( ~x19 & x108 ) | ( ~x19 & n793 ) | ( x108 & n793 ) ;
  assign n2260 = ( x27 & ~n1151 ) | ( x27 & n2259 ) | ( ~n1151 & n2259 ) ;
  assign n2265 = n2264 ^ n2262 ^ n2260 ;
  assign n2266 = n2265 ^ n661 ^ x254 ;
  assign n2267 = n540 ^ n257 ^ 1'b0 ;
  assign n2268 = n421 & n2267 ;
  assign n2269 = n2268 ^ n783 ^ 1'b0 ;
  assign n2270 = ~n1184 & n2269 ;
  assign n2271 = n2270 ^ n1642 ^ n970 ;
  assign n2276 = n1121 & ~n1670 ;
  assign n2277 = n2276 ^ n857 ^ 1'b0 ;
  assign n2278 = n2277 ^ n2268 ^ n631 ;
  assign n2272 = n1186 ^ x217 ^ x173 ;
  assign n2273 = n1899 ^ n917 ^ 1'b0 ;
  assign n2274 = n700 & ~n2273 ;
  assign n2275 = n2272 & n2274 ;
  assign n2279 = n2278 ^ n2275 ^ 1'b0 ;
  assign n2280 = x30 & ~n2279 ;
  assign n2281 = n1172 ^ x202 ^ 1'b0 ;
  assign n2282 = ( ~n1186 & n1655 ) | ( ~n1186 & n2281 ) | ( n1655 & n2281 ) ;
  assign n2283 = n332 ^ x78 ^ x16 ;
  assign n2284 = n2283 ^ n1537 ^ 1'b0 ;
  assign n2285 = x26 & ~n2284 ;
  assign n2286 = ( x215 & n1060 ) | ( x215 & ~n2285 ) | ( n1060 & ~n2285 ) ;
  assign n2287 = x171 & ~n2286 ;
  assign n2288 = ~n2257 & n2287 ;
  assign n2289 = n2288 ^ n1803 ^ n1151 ;
  assign n2290 = ( ~n544 & n2282 ) | ( ~n544 & n2289 ) | ( n2282 & n2289 ) ;
  assign n2291 = x17 & x96 ;
  assign n2292 = n2291 ^ n1048 ^ 1'b0 ;
  assign n2293 = n760 & ~n2292 ;
  assign n2294 = n961 & n2293 ;
  assign n2295 = ( n952 & n995 ) | ( n952 & n2294 ) | ( n995 & n2294 ) ;
  assign n2296 = n950 ^ n687 ^ n310 ;
  assign n2297 = x14 & x177 ;
  assign n2298 = n1042 & n2297 ;
  assign n2299 = ( ~n1661 & n2110 ) | ( ~n1661 & n2298 ) | ( n2110 & n2298 ) ;
  assign n2300 = ( ~n1793 & n2296 ) | ( ~n1793 & n2299 ) | ( n2296 & n2299 ) ;
  assign n2301 = ( n1320 & n1618 ) | ( n1320 & ~n2300 ) | ( n1618 & ~n2300 ) ;
  assign n2302 = ( x34 & n1054 ) | ( x34 & ~n2060 ) | ( n1054 & ~n2060 ) ;
  assign n2303 = ( ~n585 & n987 ) | ( ~n585 & n1258 ) | ( n987 & n1258 ) ;
  assign n2304 = n1380 & ~n2303 ;
  assign n2305 = n1822 & n2304 ;
  assign n2306 = ( n700 & ~n1871 ) | ( n700 & n2305 ) | ( ~n1871 & n2305 ) ;
  assign n2307 = x5 & x14 ;
  assign n2308 = n2307 ^ x204 ^ 1'b0 ;
  assign n2309 = ( ~n799 & n2150 ) | ( ~n799 & n2308 ) | ( n2150 & n2308 ) ;
  assign n2310 = ( x73 & ~n452 ) | ( x73 & n2309 ) | ( ~n452 & n2309 ) ;
  assign n2311 = ~n1401 & n2310 ;
  assign n2324 = n750 ^ n639 ^ n376 ;
  assign n2325 = n2324 ^ n1604 ^ n375 ;
  assign n2319 = ( ~x198 & n271 ) | ( ~x198 & n490 ) | ( n271 & n490 ) ;
  assign n2320 = x52 & n2319 ;
  assign n2321 = ~n1850 & n2320 ;
  assign n2313 = n1119 & ~n1423 ;
  assign n2314 = n1003 & ~n2313 ;
  assign n2315 = ~n1797 & n2314 ;
  assign n2316 = n599 | n2315 ;
  assign n2317 = n1274 | n2316 ;
  assign n2312 = ~n488 & n1576 ;
  assign n2318 = n2317 ^ n2312 ^ 1'b0 ;
  assign n2322 = n2321 ^ n2318 ^ 1'b0 ;
  assign n2323 = ~n409 & n2322 ;
  assign n2326 = n2325 ^ n2323 ^ n520 ;
  assign n2327 = n2326 ^ n1266 ^ 1'b0 ;
  assign n2328 = x174 & n2327 ;
  assign n2329 = ( ~n1110 & n1312 ) | ( ~n1110 & n1585 ) | ( n1312 & n1585 ) ;
  assign n2330 = ~n982 & n1574 ;
  assign n2331 = n1565 & n2330 ;
  assign n2332 = ( ~n2286 & n2329 ) | ( ~n2286 & n2331 ) | ( n2329 & n2331 ) ;
  assign n2333 = n2332 ^ n1031 ^ 1'b0 ;
  assign n2338 = x113 & ~n539 ;
  assign n2339 = ~n1466 & n2338 ;
  assign n2340 = n2190 | n2339 ;
  assign n2341 = x45 | n2340 ;
  assign n2342 = n2341 ^ n456 ^ x239 ;
  assign n2334 = n1853 ^ n1546 ^ n372 ;
  assign n2335 = n795 & n2334 ;
  assign n2336 = n2335 ^ n1945 ^ 1'b0 ;
  assign n2337 = ~n1456 & n2336 ;
  assign n2343 = n2342 ^ n2337 ^ 1'b0 ;
  assign n2352 = n1766 | n1836 ;
  assign n2344 = n616 ^ n419 ^ 1'b0 ;
  assign n2345 = x159 & n2344 ;
  assign n2347 = ( ~x122 & x153 ) | ( ~x122 & n480 ) | ( x153 & n480 ) ;
  assign n2346 = ~n775 & n1312 ;
  assign n2348 = n2347 ^ n2346 ^ n2089 ;
  assign n2349 = n1097 & ~n2348 ;
  assign n2350 = n2349 ^ n504 ^ 1'b0 ;
  assign n2351 = n2345 & ~n2350 ;
  assign n2353 = n2352 ^ n2351 ^ 1'b0 ;
  assign n2354 = x229 & n475 ;
  assign n2355 = ~n351 & n2354 ;
  assign n2356 = x18 & n2355 ;
  assign n2357 = ( x202 & n814 ) | ( x202 & n2356 ) | ( n814 & n2356 ) ;
  assign n2359 = x224 & ~n614 ;
  assign n2360 = n2359 ^ n581 ^ 1'b0 ;
  assign n2358 = n537 | n794 ;
  assign n2361 = n2360 ^ n2358 ^ 1'b0 ;
  assign n2362 = ~n919 & n2361 ;
  assign n2363 = ~n343 & n2362 ;
  assign n2364 = ( n1882 & n2357 ) | ( n1882 & ~n2363 ) | ( n2357 & ~n2363 ) ;
  assign n2368 = ~n2022 & n2148 ;
  assign n2369 = n2368 ^ n277 ^ 1'b0 ;
  assign n2365 = x197 & n1745 ;
  assign n2366 = n438 | n2365 ;
  assign n2367 = n2366 ^ n890 ^ 1'b0 ;
  assign n2370 = n2369 ^ n2367 ^ n1876 ;
  assign n2371 = n2230 ^ n1747 ^ n1189 ;
  assign n2375 = n738 & ~n770 ;
  assign n2376 = n2375 ^ x86 ^ 1'b0 ;
  assign n2377 = n2376 ^ n1507 ^ n1139 ;
  assign n2378 = ~n385 & n2377 ;
  assign n2372 = n1161 ^ n747 ^ 1'b0 ;
  assign n2373 = n2372 ^ n1896 ^ n1476 ;
  assign n2374 = n603 | n2373 ;
  assign n2379 = n2378 ^ n2374 ^ 1'b0 ;
  assign n2382 = ( n359 & ~n397 ) | ( n359 & n565 ) | ( ~n397 & n565 ) ;
  assign n2381 = ( x249 & ~n298 ) | ( x249 & n858 ) | ( ~n298 & n858 ) ;
  assign n2380 = n2101 ^ n999 ^ n407 ;
  assign n2383 = n2382 ^ n2381 ^ n2380 ;
  assign n2384 = n2383 ^ x109 ^ 1'b0 ;
  assign n2385 = n1205 & ~n2384 ;
  assign n2387 = x251 & ~n598 ;
  assign n2388 = ~x135 & n2387 ;
  assign n2389 = n1096 ^ n653 ^ n578 ;
  assign n2390 = ( ~n1292 & n2388 ) | ( ~n1292 & n2389 ) | ( n2388 & n2389 ) ;
  assign n2391 = n2390 ^ n748 ^ 1'b0 ;
  assign n2392 = ~n1694 & n2391 ;
  assign n2386 = ~n295 & n1200 ;
  assign n2393 = n2392 ^ n2386 ^ 1'b0 ;
  assign n2394 = n2393 ^ n1582 ^ 1'b0 ;
  assign n2395 = n2394 ^ n2319 ^ n1601 ;
  assign n2396 = x45 & x172 ;
  assign n2397 = n2395 & n2396 ;
  assign n2398 = n961 ^ n289 ^ 1'b0 ;
  assign n2399 = n496 | n2398 ;
  assign n2400 = n1491 ^ n471 ^ 1'b0 ;
  assign n2401 = ( ~x10 & n706 ) | ( ~x10 & n1153 ) | ( n706 & n1153 ) ;
  assign n2402 = n2401 ^ n1618 ^ 1'b0 ;
  assign n2403 = n1028 & n2402 ;
  assign n2404 = ( n1465 & ~n2400 ) | ( n1465 & n2403 ) | ( ~n2400 & n2403 ) ;
  assign n2405 = n2404 ^ n1131 ^ 1'b0 ;
  assign n2406 = n1371 | n2405 ;
  assign n2407 = ~n1527 & n1842 ;
  assign n2408 = n2407 ^ n1096 ^ 1'b0 ;
  assign n2412 = n1569 ^ n1477 ^ 1'b0 ;
  assign n2410 = n1055 ^ n825 ^ n501 ;
  assign n2409 = ~n329 & n823 ;
  assign n2411 = n2410 ^ n2409 ^ 1'b0 ;
  assign n2413 = n2412 ^ n2411 ^ x186 ;
  assign n2414 = ( ~n1018 & n1477 ) | ( ~n1018 & n2413 ) | ( n1477 & n2413 ) ;
  assign n2415 = ( ~n1028 & n2408 ) | ( ~n1028 & n2414 ) | ( n2408 & n2414 ) ;
  assign n2416 = n639 | n2415 ;
  assign n2417 = n1155 & ~n2416 ;
  assign n2418 = n635 ^ x23 ^ 1'b0 ;
  assign n2419 = ~n885 & n2418 ;
  assign n2420 = n2419 ^ n612 ^ 1'b0 ;
  assign n2421 = n2420 ^ n1423 ^ 1'b0 ;
  assign n2422 = n2417 | n2421 ;
  assign n2423 = n2406 | n2422 ;
  assign n2424 = n2399 & ~n2423 ;
  assign n2426 = n1201 ^ n327 ^ 1'b0 ;
  assign n2425 = ~n495 & n1633 ;
  assign n2427 = n2426 ^ n2425 ^ n786 ;
  assign n2428 = x75 & ~n1577 ;
  assign n2429 = n1381 ^ x245 ^ 1'b0 ;
  assign n2430 = n1279 ^ n599 ^ n414 ;
  assign n2431 = x109 & n830 ;
  assign n2432 = n2431 ^ n639 ^ 1'b0 ;
  assign n2433 = ( n1062 & n2288 ) | ( n1062 & n2432 ) | ( n2288 & n2432 ) ;
  assign n2434 = n1226 & ~n2433 ;
  assign n2435 = ( n405 & n1602 ) | ( n405 & n2434 ) | ( n1602 & n2434 ) ;
  assign n2436 = n2132 ^ n1365 ^ x113 ;
  assign n2437 = n2068 ^ n1477 ^ 1'b0 ;
  assign n2442 = n2057 ^ n702 ^ 1'b0 ;
  assign n2439 = n529 & n1573 ;
  assign n2440 = n2439 ^ n1257 ^ 1'b0 ;
  assign n2438 = n1575 ^ n399 ^ x150 ;
  assign n2441 = n2440 ^ n2438 ^ 1'b0 ;
  assign n2443 = n2442 ^ n2441 ^ n268 ;
  assign n2444 = ( n2436 & ~n2437 ) | ( n2436 & n2443 ) | ( ~n2437 & n2443 ) ;
  assign n2445 = n731 ^ n494 ^ 1'b0 ;
  assign n2446 = x122 & ~n1467 ;
  assign n2447 = ~n2445 & n2446 ;
  assign n2448 = n2447 ^ n1024 ^ 1'b0 ;
  assign n2449 = n2448 ^ n1597 ^ 1'b0 ;
  assign n2450 = ( ~n274 & n308 ) | ( ~n274 & n1177 ) | ( n308 & n1177 ) ;
  assign n2451 = n2450 ^ n2057 ^ n1168 ;
  assign n2461 = n1674 ^ n1189 ^ n1154 ;
  assign n2462 = n2179 & n2461 ;
  assign n2463 = ( x39 & n830 ) | ( x39 & ~n2462 ) | ( n830 & ~n2462 ) ;
  assign n2464 = n2388 ^ n1795 ^ 1'b0 ;
  assign n2465 = n2463 & ~n2464 ;
  assign n2466 = ( x111 & n329 ) | ( x111 & n340 ) | ( n329 & n340 ) ;
  assign n2467 = n710 & n2466 ;
  assign n2468 = n2467 ^ n467 ^ 1'b0 ;
  assign n2469 = n287 & n336 ;
  assign n2470 = n2468 & n2469 ;
  assign n2471 = ( x39 & ~n2465 ) | ( x39 & n2470 ) | ( ~n2465 & n2470 ) ;
  assign n2452 = n2084 ^ n822 ^ x58 ;
  assign n2453 = x149 & ~n2452 ;
  assign n2454 = ( x94 & n277 ) | ( x94 & ~n334 ) | ( n277 & ~n334 ) ;
  assign n2455 = ( ~x195 & n2254 ) | ( ~x195 & n2454 ) | ( n2254 & n2454 ) ;
  assign n2456 = ( ~n396 & n1601 ) | ( ~n396 & n2455 ) | ( n1601 & n2455 ) ;
  assign n2457 = n2456 ^ n1603 ^ n1164 ;
  assign n2458 = ~n431 & n2456 ;
  assign n2459 = n2457 & n2458 ;
  assign n2460 = n2453 | n2459 ;
  assign n2472 = n2471 ^ n2460 ^ 1'b0 ;
  assign n2473 = n2133 ^ n831 ^ n608 ;
  assign n2474 = n1853 ^ n674 ^ n578 ;
  assign n2475 = n2474 ^ n1632 ^ 1'b0 ;
  assign n2476 = ( x110 & ~n2473 ) | ( x110 & n2475 ) | ( ~n2473 & n2475 ) ;
  assign n2477 = n1884 ^ n1091 ^ 1'b0 ;
  assign n2478 = ~n1155 & n2477 ;
  assign n2479 = n2476 & n2478 ;
  assign n2480 = ~n809 & n1635 ;
  assign n2481 = ( n363 & n1121 ) | ( n363 & ~n2455 ) | ( n1121 & ~n2455 ) ;
  assign n2482 = ( n557 & n1676 ) | ( n557 & n2481 ) | ( n1676 & n2481 ) ;
  assign n2483 = n2482 ^ n1230 ^ 1'b0 ;
  assign n2484 = n367 & n2483 ;
  assign n2485 = n2484 ^ n1824 ^ x158 ;
  assign n2486 = ( ~n352 & n1502 ) | ( ~n352 & n2485 ) | ( n1502 & n2485 ) ;
  assign n2487 = ~n1015 & n1561 ;
  assign n2488 = n2487 ^ n897 ^ 1'b0 ;
  assign n2489 = n2248 & n2488 ;
  assign n2490 = n1302 ^ n1214 ^ n803 ;
  assign n2491 = ( n1457 & n2489 ) | ( n1457 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = n819 ^ n790 ^ n393 ;
  assign n2493 = x37 & ~n2492 ;
  assign n2494 = n2493 ^ n2339 ^ 1'b0 ;
  assign n2495 = ~n548 & n1573 ;
  assign n2496 = ( x251 & ~n2494 ) | ( x251 & n2495 ) | ( ~n2494 & n2495 ) ;
  assign n2500 = n1423 ^ x29 ^ 1'b0 ;
  assign n2501 = n912 & ~n2500 ;
  assign n2497 = n538 ^ n287 ^ 1'b0 ;
  assign n2498 = ~n1657 & n2497 ;
  assign n2499 = n2498 ^ n2263 ^ 1'b0 ;
  assign n2502 = n2501 ^ n2499 ^ n1384 ;
  assign n2503 = n1816 ^ n963 ^ 1'b0 ;
  assign n2504 = ~n2502 & n2503 ;
  assign n2505 = n1346 ^ n461 ^ 1'b0 ;
  assign n2506 = n1200 | n2505 ;
  assign n2507 = ( n414 & n1287 ) | ( n414 & ~n2071 ) | ( n1287 & ~n2071 ) ;
  assign n2508 = n2507 ^ n1843 ^ n396 ;
  assign n2509 = ( n326 & n519 ) | ( n326 & n1122 ) | ( n519 & n1122 ) ;
  assign n2510 = ( ~n841 & n1417 ) | ( ~n841 & n2509 ) | ( n1417 & n2509 ) ;
  assign n2511 = n2508 & n2510 ;
  assign n2512 = ~n1245 & n2511 ;
  assign n2513 = n2506 | n2512 ;
  assign n2514 = n1420 | n2513 ;
  assign n2515 = ( n376 & n2504 ) | ( n376 & ~n2514 ) | ( n2504 & ~n2514 ) ;
  assign n2516 = n1440 ^ n1142 ^ 1'b0 ;
  assign n2517 = ( n966 & n1230 ) | ( n966 & ~n1955 ) | ( n1230 & ~n1955 ) ;
  assign n2520 = x241 ^ x195 ^ x21 ;
  assign n2518 = n649 ^ x88 ^ 1'b0 ;
  assign n2519 = x180 & n2518 ;
  assign n2521 = n2520 ^ n2519 ^ n308 ;
  assign n2522 = ( ~n2205 & n2517 ) | ( ~n2205 & n2521 ) | ( n2517 & n2521 ) ;
  assign n2523 = ( n1188 & n2321 ) | ( n1188 & ~n2522 ) | ( n2321 & ~n2522 ) ;
  assign n2524 = ( x226 & n1341 ) | ( x226 & ~n1943 ) | ( n1341 & ~n1943 ) ;
  assign n2525 = ~n2190 & n2524 ;
  assign n2528 = n1686 ^ n365 ^ x207 ;
  assign n2529 = ( n859 & n1334 ) | ( n859 & ~n2528 ) | ( n1334 & ~n2528 ) ;
  assign n2526 = n495 ^ n402 ^ 1'b0 ;
  assign n2527 = n2526 ^ n1046 ^ 1'b0 ;
  assign n2530 = n2529 ^ n2527 ^ 1'b0 ;
  assign n2531 = ( x40 & n2217 ) | ( x40 & ~n2451 ) | ( n2217 & ~n2451 ) ;
  assign n2532 = n1077 ^ n704 ^ 1'b0 ;
  assign n2533 = ~n1707 & n2532 ;
  assign n2538 = n2160 ^ n715 ^ n481 ;
  assign n2534 = n1616 ^ n1371 ^ 1'b0 ;
  assign n2535 = n628 | n2534 ;
  assign n2536 = ( x9 & n1355 ) | ( x9 & ~n2535 ) | ( n1355 & ~n2535 ) ;
  assign n2537 = x183 & n2536 ;
  assign n2539 = n2538 ^ n2537 ^ 1'b0 ;
  assign n2540 = n2010 ^ n1155 ^ n912 ;
  assign n2541 = n355 | n589 ;
  assign n2542 = x147 | n2541 ;
  assign n2543 = ~n989 & n2542 ;
  assign n2544 = ~n2540 & n2543 ;
  assign n2545 = ( ~x223 & n2195 ) | ( ~x223 & n2544 ) | ( n2195 & n2544 ) ;
  assign n2546 = ( n2533 & ~n2539 ) | ( n2533 & n2545 ) | ( ~n2539 & n2545 ) ;
  assign n2549 = n1689 ^ n906 ^ x245 ;
  assign n2547 = ( n582 & n740 ) | ( n582 & ~n2050 ) | ( n740 & ~n2050 ) ;
  assign n2548 = n2547 ^ n2007 ^ n1682 ;
  assign n2550 = n2549 ^ n2548 ^ n325 ;
  assign n2554 = x234 & n795 ;
  assign n2555 = n961 & n2554 ;
  assign n2553 = ~n1819 & n2156 ;
  assign n2551 = ~n799 & n2074 ;
  assign n2552 = n2186 & n2551 ;
  assign n2556 = n2555 ^ n2553 ^ n2552 ;
  assign n2557 = ( n1071 & ~n1196 ) | ( n1071 & n1398 ) | ( ~n1196 & n1398 ) ;
  assign n2558 = n2557 ^ n2108 ^ n1901 ;
  assign n2559 = ~n264 & n582 ;
  assign n2560 = ( ~n1023 & n1418 ) | ( ~n1023 & n2559 ) | ( n1418 & n2559 ) ;
  assign n2561 = ( x235 & ~n558 ) | ( x235 & n966 ) | ( ~n558 & n966 ) ;
  assign n2563 = n306 & ~n684 ;
  assign n2564 = n2563 ^ x43 ^ 1'b0 ;
  assign n2562 = n1210 ^ n692 ^ x79 ;
  assign n2565 = n2564 ^ n2562 ^ n2263 ;
  assign n2566 = n2565 ^ n713 ^ 1'b0 ;
  assign n2567 = n2053 | n2566 ;
  assign n2568 = n2561 & ~n2567 ;
  assign n2569 = ( n499 & ~n1212 ) | ( n499 & n2568 ) | ( ~n1212 & n2568 ) ;
  assign n2570 = n2098 ^ n1750 ^ 1'b0 ;
  assign n2577 = ~n370 & n1645 ;
  assign n2571 = x123 & ~n414 ;
  assign n2572 = ~n1365 & n2571 ;
  assign n2573 = ( ~n545 & n978 ) | ( ~n545 & n2572 ) | ( n978 & n2572 ) ;
  assign n2574 = n257 & n552 ;
  assign n2575 = n2574 ^ n693 ^ 1'b0 ;
  assign n2576 = ( n1612 & ~n2573 ) | ( n1612 & n2575 ) | ( ~n2573 & n2575 ) ;
  assign n2578 = n2577 ^ n2576 ^ 1'b0 ;
  assign n2579 = n1366 | n2578 ;
  assign n2583 = ( n899 & ~n1133 ) | ( n899 & n1466 ) | ( ~n1133 & n1466 ) ;
  assign n2584 = n2583 ^ x202 ^ 1'b0 ;
  assign n2585 = ( x28 & ~x59 ) | ( x28 & n2584 ) | ( ~x59 & n2584 ) ;
  assign n2580 = ( n440 & n772 ) | ( n440 & n1883 ) | ( n772 & n1883 ) ;
  assign n2581 = ( n367 & ~n526 ) | ( n367 & n2580 ) | ( ~n526 & n2580 ) ;
  assign n2582 = n450 & n2581 ;
  assign n2586 = n2585 ^ n2582 ^ 1'b0 ;
  assign n2587 = n2411 ^ n908 ^ 1'b0 ;
  assign n2588 = x171 & ~n2587 ;
  assign n2589 = x161 ^ x146 ^ x85 ;
  assign n2590 = n2589 ^ n1817 ^ n1693 ;
  assign n2596 = n871 & ~n919 ;
  assign n2597 = n2596 ^ n1288 ^ 1'b0 ;
  assign n2592 = n1402 ^ n1015 ^ x120 ;
  assign n2591 = ( ~x217 & n291 ) | ( ~x217 & n935 ) | ( n291 & n935 ) ;
  assign n2593 = n2592 ^ n2591 ^ n950 ;
  assign n2594 = n978 ^ n534 ^ 1'b0 ;
  assign n2595 = n2593 | n2594 ;
  assign n2598 = n2597 ^ n2595 ^ 1'b0 ;
  assign n2599 = ( ~n2588 & n2590 ) | ( ~n2588 & n2598 ) | ( n2590 & n2598 ) ;
  assign n2604 = x141 & n817 ;
  assign n2605 = ~n2518 & n2604 ;
  assign n2606 = ( n300 & n1851 ) | ( n300 & n2605 ) | ( n1851 & n2605 ) ;
  assign n2607 = n2606 ^ n573 ^ n528 ;
  assign n2600 = n1801 ^ x32 ^ 1'b0 ;
  assign n2601 = n1147 & n2600 ;
  assign n2602 = n2035 & n2212 ;
  assign n2603 = ~n2601 & n2602 ;
  assign n2608 = n2607 ^ n2603 ^ 1'b0 ;
  assign n2609 = n667 ^ x6 ^ 1'b0 ;
  assign n2610 = ~n1141 & n2609 ;
  assign n2611 = n1879 & ~n1914 ;
  assign n2612 = ~n1674 & n2611 ;
  assign n2613 = ( x222 & n856 ) | ( x222 & ~n1413 ) | ( n856 & ~n1413 ) ;
  assign n2614 = n455 ^ n315 ^ x128 ;
  assign n2615 = ( n380 & n487 ) | ( n380 & n2614 ) | ( n487 & n2614 ) ;
  assign n2616 = n2615 ^ n896 ^ 1'b0 ;
  assign n2617 = n2613 & ~n2616 ;
  assign n2618 = ( n1622 & ~n2612 ) | ( n1622 & n2617 ) | ( ~n2612 & n2617 ) ;
  assign n2619 = ( n848 & n1298 ) | ( n848 & n2156 ) | ( n1298 & n2156 ) ;
  assign n2620 = n2619 ^ n1844 ^ n350 ;
  assign n2621 = ( x15 & n1410 ) | ( x15 & ~n1944 ) | ( n1410 & ~n1944 ) ;
  assign n2622 = ( ~n677 & n1618 ) | ( ~n677 & n2621 ) | ( n1618 & n2621 ) ;
  assign n2623 = n300 | n1310 ;
  assign n2624 = n2623 ^ n1488 ^ 1'b0 ;
  assign n2625 = n758 ^ x156 ^ x126 ;
  assign n2626 = n2625 ^ n2366 ^ n1894 ;
  assign n2627 = n2626 ^ n1330 ^ n822 ;
  assign n2628 = x200 ^ x155 ^ 1'b0 ;
  assign n2629 = n422 & n2628 ;
  assign n2630 = ( n446 & ~n2305 ) | ( n446 & n2629 ) | ( ~n2305 & n2629 ) ;
  assign n2631 = ( n1012 & n1979 ) | ( n1012 & n2474 ) | ( n1979 & n2474 ) ;
  assign n2632 = n1980 ^ n1670 ^ n1140 ;
  assign n2633 = ( n594 & n2631 ) | ( n594 & ~n2632 ) | ( n2631 & ~n2632 ) ;
  assign n2634 = n2630 & ~n2633 ;
  assign n2643 = n2032 ^ n1568 ^ n1412 ;
  assign n2635 = n835 ^ n656 ^ 1'b0 ;
  assign n2636 = n2559 ^ n1217 ^ n507 ;
  assign n2637 = n2636 ^ n1420 ^ 1'b0 ;
  assign n2638 = n295 | n2637 ;
  assign n2639 = n1438 ^ n469 ^ 1'b0 ;
  assign n2640 = n326 & ~n2639 ;
  assign n2641 = ( ~n615 & n2638 ) | ( ~n615 & n2640 ) | ( n2638 & n2640 ) ;
  assign n2642 = n2635 & ~n2641 ;
  assign n2644 = n2643 ^ n2642 ^ 1'b0 ;
  assign n2645 = n1005 ^ n802 ^ n668 ;
  assign n2646 = n2645 ^ n1747 ^ n605 ;
  assign n2647 = n2646 ^ n1455 ^ 1'b0 ;
  assign n2648 = n2644 & ~n2647 ;
  assign n2649 = n2638 ^ n841 ^ n502 ;
  assign n2650 = x9 & n1701 ;
  assign n2651 = n2193 ^ n764 ^ x239 ;
  assign n2654 = n2080 ^ n801 ^ x130 ;
  assign n2652 = n1464 | n1757 ;
  assign n2653 = ~n1894 & n2652 ;
  assign n2655 = n2654 ^ n2653 ^ 1'b0 ;
  assign n2656 = ~n366 & n2655 ;
  assign n2657 = ( n1862 & ~n2545 ) | ( n1862 & n2656 ) | ( ~n2545 & n2656 ) ;
  assign n2658 = ( ~x104 & n378 ) | ( ~x104 & n634 ) | ( n378 & n634 ) ;
  assign n2659 = n2658 ^ n1979 ^ x160 ;
  assign n2660 = n2659 ^ n1391 ^ n838 ;
  assign n2661 = n1399 ^ n921 ^ x38 ;
  assign n2662 = ( ~n2631 & n2660 ) | ( ~n2631 & n2661 ) | ( n2660 & n2661 ) ;
  assign n2663 = x159 | n876 ;
  assign n2664 = ( n423 & ~n1012 ) | ( n423 & n2663 ) | ( ~n1012 & n2663 ) ;
  assign n2679 = ( n975 & ~n1091 ) | ( n975 & n1536 ) | ( ~n1091 & n1536 ) ;
  assign n2678 = ( ~n429 & n489 ) | ( ~n429 & n1670 ) | ( n489 & n1670 ) ;
  assign n2665 = n1397 ^ n971 ^ n299 ;
  assign n2666 = n2506 ^ n1689 ^ 1'b0 ;
  assign n2667 = x34 & ~n1842 ;
  assign n2668 = n2667 ^ n1697 ^ n1421 ;
  assign n2669 = n2615 | n2668 ;
  assign n2670 = n2669 ^ n1248 ^ 1'b0 ;
  assign n2672 = ~n379 & n2452 ;
  assign n2673 = ~x134 & n2672 ;
  assign n2674 = ( n1063 & n1246 ) | ( n1063 & ~n2673 ) | ( n1246 & ~n2673 ) ;
  assign n2671 = ~n371 & n1942 ;
  assign n2675 = n2674 ^ n2671 ^ 1'b0 ;
  assign n2676 = ( ~n2666 & n2670 ) | ( ~n2666 & n2675 ) | ( n2670 & n2675 ) ;
  assign n2677 = n2665 & ~n2676 ;
  assign n2680 = n2679 ^ n2678 ^ n2677 ;
  assign n2691 = n1244 ^ x206 ^ x11 ;
  assign n2692 = n2691 ^ n1266 ^ n320 ;
  assign n2688 = n890 ^ n886 ^ n624 ;
  assign n2687 = n1972 ^ n476 ^ x29 ;
  assign n2686 = x51 & ~n1846 ;
  assign n2689 = n2688 ^ n2687 ^ n2686 ;
  assign n2681 = ( x8 & n809 ) | ( x8 & n1670 ) | ( n809 & n1670 ) ;
  assign n2682 = n1402 | n2681 ;
  assign n2683 = n2535 & ~n2682 ;
  assign n2684 = ( ~n1972 & n2227 ) | ( ~n1972 & n2683 ) | ( n2227 & n2683 ) ;
  assign n2685 = ( n2251 & n2318 ) | ( n2251 & n2684 ) | ( n2318 & n2684 ) ;
  assign n2690 = n2689 ^ n2685 ^ n2565 ;
  assign n2693 = n2692 ^ n2690 ^ n492 ;
  assign n2694 = n1395 ^ n994 ^ x171 ;
  assign n2695 = ( x114 & n325 ) | ( x114 & n498 ) | ( n325 & n498 ) ;
  assign n2696 = n2695 ^ n2425 ^ 1'b0 ;
  assign n2697 = n2696 ^ n2355 ^ n1310 ;
  assign n2698 = n2694 & ~n2697 ;
  assign n2699 = n2698 ^ n2610 ^ 1'b0 ;
  assign n2704 = ~n1702 & n1869 ;
  assign n2702 = x253 & ~n2051 ;
  assign n2703 = n2702 ^ n492 ^ 1'b0 ;
  assign n2705 = n2704 ^ n2703 ^ n1215 ;
  assign n2700 = x3 & x24 ;
  assign n2701 = ~n1230 & n2700 ;
  assign n2706 = n2705 ^ n2701 ^ n1928 ;
  assign n2707 = n1604 ^ n1467 ^ n332 ;
  assign n2708 = n2502 ^ n1524 ^ n459 ;
  assign n2709 = n2707 & ~n2708 ;
  assign n2710 = ~n1408 & n2709 ;
  assign n2711 = n721 ^ n344 ^ n269 ;
  assign n2712 = ~n1511 & n2711 ;
  assign n2727 = n501 & n1164 ;
  assign n2728 = n1155 & n2727 ;
  assign n2724 = ( n653 & ~n894 ) | ( n653 & n1258 ) | ( ~n894 & n1258 ) ;
  assign n2725 = n2724 ^ n1728 ^ n1154 ;
  assign n2726 = n2725 ^ n264 ^ 1'b0 ;
  assign n2729 = n2728 ^ n2726 ^ n1564 ;
  assign n2714 = ( x152 & n257 ) | ( x152 & ~n812 ) | ( n257 & ~n812 ) ;
  assign n2713 = n1537 & n1668 ;
  assign n2715 = n2714 ^ n2713 ^ 1'b0 ;
  assign n2716 = n1616 ^ n904 ^ 1'b0 ;
  assign n2717 = ~n621 & n2716 ;
  assign n2718 = ( ~n1206 & n1343 ) | ( ~n1206 & n2717 ) | ( n1343 & n2717 ) ;
  assign n2719 = ( n485 & ~n868 ) | ( n485 & n2036 ) | ( ~n868 & n2036 ) ;
  assign n2720 = ( x169 & n2718 ) | ( x169 & n2719 ) | ( n2718 & n2719 ) ;
  assign n2721 = n2720 ^ n2334 ^ 1'b0 ;
  assign n2722 = ~n984 & n2721 ;
  assign n2723 = ~n2715 & n2722 ;
  assign n2730 = n2729 ^ n2723 ^ 1'b0 ;
  assign n2736 = n1382 ^ n667 ^ 1'b0 ;
  assign n2737 = n2736 ^ n2130 ^ 1'b0 ;
  assign n2731 = n1009 | n1504 ;
  assign n2732 = n2731 ^ n907 ^ 1'b0 ;
  assign n2733 = n2466 ^ n1290 ^ n795 ;
  assign n2734 = ~n2732 & n2733 ;
  assign n2735 = n2734 ^ n995 ^ 1'b0 ;
  assign n2738 = n2737 ^ n2735 ^ 1'b0 ;
  assign n2739 = x191 & ~n1206 ;
  assign n2741 = ( n278 & ~n944 ) | ( n278 & n1265 ) | ( ~n944 & n1265 ) ;
  assign n2740 = ( ~n295 & n1371 ) | ( ~n295 & n1873 ) | ( n1371 & n1873 ) ;
  assign n2742 = n2741 ^ n2740 ^ n2358 ;
  assign n2743 = n1412 ^ n984 ^ n576 ;
  assign n2744 = n1265 ^ n791 ^ 1'b0 ;
  assign n2745 = x93 & ~n2744 ;
  assign n2746 = ( n2737 & n2743 ) | ( n2737 & n2745 ) | ( n2743 & n2745 ) ;
  assign n2747 = n1243 ^ x77 ^ 1'b0 ;
  assign n2749 = ( ~n711 & n1338 ) | ( ~n711 & n2325 ) | ( n1338 & n2325 ) ;
  assign n2748 = x66 & n2499 ;
  assign n2750 = n2749 ^ n2748 ^ 1'b0 ;
  assign n2751 = n2750 ^ n2674 ^ 1'b0 ;
  assign n2754 = n2050 ^ x171 ^ 1'b0 ;
  assign n2752 = ( n415 & n1766 ) | ( n415 & ~n2182 ) | ( n1766 & ~n2182 ) ;
  assign n2753 = ( n759 & n1816 ) | ( n759 & n2752 ) | ( n1816 & n2752 ) ;
  assign n2755 = n2754 ^ n2753 ^ n2678 ;
  assign n2756 = ( ~n2747 & n2751 ) | ( ~n2747 & n2755 ) | ( n2751 & n2755 ) ;
  assign n2757 = n1191 ^ n505 ^ 1'b0 ;
  assign n2758 = ( x253 & n2397 ) | ( x253 & ~n2757 ) | ( n2397 & ~n2757 ) ;
  assign n2759 = n2323 ^ n652 ^ n529 ;
  assign n2760 = ( n458 & n825 ) | ( n458 & ~n2625 ) | ( n825 & ~n2625 ) ;
  assign n2761 = n2760 ^ n2218 ^ 1'b0 ;
  assign n2762 = x173 | n2761 ;
  assign n2763 = n2762 ^ n2614 ^ n979 ;
  assign n2764 = n2763 ^ n634 ^ n287 ;
  assign n2765 = n2764 ^ n2329 ^ n1151 ;
  assign n2766 = n2281 ^ n1299 ^ n452 ;
  assign n2769 = n1578 ^ n1100 ^ 1'b0 ;
  assign n2770 = n2520 | n2769 ;
  assign n2771 = ( n414 & n1276 ) | ( n414 & ~n2770 ) | ( n1276 & ~n2770 ) ;
  assign n2767 = ( ~n1302 & n1404 ) | ( ~n1302 & n2658 ) | ( n1404 & n2658 ) ;
  assign n2768 = ( x17 & ~n1724 ) | ( x17 & n2767 ) | ( ~n1724 & n2767 ) ;
  assign n2772 = n2771 ^ n2768 ^ 1'b0 ;
  assign n2773 = n2766 & ~n2772 ;
  assign n2774 = ( x173 & n639 ) | ( x173 & n1497 ) | ( n639 & n1497 ) ;
  assign n2775 = ( x107 & ~x220 ) | ( x107 & n571 ) | ( ~x220 & n571 ) ;
  assign n2776 = n720 & ~n822 ;
  assign n2777 = n2776 ^ n2358 ^ 1'b0 ;
  assign n2778 = ( ~n1366 & n2775 ) | ( ~n1366 & n2777 ) | ( n2775 & n2777 ) ;
  assign n2779 = ( ~n2176 & n2774 ) | ( ~n2176 & n2778 ) | ( n2774 & n2778 ) ;
  assign n2780 = n2089 ^ n1803 ^ n516 ;
  assign n2781 = ( n491 & n2715 ) | ( n491 & ~n2780 ) | ( n2715 & ~n2780 ) ;
  assign n2782 = ~n1165 & n2781 ;
  assign n2786 = ( n455 & n748 ) | ( n455 & ~n778 ) | ( n748 & ~n778 ) ;
  assign n2783 = n2581 ^ n1516 ^ 1'b0 ;
  assign n2784 = n421 & ~n2783 ;
  assign n2785 = n2784 ^ n1493 ^ n553 ;
  assign n2787 = n2786 ^ n2785 ^ n2019 ;
  assign n2788 = n2787 ^ n2476 ^ n2099 ;
  assign n2789 = ( x134 & ~n747 ) | ( x134 & n2788 ) | ( ~n747 & n2788 ) ;
  assign n2790 = n2784 ^ n2517 ^ 1'b0 ;
  assign n2791 = n289 & ~n2790 ;
  assign n2792 = ( x229 & n2752 ) | ( x229 & ~n2754 ) | ( n2752 & ~n2754 ) ;
  assign n2793 = ( n369 & n1050 ) | ( n369 & n1883 ) | ( n1050 & n1883 ) ;
  assign n2794 = ( n1488 & n2011 ) | ( n1488 & ~n2793 ) | ( n2011 & ~n2793 ) ;
  assign n2795 = ( x245 & ~n2536 ) | ( x245 & n2794 ) | ( ~n2536 & n2794 ) ;
  assign n2796 = ~n1363 & n2795 ;
  assign n2797 = n2792 & n2796 ;
  assign n2798 = n1014 ^ x89 ^ 1'b0 ;
  assign n2799 = n1603 & n2798 ;
  assign n2800 = ~n2548 & n2799 ;
  assign n2801 = n2089 ^ n1714 ^ 1'b0 ;
  assign n2802 = ( x213 & n582 ) | ( x213 & n2801 ) | ( n582 & n2801 ) ;
  assign n2803 = ( n880 & n1499 ) | ( n880 & n2259 ) | ( n1499 & n2259 ) ;
  assign n2804 = n2803 ^ n961 ^ 1'b0 ;
  assign n2805 = ~n1947 & n2804 ;
  assign n2806 = ~n726 & n2805 ;
  assign n2807 = n1907 & ~n2806 ;
  assign n2816 = ( x94 & n1108 ) | ( x94 & n1926 ) | ( n1108 & n1926 ) ;
  assign n2817 = n748 | n2816 ;
  assign n2818 = n2817 ^ n1784 ^ 1'b0 ;
  assign n2808 = n1392 & ~n1419 ;
  assign n2809 = n2808 ^ x66 ^ 1'b0 ;
  assign n2810 = n2809 ^ n1172 ^ 1'b0 ;
  assign n2811 = ( x209 & n1473 ) | ( x209 & n2200 ) | ( n1473 & n2200 ) ;
  assign n2812 = n2811 ^ n1414 ^ 1'b0 ;
  assign n2813 = x160 & ~n2812 ;
  assign n2814 = n2813 ^ n1078 ^ 1'b0 ;
  assign n2815 = ~n2810 & n2814 ;
  assign n2819 = n2818 ^ n2815 ^ n1711 ;
  assign n2820 = n2819 ^ n2232 ^ n1507 ;
  assign n2821 = n905 ^ n898 ^ 1'b0 ;
  assign n2822 = n2412 | n2821 ;
  assign n2823 = n2822 ^ n1192 ^ 1'b0 ;
  assign n2824 = n1390 ^ n1251 ^ x134 ;
  assign n2825 = n2176 & n2824 ;
  assign n2826 = n700 ^ n427 ^ 1'b0 ;
  assign n2827 = ( n1063 & n1707 ) | ( n1063 & ~n2826 ) | ( n1707 & ~n2826 ) ;
  assign n2828 = n2827 ^ n1372 ^ 1'b0 ;
  assign n2829 = n852 & n2158 ;
  assign n2830 = n901 & n2829 ;
  assign n2834 = ~n1653 & n1785 ;
  assign n2835 = n2834 ^ n1990 ^ 1'b0 ;
  assign n2836 = ( x46 & n807 ) | ( x46 & n2410 ) | ( n807 & n2410 ) ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2838 = n1076 | n2837 ;
  assign n2831 = x16 & n1981 ;
  assign n2832 = n2831 ^ n1778 ^ 1'b0 ;
  assign n2833 = ( n708 & n1979 ) | ( n708 & ~n2832 ) | ( n1979 & ~n2832 ) ;
  assign n2839 = n2838 ^ n2833 ^ n343 ;
  assign n2840 = ~n2012 & n2839 ;
  assign n2842 = n375 ^ x202 ^ x71 ;
  assign n2841 = n2754 ^ n563 ^ n405 ;
  assign n2843 = n2842 ^ n2841 ^ n603 ;
  assign n2844 = ( x186 & x227 ) | ( x186 & ~n2843 ) | ( x227 & ~n2843 ) ;
  assign n2845 = n2162 ^ n1945 ^ n917 ;
  assign n2846 = ( n1078 & n1183 ) | ( n1078 & ~n1188 ) | ( n1183 & ~n1188 ) ;
  assign n2847 = ( n1994 & n2845 ) | ( n1994 & n2846 ) | ( n2845 & n2846 ) ;
  assign n2848 = n375 | n2004 ;
  assign n2851 = x91 & n566 ;
  assign n2852 = n1855 & n2851 ;
  assign n2849 = ( x62 & x105 ) | ( x62 & ~x185 ) | ( x105 & ~x185 ) ;
  assign n2850 = ( n1471 & ~n1515 ) | ( n1471 & n2849 ) | ( ~n1515 & n2849 ) ;
  assign n2853 = n2852 ^ n2850 ^ n1238 ;
  assign n2854 = ( n987 & n2140 ) | ( n987 & ~n2853 ) | ( n2140 & ~n2853 ) ;
  assign n2855 = n1820 ^ n847 ^ 1'b0 ;
  assign n2856 = n2854 & ~n2855 ;
  assign n2857 = n349 & n1576 ;
  assign n2858 = x134 & n2857 ;
  assign n2859 = n2858 ^ n1592 ^ n1387 ;
  assign n2860 = n1893 ^ n997 ^ n801 ;
  assign n2861 = ~n389 & n2860 ;
  assign n2862 = n2601 ^ n2017 ^ n1379 ;
  assign n2863 = ( n971 & n2720 ) | ( n971 & n2758 ) | ( n2720 & n2758 ) ;
  assign n2864 = ( n1455 & ~n2032 ) | ( n1455 & n2729 ) | ( ~n2032 & n2729 ) ;
  assign n2865 = ( ~x67 & n369 ) | ( ~x67 & n1066 ) | ( n369 & n1066 ) ;
  assign n2866 = ( x173 & n1062 ) | ( x173 & n2865 ) | ( n1062 & n2865 ) ;
  assign n2867 = x187 | n359 ;
  assign n2868 = n2867 ^ n1390 ^ n410 ;
  assign n2869 = n2868 ^ n1118 ^ n513 ;
  assign n2883 = ( ~x206 & n722 ) | ( ~x206 & n2401 ) | ( n722 & n2401 ) ;
  assign n2884 = n2883 ^ n1100 ^ n877 ;
  assign n2874 = x17 & ~n1124 ;
  assign n2875 = ~n1842 & n2874 ;
  assign n2870 = n1689 ^ x19 ^ 1'b0 ;
  assign n2871 = n1046 ^ n597 ^ n425 ;
  assign n2872 = n2871 ^ n1009 ^ n802 ;
  assign n2873 = n2870 | n2872 ;
  assign n2876 = n2875 ^ n2873 ^ 1'b0 ;
  assign n2877 = n486 ^ n438 ^ x125 ;
  assign n2878 = n1495 & ~n2877 ;
  assign n2879 = n649 | n2878 ;
  assign n2880 = n1716 & ~n2879 ;
  assign n2881 = ( ~n672 & n2876 ) | ( ~n672 & n2880 ) | ( n2876 & n2880 ) ;
  assign n2882 = ( n950 & ~n1389 ) | ( n950 & n2881 ) | ( ~n1389 & n2881 ) ;
  assign n2885 = n2884 ^ n2882 ^ n2390 ;
  assign n2896 = n2133 ^ n385 ^ x65 ;
  assign n2894 = n1962 ^ n1510 ^ 1'b0 ;
  assign n2895 = ( n1663 & n2837 ) | ( n1663 & ~n2894 ) | ( n2837 & ~n2894 ) ;
  assign n2890 = ( ~n664 & n1006 ) | ( ~n664 & n1141 ) | ( n1006 & n1141 ) ;
  assign n2886 = ( n317 & ~n462 ) | ( n317 & n778 ) | ( ~n462 & n778 ) ;
  assign n2887 = x6 & ~n2886 ;
  assign n2888 = n2887 ^ n626 ^ x184 ;
  assign n2889 = n1948 | n2888 ;
  assign n2891 = n2890 ^ n2889 ^ 1'b0 ;
  assign n2892 = n268 | n2891 ;
  assign n2893 = n1685 & ~n2892 ;
  assign n2897 = n2896 ^ n2895 ^ n2893 ;
  assign n2898 = x245 ^ x32 ^ 1'b0 ;
  assign n2899 = x114 & n2898 ;
  assign n2900 = n487 ^ x84 ^ 1'b0 ;
  assign n2901 = n676 | n2900 ;
  assign n2902 = n2901 ^ n1005 ^ 1'b0 ;
  assign n2903 = n2033 | n2902 ;
  assign n2904 = n2903 ^ n2643 ^ n2016 ;
  assign n2905 = n2899 & ~n2904 ;
  assign n2923 = x177 ^ x129 ^ 1'b0 ;
  assign n2917 = n380 | n1521 ;
  assign n2918 = n2917 ^ n498 ^ 1'b0 ;
  assign n2919 = n944 & n2360 ;
  assign n2920 = ~n2918 & n2919 ;
  assign n2921 = n2920 ^ n393 ^ 1'b0 ;
  assign n2922 = n1238 & n2921 ;
  assign n2906 = n1419 | n1808 ;
  assign n2907 = n2906 ^ n1114 ^ 1'b0 ;
  assign n2908 = x88 & ~n1627 ;
  assign n2909 = ~x157 & n2908 ;
  assign n2910 = n2909 ^ n1093 ^ 1'b0 ;
  assign n2911 = n1282 ^ n380 ^ x184 ;
  assign n2912 = ( n318 & n641 ) | ( n318 & ~n2911 ) | ( n641 & ~n2911 ) ;
  assign n2913 = n2912 ^ n1544 ^ n382 ;
  assign n2914 = ( ~n1288 & n2910 ) | ( ~n1288 & n2913 ) | ( n2910 & n2913 ) ;
  assign n2915 = n356 & ~n2914 ;
  assign n2916 = n2907 & n2915 ;
  assign n2924 = n2923 ^ n2922 ^ n2916 ;
  assign n2925 = ( n1070 & n1126 ) | ( n1070 & ~n1449 ) | ( n1126 & ~n1449 ) ;
  assign n2926 = n2925 ^ n2905 ^ x92 ;
  assign n2927 = n2922 ^ n1137 ^ n574 ;
  assign n2928 = ( ~n856 & n1456 ) | ( ~n856 & n2927 ) | ( n1456 & n2927 ) ;
  assign n2929 = n2928 ^ n2392 ^ n259 ;
  assign n2930 = ( x75 & x114 ) | ( x75 & ~n466 ) | ( x114 & ~n466 ) ;
  assign n2931 = n706 | n756 ;
  assign n2932 = n2931 ^ n579 ^ n427 ;
  assign n2933 = ( ~n2490 & n2930 ) | ( ~n2490 & n2932 ) | ( n2930 & n2932 ) ;
  assign n2934 = ( x211 & ~n461 ) | ( x211 & n966 ) | ( ~n461 & n966 ) ;
  assign n2935 = n1319 ^ n481 ^ 1'b0 ;
  assign n2936 = ~n1663 & n2935 ;
  assign n2937 = n2934 & n2936 ;
  assign n2938 = n2853 ^ n2017 ^ 1'b0 ;
  assign n2939 = n723 & n2938 ;
  assign n2944 = n781 | n948 ;
  assign n2945 = n2944 ^ n1796 ^ 1'b0 ;
  assign n2940 = ~n308 & n854 ;
  assign n2941 = n2940 ^ n376 ^ 1'b0 ;
  assign n2942 = n2941 ^ n476 ^ x36 ;
  assign n2943 = n2942 ^ n2499 ^ n2488 ;
  assign n2946 = n2945 ^ n2943 ^ 1'b0 ;
  assign n2947 = n1434 & ~n2946 ;
  assign n2948 = ( ~n871 & n1192 ) | ( ~n871 & n2277 ) | ( n1192 & n2277 ) ;
  assign n2949 = n2948 ^ n797 ^ 1'b0 ;
  assign n2950 = ( x146 & ~n1365 ) | ( x146 & n2259 ) | ( ~n1365 & n2259 ) ;
  assign n2951 = n2950 ^ n2844 ^ n368 ;
  assign n2952 = n2007 ^ n1534 ^ n374 ;
  assign n2953 = n1141 ^ n1129 ^ x157 ;
  assign n2954 = n2953 ^ n2077 ^ 1'b0 ;
  assign n2955 = n656 | n2954 ;
  assign n2956 = n2952 | n2955 ;
  assign n2959 = n605 & n1913 ;
  assign n2960 = n2959 ^ n750 ^ 1'b0 ;
  assign n2958 = n1375 & n2452 ;
  assign n2961 = n2960 ^ n2958 ^ n286 ;
  assign n2957 = ( ~n955 & n2092 ) | ( ~n955 & n2747 ) | ( n2092 & n2747 ) ;
  assign n2962 = n2961 ^ n2957 ^ n771 ;
  assign n2963 = n2962 ^ n270 ^ x89 ;
  assign n2964 = n1957 ^ n1269 ^ n890 ;
  assign n2965 = ~n2300 & n2964 ;
  assign n2966 = n1422 ^ n1070 ^ 1'b0 ;
  assign n2967 = n2074 ^ n952 ^ n795 ;
  assign n2968 = n1488 & ~n1929 ;
  assign n2969 = ~n1924 & n2968 ;
  assign n2970 = n2967 & ~n2969 ;
  assign n2971 = ~n2966 & n2970 ;
  assign n2972 = n1312 & ~n2678 ;
  assign n2973 = ~n2152 & n2972 ;
  assign n2975 = n2194 ^ x2 ^ 1'b0 ;
  assign n2974 = n747 | n2547 ;
  assign n2976 = n2975 ^ n2974 ^ x206 ;
  assign n2977 = n2399 ^ n1130 ^ n1066 ;
  assign n2978 = n672 ^ n488 ^ 1'b0 ;
  assign n2981 = n2223 ^ n1147 ^ n640 ;
  assign n2982 = n422 & n1159 ;
  assign n2983 = ~n2981 & n2982 ;
  assign n2984 = n2983 ^ n2527 ^ n1155 ;
  assign n2979 = ~n345 & n1612 ;
  assign n2980 = n2979 ^ n1951 ^ x89 ;
  assign n2985 = n2984 ^ n2980 ^ n911 ;
  assign n2986 = n2066 ^ x70 ^ 1'b0 ;
  assign n2987 = n2922 & ~n2986 ;
  assign n2995 = ( n330 & n341 ) | ( n330 & n390 ) | ( n341 & n390 ) ;
  assign n2996 = n2995 ^ n273 ^ x49 ;
  assign n2991 = n720 ^ x61 ^ 1'b0 ;
  assign n2992 = x131 & n2991 ;
  assign n2993 = ( ~n373 & n1261 ) | ( ~n373 & n2992 ) | ( n1261 & n2992 ) ;
  assign n2994 = n2993 ^ n754 ^ n500 ;
  assign n2997 = n2996 ^ n2994 ^ n408 ;
  assign n2989 = n1962 ^ n1599 ^ n866 ;
  assign n2990 = n2989 ^ n930 ^ n352 ;
  assign n2998 = n2997 ^ n2990 ^ n2482 ;
  assign n2988 = ( n641 & n726 ) | ( n641 & ~n894 ) | ( n726 & ~n894 ) ;
  assign n2999 = n2998 ^ n2988 ^ 1'b0 ;
  assign n3000 = n779 & n1534 ;
  assign n3001 = n3000 ^ n1324 ^ 1'b0 ;
  assign n3002 = ~n1426 & n3001 ;
  assign n3003 = ~n2835 & n3002 ;
  assign n3004 = n2459 & n3003 ;
  assign n3005 = n1952 ^ n566 ^ n486 ;
  assign n3006 = n3005 ^ n2326 ^ n645 ;
  assign n3007 = n3006 ^ n2989 ^ n2449 ;
  assign n3008 = n1988 ^ n1373 ^ x100 ;
  assign n3009 = ( x189 & ~n1709 ) | ( x189 & n3008 ) | ( ~n1709 & n3008 ) ;
  assign n3010 = n924 ^ n840 ^ x253 ;
  assign n3011 = n3010 ^ n2850 ^ 1'b0 ;
  assign n3012 = x122 & ~n3011 ;
  assign n3013 = ~n300 & n3012 ;
  assign n3014 = n3013 ^ n2601 ^ 1'b0 ;
  assign n3015 = ( ~x105 & n373 ) | ( ~x105 & n997 ) | ( n373 & n997 ) ;
  assign n3016 = ( n2187 & n2755 ) | ( n2187 & ~n3015 ) | ( n2755 & ~n3015 ) ;
  assign n3017 = n2217 ^ n1568 ^ 1'b0 ;
  assign n3018 = ( n488 & n1582 ) | ( n488 & n2001 ) | ( n1582 & n2001 ) ;
  assign n3019 = ( ~n552 & n3017 ) | ( ~n552 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3024 = n2466 ^ n2170 ^ n401 ;
  assign n3025 = n2794 ^ n2004 ^ x113 ;
  assign n3026 = n1074 & n2542 ;
  assign n3027 = ( ~n3024 & n3025 ) | ( ~n3024 & n3026 ) | ( n3025 & n3026 ) ;
  assign n3020 = n509 & ~n566 ;
  assign n3021 = n1061 & n3020 ;
  assign n3022 = ~n2022 & n3021 ;
  assign n3023 = n2315 & n3022 ;
  assign n3028 = n3027 ^ n3023 ^ x248 ;
  assign n3029 = n2526 ^ n866 ^ x174 ;
  assign n3030 = ( n346 & n591 ) | ( n346 & ~n3029 ) | ( n591 & ~n3029 ) ;
  assign n3031 = n275 & n605 ;
  assign n3032 = ~n632 & n3031 ;
  assign n3033 = n975 & n3032 ;
  assign n3034 = n2450 & n3033 ;
  assign n3035 = ( n327 & n3030 ) | ( n327 & n3034 ) | ( n3030 & n3034 ) ;
  assign n3036 = ~n525 & n1189 ;
  assign n3039 = n1585 ^ n742 ^ 1'b0 ;
  assign n3037 = n1210 ^ n944 ^ n364 ;
  assign n3038 = n3037 ^ n2659 ^ x107 ;
  assign n3040 = n3039 ^ n3038 ^ n1354 ;
  assign n3041 = n619 & n3040 ;
  assign n3042 = n3041 ^ n2189 ^ 1'b0 ;
  assign n3043 = n1362 ^ n1252 ^ n421 ;
  assign n3044 = ( n777 & ~n1555 ) | ( n777 & n3043 ) | ( ~n1555 & n3043 ) ;
  assign n3045 = ( x191 & n326 ) | ( x191 & ~n3044 ) | ( n326 & ~n3044 ) ;
  assign n3046 = n3045 ^ n963 ^ n527 ;
  assign n3047 = ~n1971 & n2220 ;
  assign n3048 = n3047 ^ x227 ^ 1'b0 ;
  assign n3049 = ( n1012 & n1302 ) | ( n1012 & ~n3048 ) | ( n1302 & ~n3048 ) ;
  assign n3050 = n706 | n1848 ;
  assign n3051 = ( n2427 & n3049 ) | ( n2427 & ~n3050 ) | ( n3049 & ~n3050 ) ;
  assign n3052 = n1688 ^ n636 ^ n384 ;
  assign n3053 = n1301 ^ n910 ^ n326 ;
  assign n3054 = n3053 ^ n2613 ^ n930 ;
  assign n3055 = n3054 ^ n1595 ^ 1'b0 ;
  assign n3056 = n3052 & n3055 ;
  assign n3057 = n696 & n1257 ;
  assign n3058 = n3057 ^ x90 ^ 1'b0 ;
  assign n3059 = ( n501 & ~n1472 ) | ( n501 & n3058 ) | ( ~n1472 & n3058 ) ;
  assign n3060 = n3059 ^ n1487 ^ n1295 ;
  assign n3061 = n2324 ^ n1080 ^ n471 ;
  assign n3062 = ( x245 & n1188 ) | ( x245 & ~n3061 ) | ( n1188 & ~n3061 ) ;
  assign n3063 = n3062 ^ n1674 ^ 1'b0 ;
  assign n3070 = n396 & ~n1999 ;
  assign n3071 = ~n2607 & n3070 ;
  assign n3072 = n3071 ^ x126 ^ 1'b0 ;
  assign n3065 = ~n574 & n1373 ;
  assign n3064 = ( ~x106 & n1402 ) | ( ~x106 & n1449 ) | ( n1402 & n1449 ) ;
  assign n3066 = n3065 ^ n3064 ^ n2199 ;
  assign n3067 = n3066 ^ n2803 ^ n485 ;
  assign n3068 = ~n2166 & n3067 ;
  assign n3069 = n2348 | n3068 ;
  assign n3073 = n3072 ^ n3069 ^ 1'b0 ;
  assign n3074 = x250 & n1784 ;
  assign n3075 = n1080 ^ x64 ^ 1'b0 ;
  assign n3076 = n3074 & ~n3075 ;
  assign n3077 = n2714 ^ n2280 ^ 1'b0 ;
  assign n3080 = n1344 ^ n562 ^ 1'b0 ;
  assign n3081 = n1098 & ~n3080 ;
  assign n3082 = x167 & ~n3081 ;
  assign n3083 = n805 & n3082 ;
  assign n3084 = n3083 ^ n469 ^ 1'b0 ;
  assign n3078 = n3039 ^ n2990 ^ n1774 ;
  assign n3079 = n478 | n3078 ;
  assign n3085 = n3084 ^ n3079 ^ 1'b0 ;
  assign n3086 = n2581 ^ n1898 ^ n1380 ;
  assign n3087 = n3086 ^ n2509 ^ 1'b0 ;
  assign n3088 = n2757 & ~n3087 ;
  assign n3089 = n3088 ^ n3060 ^ n1601 ;
  assign n3090 = n449 & ~n902 ;
  assign n3091 = n3090 ^ n1790 ^ x56 ;
  assign n3092 = n3091 ^ n1121 ^ n304 ;
  assign n3094 = ( ~n616 & n1434 ) | ( ~n616 & n1750 ) | ( n1434 & n1750 ) ;
  assign n3095 = ~n1891 & n3094 ;
  assign n3096 = n3095 ^ n1134 ^ 1'b0 ;
  assign n3093 = n1402 | n2113 ;
  assign n3097 = n3096 ^ n3093 ^ 1'b0 ;
  assign n3098 = n3097 ^ n2358 ^ 1'b0 ;
  assign n3099 = n2803 ^ n914 ^ n871 ;
  assign n3100 = n3099 ^ n1578 ^ 1'b0 ;
  assign n3101 = n945 | n3100 ;
  assign n3102 = ( n1155 & n1454 ) | ( n1155 & ~n3101 ) | ( n1454 & ~n3101 ) ;
  assign n3103 = n1747 ^ n929 ^ x9 ;
  assign n3104 = ( n2414 & ~n2967 ) | ( n2414 & n3103 ) | ( ~n2967 & n3103 ) ;
  assign n3105 = x129 & ~n3104 ;
  assign n3106 = n3105 ^ n1576 ^ 1'b0 ;
  assign n3107 = x219 & ~n2539 ;
  assign n3108 = ( n669 & n3078 ) | ( n669 & n3107 ) | ( n3078 & n3107 ) ;
  assign n3109 = n764 | n2875 ;
  assign n3110 = n2014 ^ n1339 ^ n409 ;
  assign n3111 = ( n513 & n876 ) | ( n513 & n3110 ) | ( n876 & n3110 ) ;
  assign n3112 = n317 & ~n3111 ;
  assign n3113 = ~n2927 & n3112 ;
  assign n3116 = ( x240 & n350 ) | ( x240 & n452 ) | ( n350 & n452 ) ;
  assign n3114 = ~n595 & n1583 ;
  assign n3115 = n3114 ^ n922 ^ 1'b0 ;
  assign n3117 = n3116 ^ n3115 ^ n1207 ;
  assign n3118 = n498 & n2867 ;
  assign n3119 = ( n3113 & ~n3117 ) | ( n3113 & n3118 ) | ( ~n3117 & n3118 ) ;
  assign n3120 = n327 | n1705 ;
  assign n3121 = n3120 ^ n2696 ^ 1'b0 ;
  assign n3122 = n2613 & n3121 ;
  assign n3123 = ~n736 & n3122 ;
  assign n3124 = n1626 & n3123 ;
  assign n3128 = n3115 ^ n2568 ^ x21 ;
  assign n3125 = ~n617 & n1250 ;
  assign n3126 = n261 & ~n3125 ;
  assign n3127 = ( n1012 & n2245 ) | ( n1012 & n3126 ) | ( n2245 & n3126 ) ;
  assign n3129 = n3128 ^ n3127 ^ 1'b0 ;
  assign n3130 = n1153 ^ x161 ^ x49 ;
  assign n3131 = n3130 ^ n1568 ^ x193 ;
  assign n3132 = n3131 ^ n2763 ^ n813 ;
  assign n3133 = n1031 ^ n962 ^ 1'b0 ;
  assign n3134 = n680 | n3133 ;
  assign n3135 = n3134 ^ n1168 ^ x167 ;
  assign n3136 = n3132 | n3135 ;
  assign n3137 = ( ~n562 & n1695 ) | ( ~n562 & n3136 ) | ( n1695 & n3136 ) ;
  assign n3138 = ( x228 & n534 ) | ( x228 & n2183 ) | ( n534 & n2183 ) ;
  assign n3139 = ( n364 & ~n458 ) | ( n364 & n882 ) | ( ~n458 & n882 ) ;
  assign n3140 = n3138 & ~n3139 ;
  assign n3141 = n3140 ^ n621 ^ 1'b0 ;
  assign n3142 = n2357 & ~n3134 ;
  assign n3143 = ( x213 & n1223 ) | ( x213 & ~n1231 ) | ( n1223 & ~n1231 ) ;
  assign n3144 = n1093 ^ x75 ^ 1'b0 ;
  assign n3145 = ( n719 & ~n3143 ) | ( n719 & n3144 ) | ( ~n3143 & n3144 ) ;
  assign n3146 = n3145 ^ n2296 ^ n786 ;
  assign n3147 = ( ~n928 & n2436 ) | ( ~n928 & n2454 ) | ( n2436 & n2454 ) ;
  assign n3148 = n2324 ^ n526 ^ 1'b0 ;
  assign n3149 = n3147 & n3148 ;
  assign n3150 = n283 ^ x244 ^ x34 ;
  assign n3151 = ( ~x164 & n478 ) | ( ~x164 & n3150 ) | ( n478 & n3150 ) ;
  assign n3152 = n3151 ^ x220 ^ x212 ;
  assign n3154 = n550 ^ x163 ^ x91 ;
  assign n3153 = x232 & n1869 ;
  assign n3155 = n3154 ^ n3153 ^ 1'b0 ;
  assign n3156 = n3155 ^ n3117 ^ 1'b0 ;
  assign n3157 = ( n833 & n3152 ) | ( n833 & n3156 ) | ( n3152 & n3156 ) ;
  assign n3158 = n1523 ^ n416 ^ x200 ;
  assign n3159 = ~n1564 & n1728 ;
  assign n3160 = n505 & n3159 ;
  assign n3161 = ( n2214 & ~n3158 ) | ( n2214 & n3160 ) | ( ~n3158 & n3160 ) ;
  assign n3162 = n3049 ^ n2157 ^ n1976 ;
  assign n3163 = ( ~n279 & n1381 ) | ( ~n279 & n2064 ) | ( n1381 & n2064 ) ;
  assign n3164 = n973 ^ n856 ^ n631 ;
  assign n3165 = x114 & n1108 ;
  assign n3166 = n3165 ^ n1336 ^ 1'b0 ;
  assign n3167 = n3166 ^ n2922 ^ n993 ;
  assign n3168 = n3167 ^ n1693 ^ 1'b0 ;
  assign n3169 = ~n3164 & n3168 ;
  assign n3170 = n3169 ^ n2213 ^ n1141 ;
  assign n3171 = ( n2011 & ~n3163 ) | ( n2011 & n3170 ) | ( ~n3163 & n3170 ) ;
  assign n3172 = n604 ^ n373 ^ 1'b0 ;
  assign n3173 = x56 & ~n3172 ;
  assign n3174 = n3173 ^ x98 ^ 1'b0 ;
  assign n3175 = n3171 & n3174 ;
  assign n3176 = n1321 ^ n770 ^ 1'b0 ;
  assign n3177 = n1016 | n2774 ;
  assign n3178 = n3177 ^ n1366 ^ 1'b0 ;
  assign n3179 = n1893 | n3178 ;
  assign n3180 = n2017 | n3179 ;
  assign n3181 = n3180 ^ n2355 ^ 1'b0 ;
  assign n3182 = ( ~n444 & n790 ) | ( ~n444 & n3181 ) | ( n790 & n3181 ) ;
  assign n3187 = n2285 ^ n864 ^ 1'b0 ;
  assign n3188 = n522 & n3187 ;
  assign n3183 = n2992 & n3150 ;
  assign n3184 = n3183 ^ n503 ^ 1'b0 ;
  assign n3185 = n3184 ^ n2836 ^ n2594 ;
  assign n3186 = n501 | n3185 ;
  assign n3189 = n3188 ^ n3186 ^ 1'b0 ;
  assign n3190 = n2057 ^ n815 ^ n326 ;
  assign n3191 = x34 | n259 ;
  assign n3192 = ~n706 & n3191 ;
  assign n3193 = ( ~n818 & n1655 ) | ( ~n818 & n3192 ) | ( n1655 & n3192 ) ;
  assign n3194 = x109 & ~n3193 ;
  assign n3195 = n3194 ^ n534 ^ 1'b0 ;
  assign n3207 = n2151 ^ n1457 ^ 1'b0 ;
  assign n3203 = n1735 ^ n1194 ^ x219 ;
  assign n3204 = n3203 ^ n344 ^ 1'b0 ;
  assign n3205 = n3204 ^ n422 ^ n290 ;
  assign n3206 = ( ~n774 & n1222 ) | ( ~n774 & n3205 ) | ( n1222 & n3205 ) ;
  assign n3196 = n983 ^ n640 ^ x113 ;
  assign n3197 = n2993 & n3002 ;
  assign n3198 = n3196 & n3197 ;
  assign n3199 = ~n1709 & n2711 ;
  assign n3200 = n825 & n3199 ;
  assign n3201 = n3200 ^ n2684 ^ 1'b0 ;
  assign n3202 = n3198 | n3201 ;
  assign n3208 = n3207 ^ n3206 ^ n3202 ;
  assign n3217 = n2190 ^ n1591 ^ n353 ;
  assign n3210 = ( x54 & ~n594 ) | ( x54 & n628 ) | ( ~n594 & n628 ) ;
  assign n3211 = n3210 ^ n1267 ^ n324 ;
  assign n3212 = n1357 | n2123 ;
  assign n3213 = ( n759 & n3039 ) | ( n759 & ~n3212 ) | ( n3039 & ~n3212 ) ;
  assign n3214 = n1921 | n3213 ;
  assign n3215 = n3211 & n3214 ;
  assign n3216 = n1925 & n3215 ;
  assign n3209 = n2722 ^ x227 ^ x0 ;
  assign n3218 = n3217 ^ n3216 ^ n3209 ;
  assign n3219 = ( ~x0 & n572 ) | ( ~x0 & n1883 ) | ( n572 & n1883 ) ;
  assign n3220 = n2927 ^ n2244 ^ 1'b0 ;
  assign n3222 = n1855 & ~n2358 ;
  assign n3221 = n1162 & n3196 ;
  assign n3223 = n3222 ^ n3221 ^ 1'b0 ;
  assign n3224 = n2185 ^ n1612 ^ 1'b0 ;
  assign n3225 = n2614 & n3224 ;
  assign n3226 = n3188 ^ n1282 ^ n455 ;
  assign n3227 = n919 & ~n1378 ;
  assign n3228 = ( ~n883 & n1434 ) | ( ~n883 & n3227 ) | ( n1434 & n3227 ) ;
  assign n3229 = ( n2461 & n3226 ) | ( n2461 & n3228 ) | ( n3226 & n3228 ) ;
  assign n3230 = ( n1331 & ~n3225 ) | ( n1331 & n3229 ) | ( ~n3225 & n3229 ) ;
  assign n3231 = ( n846 & n1894 ) | ( n846 & n3230 ) | ( n1894 & n3230 ) ;
  assign n3235 = n505 ^ n296 ^ x111 ;
  assign n3236 = n2032 ^ x111 ^ 1'b0 ;
  assign n3237 = n3236 ^ n1592 ^ 1'b0 ;
  assign n3238 = n3235 & n3237 ;
  assign n3239 = n784 ^ n456 ^ 1'b0 ;
  assign n3240 = ~n3238 & n3239 ;
  assign n3232 = n1332 ^ x141 ^ 1'b0 ;
  assign n3233 = n3232 ^ n1463 ^ 1'b0 ;
  assign n3234 = n1012 & n3233 ;
  assign n3241 = n3240 ^ n3234 ^ 1'b0 ;
  assign n3242 = n2137 & ~n2466 ;
  assign n3252 = x143 & ~n495 ;
  assign n3253 = n3252 ^ n894 ^ 1'b0 ;
  assign n3254 = ~n2466 & n3253 ;
  assign n3249 = ( x218 & n496 ) | ( x218 & n794 ) | ( n496 & n794 ) ;
  assign n3248 = n396 & ~n758 ;
  assign n3243 = x137 & ~n1437 ;
  assign n3244 = n3243 ^ x182 ^ 1'b0 ;
  assign n3245 = n1570 | n2760 ;
  assign n3246 = n3244 | n3245 ;
  assign n3247 = n3246 ^ n1456 ^ 1'b0 ;
  assign n3250 = n3249 ^ n3248 ^ n3247 ;
  assign n3251 = n1212 & ~n3250 ;
  assign n3255 = n3254 ^ n3251 ^ n3192 ;
  assign n3257 = ( ~x40 & n538 ) | ( ~x40 & n2841 ) | ( n538 & n2841 ) ;
  assign n3256 = n393 | n2272 ;
  assign n3258 = n3257 ^ n3256 ^ 1'b0 ;
  assign n3259 = x204 & n3258 ;
  assign n3260 = n1853 ^ x245 ^ x29 ;
  assign n3261 = n3260 ^ n1663 ^ n1269 ;
  assign n3262 = ( x146 & x252 ) | ( x146 & ~n275 ) | ( x252 & ~n275 ) ;
  assign n3263 = x37 & n3262 ;
  assign n3264 = ( ~n2718 & n3261 ) | ( ~n2718 & n3263 ) | ( n3261 & n3263 ) ;
  assign n3269 = n924 & n1524 ;
  assign n3265 = x155 & ~n1485 ;
  assign n3266 = n818 & n1896 ;
  assign n3267 = n3266 ^ n2743 ^ n1019 ;
  assign n3268 = ( n1358 & ~n3265 ) | ( n1358 & n3267 ) | ( ~n3265 & n3267 ) ;
  assign n3270 = n3269 ^ n3268 ^ n825 ;
  assign n3271 = ( x42 & n471 ) | ( x42 & n3144 ) | ( n471 & n3144 ) ;
  assign n3272 = n3271 ^ n1177 ^ x111 ;
  assign n3273 = n3272 ^ n1214 ^ 1'b0 ;
  assign n3274 = ~n3270 & n3273 ;
  assign n3275 = n2937 ^ n2579 ^ n1920 ;
  assign n3276 = ( ~x124 & n1481 ) | ( ~x124 & n1734 ) | ( n1481 & n1734 ) ;
  assign n3277 = x113 & ~n849 ;
  assign n3278 = n3276 & n3277 ;
  assign n3279 = ( x42 & ~n2666 ) | ( x42 & n2777 ) | ( ~n2666 & n2777 ) ;
  assign n3280 = ( x21 & ~n357 ) | ( x21 & n1544 ) | ( ~n357 & n1544 ) ;
  assign n3281 = n3280 ^ n2125 ^ x135 ;
  assign n3285 = ( n677 & n1359 ) | ( n677 & n1740 ) | ( n1359 & n1740 ) ;
  assign n3282 = n2533 ^ n2113 ^ n1080 ;
  assign n3283 = n2256 | n3282 ;
  assign n3284 = n3283 ^ n1753 ^ 1'b0 ;
  assign n3286 = n3285 ^ n3284 ^ n2822 ;
  assign n3288 = n3167 ^ n1120 ^ x176 ;
  assign n3289 = ~n1948 & n2967 ;
  assign n3290 = n3288 & n3289 ;
  assign n3287 = ( n578 & n1155 ) | ( n578 & n1981 ) | ( n1155 & n1981 ) ;
  assign n3291 = n3290 ^ n3287 ^ 1'b0 ;
  assign n3292 = ( ~n430 & n930 ) | ( ~n430 & n2909 ) | ( n930 & n2909 ) ;
  assign n3293 = ( n326 & n877 ) | ( n326 & n942 ) | ( n877 & n942 ) ;
  assign n3294 = ( n2079 & n3292 ) | ( n2079 & n3293 ) | ( n3292 & n3293 ) ;
  assign n3306 = ( n1395 & n1498 ) | ( n1395 & n1892 ) | ( n1498 & n1892 ) ;
  assign n3295 = x178 & ~n1240 ;
  assign n3296 = ~x210 & n3295 ;
  assign n3297 = n1730 ^ n476 ^ 1'b0 ;
  assign n3298 = x188 & n3297 ;
  assign n3299 = ( n345 & ~n1151 ) | ( n345 & n1358 ) | ( ~n1151 & n1358 ) ;
  assign n3300 = ( n3296 & n3298 ) | ( n3296 & ~n3299 ) | ( n3298 & ~n3299 ) ;
  assign n3301 = ( n906 & n2708 ) | ( n906 & ~n3300 ) | ( n2708 & ~n3300 ) ;
  assign n3302 = x113 & ~n527 ;
  assign n3303 = n3302 ^ x38 ^ 1'b0 ;
  assign n3304 = n3303 ^ n1276 ^ 1'b0 ;
  assign n3305 = ~n3301 & n3304 ;
  assign n3307 = n3306 ^ n3305 ^ 1'b0 ;
  assign n3308 = ( ~x12 & x115 ) | ( ~x12 & n719 ) | ( x115 & n719 ) ;
  assign n3309 = n3308 ^ n1108 ^ n885 ;
  assign n3310 = ( n702 & n1236 ) | ( n702 & n3309 ) | ( n1236 & n3309 ) ;
  assign n3311 = ( x61 & n2857 ) | ( x61 & n2905 ) | ( n2857 & n2905 ) ;
  assign n3312 = n2774 ^ n626 ^ x57 ;
  assign n3313 = n3312 ^ n1868 ^ x221 ;
  assign n3314 = n2268 & ~n3313 ;
  assign n3315 = n2475 & n3314 ;
  assign n3316 = n1899 ^ n1399 ^ x222 ;
  assign n3321 = n2235 | n3303 ;
  assign n3322 = n3321 ^ n1603 ^ 1'b0 ;
  assign n3323 = n3322 ^ n2352 ^ n498 ;
  assign n3319 = ( ~n407 & n859 ) | ( ~n407 & n2163 ) | ( n859 & n2163 ) ;
  assign n3320 = n3319 ^ n2849 ^ n1200 ;
  assign n3324 = n3323 ^ n3320 ^ 1'b0 ;
  assign n3325 = n1034 & n3324 ;
  assign n3326 = n3325 ^ n820 ^ 1'b0 ;
  assign n3317 = n1276 | n3130 ;
  assign n3318 = ( n2143 & ~n2557 ) | ( n2143 & n3317 ) | ( ~n2557 & n3317 ) ;
  assign n3327 = n3326 ^ n3318 ^ n1188 ;
  assign n3332 = n2372 ^ n748 ^ n323 ;
  assign n3333 = ( x121 & n549 ) | ( x121 & n3332 ) | ( n549 & n3332 ) ;
  assign n3329 = n747 & n1794 ;
  assign n3330 = ~n394 & n3329 ;
  assign n3328 = n1758 ^ n789 ^ n664 ;
  assign n3331 = n3330 ^ n3328 ^ n2980 ;
  assign n3334 = n3333 ^ n3331 ^ n1726 ;
  assign n3335 = ( ~n788 & n1948 ) | ( ~n788 & n3334 ) | ( n1948 & n3334 ) ;
  assign n3336 = ( n526 & n1839 ) | ( n526 & n2989 ) | ( n1839 & n2989 ) ;
  assign n3337 = ( ~n1123 & n1156 ) | ( ~n1123 & n2084 ) | ( n1156 & n2084 ) ;
  assign n3338 = n3337 ^ n1819 ^ 1'b0 ;
  assign n3339 = ~n1816 & n2401 ;
  assign n3340 = n3339 ^ n2401 ^ 1'b0 ;
  assign n3341 = n3340 ^ n997 ^ n798 ;
  assign n3342 = n1243 ^ n986 ^ 1'b0 ;
  assign n3343 = ( n415 & n1350 ) | ( n415 & ~n3342 ) | ( n1350 & ~n3342 ) ;
  assign n3344 = n3343 ^ n2245 ^ 1'b0 ;
  assign n3345 = n1400 & ~n3344 ;
  assign n3346 = n3341 & n3345 ;
  assign n3347 = ~n3338 & n3346 ;
  assign n3348 = n1520 | n3347 ;
  assign n3349 = n3348 ^ n2832 ^ 1'b0 ;
  assign n3350 = n3144 ^ n686 ^ n465 ;
  assign n3351 = ( n670 & n1252 ) | ( n670 & ~n3350 ) | ( n1252 & ~n3350 ) ;
  assign n3352 = n3351 ^ n2993 ^ n1676 ;
  assign n3353 = ( x189 & n3228 ) | ( x189 & n3352 ) | ( n3228 & n3352 ) ;
  assign n3354 = n2326 ^ n1472 ^ 1'b0 ;
  assign n3355 = n3005 | n3354 ;
  assign n3356 = n2406 | n3355 ;
  assign n3357 = n2495 ^ n2282 ^ 1'b0 ;
  assign n3358 = x31 & n3357 ;
  assign n3359 = ( ~n1061 & n2861 ) | ( ~n1061 & n3306 ) | ( n2861 & n3306 ) ;
  assign n3364 = x97 & ~n595 ;
  assign n3365 = ~n1077 & n3364 ;
  assign n3366 = ( ~x157 & n2918 ) | ( ~x157 & n3365 ) | ( n2918 & n3365 ) ;
  assign n3361 = ( x221 & ~n458 ) | ( x221 & n691 ) | ( ~n458 & n691 ) ;
  assign n3360 = ( n508 & ~n523 ) | ( n508 & n705 ) | ( ~n523 & n705 ) ;
  assign n3362 = n3361 ^ n3360 ^ n1054 ;
  assign n3363 = n3362 ^ n1405 ^ n558 ;
  assign n3367 = n3366 ^ n3363 ^ n2461 ;
  assign n3377 = ( n993 & n1927 ) | ( n993 & n2445 ) | ( n1927 & n2445 ) ;
  assign n3368 = n869 ^ x249 ^ 1'b0 ;
  assign n3369 = n3368 ^ n794 ^ n289 ;
  assign n3370 = n903 ^ n503 ^ 1'b0 ;
  assign n3371 = ~n3369 & n3370 ;
  assign n3372 = n1570 & n3371 ;
  assign n3373 = n3372 ^ n711 ^ 1'b0 ;
  assign n3374 = ~n748 & n3373 ;
  assign n3375 = n3374 ^ x90 ^ 1'b0 ;
  assign n3376 = ~n1214 & n3375 ;
  assign n3378 = n3377 ^ n3376 ^ n438 ;
  assign n3379 = n1269 & ~n3378 ;
  assign n3380 = x154 & n1902 ;
  assign n3381 = n3380 ^ n1649 ^ 1'b0 ;
  assign n3382 = n597 & ~n1292 ;
  assign n3383 = ~n1381 & n3382 ;
  assign n3384 = n3276 & ~n3383 ;
  assign n3385 = n3384 ^ n2210 ^ 1'b0 ;
  assign n3386 = ( n3296 & ~n3381 ) | ( n3296 & n3385 ) | ( ~n3381 & n3385 ) ;
  assign n3387 = n381 & ~n2606 ;
  assign n3388 = n3387 ^ n419 ^ 1'b0 ;
  assign n3389 = x79 & ~n3388 ;
  assign n3390 = n2564 ^ n1029 ^ n535 ;
  assign n3391 = n3390 ^ n3245 ^ n1154 ;
  assign n3400 = n357 & ~n2318 ;
  assign n3401 = n3400 ^ x120 ^ 1'b0 ;
  assign n3394 = ~n1191 & n2277 ;
  assign n3395 = ~n1146 & n3394 ;
  assign n3396 = n3395 ^ n1394 ^ 1'b0 ;
  assign n3397 = ~n1870 & n3396 ;
  assign n3398 = ( x129 & n389 ) | ( x129 & n3397 ) | ( n389 & n3397 ) ;
  assign n3399 = n3398 ^ n1108 ^ n293 ;
  assign n3402 = n3401 ^ n3399 ^ n1991 ;
  assign n3403 = n2913 ^ n1546 ^ 1'b0 ;
  assign n3404 = n3402 | n3403 ;
  assign n3392 = n739 ^ n585 ^ 1'b0 ;
  assign n3393 = ~n3240 & n3392 ;
  assign n3405 = n3404 ^ n3393 ^ n3304 ;
  assign n3406 = n2519 ^ n1729 ^ n557 ;
  assign n3407 = n269 & ~n3406 ;
  assign n3413 = n793 ^ n287 ^ 1'b0 ;
  assign n3414 = ~n566 & n3413 ;
  assign n3415 = ~n794 & n3414 ;
  assign n3408 = x181 ^ x42 ^ 1'b0 ;
  assign n3409 = ~n1706 & n2504 ;
  assign n3410 = n612 & n3409 ;
  assign n3411 = n3410 ^ x208 ^ x134 ;
  assign n3412 = ( n480 & n3408 ) | ( n480 & n3411 ) | ( n3408 & n3411 ) ;
  assign n3416 = n3415 ^ n3412 ^ n639 ;
  assign n3417 = ( ~x88 & n887 ) | ( ~x88 & n1787 ) | ( n887 & n1787 ) ;
  assign n3418 = n3417 ^ n2793 ^ n1809 ;
  assign n3419 = n3418 ^ n3094 ^ 1'b0 ;
  assign n3420 = x111 & ~n3419 ;
  assign n3422 = ~x22 & n1340 ;
  assign n3421 = x223 & n420 ;
  assign n3423 = n3422 ^ n3421 ^ 1'b0 ;
  assign n3429 = n1836 & ~n2519 ;
  assign n3424 = ( n310 & ~n446 ) | ( n310 & n733 ) | ( ~n446 & n733 ) ;
  assign n3425 = ~n811 & n3424 ;
  assign n3426 = n3425 ^ n1133 ^ 1'b0 ;
  assign n3427 = ( n431 & ~n1017 ) | ( n431 & n3426 ) | ( ~n1017 & n3426 ) ;
  assign n3428 = n3427 ^ n1423 ^ n1019 ;
  assign n3430 = n3429 ^ n3428 ^ n1164 ;
  assign n3431 = n1254 | n2853 ;
  assign n3432 = ( n2257 & n2607 ) | ( n2257 & ~n3431 ) | ( n2607 & ~n3431 ) ;
  assign n3433 = n951 | n3288 ;
  assign n3434 = n3432 & ~n3433 ;
  assign n3435 = ~n311 & n3434 ;
  assign n3442 = n390 ^ x228 ^ 1'b0 ;
  assign n3443 = n1090 & n3442 ;
  assign n3444 = n3443 ^ n1269 ^ n608 ;
  assign n3436 = n1003 ^ x65 ^ 1'b0 ;
  assign n3437 = x221 & n3436 ;
  assign n3438 = n3437 ^ n1246 ^ n1224 ;
  assign n3439 = n2868 & n3438 ;
  assign n3440 = n1646 | n3439 ;
  assign n3441 = n2925 & ~n3440 ;
  assign n3445 = n3444 ^ n3441 ^ n621 ;
  assign n3446 = ( ~n1090 & n3332 ) | ( ~n1090 & n3445 ) | ( n3332 & n3445 ) ;
  assign n3447 = n2864 ^ n399 ^ n387 ;
  assign n3448 = ( n895 & ~n1573 ) | ( n895 & n1948 ) | ( ~n1573 & n1948 ) ;
  assign n3450 = n1670 ^ n1130 ^ x188 ;
  assign n3451 = n3450 ^ n1018 ^ 1'b0 ;
  assign n3452 = n677 & n3451 ;
  assign n3449 = n3115 ^ n420 ^ 1'b0 ;
  assign n3453 = n3452 ^ n3449 ^ 1'b0 ;
  assign n3454 = ( n1907 & n2230 ) | ( n1907 & n2599 ) | ( n2230 & n2599 ) ;
  assign n3455 = ( n1144 & n2214 ) | ( n1144 & n3139 ) | ( n2214 & n3139 ) ;
  assign n3456 = n3135 ^ n561 ^ 1'b0 ;
  assign n3457 = ( n1325 & ~n1813 ) | ( n1325 & n3456 ) | ( ~n1813 & n3456 ) ;
  assign n3458 = n3457 ^ n2011 ^ 1'b0 ;
  assign n3463 = n3322 ^ n1758 ^ x7 ;
  assign n3459 = n779 & ~n1948 ;
  assign n3460 = n3459 ^ n2420 ^ n449 ;
  assign n3461 = n3460 ^ n1235 ^ x16 ;
  assign n3462 = n3461 ^ n2662 ^ 1'b0 ;
  assign n3464 = n3463 ^ n3462 ^ 1'b0 ;
  assign n3465 = n2715 | n3464 ;
  assign n3466 = n1155 ^ x89 ^ 1'b0 ;
  assign n3467 = n1870 | n3466 ;
  assign n3468 = n1433 & ~n3467 ;
  assign n3469 = ( n325 & n1302 ) | ( n325 & n1905 ) | ( n1302 & n1905 ) ;
  assign n3470 = n896 & n1018 ;
  assign n3471 = n3470 ^ n2732 ^ 1'b0 ;
  assign n3472 = ( n429 & ~n846 ) | ( n429 & n1246 ) | ( ~n846 & n1246 ) ;
  assign n3473 = n3472 ^ n2457 ^ n771 ;
  assign n3474 = n1926 ^ n994 ^ x237 ;
  assign n3475 = n2360 & n3474 ;
  assign n3476 = ~n1672 & n3475 ;
  assign n3477 = n2408 | n2893 ;
  assign n3478 = n3476 & ~n3477 ;
  assign n3479 = ( n449 & ~n1024 ) | ( n449 & n2961 ) | ( ~n1024 & n2961 ) ;
  assign n3480 = ~n1822 & n3155 ;
  assign n3481 = n987 & n3480 ;
  assign n3482 = n1503 & ~n3481 ;
  assign n3483 = n825 & ~n3482 ;
  assign n3484 = ( x233 & n1292 ) | ( x233 & ~n2051 ) | ( n1292 & ~n2051 ) ;
  assign n3485 = n3484 ^ n1363 ^ n1162 ;
  assign n3486 = ( x3 & n1446 ) | ( x3 & n2754 ) | ( n1446 & n2754 ) ;
  assign n3487 = n3486 ^ n1116 ^ n1037 ;
  assign n3488 = ( ~n2059 & n3485 ) | ( ~n2059 & n3487 ) | ( n3485 & n3487 ) ;
  assign n3491 = ~n291 & n1252 ;
  assign n3492 = n894 & n3491 ;
  assign n3489 = ( n414 & ~n899 ) | ( n414 & n2382 ) | ( ~n899 & n2382 ) ;
  assign n3490 = n3489 ^ n1616 ^ x14 ;
  assign n3493 = n3492 ^ n3490 ^ x53 ;
  assign n3494 = n3493 ^ n868 ^ n725 ;
  assign n3495 = ( n568 & n1982 ) | ( n568 & n3494 ) | ( n1982 & n3494 ) ;
  assign n3497 = n1172 ^ n801 ^ n524 ;
  assign n3498 = ( n2209 & ~n3296 ) | ( n2209 & n3497 ) | ( ~n3296 & n3497 ) ;
  assign n3499 = n3498 ^ x135 ^ 1'b0 ;
  assign n3500 = ~n2667 & n3499 ;
  assign n3501 = n3500 ^ n3337 ^ x177 ;
  assign n3496 = ( n640 & ~n1884 ) | ( n640 & n2877 ) | ( ~n1884 & n2877 ) ;
  assign n3502 = n3501 ^ n3496 ^ n1408 ;
  assign n3503 = n515 | n3502 ;
  assign n3504 = n3495 & ~n3503 ;
  assign n3508 = n924 | n1211 ;
  assign n3509 = n3508 ^ n1631 ^ n594 ;
  assign n3505 = n2239 ^ n1754 ^ n1677 ;
  assign n3506 = n3493 ^ n2635 ^ n1264 ;
  assign n3507 = ( n2128 & n3505 ) | ( n2128 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3510 = n3509 ^ n3507 ^ 1'b0 ;
  assign n3511 = ( n3488 & ~n3504 ) | ( n3488 & n3510 ) | ( ~n3504 & n3510 ) ;
  assign n3512 = ( ~n1672 & n2086 ) | ( ~n1672 & n2785 ) | ( n2086 & n2785 ) ;
  assign n3515 = ( n873 & n1146 ) | ( n873 & n2166 ) | ( n1146 & n2166 ) ;
  assign n3513 = ~n379 & n470 ;
  assign n3514 = n2183 & n3513 ;
  assign n3516 = n3515 ^ n3514 ^ n1144 ;
  assign n3517 = n2141 & ~n3516 ;
  assign n3518 = ( ~n574 & n1251 ) | ( ~n574 & n3517 ) | ( n1251 & n3517 ) ;
  assign n3519 = ( n289 & ~n401 ) | ( n289 & n3266 ) | ( ~n401 & n3266 ) ;
  assign n3520 = ( ~x141 & n1535 ) | ( ~x141 & n3164 ) | ( n1535 & n3164 ) ;
  assign n3521 = n3520 ^ n2410 ^ 1'b0 ;
  assign n3522 = n3519 & n3521 ;
  assign n3524 = n1306 ^ n1007 ^ n664 ;
  assign n3523 = n1561 ^ n1444 ^ n313 ;
  assign n3525 = n3524 ^ n3523 ^ x21 ;
  assign n3526 = n1728 ^ n1596 ^ 1'b0 ;
  assign n3527 = ~n304 & n795 ;
  assign n3528 = n3527 ^ n2527 ^ 1'b0 ;
  assign n3529 = ( ~n683 & n3526 ) | ( ~n683 & n3528 ) | ( n3526 & n3528 ) ;
  assign n3530 = n3529 ^ n1304 ^ 1'b0 ;
  assign n3531 = n1142 & n1573 ;
  assign n3532 = n3531 ^ n3022 ^ 1'b0 ;
  assign n3533 = ~n3290 & n3532 ;
  assign n3534 = n3530 & n3533 ;
  assign n3535 = ( x7 & ~n3525 ) | ( x7 & n3534 ) | ( ~n3525 & n3534 ) ;
  assign n3536 = n3402 ^ n2373 ^ n1295 ;
  assign n3537 = ( ~x16 & n3053 ) | ( ~x16 & n3536 ) | ( n3053 & n3536 ) ;
  assign n3538 = n2992 ^ n2027 ^ n1154 ;
  assign n3539 = n3538 ^ n3326 ^ n1315 ;
  assign n3540 = n2182 | n3539 ;
  assign n3541 = n3160 ^ n924 ^ n301 ;
  assign n3542 = ( ~n1488 & n2392 ) | ( ~n1488 & n3541 ) | ( n2392 & n3541 ) ;
  assign n3543 = n3542 ^ n2840 ^ 1'b0 ;
  assign n3544 = n291 | n3543 ;
  assign n3545 = n3544 ^ n1728 ^ 1'b0 ;
  assign n3548 = n382 ^ n302 ^ n288 ;
  assign n3549 = n3548 ^ n1011 ^ n461 ;
  assign n3550 = n3549 ^ x107 ^ x24 ;
  assign n3546 = ( x58 & n274 ) | ( x58 & ~n3365 ) | ( n274 & ~n3365 ) ;
  assign n3547 = n3546 ^ n2456 ^ n1440 ;
  assign n3551 = n3550 ^ n3547 ^ n608 ;
  assign n3552 = n1697 ^ n1378 ^ 1'b0 ;
  assign n3553 = x153 & ~n3552 ;
  assign n3563 = n799 | n2076 ;
  assign n3564 = n2606 & ~n3563 ;
  assign n3560 = n466 & ~n575 ;
  assign n3561 = n3560 ^ n1369 ^ 1'b0 ;
  assign n3559 = ~n579 & n1028 ;
  assign n3562 = n3561 ^ n3559 ^ 1'b0 ;
  assign n3565 = n3564 ^ n3562 ^ 1'b0 ;
  assign n3566 = n1930 & n3565 ;
  assign n3567 = n1747 & n3566 ;
  assign n3554 = n1755 ^ x213 ^ 1'b0 ;
  assign n3555 = ( ~n589 & n1788 ) | ( ~n589 & n3554 ) | ( n1788 & n3554 ) ;
  assign n3556 = n3555 ^ n2116 ^ n293 ;
  assign n3557 = ( n1529 & n1803 ) | ( n1529 & n3556 ) | ( n1803 & n3556 ) ;
  assign n3558 = x48 & ~n3557 ;
  assign n3568 = n3567 ^ n3558 ^ 1'b0 ;
  assign n3569 = n3271 ^ n2746 ^ n578 ;
  assign n3570 = ~n2755 & n3569 ;
  assign n3571 = n3500 & n3570 ;
  assign n3572 = n3571 ^ n1853 ^ n1207 ;
  assign n3573 = n3572 ^ n1828 ^ 1'b0 ;
  assign n3574 = n3568 & ~n3573 ;
  assign n3577 = ( x243 & n2084 ) | ( x243 & ~n3191 ) | ( n2084 & ~n3191 ) ;
  assign n3575 = n966 | n1729 ;
  assign n3576 = ~n452 & n3575 ;
  assign n3578 = n3577 ^ n3576 ^ 1'b0 ;
  assign n3579 = n1756 ^ n1111 ^ x59 ;
  assign n3580 = ~n460 & n3579 ;
  assign n3581 = ( n387 & n2521 ) | ( n387 & n3580 ) | ( n2521 & n3580 ) ;
  assign n3585 = ( n325 & n490 ) | ( n325 & ~n2050 ) | ( n490 & ~n2050 ) ;
  assign n3586 = n2360 & ~n3585 ;
  assign n3587 = n3586 ^ n1877 ^ 1'b0 ;
  assign n3582 = ~n1467 & n1883 ;
  assign n3583 = n3582 ^ n1799 ^ 1'b0 ;
  assign n3584 = n3450 & ~n3583 ;
  assign n3588 = n3587 ^ n3584 ^ n3185 ;
  assign n3589 = n3024 ^ n2342 ^ n348 ;
  assign n3591 = ( n511 & n857 ) | ( n511 & n3163 ) | ( n857 & n3163 ) ;
  assign n3590 = n969 & n2230 ;
  assign n3592 = n3591 ^ n3590 ^ 1'b0 ;
  assign n3593 = ( n829 & n3589 ) | ( n829 & n3592 ) | ( n3589 & n3592 ) ;
  assign n3594 = ( n2152 & ~n2629 ) | ( n2152 & n3584 ) | ( ~n2629 & n3584 ) ;
  assign n3595 = n2710 ^ n1516 ^ n633 ;
  assign n3596 = n3369 ^ n606 ^ x193 ;
  assign n3597 = n3596 ^ n3474 ^ 1'b0 ;
  assign n3598 = ( ~n1242 & n1855 ) | ( ~n1242 & n2920 ) | ( n1855 & n2920 ) ;
  assign n3599 = n1959 ^ n1850 ^ n1186 ;
  assign n3600 = ( n1200 & ~n3598 ) | ( n1200 & n3599 ) | ( ~n3598 & n3599 ) ;
  assign n3601 = ( n967 & ~n2346 ) | ( n967 & n3600 ) | ( ~n2346 & n3600 ) ;
  assign n3602 = n3601 ^ x42 ^ 1'b0 ;
  assign n3603 = ~n3597 & n3602 ;
  assign n3604 = n3228 ^ n379 ^ 1'b0 ;
  assign n3605 = ~n809 & n3604 ;
  assign n3606 = n3605 ^ n431 ^ 1'b0 ;
  assign n3607 = n3606 ^ x207 ^ 1'b0 ;
  assign n3608 = ( n361 & n1763 ) | ( n361 & ~n2643 ) | ( n1763 & ~n2643 ) ;
  assign n3609 = ( ~n1046 & n2750 ) | ( ~n1046 & n3608 ) | ( n2750 & n3608 ) ;
  assign n3610 = ~n1896 & n2277 ;
  assign n3611 = n1293 & n3610 ;
  assign n3612 = n3210 ^ n1293 ^ n461 ;
  assign n3613 = n3612 ^ n2777 ^ n1433 ;
  assign n3614 = ( n300 & n808 ) | ( n300 & ~n2240 ) | ( n808 & ~n2240 ) ;
  assign n3615 = ~n708 & n3614 ;
  assign n3616 = n1875 ^ n944 ^ n382 ;
  assign n3617 = n3616 ^ n2606 ^ 1'b0 ;
  assign n3618 = n1207 ^ n849 ^ 1'b0 ;
  assign n3619 = n563 & ~n3618 ;
  assign n3620 = n3619 ^ n499 ^ n275 ;
  assign n3621 = ( ~n1645 & n3617 ) | ( ~n1645 & n3620 ) | ( n3617 & n3620 ) ;
  assign n3622 = n3621 ^ n1971 ^ n540 ;
  assign n3623 = n3298 ^ n3111 ^ n1724 ;
  assign n3624 = ( ~n538 & n784 ) | ( ~n538 & n2412 ) | ( n784 & n2412 ) ;
  assign n3625 = n1392 & n3624 ;
  assign n3626 = n3625 ^ n375 ^ 1'b0 ;
  assign n3627 = n3626 ^ n2031 ^ 1'b0 ;
  assign n3628 = ~n1762 & n3627 ;
  assign n3629 = n3628 ^ n2715 ^ 1'b0 ;
  assign n3630 = ( n1929 & n3623 ) | ( n1929 & ~n3629 ) | ( n3623 & ~n3629 ) ;
  assign n3631 = ( n351 & n777 ) | ( n351 & ~n3266 ) | ( n777 & ~n3266 ) ;
  assign n3632 = n3631 ^ n903 ^ n858 ;
  assign n3638 = n332 & ~n538 ;
  assign n3639 = ( n815 & n1122 ) | ( n815 & ~n3638 ) | ( n1122 & ~n3638 ) ;
  assign n3640 = n3639 ^ n1294 ^ 1'b0 ;
  assign n3641 = x104 & n3640 ;
  assign n3633 = n3244 ^ n1212 ^ x4 ;
  assign n3634 = n890 ^ n555 ^ 1'b0 ;
  assign n3635 = n974 & n3634 ;
  assign n3636 = ( n2083 & ~n2694 ) | ( n2083 & n3635 ) | ( ~n2694 & n3635 ) ;
  assign n3637 = n3633 & ~n3636 ;
  assign n3642 = n3641 ^ n3637 ^ 1'b0 ;
  assign n3643 = n3642 ^ n2451 ^ n1408 ;
  assign n3644 = n3484 ^ x175 ^ 1'b0 ;
  assign n3645 = ( x106 & n1280 ) | ( x106 & n3644 ) | ( n1280 & n3644 ) ;
  assign n3646 = ~n2070 & n3645 ;
  assign n3647 = n2256 ^ n1638 ^ n1064 ;
  assign n3648 = ~n3272 & n3647 ;
  assign n3651 = n1295 & n1673 ;
  assign n3652 = n3303 ^ n2372 ^ 1'b0 ;
  assign n3653 = ~n3651 & n3652 ;
  assign n3649 = ( n2380 & n2490 ) | ( n2380 & ~n3269 ) | ( n2490 & ~n3269 ) ;
  assign n3650 = n348 & ~n3649 ;
  assign n3654 = n3653 ^ n3650 ^ 1'b0 ;
  assign n3655 = n2512 ^ n1291 ^ 1'b0 ;
  assign n3656 = n3654 | n3655 ;
  assign n3657 = n3432 ^ n2283 ^ n372 ;
  assign n3658 = ( n1181 & n2863 ) | ( n1181 & n3657 ) | ( n2863 & n3657 ) ;
  assign n3673 = n1172 & ~n1827 ;
  assign n3666 = n2715 ^ n1943 ^ 1'b0 ;
  assign n3667 = n1759 & ~n3666 ;
  assign n3668 = n3247 ^ n476 ^ 1'b0 ;
  assign n3669 = ( n1164 & n2816 ) | ( n1164 & ~n3668 ) | ( n2816 & ~n3668 ) ;
  assign n3670 = n3399 ^ n2376 ^ n1219 ;
  assign n3671 = ( n3667 & ~n3669 ) | ( n3667 & n3670 ) | ( ~n3669 & n3670 ) ;
  assign n3659 = ( x45 & ~n283 ) | ( x45 & n313 ) | ( ~n283 & n313 ) ;
  assign n3660 = n1189 & n3659 ;
  assign n3661 = ~x130 & n3660 ;
  assign n3662 = n1629 ^ x130 ^ 1'b0 ;
  assign n3663 = n1308 & n3662 ;
  assign n3664 = n3663 ^ n3644 ^ n2277 ;
  assign n3665 = n3661 | n3664 ;
  assign n3672 = n3671 ^ n3665 ^ 1'b0 ;
  assign n3674 = n3673 ^ n3672 ^ n3614 ;
  assign n3675 = n3674 ^ n507 ^ x78 ;
  assign n3676 = ( ~n313 & n505 ) | ( ~n313 & n1141 ) | ( n505 & n1141 ) ;
  assign n3677 = n3676 ^ n3365 ^ n2641 ;
  assign n3678 = ( ~n1676 & n1702 ) | ( ~n1676 & n2041 ) | ( n1702 & n2041 ) ;
  assign n3679 = ( ~n2272 & n3677 ) | ( ~n2272 & n3678 ) | ( n3677 & n3678 ) ;
  assign n3687 = n2259 ^ n688 ^ 1'b0 ;
  assign n3688 = n573 | n3687 ;
  assign n3689 = x219 | n3688 ;
  assign n3680 = ~n325 & n1928 ;
  assign n3681 = ( x62 & n433 ) | ( x62 & ~n3680 ) | ( n433 & ~n3680 ) ;
  assign n3682 = ( n270 & ~n1431 ) | ( n270 & n1454 ) | ( ~n1431 & n1454 ) ;
  assign n3683 = n275 & ~n1331 ;
  assign n3684 = ~n3682 & n3683 ;
  assign n3685 = n3684 ^ n2235 ^ n467 ;
  assign n3686 = ( x158 & ~n3681 ) | ( x158 & n3685 ) | ( ~n3681 & n3685 ) ;
  assign n3690 = n3689 ^ n3686 ^ n1880 ;
  assign n3691 = n3333 ^ n1748 ^ n1714 ;
  assign n3693 = n398 ^ x218 ^ x112 ;
  assign n3692 = x197 & ~n2064 ;
  assign n3694 = n3693 ^ n3692 ^ 1'b0 ;
  assign n3695 = ( n801 & ~n1813 ) | ( n801 & n2473 ) | ( ~n1813 & n2473 ) ;
  assign n3696 = ( ~n1029 & n3694 ) | ( ~n1029 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3697 = n2336 ^ x178 ^ 1'b0 ;
  assign n3698 = n1232 & ~n3697 ;
  assign n3699 = ~n3696 & n3698 ;
  assign n3700 = ( n2929 & ~n3691 ) | ( n2929 & n3699 ) | ( ~n3691 & n3699 ) ;
  assign n3701 = ( n1392 & n1451 ) | ( n1392 & ~n2317 ) | ( n1451 & ~n2317 ) ;
  assign n3702 = n3701 ^ n1958 ^ 1'b0 ;
  assign n3703 = ~n1424 & n3702 ;
  assign n3704 = ( n1269 & ~n2313 ) | ( n1269 & n3703 ) | ( ~n2313 & n3703 ) ;
  assign n3705 = n3704 ^ n2468 ^ 1'b0 ;
  assign n3706 = n3700 | n3705 ;
  assign n3707 = n3115 ^ n2029 ^ 1'b0 ;
  assign n3708 = ( n2088 & ~n2468 ) | ( n2088 & n3538 ) | ( ~n2468 & n3538 ) ;
  assign n3710 = n585 ^ n280 ^ x87 ;
  assign n3709 = n293 | n1916 ;
  assign n3711 = n3710 ^ n3709 ^ 1'b0 ;
  assign n3712 = x220 & ~n1513 ;
  assign n3713 = ~n1737 & n3712 ;
  assign n3714 = n2629 ^ x212 ^ 1'b0 ;
  assign n3715 = n650 & n3714 ;
  assign n3716 = ( n2556 & n2787 ) | ( n2556 & n3715 ) | ( n2787 & n3715 ) ;
  assign n3717 = ( ~n2755 & n3713 ) | ( ~n2755 & n3716 ) | ( n3713 & n3716 ) ;
  assign n3718 = n2106 | n2824 ;
  assign n3719 = x249 | n3718 ;
  assign n3720 = n3719 ^ n2784 ^ 1'b0 ;
  assign n3721 = n1208 ^ n1164 ^ 1'b0 ;
  assign n3730 = n3663 ^ n2638 ^ n1503 ;
  assign n3727 = n872 ^ n273 ^ 1'b0 ;
  assign n3722 = ( n269 & ~n537 ) | ( n269 & n649 ) | ( ~n537 & n649 ) ;
  assign n3723 = n3722 ^ n1762 ^ n1256 ;
  assign n3724 = n2313 ^ n1952 ^ n1186 ;
  assign n3725 = ( n2050 & n3723 ) | ( n2050 & n3724 ) | ( n3723 & n3724 ) ;
  assign n3726 = ( n1676 & ~n1773 ) | ( n1676 & n3725 ) | ( ~n1773 & n3725 ) ;
  assign n3728 = n3727 ^ n3726 ^ n352 ;
  assign n3729 = n3728 ^ x94 ^ 1'b0 ;
  assign n3731 = n3730 ^ n3729 ^ n786 ;
  assign n3732 = n3548 ^ n720 ^ x33 ;
  assign n3733 = n3732 ^ n3691 ^ 1'b0 ;
  assign n3734 = ( n2275 & n3731 ) | ( n2275 & n3733 ) | ( n3731 & n3733 ) ;
  assign n3735 = n2992 ^ n1740 ^ 1'b0 ;
  assign n3736 = n2101 ^ n1088 ^ x85 ;
  assign n3737 = n3736 ^ n2948 ^ n1645 ;
  assign n3738 = ( n1737 & n2479 ) | ( n1737 & n3737 ) | ( n2479 & n3737 ) ;
  assign n3739 = n1218 ^ n522 ^ n450 ;
  assign n3740 = n3739 ^ n1455 ^ 1'b0 ;
  assign n3741 = n3086 ^ n2763 ^ 1'b0 ;
  assign n3742 = n3157 ^ n969 ^ 1'b0 ;
  assign n3743 = ( n1167 & n1431 ) | ( n1167 & n2953 ) | ( n1431 & n2953 ) ;
  assign n3744 = ( n944 & n1925 ) | ( n944 & ~n3715 ) | ( n1925 & ~n3715 ) ;
  assign n3745 = ( n336 & n3743 ) | ( n336 & ~n3744 ) | ( n3743 & ~n3744 ) ;
  assign n3746 = n963 | n3502 ;
  assign n3749 = n263 & n1317 ;
  assign n3747 = ( ~n642 & n1332 ) | ( ~n642 & n3417 ) | ( n1332 & n3417 ) ;
  assign n3748 = ( n1716 & ~n2366 ) | ( n1716 & n3747 ) | ( ~n2366 & n3747 ) ;
  assign n3750 = n3749 ^ n3748 ^ n1974 ;
  assign n3751 = n1587 | n1868 ;
  assign n3752 = n906 ^ n364 ^ n293 ;
  assign n3753 = n2810 ^ n1495 ^ n579 ;
  assign n3754 = n2189 ^ x40 ^ 1'b0 ;
  assign n3755 = n2559 ^ n2026 ^ 1'b0 ;
  assign n3756 = ~n3754 & n3755 ;
  assign n3757 = ( n1136 & ~n3753 ) | ( n1136 & n3756 ) | ( ~n3753 & n3756 ) ;
  assign n3758 = ( n999 & n3752 ) | ( n999 & n3757 ) | ( n3752 & n3757 ) ;
  assign n3759 = n2084 ^ x249 ^ x113 ;
  assign n3760 = n2319 & ~n3759 ;
  assign n3761 = n3760 ^ n3267 ^ 1'b0 ;
  assign n3762 = ~n3758 & n3761 ;
  assign n3763 = n3762 ^ n3612 ^ 1'b0 ;
  assign n3764 = n3710 ^ n2882 ^ x211 ;
  assign n3767 = n2139 ^ n1983 ^ n1292 ;
  assign n3766 = x252 & n1090 ;
  assign n3765 = ~n869 & n1294 ;
  assign n3768 = n3767 ^ n3766 ^ n3765 ;
  assign n3769 = n3377 ^ n1421 ^ n766 ;
  assign n3770 = ~n1287 & n3561 ;
  assign n3771 = ( n2091 & ~n3769 ) | ( n2091 & n3770 ) | ( ~n3769 & n3770 ) ;
  assign n3772 = n1200 ^ x90 ^ 1'b0 ;
  assign n3773 = ( n711 & ~n3726 ) | ( n711 & n3772 ) | ( ~n3726 & n3772 ) ;
  assign n3774 = ( x248 & n3771 ) | ( x248 & ~n3773 ) | ( n3771 & ~n3773 ) ;
  assign n3775 = n2880 ^ n2110 ^ 1'b0 ;
  assign n3776 = ( ~n312 & n3736 ) | ( ~n312 & n3775 ) | ( n3736 & n3775 ) ;
  assign n3777 = n3776 ^ n2912 ^ n1561 ;
  assign n3778 = n1067 & ~n2129 ;
  assign n3779 = n3777 & n3778 ;
  assign n3780 = x230 & ~n3703 ;
  assign n3781 = n2187 ^ n1718 ^ n560 ;
  assign n3782 = ( x176 & ~n3780 ) | ( x176 & n3781 ) | ( ~n3780 & n3781 ) ;
  assign n3783 = n1579 & n2197 ;
  assign n3784 = n1273 & n3783 ;
  assign n3785 = ( ~n1440 & n1758 ) | ( ~n1440 & n3784 ) | ( n1758 & n3784 ) ;
  assign n3786 = n327 & n3548 ;
  assign n3788 = n1042 | n3203 ;
  assign n3789 = n3788 ^ x173 ^ 1'b0 ;
  assign n3787 = n3686 ^ n2928 ^ 1'b0 ;
  assign n3790 = n3789 ^ n3787 ^ 1'b0 ;
  assign n3791 = ~n1106 & n3790 ;
  assign n3792 = ( x26 & n2515 ) | ( x26 & ~n2858 ) | ( n2515 & ~n2858 ) ;
  assign n3793 = n1440 | n2160 ;
  assign n3794 = n603 | n817 ;
  assign n3795 = n736 | n1761 ;
  assign n3796 = n3795 ^ n2706 ^ 1'b0 ;
  assign n3797 = n3794 & ~n3796 ;
  assign n3798 = n3797 ^ n2383 ^ n1392 ;
  assign n3807 = n1027 | n1469 ;
  assign n3808 = n324 | n3807 ;
  assign n3803 = ( n513 & n2133 ) | ( n513 & n2654 ) | ( n2133 & n2654 ) ;
  assign n3802 = n834 ^ x151 ^ 1'b0 ;
  assign n3804 = n3803 ^ n3802 ^ n3160 ;
  assign n3805 = ~n1712 & n3689 ;
  assign n3806 = n3804 & n3805 ;
  assign n3809 = n3808 ^ n3806 ^ 1'b0 ;
  assign n3799 = n2754 ^ n993 ^ x194 ;
  assign n3800 = n3799 ^ n3497 ^ x173 ;
  assign n3801 = ( ~n2592 & n3447 ) | ( ~n2592 & n3800 ) | ( n3447 & n3800 ) ;
  assign n3810 = n3809 ^ n3801 ^ n1632 ;
  assign n3811 = ( n1327 & ~n1677 ) | ( n1327 & n3021 ) | ( ~n1677 & n3021 ) ;
  assign n3812 = n2012 ^ n1307 ^ n688 ;
  assign n3813 = ( n536 & n3811 ) | ( n536 & n3812 ) | ( n3811 & n3812 ) ;
  assign n3814 = ( x123 & n3730 ) | ( x123 & n3813 ) | ( n3730 & n3813 ) ;
  assign n3815 = n2453 ^ n925 ^ 1'b0 ;
  assign n3816 = n2323 & ~n3815 ;
  assign n3817 = n721 & ~n1085 ;
  assign n3818 = n3817 ^ n781 ^ 1'b0 ;
  assign n3819 = n2853 & n3818 ;
  assign n3820 = n2217 ^ n1943 ^ 1'b0 ;
  assign n3821 = n2777 | n3820 ;
  assign n3822 = n1375 & ~n3821 ;
  assign n3823 = n907 ^ n857 ^ 1'b0 ;
  assign n3824 = ~n1832 & n3823 ;
  assign n3825 = ~n1180 & n3824 ;
  assign n3826 = ~n1208 & n3825 ;
  assign n3827 = n971 & ~n1747 ;
  assign n3828 = ~x246 & n3827 ;
  assign n3829 = ( n875 & n3826 ) | ( n875 & ~n3828 ) | ( n3826 & ~n3828 ) ;
  assign n3830 = n876 | n3829 ;
  assign n3831 = n2152 ^ n649 ^ 1'b0 ;
  assign n3832 = x149 & ~n3831 ;
  assign n3833 = n3832 ^ n2319 ^ n1559 ;
  assign n3834 = n264 & n3833 ;
  assign n3835 = n291 & n3834 ;
  assign n3836 = n1185 & ~n3835 ;
  assign n3837 = n861 & ~n1823 ;
  assign n3838 = n468 & ~n2521 ;
  assign n3840 = n2243 ^ x136 ^ 1'b0 ;
  assign n3839 = ~n1439 & n2659 ;
  assign n3841 = n3840 ^ n3839 ^ n873 ;
  assign n3842 = n3841 ^ n1580 ^ n890 ;
  assign n3843 = ~n2506 & n3842 ;
  assign n3844 = ~n1530 & n3843 ;
  assign n3845 = ( ~n866 & n3838 ) | ( ~n866 & n3844 ) | ( n3838 & n3844 ) ;
  assign n3846 = n984 & n2890 ;
  assign n3847 = n3846 ^ n326 ^ 1'b0 ;
  assign n3848 = n2029 ^ n1898 ^ 1'b0 ;
  assign n3849 = n771 ^ n390 ^ x167 ;
  assign n3850 = n1523 | n3849 ;
  assign n3851 = n2780 & ~n3850 ;
  assign n3852 = ( n756 & n2385 ) | ( n756 & n3644 ) | ( n2385 & n3644 ) ;
  assign n3853 = ~n2555 & n3852 ;
  assign n3861 = n1011 & n1139 ;
  assign n3862 = n3861 ^ n1839 ^ 1'b0 ;
  assign n3854 = n2339 ^ n1413 ^ n536 ;
  assign n3855 = n2012 ^ n1175 ^ x13 ;
  assign n3856 = ( n1167 & n3854 ) | ( n1167 & ~n3855 ) | ( n3854 & ~n3855 ) ;
  assign n3857 = n3856 ^ n2221 ^ n787 ;
  assign n3858 = x221 & n2606 ;
  assign n3859 = x143 | n3858 ;
  assign n3860 = n3857 & n3859 ;
  assign n3863 = n3862 ^ n3860 ^ 1'b0 ;
  assign n3864 = n3853 & ~n3863 ;
  assign n3865 = ( n2813 & n3851 ) | ( n2813 & ~n3864 ) | ( n3851 & ~n3864 ) ;
  assign n3877 = n3319 ^ n1722 ^ n1428 ;
  assign n3866 = n2169 ^ n732 ^ n501 ;
  assign n3867 = n3866 ^ n2173 ^ x144 ;
  assign n3868 = ( n491 & n3342 ) | ( n491 & n3867 ) | ( n3342 & n3867 ) ;
  assign n3872 = n2494 ^ n1401 ^ x97 ;
  assign n3873 = ( ~n365 & n3228 ) | ( ~n365 & n3872 ) | ( n3228 & n3872 ) ;
  assign n3869 = ( ~n524 & n1417 ) | ( ~n524 & n1853 ) | ( n1417 & n1853 ) ;
  assign n3870 = ( n619 & n1944 ) | ( n619 & n2559 ) | ( n1944 & n2559 ) ;
  assign n3871 = ( ~n2090 & n3869 ) | ( ~n2090 & n3870 ) | ( n3869 & n3870 ) ;
  assign n3874 = n3873 ^ n3871 ^ n3401 ;
  assign n3875 = ~n1656 & n3874 ;
  assign n3876 = ~n3868 & n3875 ;
  assign n3878 = n3877 ^ n3876 ^ n2643 ;
  assign n3879 = ( n284 & ~n866 ) | ( n284 & n3266 ) | ( ~n866 & n3266 ) ;
  assign n3880 = n1042 ^ n499 ^ 1'b0 ;
  assign n3881 = n2575 & ~n3880 ;
  assign n3882 = n2501 & n3881 ;
  assign n3883 = n3882 ^ n299 ^ 1'b0 ;
  assign n3884 = n3883 ^ n3134 ^ n664 ;
  assign n3885 = ( ~n2588 & n3879 ) | ( ~n2588 & n3884 ) | ( n3879 & n3884 ) ;
  assign n3886 = ~n2496 & n3253 ;
  assign n3887 = n3886 ^ n3067 ^ 1'b0 ;
  assign n3888 = n1925 ^ x153 ^ 1'b0 ;
  assign n3889 = n3888 ^ n2492 ^ n501 ;
  assign n3890 = n3889 ^ n574 ^ 1'b0 ;
  assign n3891 = ~n789 & n3890 ;
  assign n3892 = ~n3887 & n3891 ;
  assign n3893 = n1129 & ~n1718 ;
  assign n3894 = n2894 & n3893 ;
  assign n3895 = n3894 ^ n1451 ^ n1297 ;
  assign n3896 = n3895 ^ n1528 ^ n574 ;
  assign n3897 = n3896 ^ n1683 ^ 1'b0 ;
  assign n3898 = x196 & n809 ;
  assign n3899 = n3898 ^ n1473 ^ 1'b0 ;
  assign n3900 = n3899 ^ n1980 ^ n291 ;
  assign n3901 = n3900 ^ n1894 ^ n1695 ;
  assign n3905 = n329 | n3688 ;
  assign n3906 = ( x17 & n3846 ) | ( x17 & n3905 ) | ( n3846 & n3905 ) ;
  assign n3902 = n3260 ^ n2331 ^ n2223 ;
  assign n3903 = n1590 | n3902 ;
  assign n3904 = n1835 | n3903 ;
  assign n3907 = n3906 ^ n3904 ^ 1'b0 ;
  assign n3908 = n3907 ^ n2183 ^ 1'b0 ;
  assign n3909 = n1032 ^ n329 ^ 1'b0 ;
  assign n3910 = ( n1689 & n3225 ) | ( n1689 & n3909 ) | ( n3225 & n3909 ) ;
  assign n3911 = n3317 ^ n1616 ^ n587 ;
  assign n3912 = ( ~n3135 & n3910 ) | ( ~n3135 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3913 = ~n505 & n694 ;
  assign n3914 = ~n1237 & n3913 ;
  assign n3915 = ( ~n1114 & n2281 ) | ( ~n1114 & n3914 ) | ( n2281 & n3914 ) ;
  assign n3916 = n738 & ~n3915 ;
  assign n3917 = n3497 ^ n1591 ^ n1556 ;
  assign n3918 = ( ~n666 & n1108 ) | ( ~n666 & n3308 ) | ( n1108 & n3308 ) ;
  assign n3919 = n3869 & ~n3918 ;
  assign n3920 = n3919 ^ n3841 ^ n3427 ;
  assign n3921 = n3917 & ~n3920 ;
  assign n3922 = ( n1200 & n1226 ) | ( n1200 & ~n2402 ) | ( n1226 & ~n2402 ) ;
  assign n3923 = n3922 ^ n2134 ^ n1285 ;
  assign n3926 = n589 ^ x156 ^ x89 ;
  assign n3927 = ~n3067 & n3926 ;
  assign n3924 = n702 & ~n2245 ;
  assign n3925 = n3924 ^ x210 ^ 1'b0 ;
  assign n3928 = n3927 ^ n3925 ^ 1'b0 ;
  assign n3929 = n1843 & ~n3928 ;
  assign n3933 = n2133 ^ n1334 ^ n835 ;
  assign n3934 = ( n1317 & ~n3260 ) | ( n1317 & n3933 ) | ( ~n3260 & n3933 ) ;
  assign n3935 = n3934 ^ n1088 ^ 1'b0 ;
  assign n3936 = ~n455 & n3935 ;
  assign n3937 = n545 ^ n486 ^ x215 ;
  assign n3938 = ( n1593 & ~n3936 ) | ( n1593 & n3937 ) | ( ~n3936 & n3937 ) ;
  assign n3930 = n1345 ^ n1106 ^ 1'b0 ;
  assign n3931 = ~n932 & n3930 ;
  assign n3932 = ( n2865 & ~n3073 ) | ( n2865 & n3931 ) | ( ~n3073 & n3931 ) ;
  assign n3939 = n3938 ^ n3932 ^ 1'b0 ;
  assign n3940 = n3939 ^ n3522 ^ n2606 ;
  assign n3941 = n2388 ^ x144 ^ 1'b0 ;
  assign n3942 = n1167 & ~n3941 ;
  assign n3943 = n3942 ^ n556 ^ n399 ;
  assign n3944 = ( n463 & n877 ) | ( n463 & ~n3181 ) | ( n877 & ~n3181 ) ;
  assign n3952 = n3873 ^ n801 ^ n498 ;
  assign n3947 = n1403 ^ n1384 ^ n649 ;
  assign n3945 = n1795 ^ n1107 ^ n774 ;
  assign n3946 = ~n1853 & n3945 ;
  assign n3948 = n3947 ^ n3946 ^ 1'b0 ;
  assign n3949 = ( ~n331 & n1623 ) | ( ~n331 & n3828 ) | ( n1623 & n3828 ) ;
  assign n3950 = n3949 ^ n1759 ^ x119 ;
  assign n3951 = ( n606 & n3948 ) | ( n606 & ~n3950 ) | ( n3948 & ~n3950 ) ;
  assign n3953 = n3952 ^ n3951 ^ 1'b0 ;
  assign n3954 = ( n942 & n2766 ) | ( n942 & ~n3953 ) | ( n2766 & ~n3953 ) ;
  assign n3958 = ( ~n329 & n766 ) | ( ~n329 & n2544 ) | ( n766 & n2544 ) ;
  assign n3959 = n3958 ^ n3235 ^ n1085 ;
  assign n3960 = n3959 ^ n786 ^ x108 ;
  assign n3955 = ( x68 & n1469 ) | ( x68 & n2994 ) | ( n1469 & n2994 ) ;
  assign n3956 = n2872 | n3955 ;
  assign n3957 = n1523 | n3956 ;
  assign n3961 = n3960 ^ n3957 ^ 1'b0 ;
  assign n3962 = n3211 ^ n3154 ^ 1'b0 ;
  assign n3963 = n3753 ^ n1726 ^ n819 ;
  assign n3964 = ( n414 & n3962 ) | ( n414 & n3963 ) | ( n3962 & n3963 ) ;
  assign n3971 = x198 & n1181 ;
  assign n3972 = n592 & n3971 ;
  assign n3973 = ~x136 & n3972 ;
  assign n3974 = ( x37 & ~x230 ) | ( x37 & n3973 ) | ( ~x230 & n3973 ) ;
  assign n3965 = n2925 ^ n992 ^ x42 ;
  assign n3966 = n3965 ^ n321 ^ x79 ;
  assign n3967 = ( x162 & ~n2072 ) | ( x162 & n3966 ) | ( ~n2072 & n3966 ) ;
  assign n3968 = n527 | n1685 ;
  assign n3969 = n3968 ^ n1323 ^ 1'b0 ;
  assign n3970 = ( n540 & n3967 ) | ( n540 & n3969 ) | ( n3967 & n3969 ) ;
  assign n3975 = n3974 ^ n3970 ^ n1539 ;
  assign n3976 = n3575 ^ n1690 ^ n1027 ;
  assign n3978 = ( n1026 & n1340 ) | ( n1026 & ~n1609 ) | ( n1340 & ~n1609 ) ;
  assign n3977 = n2724 ^ n1945 ^ n1248 ;
  assign n3979 = n3978 ^ n3977 ^ n1769 ;
  assign n3980 = ( n2536 & ~n3976 ) | ( n2536 & n3979 ) | ( ~n3976 & n3979 ) ;
  assign n3981 = n3651 ^ n2484 ^ x39 ;
  assign n3982 = n3981 ^ n2638 ^ 1'b0 ;
  assign n3983 = n3980 & ~n3982 ;
  assign n3984 = n3983 ^ n3931 ^ 1'b0 ;
  assign n3985 = n1882 & n3984 ;
  assign n3986 = n1898 ^ n1509 ^ n1265 ;
  assign n3987 = n3986 ^ n3979 ^ 1'b0 ;
  assign n3988 = n3987 ^ n3629 ^ n760 ;
  assign n3989 = n401 | n1544 ;
  assign n3990 = n3134 & n3989 ;
  assign n3995 = n2452 ^ n2392 ^ n735 ;
  assign n3991 = n1898 ^ n1437 ^ n896 ;
  assign n3992 = n2889 | n3991 ;
  assign n3993 = n3992 ^ n1316 ^ 1'b0 ;
  assign n3994 = n1181 & n3993 ;
  assign n3996 = n3995 ^ n3994 ^ 1'b0 ;
  assign n3997 = ( x69 & n626 ) | ( x69 & n1296 ) | ( n626 & n1296 ) ;
  assign n3998 = n2054 ^ n856 ^ 1'b0 ;
  assign n3999 = n3998 ^ n3967 ^ n1994 ;
  assign n4001 = n2714 ^ n2081 ^ n1060 ;
  assign n4000 = n3854 ^ n987 ^ n340 ;
  assign n4002 = n4001 ^ n4000 ^ n1920 ;
  assign n4003 = n2988 ^ n1778 ^ n1457 ;
  assign n4004 = n4003 ^ n1179 ^ 1'b0 ;
  assign n4005 = n1719 ^ n1131 ^ x210 ;
  assign n4006 = n2070 & ~n4005 ;
  assign n4007 = n4004 & n4006 ;
  assign n4008 = n4002 & n4007 ;
  assign n4009 = ( ~n418 & n3864 ) | ( ~n418 & n4008 ) | ( n3864 & n4008 ) ;
  assign n4010 = ( ~x239 & n1466 ) | ( ~x239 & n1530 ) | ( n1466 & n1530 ) ;
  assign n4011 = n4010 ^ n2905 ^ n1320 ;
  assign n4012 = n3975 | n4011 ;
  assign n4013 = ( n1449 & n2455 ) | ( n1449 & n2786 ) | ( n2455 & n2786 ) ;
  assign n4014 = n4013 ^ n2206 ^ x149 ;
  assign n4015 = n2052 ^ n1880 ^ n284 ;
  assign n4016 = n4015 ^ n3934 ^ n3482 ;
  assign n4021 = n559 & ~n1204 ;
  assign n4022 = ~n1876 & n4021 ;
  assign n4017 = n2341 ^ n1368 ^ n1201 ;
  assign n4018 = n1679 ^ n825 ^ n580 ;
  assign n4019 = n4018 ^ n562 ^ x52 ;
  assign n4020 = n4017 & n4019 ;
  assign n4023 = n4022 ^ n4020 ^ 1'b0 ;
  assign n4024 = n762 | n4023 ;
  assign n4025 = n2943 & n3492 ;
  assign n4026 = ( x29 & n2894 ) | ( x29 & ~n3868 ) | ( n2894 & ~n3868 ) ;
  assign n4027 = ( n438 & n1679 ) | ( n438 & ~n4026 ) | ( n1679 & ~n4026 ) ;
  assign n4029 = n2794 & n2835 ;
  assign n4028 = n1569 | n1722 ;
  assign n4030 = n4029 ^ n4028 ^ 1'b0 ;
  assign n4032 = ( n453 & n1101 ) | ( n453 & ~n2809 ) | ( n1101 & ~n2809 ) ;
  assign n4033 = n1929 & n4032 ;
  assign n4034 = ( n643 & ~n2562 ) | ( n643 & n4033 ) | ( ~n2562 & n4033 ) ;
  assign n4035 = n4034 ^ n3323 ^ 1'b0 ;
  assign n4036 = ( n674 & n2950 ) | ( n674 & ~n4035 ) | ( n2950 & ~n4035 ) ;
  assign n4031 = n916 & n2854 ;
  assign n4037 = n4036 ^ n4031 ^ 1'b0 ;
  assign n4038 = ~n4030 & n4037 ;
  assign n4039 = ( n368 & n2109 ) | ( n368 & ~n2691 ) | ( n2109 & ~n2691 ) ;
  assign n4040 = n4039 ^ x159 ^ 1'b0 ;
  assign n4041 = ~n836 & n2664 ;
  assign n4042 = n4040 & n4041 ;
  assign n4043 = n2148 ^ n1659 ^ 1'b0 ;
  assign n4044 = n2641 ^ n1516 ^ n1320 ;
  assign n4045 = n1643 | n4044 ;
  assign n4046 = ~n2909 & n3163 ;
  assign n4049 = ( n2197 & n2216 ) | ( n2197 & n2254 ) | ( n2216 & n2254 ) ;
  assign n4050 = ( ~n526 & n945 ) | ( ~n526 & n4049 ) | ( n945 & n4049 ) ;
  assign n4047 = n1544 ^ n811 ^ n347 ;
  assign n4048 = ( ~x160 & n3171 ) | ( ~x160 & n4047 ) | ( n3171 & n4047 ) ;
  assign n4051 = n4050 ^ n4048 ^ n572 ;
  assign n4052 = n3849 ^ n331 ^ x135 ;
  assign n4053 = n4052 ^ n3222 ^ 1'b0 ;
  assign n4054 = ~n3303 & n4053 ;
  assign n4055 = ~n520 & n4054 ;
  assign n4056 = n4055 ^ n3240 ^ 1'b0 ;
  assign n4057 = n2232 ^ n637 ^ 1'b0 ;
  assign n4058 = ~n688 & n3765 ;
  assign n4059 = n2298 & n4058 ;
  assign n4060 = ( ~n1420 & n1485 ) | ( ~n1420 & n4059 ) | ( n1485 & n4059 ) ;
  assign n4061 = n865 & ~n1391 ;
  assign n4062 = n4061 ^ n1093 ^ 1'b0 ;
  assign n4063 = ( ~n845 & n2433 ) | ( ~n845 & n4062 ) | ( n2433 & n4062 ) ;
  assign n4064 = n4063 ^ n1661 ^ 1'b0 ;
  assign n4065 = n3948 ^ n1736 ^ 1'b0 ;
  assign n4066 = n1113 & n4065 ;
  assign n4067 = n1217 | n3007 ;
  assign n4068 = n1392 ^ n447 ^ n269 ;
  assign n4069 = n4068 ^ n2203 ^ n1301 ;
  assign n4070 = ~n1419 & n4069 ;
  assign n4071 = n447 & ~n1106 ;
  assign n4072 = n310 & n4071 ;
  assign n4073 = n4070 | n4072 ;
  assign n4074 = n4073 ^ x58 ^ 1'b0 ;
  assign n4075 = n4074 ^ n1880 ^ n830 ;
  assign n4076 = n2910 ^ n1392 ^ 1'b0 ;
  assign n4077 = n2526 & ~n4076 ;
  assign n4078 = ( ~n1003 & n3515 ) | ( ~n1003 & n4077 ) | ( n3515 & n4077 ) ;
  assign n4079 = ( n2300 & ~n2531 ) | ( n2300 & n4078 ) | ( ~n2531 & n4078 ) ;
  assign n4080 = ( ~x245 & n406 ) | ( ~x245 & n1242 ) | ( n406 & n1242 ) ;
  assign n4081 = ( n766 & ~n2720 ) | ( n766 & n4080 ) | ( ~n2720 & n4080 ) ;
  assign n4082 = n3443 & ~n3828 ;
  assign n4083 = ~n2432 & n4082 ;
  assign n4084 = ( ~n933 & n1325 ) | ( ~n933 & n1554 ) | ( n1325 & n1554 ) ;
  assign n4085 = n4084 ^ n1795 ^ 1'b0 ;
  assign n4086 = n503 & ~n4085 ;
  assign n4087 = ( ~x144 & x198 ) | ( ~x144 & n2887 ) | ( x198 & n2887 ) ;
  assign n4088 = n4086 & ~n4087 ;
  assign n4089 = n4088 ^ x126 ^ 1'b0 ;
  assign n4090 = n4089 ^ n1292 ^ n471 ;
  assign n4091 = ( n4081 & n4083 ) | ( n4081 & n4090 ) | ( n4083 & n4090 ) ;
  assign n4092 = n3360 ^ n2016 ^ x233 ;
  assign n4093 = ( n988 & n1855 ) | ( n988 & ~n4092 ) | ( n1855 & ~n4092 ) ;
  assign n4095 = ~n581 & n2160 ;
  assign n4096 = n4095 ^ n366 ^ 1'b0 ;
  assign n4094 = n2684 ^ n2080 ^ 1'b0 ;
  assign n4097 = n4096 ^ n4094 ^ n398 ;
  assign n4098 = n1906 ^ n719 ^ 1'b0 ;
  assign n4099 = x228 & ~n4098 ;
  assign n4100 = n4099 ^ n2519 ^ n2162 ;
  assign n4101 = n1537 & n1803 ;
  assign n4102 = ( ~x24 & n4100 ) | ( ~x24 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = n1758 & ~n4102 ;
  assign n4104 = ~n1661 & n4103 ;
  assign n4108 = n1147 ^ n747 ^ 1'b0 ;
  assign n4105 = n353 & ~n2934 ;
  assign n4106 = n4105 ^ n3616 ^ 1'b0 ;
  assign n4107 = ~n3104 & n4106 ;
  assign n4109 = n4108 ^ n4107 ^ 1'b0 ;
  assign n4111 = n1096 & n1452 ;
  assign n4112 = n4111 ^ n620 ^ 1'b0 ;
  assign n4110 = n1323 & ~n2355 ;
  assign n4113 = n4112 ^ n4110 ^ n3779 ;
  assign n4114 = n3433 ^ n3160 ^ 1'b0 ;
  assign n4115 = n2950 & n4114 ;
  assign n4116 = n4115 ^ n3371 ^ x198 ;
  assign n4117 = ~n958 & n2278 ;
  assign n4118 = n4117 ^ n823 ^ 1'b0 ;
  assign n4119 = n3701 ^ n2547 ^ x92 ;
  assign n4120 = x118 & ~n3341 ;
  assign n4121 = n4120 ^ n1291 ^ 1'b0 ;
  assign n4122 = n2659 & ~n4121 ;
  assign n4123 = ( n870 & ~n1200 ) | ( n870 & n2146 ) | ( ~n1200 & n2146 ) ;
  assign n4124 = ~n4122 & n4123 ;
  assign n4135 = n1763 ^ n1118 ^ 1'b0 ;
  assign n4125 = n2960 ^ n886 ^ 1'b0 ;
  assign n4126 = n1093 & n4125 ;
  assign n4127 = n1339 ^ n633 ^ 1'b0 ;
  assign n4128 = ~n2605 & n4127 ;
  assign n4129 = n4128 ^ n2317 ^ 1'b0 ;
  assign n4130 = n4126 & n4129 ;
  assign n4131 = ( ~n655 & n1554 ) | ( ~n655 & n4130 ) | ( n1554 & n4130 ) ;
  assign n4132 = n373 & ~n2935 ;
  assign n4133 = n2187 | n4132 ;
  assign n4134 = n4131 | n4133 ;
  assign n4136 = n4135 ^ n4134 ^ n2540 ;
  assign n4137 = n3469 ^ n2309 ^ 1'b0 ;
  assign n4138 = ( n653 & n1180 ) | ( n653 & n4137 ) | ( n1180 & n4137 ) ;
  assign n4139 = ( ~n461 & n833 ) | ( ~n461 & n2178 ) | ( n833 & n2178 ) ;
  assign n4140 = n3844 ^ n1244 ^ 1'b0 ;
  assign n4141 = n2459 | n4140 ;
  assign n4142 = ( n544 & ~n4139 ) | ( n544 & n4141 ) | ( ~n4139 & n4141 ) ;
  assign n4143 = x210 & ~n4025 ;
  assign n4144 = n1977 & n3961 ;
  assign n4145 = ( ~n1703 & n4143 ) | ( ~n1703 & n4144 ) | ( n4143 & n4144 ) ;
  assign n4152 = n2849 ^ n616 ^ 1'b0 ;
  assign n4153 = n4152 ^ n1500 ^ 1'b0 ;
  assign n4154 = ~n2740 & n4153 ;
  assign n4146 = n525 & n981 ;
  assign n4147 = ~n416 & n4146 ;
  assign n4148 = ~n528 & n4147 ;
  assign n4149 = n4148 ^ x120 ^ 1'b0 ;
  assign n4150 = n4149 ^ n1759 ^ 1'b0 ;
  assign n4151 = n4150 ^ n4005 ^ n814 ;
  assign n4155 = n4154 ^ n4151 ^ 1'b0 ;
  assign n4156 = n2728 ^ x174 ^ 1'b0 ;
  assign n4157 = ~n308 & n3493 ;
  assign n4158 = n4157 ^ x68 ^ 1'b0 ;
  assign n4159 = n3889 & ~n4158 ;
  assign n4160 = n4159 ^ n3137 ^ n1052 ;
  assign n4161 = ( n2507 & ~n4156 ) | ( n2507 & n4160 ) | ( ~n4156 & n4160 ) ;
  assign n4170 = n3959 ^ n936 ^ 1'b0 ;
  assign n4168 = ( n541 & ~n1449 ) | ( n541 & n2103 ) | ( ~n1449 & n2103 ) ;
  assign n4169 = ( n1514 & ~n1999 ) | ( n1514 & n4168 ) | ( ~n1999 & n4168 ) ;
  assign n4171 = n4170 ^ n4169 ^ n264 ;
  assign n4165 = n2704 ^ n678 ^ n480 ;
  assign n4163 = n2763 ^ n2621 ^ n1464 ;
  assign n4162 = n1741 & n1879 ;
  assign n4164 = n4163 ^ n4162 ^ 1'b0 ;
  assign n4166 = n4165 ^ n4164 ^ 1'b0 ;
  assign n4167 = n1835 & n4166 ;
  assign n4172 = n4171 ^ n4167 ^ 1'b0 ;
  assign n4173 = n394 & n1406 ;
  assign n4174 = ~n3027 & n4173 ;
  assign n4175 = n3485 ^ n2770 ^ 1'b0 ;
  assign n4176 = n4175 ^ n3767 ^ n1820 ;
  assign n4177 = n4176 ^ n898 ^ n350 ;
  assign n4178 = n4177 ^ n4056 ^ n2321 ;
  assign n4179 = n579 | n947 ;
  assign n4180 = ( x128 & n930 ) | ( x128 & ~n1716 ) | ( n930 & ~n1716 ) ;
  assign n4181 = ( x228 & ~n1091 ) | ( x228 & n1571 ) | ( ~n1091 & n1571 ) ;
  assign n4182 = n4180 & n4181 ;
  assign n4183 = n950 & n4182 ;
  assign n4184 = ~n4179 & n4183 ;
  assign n4185 = x91 & ~n2901 ;
  assign n4186 = ~x21 & n4185 ;
  assign n4188 = n450 ^ x126 ^ 1'b0 ;
  assign n4189 = ( ~n490 & n1897 ) | ( ~n490 & n4188 ) | ( n1897 & n4188 ) ;
  assign n4190 = ( n352 & n974 ) | ( n352 & ~n4189 ) | ( n974 & ~n4189 ) ;
  assign n4187 = x22 & ~n1905 ;
  assign n4191 = n4190 ^ n4187 ^ 1'b0 ;
  assign n4192 = ( n2318 & ~n4186 ) | ( n2318 & n4191 ) | ( ~n4186 & n4191 ) ;
  assign n4193 = n745 & n1535 ;
  assign n4194 = n4193 ^ n534 ^ 1'b0 ;
  assign n4196 = ( x30 & n684 ) | ( x30 & ~n1031 ) | ( n684 & ~n1031 ) ;
  assign n4195 = ~n1307 & n1477 ;
  assign n4197 = n4196 ^ n4195 ^ 1'b0 ;
  assign n4198 = ( n1546 & ~n3441 ) | ( n1546 & n4197 ) | ( ~n3441 & n4197 ) ;
  assign n4199 = n4198 ^ n751 ^ 1'b0 ;
  assign n4200 = ~n4194 & n4199 ;
  assign n4201 = ( ~n1705 & n1852 ) | ( ~n1705 & n3574 ) | ( n1852 & n3574 ) ;
  assign n4202 = n3611 | n4201 ;
  assign n4203 = n1576 ^ n334 ^ 1'b0 ;
  assign n4204 = n4203 ^ n619 ^ n545 ;
  assign n4205 = n1271 ^ n1241 ^ n270 ;
  assign n4206 = n4205 ^ n958 ^ 1'b0 ;
  assign n4207 = n4206 ^ n3654 ^ n798 ;
  assign n4208 = ~n3727 & n4207 ;
  assign n4209 = n597 | n2399 ;
  assign n4210 = n1784 & ~n2718 ;
  assign n4211 = ~n4209 & n4210 ;
  assign n4212 = n1603 | n4211 ;
  assign n4213 = n2070 ^ n1787 ^ n1421 ;
  assign n4214 = n1093 & n2266 ;
  assign n4215 = ~n509 & n4214 ;
  assign n4216 = ( x92 & n1544 ) | ( x92 & ~n2540 ) | ( n1544 & ~n2540 ) ;
  assign n4217 = ( x17 & ~n1710 ) | ( x17 & n1965 ) | ( ~n1710 & n1965 ) ;
  assign n4218 = n4175 ^ n2377 ^ 1'b0 ;
  assign n4219 = n4217 & n4218 ;
  assign n4225 = n1988 ^ n1761 ^ n1099 ;
  assign n4220 = x224 & n1070 ;
  assign n4221 = n4220 ^ n507 ^ 1'b0 ;
  assign n4222 = n1980 ^ x185 ^ 1'b0 ;
  assign n4223 = n4221 | n4222 ;
  assign n4224 = ( n568 & ~n2754 ) | ( n568 & n4223 ) | ( ~n2754 & n4223 ) ;
  assign n4226 = n4225 ^ n4224 ^ n330 ;
  assign n4227 = n4226 ^ n841 ^ 1'b0 ;
  assign n4228 = x192 & ~n4227 ;
  assign n4229 = ( x0 & n3139 ) | ( x0 & n4228 ) | ( n3139 & n4228 ) ;
  assign n4230 = ( n898 & n3465 ) | ( n898 & n4229 ) | ( n3465 & n4229 ) ;
  assign n4231 = n4219 & n4230 ;
  assign n4232 = n4216 & n4231 ;
  assign n4233 = n1033 ^ n943 ^ 1'b0 ;
  assign n4234 = n1294 | n4233 ;
  assign n4235 = n4234 ^ n3767 ^ 1'b0 ;
  assign n4236 = n3065 | n4235 ;
  assign n4237 = n3632 ^ x233 ^ 1'b0 ;
  assign n4238 = ( n458 & n2553 ) | ( n458 & ~n3980 ) | ( n2553 & ~n3980 ) ;
  assign n4239 = n3888 ^ n3551 ^ n3130 ;
  assign n4240 = n1431 ^ n592 ^ 1'b0 ;
  assign n4241 = n4240 ^ n1400 ^ n1376 ;
  assign n4242 = x130 & ~n3481 ;
  assign n4243 = n4242 ^ n1305 ^ 1'b0 ;
  assign n4244 = ~n1933 & n2726 ;
  assign n4245 = ~n4243 & n4244 ;
  assign n4246 = n4245 ^ n2614 ^ 1'b0 ;
  assign n4247 = n4241 & ~n4246 ;
  assign n4248 = n3244 ^ n1418 ^ x44 ;
  assign n4249 = n4248 ^ n3877 ^ n455 ;
  assign n4250 = n4249 ^ n3261 ^ 1'b0 ;
  assign n4251 = n408 | n1655 ;
  assign n4252 = n2432 | n4251 ;
  assign n4253 = n4250 & n4252 ;
  assign n4254 = ~x137 & n4253 ;
  assign n4259 = n4068 ^ n2425 ^ 1'b0 ;
  assign n4260 = n1631 | n4259 ;
  assign n4257 = n1127 ^ n331 ^ 1'b0 ;
  assign n4256 = ( ~n2406 & n3967 ) | ( ~n2406 & n4148 ) | ( n3967 & n4148 ) ;
  assign n4255 = n2613 | n3359 ;
  assign n4258 = n4257 ^ n4256 ^ n4255 ;
  assign n4261 = n4260 ^ n4258 ^ n3894 ;
  assign n4262 = n2953 & ~n3514 ;
  assign n4263 = n2515 ^ n2241 ^ n1406 ;
  assign n4264 = n4263 ^ n1785 ^ n983 ;
  assign n4266 = n2791 ^ x250 ^ 1'b0 ;
  assign n4267 = ~n680 & n4266 ;
  assign n4265 = ( n904 & ~n1181 ) | ( n904 & n2488 ) | ( ~n1181 & n2488 ) ;
  assign n4268 = n4267 ^ n4265 ^ n1930 ;
  assign n4269 = n1520 & ~n2058 ;
  assign n4273 = n4180 ^ n559 ^ x30 ;
  assign n4270 = n723 & n846 ;
  assign n4271 = ~n585 & n4270 ;
  assign n4272 = ( n2388 & ~n3101 ) | ( n2388 & n4271 ) | ( ~n3101 & n4271 ) ;
  assign n4274 = n4273 ^ n4272 ^ 1'b0 ;
  assign n4275 = n2546 & n4274 ;
  assign n4276 = ~n1054 & n4275 ;
  assign n4277 = n2646 & n4276 ;
  assign n4278 = n4277 ^ n903 ^ n550 ;
  assign n4283 = n1261 ^ n1046 ^ n494 ;
  assign n4284 = n4283 ^ n2021 ^ n1091 ;
  assign n4281 = ( x68 & ~n580 ) | ( x68 & n827 ) | ( ~n580 & n827 ) ;
  assign n4279 = ~x187 & n2836 ;
  assign n4280 = n704 & ~n4279 ;
  assign n4282 = n4281 ^ n4280 ^ 1'b0 ;
  assign n4285 = n4284 ^ n4282 ^ n1856 ;
  assign n4286 = ( n503 & n1268 ) | ( n503 & ~n1502 ) | ( n1268 & ~n1502 ) ;
  assign n4287 = n296 & n4286 ;
  assign n4288 = ~n3497 & n4287 ;
  assign n4289 = ( n2283 & n3732 ) | ( n2283 & ~n4288 ) | ( n3732 & ~n4288 ) ;
  assign n4290 = n293 | n581 ;
  assign n4291 = n371 & ~n4290 ;
  assign n4292 = n4291 ^ n1625 ^ 1'b0 ;
  assign n4295 = ( n257 & ~n557 ) | ( n257 & n1248 ) | ( ~n557 & n1248 ) ;
  assign n4296 = n4295 ^ n1620 ^ 1'b0 ;
  assign n4297 = n4296 ^ n1173 ^ 1'b0 ;
  assign n4293 = ( n1507 & n1585 ) | ( n1507 & n3155 ) | ( n1585 & n3155 ) ;
  assign n4294 = n4293 ^ x80 ^ 1'b0 ;
  assign n4298 = n4297 ^ n4294 ^ 1'b0 ;
  assign n4305 = ( n781 & n2068 ) | ( n781 & n3340 ) | ( n2068 & n3340 ) ;
  assign n4306 = n4305 ^ n1747 ^ 1'b0 ;
  assign n4303 = n2089 ^ n1449 ^ n733 ;
  assign n4302 = ( x40 & ~n943 ) | ( x40 & n999 ) | ( ~n943 & n999 ) ;
  assign n4301 = ~n3516 & n4180 ;
  assign n4304 = n4303 ^ n4302 ^ n4301 ;
  assign n4299 = n2820 & n3644 ;
  assign n4300 = ( x114 & n1602 ) | ( x114 & n4299 ) | ( n1602 & n4299 ) ;
  assign n4307 = n4306 ^ n4304 ^ n4300 ;
  assign n4308 = n2593 ^ n2086 ^ 1'b0 ;
  assign n4309 = n3061 | n4308 ;
  assign n4310 = n4249 | n4309 ;
  assign n4311 = n578 | n796 ;
  assign n4312 = n4311 ^ n1267 ^ n562 ;
  assign n4313 = n261 | n444 ;
  assign n4314 = n4312 | n4313 ;
  assign n4315 = ~n4310 & n4314 ;
  assign n4316 = n4315 ^ n419 ^ 1'b0 ;
  assign n4317 = ~n2147 & n3965 ;
  assign n4318 = n4317 ^ n938 ^ 1'b0 ;
  assign n4319 = n4318 ^ n2819 ^ 1'b0 ;
  assign n4323 = n3450 ^ n729 ^ 1'b0 ;
  assign n4320 = n2108 ^ n1707 ^ 1'b0 ;
  assign n4321 = x33 & ~n813 ;
  assign n4322 = ~n4320 & n4321 ;
  assign n4324 = n4323 ^ n4322 ^ n1305 ;
  assign n4325 = n3189 ^ n580 ^ 1'b0 ;
  assign n4326 = n4325 ^ n3461 ^ n441 ;
  assign n4327 = n491 & ~n4326 ;
  assign n4328 = n2945 ^ n2683 ^ 1'b0 ;
  assign n4329 = x2 & n4328 ;
  assign n4332 = ( n1447 & ~n3143 ) | ( n1447 & n3438 ) | ( ~n3143 & n3438 ) ;
  assign n4333 = n4332 ^ n3524 ^ n2081 ;
  assign n4331 = n2169 ^ n1643 ^ n692 ;
  assign n4330 = n3817 ^ n407 ^ n367 ;
  assign n4334 = n4333 ^ n4331 ^ n4330 ;
  assign n4335 = n4334 ^ n3567 ^ n2666 ;
  assign n4336 = n1804 | n4206 ;
  assign n4337 = n1916 & n4336 ;
  assign n4338 = ~n773 & n1360 ;
  assign n4339 = ( n480 & n1737 ) | ( n480 & n2866 ) | ( n1737 & n2866 ) ;
  assign n4340 = ( n1196 & ~n1605 ) | ( n1196 & n1635 ) | ( ~n1605 & n1635 ) ;
  assign n4341 = n1728 ^ n634 ^ 1'b0 ;
  assign n4342 = n2581 ^ n552 ^ 1'b0 ;
  assign n4343 = n3583 ^ x89 ^ 1'b0 ;
  assign n4344 = n1488 & n4343 ;
  assign n4345 = ~n1032 & n4344 ;
  assign n4346 = n2512 & n4345 ;
  assign n4347 = ~n1486 & n4346 ;
  assign n4348 = ( n4341 & n4342 ) | ( n4341 & ~n4347 ) | ( n4342 & ~n4347 ) ;
  assign n4349 = n4348 ^ n3624 ^ n1553 ;
  assign n4350 = ( ~n3528 & n4340 ) | ( ~n3528 & n4349 ) | ( n4340 & n4349 ) ;
  assign n4351 = n2750 ^ n1106 ^ 1'b0 ;
  assign n4352 = ( n2123 & ~n2884 ) | ( n2123 & n3363 ) | ( ~n2884 & n3363 ) ;
  assign n4353 = n2945 ^ n920 ^ 1'b0 ;
  assign n4354 = n2451 | n4353 ;
  assign n4355 = n4354 ^ n1968 ^ n1933 ;
  assign n4356 = n1776 & ~n4355 ;
  assign n4357 = n3501 & n4356 ;
  assign n4358 = n3082 | n4357 ;
  assign n4359 = n3619 ^ n1725 ^ n808 ;
  assign n4360 = n4359 ^ n3247 ^ 1'b0 ;
  assign n4361 = x146 | n4360 ;
  assign n4363 = ( x72 & ~n1377 ) | ( x72 & n1446 ) | ( ~n1377 & n1446 ) ;
  assign n4364 = n2085 | n4363 ;
  assign n4365 = n1424 & ~n4364 ;
  assign n4366 = ( x65 & n1567 ) | ( x65 & ~n4365 ) | ( n1567 & ~n4365 ) ;
  assign n4367 = n4366 ^ n1546 ^ 1'b0 ;
  assign n4368 = n818 & ~n4367 ;
  assign n4362 = n2904 ^ n2793 ^ n1629 ;
  assign n4369 = n4368 ^ n4362 ^ n4087 ;
  assign n4370 = n3967 ^ n1505 ^ 1'b0 ;
  assign n4371 = ~n920 & n4370 ;
  assign n4372 = n4371 ^ n3696 ^ n1358 ;
  assign n4373 = n3963 ^ n3376 ^ n2185 ;
  assign n4378 = n842 ^ x225 ^ 1'b0 ;
  assign n4379 = n635 & n4378 ;
  assign n4374 = n3670 ^ n349 ^ 1'b0 ;
  assign n4375 = n1298 & n4374 ;
  assign n4376 = n4375 ^ n2494 ^ n2438 ;
  assign n4377 = n2859 | n4376 ;
  assign n4380 = n4379 ^ n4377 ^ 1'b0 ;
  assign n4398 = n3969 ^ n870 ^ n368 ;
  assign n4399 = ( n1548 & ~n3724 ) | ( n1548 & n4398 ) | ( ~n3724 & n4398 ) ;
  assign n4393 = n1261 & n2581 ;
  assign n4394 = n4393 ^ x250 ^ 1'b0 ;
  assign n4395 = n4394 ^ x143 ^ 1'b0 ;
  assign n4396 = n1317 | n4395 ;
  assign n4386 = n1890 & ~n1947 ;
  assign n4387 = n1928 & n2935 ;
  assign n4388 = ~n1850 & n4387 ;
  assign n4389 = n4388 ^ n1546 ^ n459 ;
  assign n4390 = ~n4386 & n4389 ;
  assign n4391 = n4390 ^ n1475 ^ 1'b0 ;
  assign n4381 = ~n466 & n2890 ;
  assign n4382 = n3811 ^ n486 ^ 1'b0 ;
  assign n4383 = ~n4381 & n4382 ;
  assign n4384 = ( n355 & ~n3254 ) | ( n355 & n4383 ) | ( ~n3254 & n4383 ) ;
  assign n4385 = n1784 & n4384 ;
  assign n4392 = n4391 ^ n4385 ^ 1'b0 ;
  assign n4397 = n4396 ^ n4392 ^ n1980 ;
  assign n4400 = n4399 ^ n4397 ^ n3541 ;
  assign n4401 = n2477 ^ n1711 ^ x168 ;
  assign n4402 = ~n1527 & n2200 ;
  assign n4403 = n2923 & n4402 ;
  assign n4404 = n2113 & n4403 ;
  assign n4405 = ( x19 & n1262 ) | ( x19 & ~n4404 ) | ( n1262 & ~n4404 ) ;
  assign n4406 = n3601 ^ n2033 ^ n1976 ;
  assign n4407 = n2890 ^ n2321 ^ 1'b0 ;
  assign n4408 = n4407 ^ n2073 ^ n1447 ;
  assign n4409 = n4408 ^ n4396 ^ 1'b0 ;
  assign n4410 = ~n1714 & n4409 ;
  assign n4411 = n773 & ~n1487 ;
  assign n4412 = n4410 & ~n4411 ;
  assign n4413 = n4412 ^ n2689 ^ 1'b0 ;
  assign n4414 = ( n1843 & n1931 ) | ( n1843 & n3872 ) | ( n1931 & n3872 ) ;
  assign n4415 = n3286 ^ n2066 ^ 1'b0 ;
  assign n4419 = n4164 ^ n2918 ^ n2508 ;
  assign n4420 = n2925 ^ x254 ^ 1'b0 ;
  assign n4421 = n1616 & ~n4420 ;
  assign n4422 = ( n3239 & n4419 ) | ( n3239 & n4421 ) | ( n4419 & n4421 ) ;
  assign n4416 = n501 & n592 ;
  assign n4417 = n3071 & n4416 ;
  assign n4418 = ( n1870 & n2381 ) | ( n1870 & n4417 ) | ( n2381 & n4417 ) ;
  assign n4423 = n4422 ^ n4418 ^ n4123 ;
  assign n4424 = n2800 ^ x45 ^ x9 ;
  assign n4425 = n3061 ^ n2491 ^ 1'b0 ;
  assign n4426 = ( ~n563 & n3025 ) | ( ~n563 & n3350 ) | ( n3025 & n3350 ) ;
  assign n4427 = n3772 ^ n3120 ^ n1204 ;
  assign n4428 = ( n337 & n4426 ) | ( n337 & n4427 ) | ( n4426 & n4427 ) ;
  assign n4430 = n1759 ^ n453 ^ 1'b0 ;
  assign n4431 = n3226 & ~n4430 ;
  assign n4432 = ( n1207 & n1349 ) | ( n1207 & n4431 ) | ( n1349 & n4431 ) ;
  assign n4429 = ( n859 & n2443 ) | ( n859 & n3399 ) | ( n2443 & n3399 ) ;
  assign n4433 = n4432 ^ n4429 ^ n3192 ;
  assign n4434 = n4433 ^ n4235 ^ n993 ;
  assign n4438 = n3368 ^ n1754 ^ n1404 ;
  assign n4435 = n2009 ^ n1824 ^ 1'b0 ;
  assign n4436 = n4005 | n4435 ;
  assign n4437 = n4436 ^ n3651 ^ 1'b0 ;
  assign n4439 = n4438 ^ n4437 ^ n4275 ;
  assign n4440 = ( n1570 & n3049 ) | ( n1570 & n4029 ) | ( n3049 & n4029 ) ;
  assign n4441 = ( n293 & ~n1766 ) | ( n293 & n2786 ) | ( ~n1766 & n2786 ) ;
  assign n4442 = n4441 ^ n2901 ^ n1634 ;
  assign n4443 = x3 & n4442 ;
  assign n4444 = n4443 ^ n2348 ^ 1'b0 ;
  assign n4445 = n2345 ^ n1378 ^ 1'b0 ;
  assign n4446 = n4445 ^ n3299 ^ n3082 ;
  assign n4447 = ( n2382 & ~n4444 ) | ( n2382 & n4446 ) | ( ~n4444 & n4446 ) ;
  assign n4448 = ( n2336 & ~n4070 ) | ( n2336 & n4447 ) | ( ~n4070 & n4447 ) ;
  assign n4449 = ( n1067 & n1232 ) | ( n1067 & ~n2400 ) | ( n1232 & ~n2400 ) ;
  assign n4450 = ( n2441 & ~n3278 ) | ( n2441 & n4449 ) | ( ~n3278 & n4449 ) ;
  assign n4451 = n2108 ^ n956 ^ 1'b0 ;
  assign n4452 = ~n3715 & n4451 ;
  assign n4453 = ( n3189 & n4152 ) | ( n3189 & ~n4452 ) | ( n4152 & ~n4452 ) ;
  assign n4454 = n2436 | n3548 ;
  assign n4455 = n3149 ^ n936 ^ 1'b0 ;
  assign n4456 = ~n2184 & n4455 ;
  assign n4457 = ( n751 & n1530 ) | ( n751 & n2468 ) | ( n1530 & n2468 ) ;
  assign n4458 = x231 & n4457 ;
  assign n4459 = ~x70 & n4458 ;
  assign n4460 = n3849 ^ n2006 ^ n1206 ;
  assign n4461 = n352 | n4460 ;
  assign n4462 = n2254 | n4461 ;
  assign n4463 = ( n3894 & ~n4459 ) | ( n3894 & n4462 ) | ( ~n4459 & n4462 ) ;
  assign n4464 = ( n1471 & n2333 ) | ( n1471 & n4063 ) | ( n2333 & n4063 ) ;
  assign n4466 = n735 ^ x245 ^ 1'b0 ;
  assign n4465 = n681 & n2886 ;
  assign n4467 = n4466 ^ n4465 ^ n2953 ;
  assign n4468 = ( n2560 & ~n3299 ) | ( n2560 & n3907 ) | ( ~n3299 & n3907 ) ;
  assign n4469 = n4468 ^ n2235 ^ n861 ;
  assign n4474 = ( x220 & n942 ) | ( x220 & ~n4295 ) | ( n942 & ~n4295 ) ;
  assign n4471 = ( ~n396 & n446 ) | ( ~n396 & n490 ) | ( n446 & n490 ) ;
  assign n4472 = n4471 ^ n261 ^ 1'b0 ;
  assign n4473 = n3232 & n4472 ;
  assign n4475 = n4474 ^ n4473 ^ 1'b0 ;
  assign n4470 = ( ~n2002 & n2334 ) | ( ~n2002 & n2771 ) | ( n2334 & n2771 ) ;
  assign n4476 = n4475 ^ n4470 ^ 1'b0 ;
  assign n4477 = ( n751 & n1101 ) | ( n751 & n1707 ) | ( n1101 & n1707 ) ;
  assign n4478 = ( x138 & ~n526 ) | ( x138 & n1499 ) | ( ~n526 & n1499 ) ;
  assign n4479 = ( n405 & n1475 ) | ( n405 & ~n4478 ) | ( n1475 & ~n4478 ) ;
  assign n4480 = n4477 & n4479 ;
  assign n4481 = n2470 ^ n1991 ^ n295 ;
  assign n4482 = ( n2105 & n2231 ) | ( n2105 & n4481 ) | ( n2231 & n4481 ) ;
  assign n4483 = n4480 & ~n4482 ;
  assign n4484 = ~n1209 & n4483 ;
  assign n4491 = x215 & n3680 ;
  assign n4492 = n4491 ^ n2845 ^ 1'b0 ;
  assign n4493 = ~n315 & n1158 ;
  assign n4494 = ~n1473 & n4493 ;
  assign n4495 = n4494 ^ x226 ^ 1'b0 ;
  assign n4496 = n4492 & ~n4495 ;
  assign n4485 = n1814 ^ n987 ^ n526 ;
  assign n4486 = n4485 ^ n2310 ^ n369 ;
  assign n4487 = ( x10 & n1394 ) | ( x10 & ~n2360 ) | ( n1394 & ~n2360 ) ;
  assign n4488 = n3097 & ~n4487 ;
  assign n4489 = n4488 ^ n3803 ^ 1'b0 ;
  assign n4490 = ~n4486 & n4489 ;
  assign n4497 = n4496 ^ n4490 ^ 1'b0 ;
  assign n4498 = n993 ^ x37 ^ 1'b0 ;
  assign n4499 = n4498 ^ n2068 ^ n1679 ;
  assign n4500 = n4499 ^ n3091 ^ 1'b0 ;
  assign n4501 = ~n740 & n4500 ;
  assign n4505 = n312 & ~n1493 ;
  assign n4506 = n627 & n4505 ;
  assign n4502 = ( ~n459 & n3293 ) | ( ~n459 & n3514 ) | ( n3293 & n3514 ) ;
  assign n4503 = ( n2213 & n2512 ) | ( n2213 & n3068 ) | ( n2512 & n3068 ) ;
  assign n4504 = n4502 & ~n4503 ;
  assign n4507 = n4506 ^ n4504 ^ 1'b0 ;
  assign n4508 = n4507 ^ n2070 ^ 1'b0 ;
  assign n4509 = n1097 & n4508 ;
  assign n4510 = n1028 ^ n716 ^ n290 ;
  assign n4511 = n4510 ^ n4181 ^ n3381 ;
  assign n4518 = n2115 | n3323 ;
  assign n4513 = n2751 ^ n391 ^ 1'b0 ;
  assign n4514 = ~n2321 & n4513 ;
  assign n4515 = n4514 ^ n2646 ^ n2174 ;
  assign n4516 = n4515 ^ n2545 ^ n1683 ;
  assign n4517 = n4516 ^ n1538 ^ x89 ;
  assign n4512 = n3031 ^ n2894 ^ n511 ;
  assign n4519 = n4518 ^ n4517 ^ n4512 ;
  assign n4520 = n2011 | n3888 ;
  assign n4521 = ~n3433 & n4520 ;
  assign n4523 = ( x227 & n290 ) | ( x227 & ~n1740 ) | ( n290 & ~n1740 ) ;
  assign n4524 = ( ~n523 & n2432 ) | ( ~n523 & n4523 ) | ( n2432 & n4523 ) ;
  assign n4522 = n798 & ~n3920 ;
  assign n4525 = n4524 ^ n4522 ^ 1'b0 ;
  assign n4526 = ( ~x16 & n1327 ) | ( ~x16 & n1697 ) | ( n1327 & n1697 ) ;
  assign n4527 = n1112 & ~n4526 ;
  assign n4528 = n4527 ^ n3270 ^ 1'b0 ;
  assign n4529 = n4410 & ~n4528 ;
  assign n4530 = ( ~n883 & n1747 ) | ( ~n883 & n4529 ) | ( n1747 & n4529 ) ;
  assign n4531 = ( ~x153 & n383 ) | ( ~x153 & n1385 ) | ( n383 & n1385 ) ;
  assign n4532 = n2394 & n3515 ;
  assign n4533 = ~n4531 & n4532 ;
  assign n4534 = n1391 ^ n412 ^ x249 ;
  assign n4535 = ( n1121 & n4533 ) | ( n1121 & n4534 ) | ( n4533 & n4534 ) ;
  assign n4536 = n3824 ^ n2693 ^ n2197 ;
  assign n4537 = n345 ^ x22 ^ 1'b0 ;
  assign n4538 = ( ~x126 & x174 ) | ( ~x126 & n1564 ) | ( x174 & n1564 ) ;
  assign n4539 = ( n405 & n1401 ) | ( n405 & n4538 ) | ( n1401 & n4538 ) ;
  assign n4540 = n4537 | n4539 ;
  assign n4541 = n528 | n1182 ;
  assign n4542 = x27 & n267 ;
  assign n4543 = n4542 ^ n3996 ^ 1'b0 ;
  assign n4544 = n4543 ^ n544 ^ 1'b0 ;
  assign n4545 = n4544 ^ n4388 ^ n4164 ;
  assign n4546 = n4541 & n4545 ;
  assign n4547 = ~n3864 & n4546 ;
  assign n4548 = n2160 ^ n1647 ^ n1629 ;
  assign n4549 = ( n1819 & ~n4438 ) | ( n1819 & n4548 ) | ( ~n4438 & n4548 ) ;
  assign n4550 = n4549 ^ n3866 ^ n929 ;
  assign n4551 = ( x32 & n1251 ) | ( x32 & n4550 ) | ( n1251 & n4550 ) ;
  assign n4552 = n4551 ^ n4112 ^ 1'b0 ;
  assign n4553 = n3181 & ~n4552 ;
  assign n4557 = n3822 ^ x168 ^ 1'b0 ;
  assign n4554 = n4096 ^ n1426 ^ n943 ;
  assign n4555 = n4554 ^ n2993 ^ 1'b0 ;
  assign n4556 = n3562 | n4555 ;
  assign n4558 = n4557 ^ n4556 ^ 1'b0 ;
  assign n4559 = n2833 & n4558 ;
  assign n4560 = ( n1137 & n2778 ) | ( n1137 & ~n3839 ) | ( n2778 & ~n3839 ) ;
  assign n4561 = n3441 | n4560 ;
  assign n4562 = n1967 | n4561 ;
  assign n4563 = ( ~n1232 & n3991 ) | ( ~n1232 & n4526 ) | ( n3991 & n4526 ) ;
  assign n4564 = ( n1419 & n3912 ) | ( n1419 & ~n4470 ) | ( n3912 & ~n4470 ) ;
  assign n4565 = n4563 | n4564 ;
  assign n4566 = n4562 | n4565 ;
  assign n4567 = ( x235 & n1338 ) | ( x235 & ~n4205 ) | ( n1338 & ~n4205 ) ;
  assign n4568 = ( n2185 & ~n2331 ) | ( n2185 & n4567 ) | ( ~n2331 & n4567 ) ;
  assign n4569 = n1299 & n1679 ;
  assign n4570 = x173 & n4569 ;
  assign n4571 = n3695 ^ x168 ^ 1'b0 ;
  assign n4572 = x69 | n4571 ;
  assign n4573 = ~n4570 & n4572 ;
  assign n4574 = ~n332 & n4573 ;
  assign n4575 = n4574 ^ n2132 ^ n1787 ;
  assign n4576 = n2777 ^ n1140 ^ 1'b0 ;
  assign n4577 = n2887 ^ n369 ^ 1'b0 ;
  assign n4578 = n381 & n4577 ;
  assign n4579 = ( n358 & n1498 ) | ( n358 & ~n3360 ) | ( n1498 & ~n3360 ) ;
  assign n4580 = n1697 & n4579 ;
  assign n4581 = n1111 & n4580 ;
  assign n4582 = ( n4576 & n4578 ) | ( n4576 & n4581 ) | ( n4578 & n4581 ) ;
  assign n4583 = n467 & ~n2586 ;
  assign n4584 = ( n2960 & n4582 ) | ( n2960 & n4583 ) | ( n4582 & n4583 ) ;
  assign n4585 = ( ~n425 & n1868 ) | ( ~n425 & n2062 ) | ( n1868 & n2062 ) ;
  assign n4588 = n2283 ^ n1271 ^ 1'b0 ;
  assign n4586 = n2162 ^ n538 ^ x82 ;
  assign n4587 = n1350 & ~n4586 ;
  assign n4589 = n4588 ^ n4587 ^ 1'b0 ;
  assign n4593 = n1423 | n1774 ;
  assign n4590 = ( ~n1161 & n1686 ) | ( ~n1161 & n2901 ) | ( n1686 & n2901 ) ;
  assign n4591 = n4590 ^ n2993 ^ n1632 ;
  assign n4592 = n4591 ^ n947 ^ 1'b0 ;
  assign n4594 = n4593 ^ n4592 ^ 1'b0 ;
  assign n4595 = ( n3453 & n4589 ) | ( n3453 & ~n4594 ) | ( n4589 & ~n4594 ) ;
  assign n4596 = ~n758 & n2345 ;
  assign n4597 = n3366 & n4596 ;
  assign n4598 = n1218 ^ x46 ^ 1'b0 ;
  assign n4599 = n1612 ^ n442 ^ 1'b0 ;
  assign n4600 = ( n2019 & ~n3902 ) | ( n2019 & n4599 ) | ( ~n3902 & n4599 ) ;
  assign n4601 = n4600 ^ n2894 ^ n1747 ;
  assign n4602 = ~n4598 & n4601 ;
  assign n4603 = n4602 ^ n2626 ^ 1'b0 ;
  assign n4604 = n2178 & ~n4603 ;
  assign n4605 = n4604 ^ n773 ^ 1'b0 ;
  assign n4606 = ( n2489 & n4597 ) | ( n2489 & n4605 ) | ( n4597 & n4605 ) ;
  assign n4607 = n4606 ^ n2980 ^ n2674 ;
  assign n4608 = n1012 ^ n731 ^ 1'b0 ;
  assign n4609 = n4608 ^ x227 ^ 1'b0 ;
  assign n4610 = ( n517 & n3668 ) | ( n517 & ~n4609 ) | ( n3668 & ~n4609 ) ;
  assign n4611 = ( n1668 & n2572 ) | ( n1668 & ~n4610 ) | ( n2572 & ~n4610 ) ;
  assign n4612 = ( x206 & n1935 ) | ( x206 & ~n2663 ) | ( n1935 & ~n2663 ) ;
  assign n4617 = x240 & ~n2309 ;
  assign n4618 = ~x60 & n4617 ;
  assign n4619 = n4618 ^ n3731 ^ n2476 ;
  assign n4613 = n3395 ^ n3091 ^ n628 ;
  assign n4614 = ( n1162 & n1758 ) | ( n1162 & n4613 ) | ( n1758 & n4613 ) ;
  assign n4615 = x59 | n885 ;
  assign n4616 = ( n3038 & n4614 ) | ( n3038 & ~n4615 ) | ( n4614 & ~n4615 ) ;
  assign n4620 = n4619 ^ n4616 ^ n3479 ;
  assign n4621 = n3009 ^ n1511 ^ x144 ;
  assign n4622 = n1412 ^ n877 ^ 1'b0 ;
  assign n4623 = n838 & n4622 ;
  assign n4624 = x146 & ~n2605 ;
  assign n4625 = ~n4623 & n4624 ;
  assign n4626 = n4625 ^ n3101 ^ n2332 ;
  assign n4627 = ( x194 & n2514 ) | ( x194 & ~n4626 ) | ( n2514 & ~n4626 ) ;
  assign n4628 = n4627 ^ n2928 ^ n271 ;
  assign n4629 = ( n3614 & n4621 ) | ( n3614 & ~n4628 ) | ( n4621 & ~n4628 ) ;
  assign n4634 = n3332 ^ n1395 ^ x223 ;
  assign n4630 = n1783 ^ n1544 ^ n778 ;
  assign n4631 = n4630 ^ n664 ^ 1'b0 ;
  assign n4632 = n4631 ^ n1085 ^ 1'b0 ;
  assign n4633 = n2619 & ~n4632 ;
  assign n4635 = n4634 ^ n4633 ^ n1718 ;
  assign n4636 = ( ~n2784 & n3244 ) | ( ~n2784 & n4635 ) | ( n3244 & n4635 ) ;
  assign n4637 = n1691 & ~n4636 ;
  assign n4638 = ~n4164 & n4637 ;
  assign n4639 = n3579 | n4638 ;
  assign n4640 = n3306 ^ n2896 ^ 1'b0 ;
  assign n4641 = n771 ^ n519 ^ 1'b0 ;
  assign n4642 = ( n499 & n1246 ) | ( n499 & ~n3963 ) | ( n1246 & ~n3963 ) ;
  assign n4643 = n3638 & n4642 ;
  assign n4644 = n4643 ^ n2410 ^ 1'b0 ;
  assign n4645 = n4644 ^ n3325 ^ n1184 ;
  assign n4646 = ~n4641 & n4645 ;
  assign n4647 = ~n4640 & n4646 ;
  assign n4648 = ~n1504 & n1588 ;
  assign n4649 = ~n3936 & n4648 ;
  assign n4650 = n3776 ^ n803 ^ n571 ;
  assign n4651 = n1056 ^ n1015 ^ x225 ;
  assign n4652 = n4651 ^ n4052 ^ n3267 ;
  assign n4653 = n779 & ~n4652 ;
  assign n4654 = n2286 ^ n1440 ^ n407 ;
  assign n4655 = n4001 ^ n704 ^ 1'b0 ;
  assign n4656 = n899 | n4655 ;
  assign n4657 = n2088 | n4656 ;
  assign n4658 = ( n453 & n2813 ) | ( n453 & n4657 ) | ( n2813 & n4657 ) ;
  assign n4659 = n4654 | n4658 ;
  assign n4660 = n1754 ^ n1241 ^ 1'b0 ;
  assign n4661 = n622 & ~n4660 ;
  assign n4662 = ~x227 & n500 ;
  assign n4663 = ~n783 & n4662 ;
  assign n4664 = n4663 ^ x227 ^ x199 ;
  assign n4665 = n1391 ^ n1209 ^ n430 ;
  assign n4666 = n4665 ^ n2308 ^ n1894 ;
  assign n4667 = ( n4661 & n4664 ) | ( n4661 & ~n4666 ) | ( n4664 & ~n4666 ) ;
  assign n4668 = ( ~n3879 & n4034 ) | ( ~n3879 & n4479 ) | ( n4034 & n4479 ) ;
  assign n4669 = ~n1379 & n4668 ;
  assign n4671 = n1394 | n3198 ;
  assign n4670 = ( ~n2080 & n2325 ) | ( ~n2080 & n2931 ) | ( n2325 & n2931 ) ;
  assign n4672 = n4671 ^ n4670 ^ n3837 ;
  assign n4673 = ( n1466 & ~n3474 ) | ( n1466 & n3772 ) | ( ~n3474 & n3772 ) ;
  assign n4675 = n1746 ^ x233 ^ 1'b0 ;
  assign n4674 = n672 | n4446 ;
  assign n4676 = n4675 ^ n4674 ^ n3889 ;
  assign n4677 = n4676 ^ n4503 ^ n2343 ;
  assign n4678 = ( ~n919 & n4673 ) | ( ~n919 & n4677 ) | ( n4673 & n4677 ) ;
  assign n4679 = n2605 ^ x213 ^ x53 ;
  assign n4680 = n3299 ^ n2055 ^ x238 ;
  assign n4681 = n4680 ^ n394 ^ x80 ;
  assign n4712 = ~n2144 & n2526 ;
  assign n4708 = x187 & n2218 ;
  assign n4709 = n4708 ^ n2092 ^ 1'b0 ;
  assign n4702 = ( ~n868 & n2360 ) | ( ~n868 & n3288 ) | ( n2360 & n3288 ) ;
  assign n4703 = ( ~n3180 & n3333 ) | ( ~n3180 & n4702 ) | ( n3333 & n4702 ) ;
  assign n4704 = ( ~x148 & n1385 ) | ( ~x148 & n3088 ) | ( n1385 & n3088 ) ;
  assign n4705 = ( ~n1555 & n4703 ) | ( ~n1555 & n4704 ) | ( n4703 & n4704 ) ;
  assign n4706 = ~n341 & n4705 ;
  assign n4699 = n3096 ^ n1367 ^ 1'b0 ;
  assign n4700 = n1327 & n4699 ;
  assign n4701 = n4700 ^ n4628 ^ n1950 ;
  assign n4707 = n4706 ^ n4701 ^ n1334 ;
  assign n4696 = ~n283 & n537 ;
  assign n4697 = n4696 ^ n598 ^ 1'b0 ;
  assign n4682 = n3854 ^ n3192 ^ x230 ;
  assign n4683 = n4682 ^ n3260 ^ 1'b0 ;
  assign n4684 = n3644 & n4683 ;
  assign n4689 = n4062 ^ n927 ^ n603 ;
  assign n4690 = n4689 ^ n2263 ^ 1'b0 ;
  assign n4691 = x52 & n4690 ;
  assign n4685 = n3520 ^ n1009 ^ x32 ;
  assign n4686 = n840 & ~n4001 ;
  assign n4687 = n1569 & n4686 ;
  assign n4688 = ~n4685 & n4687 ;
  assign n4692 = n4691 ^ n4688 ^ n3808 ;
  assign n4693 = ( x225 & ~n4684 ) | ( x225 & n4692 ) | ( ~n4684 & n4692 ) ;
  assign n4694 = n4139 ^ n870 ^ n667 ;
  assign n4695 = n4693 | n4694 ;
  assign n4698 = n4697 ^ n4695 ^ 1'b0 ;
  assign n4710 = n4709 ^ n4707 ^ n4698 ;
  assign n4711 = ~n3518 & n4710 ;
  assign n4713 = n4712 ^ n4711 ^ 1'b0 ;
  assign n4714 = n4205 ^ n2332 ^ 1'b0 ;
  assign n4715 = n3149 & ~n4714 ;
  assign n4716 = ~n2527 & n4715 ;
  assign n4717 = ~n4527 & n4716 ;
  assign n4718 = n4717 ^ n3313 ^ n3150 ;
  assign n4724 = n1340 ^ n1200 ^ n673 ;
  assign n4722 = n2087 ^ n1437 ^ 1'b0 ;
  assign n4719 = n1407 & n3363 ;
  assign n4720 = n4719 ^ n1827 ^ 1'b0 ;
  assign n4721 = ~n1293 & n4720 ;
  assign n4723 = n4722 ^ n4721 ^ x245 ;
  assign n4725 = n4724 ^ n4723 ^ 1'b0 ;
  assign n4726 = n3528 ^ x46 ^ 1'b0 ;
  assign n4727 = n929 | n932 ;
  assign n4728 = n4727 ^ n4417 ^ 1'b0 ;
  assign n4729 = n4728 ^ n1724 ^ n762 ;
  assign n4730 = ( ~n644 & n4726 ) | ( ~n644 & n4729 ) | ( n4726 & n4729 ) ;
  assign n4734 = ( n981 & ~n1544 ) | ( n981 & n1652 ) | ( ~n1544 & n1652 ) ;
  assign n4735 = n4734 ^ n1541 ^ n324 ;
  assign n4736 = ( ~n1641 & n3102 ) | ( ~n1641 & n4735 ) | ( n3102 & n4735 ) ;
  assign n4731 = n3722 ^ n3319 ^ n482 ;
  assign n4732 = n4731 ^ n3209 ^ 1'b0 ;
  assign n4733 = ( ~n2328 & n4150 ) | ( ~n2328 & n4732 ) | ( n4150 & n4732 ) ;
  assign n4737 = n4736 ^ n4733 ^ 1'b0 ;
  assign n4738 = n3717 & ~n4737 ;
  assign n4744 = n3296 ^ n2707 ^ n1261 ;
  assign n4741 = ( n1907 & n1977 ) | ( n1907 & ~n3529 ) | ( n1977 & ~n3529 ) ;
  assign n4739 = n1340 ^ n993 ^ 1'b0 ;
  assign n4740 = n2952 & ~n4739 ;
  assign n4742 = n4741 ^ n4740 ^ 1'b0 ;
  assign n4743 = n3633 & n4742 ;
  assign n4745 = n4744 ^ n4743 ^ 1'b0 ;
  assign n4746 = n3084 ^ n2235 ^ n711 ;
  assign n4747 = ( n2295 & ~n4288 ) | ( n2295 & n4746 ) | ( ~n4288 & n4746 ) ;
  assign n4748 = n2209 ^ x226 ^ x109 ;
  assign n4749 = n4748 ^ n2767 ^ 1'b0 ;
  assign n4750 = ( n4745 & ~n4747 ) | ( n4745 & n4749 ) | ( ~n4747 & n4749 ) ;
  assign n4751 = n4015 | n4750 ;
  assign n4753 = n2009 ^ n430 ^ 1'b0 ;
  assign n4754 = n582 & n4753 ;
  assign n4752 = n4186 ^ n3455 ^ n2651 ;
  assign n4755 = n4754 ^ n4752 ^ n4293 ;
  assign n4761 = ( x122 & ~n687 ) | ( x122 & n3770 ) | ( ~n687 & n3770 ) ;
  assign n4756 = n1475 ^ n1338 ^ 1'b0 ;
  assign n4757 = x69 & ~n4756 ;
  assign n4758 = n4757 ^ n2646 ^ n1690 ;
  assign n4759 = n4758 ^ n3937 ^ 1'b0 ;
  assign n4760 = ~n604 & n4759 ;
  assign n4762 = n4761 ^ n4760 ^ x25 ;
  assign n4764 = n1517 ^ n1111 ^ x161 ;
  assign n4763 = ~n293 & n4054 ;
  assign n4765 = n4764 ^ n4763 ^ 1'b0 ;
  assign n4766 = x235 & ~n1272 ;
  assign n4767 = n4766 ^ n2684 ^ 1'b0 ;
  assign n4768 = n2560 ^ n788 ^ 1'b0 ;
  assign n4769 = ( n666 & n673 ) | ( n666 & ~n4574 ) | ( n673 & ~n4574 ) ;
  assign n4770 = n2372 | n3444 ;
  assign n4771 = n4770 ^ n3494 ^ 1'b0 ;
  assign n4772 = ( n394 & n1305 ) | ( n394 & n4188 ) | ( n1305 & n4188 ) ;
  assign n4774 = n3596 | n4549 ;
  assign n4773 = ( ~n668 & n870 ) | ( ~n668 & n3099 ) | ( n870 & n3099 ) ;
  assign n4775 = n4774 ^ n4773 ^ 1'b0 ;
  assign n4776 = n856 & n4775 ;
  assign n4777 = n4776 ^ n2528 ^ x24 ;
  assign n4778 = ~n4772 & n4777 ;
  assign n4779 = n4771 & n4778 ;
  assign n4780 = ( n1642 & ~n3340 ) | ( n1642 & n4015 ) | ( ~n3340 & n4015 ) ;
  assign n4781 = ~n956 & n1799 ;
  assign n4782 = ( n430 & n523 ) | ( n430 & n4781 ) | ( n523 & n4781 ) ;
  assign n4783 = n4780 & n4782 ;
  assign n4784 = ~x124 & n4783 ;
  assign n4785 = ~n3731 & n3793 ;
  assign n4786 = ( ~n1201 & n2608 ) | ( ~n1201 & n3835 ) | ( n2608 & n3835 ) ;
  assign n4787 = n2732 ^ n1957 ^ n993 ;
  assign n4788 = n4787 ^ n4221 ^ n2022 ;
  assign n4789 = n3005 | n4788 ;
  assign n4790 = n4667 | n4789 ;
  assign n4791 = n4510 ^ n2652 ^ 1'b0 ;
  assign n4792 = n2960 ^ n582 ^ 1'b0 ;
  assign n4793 = ( n2875 & n4791 ) | ( n2875 & ~n4792 ) | ( n4791 & ~n4792 ) ;
  assign n4799 = n3065 ^ n2113 ^ 1'b0 ;
  assign n4800 = n1236 & n4799 ;
  assign n4794 = ~n339 & n1688 ;
  assign n4795 = n4794 ^ n1634 ^ n704 ;
  assign n4796 = ( x160 & n2793 ) | ( x160 & n4795 ) | ( n2793 & n4795 ) ;
  assign n4797 = ~n1746 & n4796 ;
  assign n4798 = n632 & n4797 ;
  assign n4801 = n4800 ^ n4798 ^ 1'b0 ;
  assign n4803 = n2988 & n3986 ;
  assign n4802 = n610 | n1264 ;
  assign n4804 = n4803 ^ n4802 ^ n4175 ;
  assign n4805 = n1003 & n2793 ;
  assign n4806 = n279 & n760 ;
  assign n4807 = n621 & n4806 ;
  assign n4808 = ( ~n681 & n1682 ) | ( ~n681 & n4807 ) | ( n1682 & n4807 ) ;
  assign n4809 = n4808 ^ n1143 ^ 1'b0 ;
  assign n4810 = ~n587 & n4809 ;
  assign n4811 = n4810 ^ n2180 ^ x87 ;
  assign n4816 = n1510 ^ n545 ^ 1'b0 ;
  assign n4817 = n698 & ~n4816 ;
  assign n4814 = n2134 ^ n2022 ^ 1'b0 ;
  assign n4815 = n494 | n4814 ;
  assign n4818 = n4817 ^ n4815 ^ n1278 ;
  assign n4812 = n971 | n4687 ;
  assign n4813 = ~n1183 & n4812 ;
  assign n4819 = n4818 ^ n4813 ^ 1'b0 ;
  assign n4820 = n1816 ^ n908 ^ n652 ;
  assign n4821 = n1668 & ~n4820 ;
  assign n4822 = n4821 ^ n1133 ^ 1'b0 ;
  assign n4823 = n4822 ^ n3722 ^ n1991 ;
  assign n4824 = n4070 | n4823 ;
  assign n4825 = n3752 ^ n2315 ^ x8 ;
  assign n4826 = n4825 ^ n3266 ^ n449 ;
  assign n4827 = n4184 | n4826 ;
  assign n4834 = ( n415 & n498 ) | ( n415 & ~n3240 ) | ( n498 & ~n3240 ) ;
  assign n4835 = ( n963 & ~n1235 ) | ( n963 & n2646 ) | ( ~n1235 & n2646 ) ;
  assign n4836 = ( ~n4363 & n4834 ) | ( ~n4363 & n4835 ) | ( n4834 & n4835 ) ;
  assign n4828 = n3752 ^ n2544 ^ 1'b0 ;
  assign n4829 = ~n1899 & n4828 ;
  assign n4830 = n4829 ^ n934 ^ 1'b0 ;
  assign n4831 = n4830 ^ n1452 ^ n1152 ;
  assign n4832 = n3567 ^ n3366 ^ n1883 ;
  assign n4833 = n4831 & ~n4832 ;
  assign n4837 = n4836 ^ n4833 ^ 1'b0 ;
  assign n4847 = n1329 ^ n771 ^ 1'b0 ;
  assign n4848 = n889 & ~n4847 ;
  assign n4845 = ~n1269 & n3212 ;
  assign n4846 = n3198 & n4845 ;
  assign n4849 = n4848 ^ n4846 ^ n735 ;
  assign n4841 = n4221 ^ n3977 ^ x214 ;
  assign n4842 = ( n890 & n2631 ) | ( n890 & n4841 ) | ( n2631 & n4841 ) ;
  assign n4840 = n4094 ^ n3397 ^ n1733 ;
  assign n4843 = n4842 ^ n4840 ^ 1'b0 ;
  assign n4844 = n4248 & ~n4843 ;
  assign n4850 = n4849 ^ n4844 ^ n3009 ;
  assign n4838 = x88 & n3952 ;
  assign n4839 = n4553 & n4838 ;
  assign n4851 = n4850 ^ n4839 ^ 1'b0 ;
  assign n4852 = ( n1055 & ~n1412 ) | ( n1055 & n1778 ) | ( ~n1412 & n1778 ) ;
  assign n4853 = n4852 ^ n1459 ^ n910 ;
  assign n4854 = n3024 | n4853 ;
  assign n4855 = n500 | n4854 ;
  assign n4856 = ( n699 & n1641 ) | ( n699 & n4855 ) | ( n1641 & n4855 ) ;
  assign n4857 = n1675 | n3309 ;
  assign n4858 = n2309 & ~n4857 ;
  assign n4859 = ( n1048 & n4856 ) | ( n1048 & n4858 ) | ( n4856 & n4858 ) ;
  assign n4860 = ( n1817 & n3757 ) | ( n1817 & n4859 ) | ( n3757 & n4859 ) ;
  assign n4861 = ~n858 & n1701 ;
  assign n4862 = n4861 ^ n2781 ^ 1'b0 ;
  assign n4863 = ( n3341 & n4466 ) | ( n3341 & n4862 ) | ( n4466 & n4862 ) ;
  assign n4864 = n927 ^ x147 ^ 1'b0 ;
  assign n4865 = ~n667 & n4864 ;
  assign n4866 = ( n463 & n2174 ) | ( n463 & n4865 ) | ( n2174 & n4865 ) ;
  assign n4867 = n2358 & n4601 ;
  assign n4868 = ~n4866 & n4867 ;
  assign n4869 = n4868 ^ n4713 ^ 1'b0 ;
  assign n4870 = n3325 ^ n657 ^ 1'b0 ;
  assign n4871 = n3490 ^ n1355 ^ 1'b0 ;
  assign n4872 = n4870 & ~n4871 ;
  assign n4876 = ( x123 & n1290 ) | ( x123 & ~n1611 ) | ( n1290 & ~n1611 ) ;
  assign n4877 = ( ~n471 & n2832 ) | ( ~n471 & n4876 ) | ( n2832 & n4876 ) ;
  assign n4878 = ( n1237 & ~n3766 ) | ( n1237 & n4877 ) | ( ~n3766 & n4877 ) ;
  assign n4874 = n1444 ^ n1351 ^ 1'b0 ;
  assign n4873 = n2557 ^ n2019 ^ n1589 ;
  assign n4875 = n4874 ^ n4873 ^ n2660 ;
  assign n4879 = n4878 ^ n4875 ^ n3534 ;
  assign n4882 = x173 & x174 ;
  assign n4883 = n4882 ^ n499 ^ 1'b0 ;
  assign n4880 = n4205 ^ n2071 ^ n1085 ;
  assign n4881 = n4880 ^ n485 ^ x143 ;
  assign n4884 = n4883 ^ n4881 ^ n4224 ;
  assign n4885 = ( n677 & ~n711 ) | ( n677 & n3933 ) | ( ~n711 & n3933 ) ;
  assign n4886 = n4885 ^ n1728 ^ n1392 ;
  assign n4887 = n2005 | n4886 ;
  assign n4888 = n508 | n4887 ;
  assign n4889 = n3406 ^ n2058 ^ n959 ;
  assign n4890 = n2465 ^ n1293 ^ n329 ;
  assign n4891 = n3286 ^ n2183 ^ x11 ;
  assign n4892 = ~n4890 & n4891 ;
  assign n4893 = n4889 & n4892 ;
  assign n4896 = n4444 ^ n2923 ^ n1037 ;
  assign n4894 = ( x213 & n1287 ) | ( x213 & ~n2489 ) | ( n1287 & ~n2489 ) ;
  assign n4895 = n4894 ^ n3264 ^ 1'b0 ;
  assign n4897 = n4896 ^ n4895 ^ n2857 ;
  assign n4900 = n378 & ~n827 ;
  assign n4901 = n4900 ^ n3977 ^ 1'b0 ;
  assign n4902 = n1860 | n4901 ;
  assign n4898 = n868 & n2867 ;
  assign n4899 = ~n1836 & n4898 ;
  assign n4903 = n4902 ^ n4899 ^ x61 ;
  assign n4904 = n3828 ^ n3049 ^ n1697 ;
  assign n4905 = n1211 & n4904 ;
  assign n4906 = n3691 ^ n643 ^ n620 ;
  assign n4907 = n4344 & ~n4906 ;
  assign n4908 = n4905 & n4907 ;
  assign n4909 = n2775 ^ n592 ^ n450 ;
  assign n4911 = n1950 | n2288 ;
  assign n4912 = n3251 & ~n4911 ;
  assign n4913 = n3249 & n4912 ;
  assign n4910 = n2521 ^ n2373 ^ 1'b0 ;
  assign n4914 = n4913 ^ n4910 ^ 1'b0 ;
  assign n4915 = n4909 | n4914 ;
  assign n4916 = n4419 ^ n2453 ^ 1'b0 ;
  assign n4917 = ( n455 & ~n4463 ) | ( n455 & n4916 ) | ( ~n4463 & n4916 ) ;
  assign n4918 = ~n1657 & n2966 ;
  assign n4919 = n4918 ^ n487 ^ 1'b0 ;
  assign n4920 = n4919 ^ n2154 ^ 1'b0 ;
  assign n4921 = ~n2932 & n4920 ;
  assign n4922 = ( n1406 & n4438 ) | ( n1406 & n4921 ) | ( n4438 & n4921 ) ;
  assign n4923 = ( n427 & ~n2939 ) | ( n427 & n4922 ) | ( ~n2939 & n4922 ) ;
  assign n4924 = n2835 ^ n1754 ^ n1339 ;
  assign n4925 = ( n944 & n961 ) | ( n944 & ~n4164 ) | ( n961 & ~n4164 ) ;
  assign n4926 = n351 & ~n1784 ;
  assign n4927 = n4925 | n4926 ;
  assign n4928 = n2762 & ~n4927 ;
  assign n4929 = n1028 & ~n4928 ;
  assign n4930 = ~n4924 & n4929 ;
  assign n4931 = n3676 ^ x133 ^ 1'b0 ;
  assign n4932 = x251 & ~n731 ;
  assign n4933 = n4932 ^ n2038 ^ 1'b0 ;
  assign n4934 = ( n553 & n1247 ) | ( n553 & n3995 ) | ( n1247 & n3995 ) ;
  assign n4935 = ( n4931 & ~n4933 ) | ( n4931 & n4934 ) | ( ~n4933 & n4934 ) ;
  assign n4936 = x171 ^ x144 ^ 1'b0 ;
  assign n4937 = x201 & n4936 ;
  assign n4938 = n1192 & n3716 ;
  assign n4939 = ~n4937 & n4938 ;
  assign n4940 = ( n379 & n812 ) | ( n379 & n1351 ) | ( n812 & n1351 ) ;
  assign n4941 = ~n1033 & n4940 ;
  assign n4942 = ~x190 & n4941 ;
  assign n4943 = n1901 | n4641 ;
  assign n4944 = n1198 | n4943 ;
  assign n4945 = n4576 ^ x19 ^ 1'b0 ;
  assign n4946 = ( n1968 & n4944 ) | ( n1968 & n4945 ) | ( n4944 & n4945 ) ;
  assign n4947 = n4946 ^ n1122 ^ x166 ;
  assign n4951 = ( n399 & ~n1605 ) | ( n399 & n3905 ) | ( ~n1605 & n3905 ) ;
  assign n4948 = n2691 ^ n644 ^ 1'b0 ;
  assign n4949 = n1377 & ~n4948 ;
  assign n4950 = ( n1152 & ~n2931 ) | ( n1152 & n4949 ) | ( ~n2931 & n4949 ) ;
  assign n4952 = n4951 ^ n4950 ^ n547 ;
  assign n4953 = n3271 ^ n2747 ^ 1'b0 ;
  assign n4954 = n711 & ~n4953 ;
  assign n4955 = ~n500 & n4954 ;
  assign n4956 = n4952 & n4955 ;
  assign n4957 = n4947 & n4956 ;
  assign n4958 = n2763 | n4957 ;
  assign n4959 = n4958 ^ n1035 ^ 1'b0 ;
  assign n4961 = n1423 ^ n1381 ^ 1'b0 ;
  assign n4962 = x159 & ~n4961 ;
  assign n4963 = n4962 ^ n2394 ^ n1352 ;
  assign n4964 = n4963 ^ n1449 ^ 1'b0 ;
  assign n4965 = n4954 & ~n4964 ;
  assign n4960 = n4175 ^ n2272 ^ n1791 ;
  assign n4966 = n4965 ^ n4960 ^ 1'b0 ;
  assign n4967 = ~n2594 & n4966 ;
  assign n4969 = n2296 ^ n481 ^ n433 ;
  assign n4970 = ( n2178 & n2472 ) | ( n2178 & ~n4969 ) | ( n2472 & ~n4969 ) ;
  assign n4971 = ( n1085 & n4081 ) | ( n1085 & n4970 ) | ( n4081 & n4970 ) ;
  assign n4972 = n4971 ^ n2654 ^ n2477 ;
  assign n4968 = n1869 & n3143 ;
  assign n4973 = n4972 ^ n4968 ^ 1'b0 ;
  assign n4974 = n865 ^ n833 ^ n371 ;
  assign n4975 = x149 & x237 ;
  assign n4976 = n361 & n4975 ;
  assign n4977 = n829 | n4976 ;
  assign n4978 = n1385 | n4977 ;
  assign n4979 = x238 & n4978 ;
  assign n4980 = ~n429 & n4979 ;
  assign n4981 = n4974 | n4980 ;
  assign n4982 = n4981 ^ n4449 ^ 1'b0 ;
  assign n4983 = ( n347 & n604 ) | ( n347 & n1373 ) | ( n604 & n1373 ) ;
  assign n4984 = n3851 & n4983 ;
  assign n4985 = ( n3519 & n4112 ) | ( n3519 & ~n4984 ) | ( n4112 & ~n4984 ) ;
  assign n4986 = ( n1091 & ~n4429 ) | ( n1091 & n4985 ) | ( ~n4429 & n4985 ) ;
  assign n4987 = ( n1156 & n1808 ) | ( n1156 & ~n2428 ) | ( n1808 & ~n2428 ) ;
  assign n4988 = ( x204 & n3947 ) | ( x204 & ~n4223 ) | ( n3947 & ~n4223 ) ;
  assign n4989 = ~n4987 & n4988 ;
  assign n4990 = n2949 & n4989 ;
  assign n4991 = ( n385 & n3635 ) | ( n385 & n4952 ) | ( n3635 & n4952 ) ;
  assign n4992 = n2777 ^ n2135 ^ n918 ;
  assign n4993 = n1570 ^ n880 ^ 1'b0 ;
  assign n4994 = ( n2169 & ~n4102 ) | ( n2169 & n4993 ) | ( ~n4102 & n4993 ) ;
  assign n4995 = ( n1233 & ~n4992 ) | ( n1233 & n4994 ) | ( ~n4992 & n4994 ) ;
  assign n4996 = n3522 ^ n453 ^ 1'b0 ;
  assign n4997 = n1799 | n4996 ;
  assign n4998 = ( ~n2115 & n2615 ) | ( ~n2115 & n3601 ) | ( n2615 & n3601 ) ;
  assign n4999 = ( n434 & ~n760 ) | ( n434 & n4967 ) | ( ~n760 & n4967 ) ;
  assign n5000 = ( n745 & n891 ) | ( n745 & ~n1336 ) | ( n891 & ~n1336 ) ;
  assign n5001 = n3942 & n5000 ;
  assign n5002 = n520 & n5001 ;
  assign n5003 = n5002 ^ n4120 ^ n2382 ;
  assign n5004 = n4015 ^ n939 ^ x209 ;
  assign n5006 = n4165 ^ n1637 ^ x250 ;
  assign n5007 = n1014 & ~n5006 ;
  assign n5008 = n993 & n5007 ;
  assign n5005 = ( n351 & n2782 ) | ( n351 & n4180 ) | ( n2782 & n4180 ) ;
  assign n5009 = n5008 ^ n5005 ^ n3164 ;
  assign n5010 = ( x240 & ~n2741 ) | ( x240 & n5009 ) | ( ~n2741 & n5009 ) ;
  assign n5011 = n1836 & n4008 ;
  assign n5012 = n3132 & n4838 ;
  assign n5013 = n5011 & n5012 ;
  assign n5019 = ( n409 & n1913 ) | ( n409 & n2183 ) | ( n1913 & n2183 ) ;
  assign n5015 = ~n1355 & n4189 ;
  assign n5016 = ( ~n999 & n2952 ) | ( ~n999 & n5015 ) | ( n2952 & n5015 ) ;
  assign n5014 = n4054 ^ n2101 ^ n1367 ;
  assign n5017 = n5016 ^ n5014 ^ n2804 ;
  assign n5018 = n5017 ^ n3083 ^ n2549 ;
  assign n5020 = n5019 ^ n5018 ^ n2441 ;
  assign n5022 = ( x90 & n310 ) | ( x90 & ~n630 ) | ( n310 & ~n630 ) ;
  assign n5023 = ( n890 & n1391 ) | ( n890 & ~n5022 ) | ( n1391 & ~n5022 ) ;
  assign n5021 = n570 | n2257 ;
  assign n5024 = n5023 ^ n5021 ^ n1467 ;
  assign n5025 = ~n545 & n3138 ;
  assign n5026 = n5025 ^ n336 ^ 1'b0 ;
  assign n5027 = n5026 ^ n1968 ^ 1'b0 ;
  assign n5028 = n4386 ^ n3956 ^ 1'b0 ;
  assign n5029 = ~n4048 & n5028 ;
  assign n5030 = n5029 ^ n4832 ^ 1'b0 ;
  assign n5031 = n2605 ^ n357 ^ 1'b0 ;
  assign n5032 = n961 | n5031 ;
  assign n5033 = n5032 ^ n4301 ^ n361 ;
  assign n5034 = n5033 ^ n4852 ^ 1'b0 ;
  assign n5035 = ( x28 & n1365 ) | ( x28 & n1732 ) | ( n1365 & n1732 ) ;
  assign n5036 = n5035 ^ n1032 ^ 1'b0 ;
  assign n5037 = n1134 | n5036 ;
  assign n5038 = n1653 ^ n763 ^ n570 ;
  assign n5039 = n4186 & ~n5038 ;
  assign n5041 = n796 ^ x136 ^ 1'b0 ;
  assign n5042 = n572 & ~n5041 ;
  assign n5040 = x186 | n3706 ;
  assign n5043 = n5042 ^ n5040 ^ 1'b0 ;
  assign n5044 = n3923 ^ n3667 ^ 1'b0 ;
  assign n5045 = ( n595 & n2530 ) | ( n595 & ~n4421 ) | ( n2530 & ~n4421 ) ;
  assign n5046 = n3113 ^ n1268 ^ 1'b0 ;
  assign n5047 = ( n4404 & n5045 ) | ( n4404 & n5046 ) | ( n5045 & n5046 ) ;
  assign n5048 = n5047 ^ n4396 ^ 1'b0 ;
  assign n5049 = n5023 ^ n3444 ^ n421 ;
  assign n5050 = ( ~n2055 & n4123 ) | ( ~n2055 & n4730 ) | ( n4123 & n4730 ) ;
  assign n5051 = n4685 ^ n2678 ^ n886 ;
  assign n5052 = ( n2350 & ~n3530 ) | ( n2350 & n5051 ) | ( ~n3530 & n5051 ) ;
  assign n5053 = n5052 ^ n3793 ^ 1'b0 ;
  assign n5054 = ( n550 & n771 ) | ( n550 & ~n4291 ) | ( n771 & ~n4291 ) ;
  assign n5055 = ( ~n834 & n2496 ) | ( ~n834 & n5054 ) | ( n2496 & n5054 ) ;
  assign n5059 = n2178 & ~n3276 ;
  assign n5060 = ~n1821 & n5059 ;
  assign n5061 = n4311 & ~n5060 ;
  assign n5062 = ~n3088 & n5061 ;
  assign n5056 = n2745 ^ x208 ^ x125 ;
  assign n5057 = n3727 & ~n5056 ;
  assign n5058 = n5057 ^ n593 ^ 1'b0 ;
  assign n5063 = n5062 ^ n5058 ^ 1'b0 ;
  assign n5064 = ~n5055 & n5063 ;
  assign n5065 = n793 & ~n1645 ;
  assign n5066 = ( n1906 & ~n1963 ) | ( n1906 & n5065 ) | ( ~n1963 & n5065 ) ;
  assign n5067 = n3192 ^ n1023 ^ x190 ;
  assign n5068 = n1305 | n2066 ;
  assign n5069 = n5068 ^ n574 ^ 1'b0 ;
  assign n5070 = ~n5067 & n5069 ;
  assign n5071 = n5070 ^ n4653 ^ 1'b0 ;
  assign n5073 = n2072 & ~n3018 ;
  assign n5074 = ~n3575 & n5073 ;
  assign n5072 = ( n423 & ~n1457 ) | ( n423 & n4498 ) | ( ~n1457 & n4498 ) ;
  assign n5075 = n5074 ^ n5072 ^ n2177 ;
  assign n5076 = n3300 ^ n1201 ^ n557 ;
  assign n5077 = ( ~n4261 & n4734 ) | ( ~n4261 & n5076 ) | ( n4734 & n5076 ) ;
  assign n5078 = n5077 ^ n2703 ^ n2241 ;
  assign n5080 = n4944 ^ n4126 ^ n1202 ;
  assign n5081 = ~n2066 & n5080 ;
  assign n5082 = n5081 ^ n359 ^ 1'b0 ;
  assign n5079 = ( n378 & ~n3769 ) | ( n378 & n4550 ) | ( ~n3769 & n4550 ) ;
  assign n5083 = n5082 ^ n5079 ^ n1142 ;
  assign n5086 = ( n699 & n845 ) | ( n699 & ~n2689 ) | ( n845 & ~n2689 ) ;
  assign n5084 = ~n3584 & n4567 ;
  assign n5085 = n5084 ^ n3218 ^ 1'b0 ;
  assign n5087 = n5086 ^ n5085 ^ 1'b0 ;
  assign n5088 = ( ~n4306 & n5083 ) | ( ~n4306 & n5087 ) | ( n5083 & n5087 ) ;
  assign n5089 = n2299 ^ n1939 ^ n1438 ;
  assign n5090 = n5089 ^ n1351 ^ n891 ;
  assign n5091 = n3770 & ~n5090 ;
  assign n5092 = n961 & n5091 ;
  assign n5095 = n1544 ^ n1365 ^ n795 ;
  assign n5096 = ( n548 & n2301 ) | ( n548 & ~n5095 ) | ( n2301 & ~n5095 ) ;
  assign n5093 = n4086 ^ n1823 ^ n1745 ;
  assign n5094 = n1455 & ~n5093 ;
  assign n5097 = n5096 ^ n5094 ^ 1'b0 ;
  assign n5098 = n5097 ^ n4503 ^ n1554 ;
  assign n5099 = n1133 & ~n4667 ;
  assign n5100 = n2016 & n5099 ;
  assign n5103 = n4460 ^ n2234 ^ n1550 ;
  assign n5101 = ~n2217 & n3086 ;
  assign n5102 = n5101 ^ n328 ^ 1'b0 ;
  assign n5104 = n5103 ^ n5102 ^ x196 ;
  assign n5105 = x227 & ~n594 ;
  assign n5106 = n5105 ^ n1988 ^ 1'b0 ;
  assign n5107 = n3039 | n5106 ;
  assign n5108 = ~n673 & n2899 ;
  assign n5109 = n5108 ^ n2771 ^ n1920 ;
  assign n5110 = ( x156 & n1352 ) | ( x156 & n1386 ) | ( n1352 & n1386 ) ;
  assign n5111 = ( ~n340 & n669 ) | ( ~n340 & n5110 ) | ( n669 & n5110 ) ;
  assign n5112 = n5111 ^ n2950 ^ n2664 ;
  assign n5113 = n2529 ^ n1327 ^ 1'b0 ;
  assign n5114 = ~x227 & n925 ;
  assign n5115 = ~n1159 & n5114 ;
  assign n5116 = n5115 ^ n4526 ^ 1'b0 ;
  assign n5117 = n5113 & ~n5116 ;
  assign n5118 = ( x195 & n3898 ) | ( x195 & n3977 ) | ( n3898 & n3977 ) ;
  assign n5119 = n5118 ^ n355 ^ x236 ;
  assign n5120 = n1691 & n2425 ;
  assign n5121 = ~n5119 & n5120 ;
  assign n5122 = n5121 ^ n4171 ^ n849 ;
  assign n5123 = n5117 & ~n5122 ;
  assign n5124 = n3253 ^ n1339 ^ 1'b0 ;
  assign n5125 = n3508 & ~n5124 ;
  assign n5126 = n5125 ^ n1068 ^ 1'b0 ;
  assign n5133 = n3253 ^ n365 ^ n334 ;
  assign n5128 = x250 & ~n1066 ;
  assign n5129 = n5128 ^ n3444 ^ 1'b0 ;
  assign n5130 = n5129 ^ n1739 ^ n284 ;
  assign n5131 = ( x244 & ~n1291 ) | ( x244 & n5130 ) | ( ~n1291 & n5130 ) ;
  assign n5127 = n1265 & ~n3615 ;
  assign n5132 = n5131 ^ n5127 ^ 1'b0 ;
  assign n5134 = n5133 ^ n5132 ^ n3107 ;
  assign n5135 = n639 ^ n585 ^ 1'b0 ;
  assign n5136 = n5135 ^ n2979 ^ 1'b0 ;
  assign n5137 = n3708 | n5136 ;
  assign n5146 = n1361 ^ n561 ^ x241 ;
  assign n5147 = n4820 ^ n1302 ^ n508 ;
  assign n5148 = n5147 ^ n1321 ^ 1'b0 ;
  assign n5149 = n1236 & n5148 ;
  assign n5150 = n5146 & n5149 ;
  assign n5151 = ~n3842 & n5150 ;
  assign n5152 = ( ~n2380 & n4046 ) | ( ~n2380 & n5151 ) | ( n4046 & n5151 ) ;
  assign n5138 = ( n1238 & n1945 ) | ( n1238 & n4974 ) | ( n1945 & n4974 ) ;
  assign n5139 = ( n802 & n4006 ) | ( n802 & n4279 ) | ( n4006 & n4279 ) ;
  assign n5140 = x24 & ~n1806 ;
  assign n5141 = n5140 ^ n393 ^ 1'b0 ;
  assign n5142 = n5141 ^ n1638 ^ 1'b0 ;
  assign n5143 = ( n1626 & n4049 ) | ( n1626 & ~n5142 ) | ( n4049 & ~n5142 ) ;
  assign n5144 = n2670 & n5143 ;
  assign n5145 = ( n5138 & ~n5139 ) | ( n5138 & n5144 ) | ( ~n5139 & n5144 ) ;
  assign n5153 = n5152 ^ n5145 ^ 1'b0 ;
  assign n5154 = n989 | n1508 ;
  assign n5155 = ( x149 & n4282 ) | ( x149 & ~n5154 ) | ( n4282 & ~n5154 ) ;
  assign n5156 = n1784 ^ n1087 ^ 1'b0 ;
  assign n5157 = n2309 | n5156 ;
  assign n5158 = n2501 ^ x79 ^ 1'b0 ;
  assign n5161 = ~n1405 & n2173 ;
  assign n5162 = n5161 ^ n4084 ^ 1'b0 ;
  assign n5168 = x180 & n2494 ;
  assign n5169 = ~n890 & n5168 ;
  assign n5170 = n1827 & ~n5169 ;
  assign n5171 = n2566 & n5170 ;
  assign n5163 = n2762 ^ n1060 ^ 1'b0 ;
  assign n5164 = n2411 ^ n592 ^ 1'b0 ;
  assign n5165 = ( n992 & ~n5163 ) | ( n992 & n5164 ) | ( ~n5163 & n5164 ) ;
  assign n5166 = n4480 ^ n4176 ^ x125 ;
  assign n5167 = n5165 & ~n5166 ;
  assign n5172 = n5171 ^ n5167 ^ 1'b0 ;
  assign n5173 = n5172 ^ n3806 ^ 1'b0 ;
  assign n5174 = n5173 ^ n3545 ^ n2965 ;
  assign n5175 = ( ~n3407 & n5162 ) | ( ~n3407 & n5174 ) | ( n5162 & n5174 ) ;
  assign n5159 = n5042 ^ n2914 ^ n324 ;
  assign n5160 = ~n5037 & n5159 ;
  assign n5176 = n5175 ^ n5160 ^ 1'b0 ;
  assign n5177 = ( n2736 & ~n5158 ) | ( n2736 & n5176 ) | ( ~n5158 & n5176 ) ;
  assign n5178 = ( ~x72 & n494 ) | ( ~x72 & n509 ) | ( n494 & n509 ) ;
  assign n5179 = n5178 ^ n2990 ^ n1294 ;
  assign n5180 = n5179 ^ n3225 ^ 1'b0 ;
  assign n5181 = n2818 ^ n1668 ^ n522 ;
  assign n5182 = n5154 ^ n4100 ^ 1'b0 ;
  assign n5183 = n693 | n5182 ;
  assign n5184 = n5183 ^ n1605 ^ 1'b0 ;
  assign n5185 = n2966 | n3914 ;
  assign n5186 = ( ~n1887 & n5184 ) | ( ~n1887 & n5185 ) | ( n5184 & n5185 ) ;
  assign n5187 = n2003 ^ n1683 ^ 1'b0 ;
  assign n5189 = n1003 | n1920 ;
  assign n5188 = ~x145 & n3500 ;
  assign n5190 = n5189 ^ n5188 ^ n2833 ;
  assign n5198 = n353 & ~n1569 ;
  assign n5199 = ~n1170 & n5198 ;
  assign n5200 = n2083 | n5199 ;
  assign n5201 = n711 | n5200 ;
  assign n5191 = n1518 | n3664 ;
  assign n5192 = n5191 ^ n4139 ^ 1'b0 ;
  assign n5193 = n5192 ^ n1610 ^ x5 ;
  assign n5194 = n1693 ^ n637 ^ n412 ;
  assign n5195 = ( n2033 & n4381 ) | ( n2033 & n5194 ) | ( n4381 & n5194 ) ;
  assign n5196 = n4776 ^ n3365 ^ x225 ;
  assign n5197 = ( ~n5193 & n5195 ) | ( ~n5193 & n5196 ) | ( n5195 & n5196 ) ;
  assign n5202 = n5201 ^ n5197 ^ n1830 ;
  assign n5203 = n4011 ^ n3288 ^ n775 ;
  assign n5204 = ( ~x140 & n917 ) | ( ~x140 & n1758 ) | ( n917 & n1758 ) ;
  assign n5206 = ( ~x3 & n747 ) | ( ~x3 & n1828 ) | ( n747 & n1828 ) ;
  assign n5207 = n5206 ^ n4780 ^ n991 ;
  assign n5205 = ~n1950 & n2920 ;
  assign n5208 = n5207 ^ n5205 ^ 1'b0 ;
  assign n5209 = ( n2871 & ~n5204 ) | ( n2871 & n5208 ) | ( ~n5204 & n5208 ) ;
  assign n5210 = n1495 ^ n945 ^ 1'b0 ;
  assign n5211 = n5210 ^ n2310 ^ 1'b0 ;
  assign n5212 = ( n2415 & ~n3600 ) | ( n2415 & n5211 ) | ( ~n3600 & n5211 ) ;
  assign n5213 = ( n456 & n3748 ) | ( n456 & n5212 ) | ( n3748 & n5212 ) ;
  assign n5214 = n2440 ^ n2004 ^ 1'b0 ;
  assign n5215 = n5214 ^ n951 ^ 1'b0 ;
  assign n5216 = n5199 | n5215 ;
  assign n5217 = n1292 | n5047 ;
  assign n5218 = n5216 & ~n5217 ;
  assign n5223 = n1341 | n3134 ;
  assign n5224 = x98 | n5223 ;
  assign n5220 = ( x141 & n624 ) | ( x141 & n836 ) | ( n624 & n836 ) ;
  assign n5219 = n3041 | n3381 ;
  assign n5221 = n5220 ^ n5219 ^ n1600 ;
  assign n5222 = n5221 ^ n3556 ^ n1119 ;
  assign n5225 = n5224 ^ n5222 ^ 1'b0 ;
  assign n5226 = n2156 ^ n466 ^ 1'b0 ;
  assign n5227 = n3680 & n5226 ;
  assign n5228 = n931 & n1542 ;
  assign n5229 = n5228 ^ n2390 ^ 1'b0 ;
  assign n5230 = ~n2447 & n5229 ;
  assign n5231 = ( n4336 & n5227 ) | ( n4336 & ~n5230 ) | ( n5227 & ~n5230 ) ;
  assign n5232 = n3725 ^ n1899 ^ n1406 ;
  assign n5237 = n482 & n650 ;
  assign n5234 = ( n374 & n722 ) | ( n374 & ~n1702 ) | ( n722 & ~n1702 ) ;
  assign n5233 = ( x157 & ~n1560 ) | ( x157 & n3116 ) | ( ~n1560 & n3116 ) ;
  assign n5235 = n5234 ^ n5233 ^ n849 ;
  assign n5236 = ( n869 & ~n3444 ) | ( n869 & n5235 ) | ( ~n3444 & n5235 ) ;
  assign n5238 = n5237 ^ n5236 ^ n656 ;
  assign n5239 = n1200 & ~n1627 ;
  assign n5240 = n5239 ^ n693 ^ 1'b0 ;
  assign n5241 = n5240 ^ n2562 ^ n1490 ;
  assign n5242 = ( x184 & ~n2492 ) | ( x184 & n4909 ) | ( ~n2492 & n4909 ) ;
  assign n5243 = n5242 ^ n4282 ^ n3734 ;
  assign n5244 = n2130 & n5243 ;
  assign n5245 = n3296 & n5244 ;
  assign n5246 = ( n450 & ~n1382 ) | ( n450 & n3824 ) | ( ~n1382 & n3824 ) ;
  assign n5247 = ( n3335 & n4265 ) | ( n3335 & n5246 ) | ( n4265 & n5246 ) ;
  assign n5250 = ( n1173 & ~n2401 ) | ( n1173 & n2867 ) | ( ~n2401 & n2867 ) ;
  assign n5251 = ( ~n505 & n1448 ) | ( ~n505 & n5250 ) | ( n1448 & n5250 ) ;
  assign n5253 = n2455 ^ n931 ^ n733 ;
  assign n5252 = n2760 ^ n324 ^ 1'b0 ;
  assign n5254 = n5253 ^ n5252 ^ 1'b0 ;
  assign n5255 = ~n2205 & n5254 ;
  assign n5256 = ( ~n2042 & n5251 ) | ( ~n2042 & n5255 ) | ( n5251 & n5255 ) ;
  assign n5248 = n2643 ^ x200 ^ 1'b0 ;
  assign n5249 = n5248 ^ n3616 ^ n365 ;
  assign n5257 = n5256 ^ n5249 ^ n1911 ;
  assign n5258 = ( n1026 & n4257 ) | ( n1026 & n5257 ) | ( n4257 & n5257 ) ;
  assign n5259 = ( ~n544 & n1339 ) | ( ~n544 & n3316 ) | ( n1339 & n3316 ) ;
  assign n5260 = n3484 & n5259 ;
  assign n5263 = n1892 ^ x227 ^ 1'b0 ;
  assign n5264 = n2526 & n5263 ;
  assign n5261 = ( n1412 & ~n1832 ) | ( n1412 & n2749 ) | ( ~n1832 & n2749 ) ;
  assign n5262 = ( ~n3144 & n4445 ) | ( ~n3144 & n5261 ) | ( n4445 & n5261 ) ;
  assign n5265 = n5264 ^ n5262 ^ n1448 ;
  assign n5266 = n3198 ^ n852 ^ 1'b0 ;
  assign n5267 = n5265 | n5266 ;
  assign n5268 = n2934 | n5138 ;
  assign n5269 = n5268 ^ x125 ^ 1'b0 ;
  assign n5270 = n5118 ^ n3794 ^ n3383 ;
  assign n5271 = ( n563 & n3700 ) | ( n563 & ~n5270 ) | ( n3700 & ~n5270 ) ;
  assign n5272 = n5269 & ~n5271 ;
  assign n5273 = n5267 & n5272 ;
  assign n5274 = ( ~n1849 & n3060 ) | ( ~n1849 & n4074 ) | ( n3060 & n4074 ) ;
  assign n5275 = n381 & ~n3881 ;
  assign n5276 = n5275 ^ n4570 ^ n3027 ;
  assign n5277 = n2444 & n4291 ;
  assign n5278 = n3027 ^ n2027 ^ 1'b0 ;
  assign n5279 = n1665 | n5278 ;
  assign n5280 = n1096 & n2411 ;
  assign n5281 = n2220 & n5280 ;
  assign n5282 = n1363 & n5281 ;
  assign n5283 = n5253 ^ x221 ^ 1'b0 ;
  assign n5284 = n1845 & ~n5283 ;
  assign n5285 = n5284 ^ n5250 ^ n3549 ;
  assign n5286 = ( ~n5279 & n5282 ) | ( ~n5279 & n5285 ) | ( n5282 & n5285 ) ;
  assign n5287 = n2656 ^ n1991 ^ n1927 ;
  assign n5298 = n2035 ^ n1336 ^ 1'b0 ;
  assign n5299 = n727 | n3131 ;
  assign n5300 = n343 & ~n5299 ;
  assign n5301 = n3575 ^ n328 ^ 1'b0 ;
  assign n5302 = ~n325 & n5301 ;
  assign n5303 = n5302 ^ n2905 ^ n817 ;
  assign n5304 = ( n1380 & n5300 ) | ( n1380 & n5303 ) | ( n5300 & n5303 ) ;
  assign n5305 = n2272 ^ n1853 ^ 1'b0 ;
  assign n5306 = n1344 & n5305 ;
  assign n5307 = n5306 ^ x239 ^ 1'b0 ;
  assign n5308 = ( n5298 & n5304 ) | ( n5298 & n5307 ) | ( n5304 & n5307 ) ;
  assign n5296 = n4452 ^ n3963 ^ n2735 ;
  assign n5297 = n5296 ^ n2975 ^ n1465 ;
  assign n5293 = ( n749 & n1402 ) | ( n749 & n5219 ) | ( n1402 & n5219 ) ;
  assign n5291 = ( ~n1783 & n1968 ) | ( ~n1783 & n2528 ) | ( n1968 & n2528 ) ;
  assign n5292 = ( x196 & n3562 ) | ( x196 & ~n5291 ) | ( n3562 & ~n5291 ) ;
  assign n5294 = n5293 ^ n5292 ^ n875 ;
  assign n5290 = n4899 ^ n1487 ^ n1444 ;
  assign n5288 = n860 & n1261 ;
  assign n5289 = n5288 ^ n3619 ^ 1'b0 ;
  assign n5295 = n5294 ^ n5290 ^ n5289 ;
  assign n5309 = n5308 ^ n5297 ^ n5295 ;
  assign n5310 = n1793 ^ n1091 ^ n813 ;
  assign n5311 = n5310 ^ n3415 ^ n2767 ;
  assign n5312 = n5311 ^ n2594 ^ x215 ;
  assign n5313 = n5312 ^ n911 ^ 1'b0 ;
  assign n5314 = n3952 ^ n2325 ^ 1'b0 ;
  assign n5315 = n5313 & n5314 ;
  assign n5316 = n2755 & n3398 ;
  assign n5317 = n5204 ^ x22 ^ 1'b0 ;
  assign n5318 = ~n5316 & n5317 ;
  assign n5319 = n3868 & n5318 ;
  assign n5320 = n4064 ^ n1433 ^ x12 ;
  assign n5321 = n1056 & ~n2674 ;
  assign n5322 = n2896 & n5321 ;
  assign n5323 = n5322 ^ n3601 ^ n2255 ;
  assign n5324 = ( ~x1 & n473 ) | ( ~x1 & n1271 ) | ( n473 & n1271 ) ;
  assign n5325 = n4515 ^ n3836 ^ 1'b0 ;
  assign n5326 = n5324 & ~n5325 ;
  assign n5327 = n2914 & ~n4881 ;
  assign n5328 = ( ~x147 & n1230 ) | ( ~x147 & n1329 ) | ( n1230 & n1329 ) ;
  assign n5329 = ~n3855 & n5328 ;
  assign n5330 = ( n1619 & ~n3773 ) | ( n1619 & n5329 ) | ( ~n3773 & n5329 ) ;
  assign n5331 = n1665 & n2055 ;
  assign n5332 = n1926 ^ n797 ^ x159 ;
  assign n5333 = x93 & ~n5332 ;
  assign n5334 = n5331 & n5333 ;
  assign n5335 = n2913 ^ n2123 ^ n973 ;
  assign n5336 = ( ~x12 & n410 ) | ( ~x12 & n1716 ) | ( n410 & n1716 ) ;
  assign n5337 = n5336 ^ n4410 ^ 1'b0 ;
  assign n5338 = n2990 & ~n5337 ;
  assign n5339 = n1447 ^ n1398 ^ 1'b0 ;
  assign n5340 = n5338 | n5339 ;
  assign n5341 = ( n899 & n1356 ) | ( n899 & n5340 ) | ( n1356 & n5340 ) ;
  assign n5342 = n2961 & n5341 ;
  assign n5343 = n3594 & n5342 ;
  assign n5344 = ( n995 & n1659 ) | ( n995 & n2058 ) | ( n1659 & n2058 ) ;
  assign n5345 = n1285 ^ n1273 ^ 1'b0 ;
  assign n5346 = n5344 & n5345 ;
  assign n5347 = ~n4841 & n5346 ;
  assign n5348 = n5347 ^ n5115 ^ n3725 ;
  assign n5349 = ( n5335 & ~n5343 ) | ( n5335 & n5348 ) | ( ~n5343 & n5348 ) ;
  assign n5350 = n3119 ^ n2756 ^ n2736 ;
  assign n5351 = ( x108 & ~n1438 ) | ( x108 & n4757 ) | ( ~n1438 & n4757 ) ;
  assign n5352 = n1727 | n3245 ;
  assign n5353 = n5352 ^ n1225 ^ x75 ;
  assign n5354 = n2122 & n5353 ;
  assign n5355 = ( ~n1484 & n2193 ) | ( ~n1484 & n5354 ) | ( n2193 & n5354 ) ;
  assign n5356 = x82 & n5355 ;
  assign n5357 = ~n5351 & n5356 ;
  assign n5358 = ( n1269 & n3150 ) | ( n1269 & ~n3211 ) | ( n3150 & ~n3211 ) ;
  assign n5359 = ( n2956 & ~n3653 ) | ( n2956 & n5358 ) | ( ~n3653 & n5358 ) ;
  assign n5360 = n5022 ^ n4744 ^ n4445 ;
  assign n5361 = n3885 & ~n5360 ;
  assign n5362 = n5359 & n5361 ;
  assign n5363 = ( n600 & n1870 ) | ( n600 & ~n2135 ) | ( n1870 & ~n2135 ) ;
  assign n5364 = ( n690 & n4029 ) | ( n690 & ~n5363 ) | ( n4029 & ~n5363 ) ;
  assign n5365 = n4863 ^ n1108 ^ 1'b0 ;
  assign n5366 = n5364 & ~n5365 ;
  assign n5367 = n1247 ^ x228 ^ x121 ;
  assign n5368 = n5367 ^ n4633 ^ n2549 ;
  assign n5369 = ~n5219 & n5240 ;
  assign n5370 = n5369 ^ n1305 ^ 1'b0 ;
  assign n5371 = n5368 & ~n5370 ;
  assign n5372 = n3748 ^ n3073 ^ n1928 ;
  assign n5373 = n5372 ^ n3917 ^ x248 ;
  assign n5374 = ~x236 & n5373 ;
  assign n5375 = ~n1423 & n3415 ;
  assign n5376 = n5375 ^ n1957 ^ 1'b0 ;
  assign n5383 = n1766 ^ n1210 ^ x174 ;
  assign n5382 = ( x25 & n516 ) | ( x25 & ~n3899 ) | ( n516 & ~n3899 ) ;
  assign n5384 = n5383 ^ n5382 ^ n4886 ;
  assign n5378 = n3432 ^ n3280 ^ n1814 ;
  assign n5379 = n5378 ^ n2613 ^ 1'b0 ;
  assign n5380 = ~n786 & n5379 ;
  assign n5377 = n1911 & ~n4925 ;
  assign n5381 = n5380 ^ n5377 ^ 1'b0 ;
  assign n5385 = n5384 ^ n5381 ^ n5060 ;
  assign n5386 = ( ~n3723 & n5376 ) | ( ~n3723 & n5385 ) | ( n5376 & n5385 ) ;
  assign n5387 = x51 & ~n3341 ;
  assign n5388 = n4923 & ~n5387 ;
  assign n5389 = ~n5386 & n5388 ;
  assign n5390 = x220 & ~n487 ;
  assign n5391 = n5390 ^ n1113 ^ n575 ;
  assign n5392 = n5391 ^ n438 ^ x57 ;
  assign n5393 = ~n2424 & n5392 ;
  assign n5398 = n2080 ^ n906 ^ 1'b0 ;
  assign n5394 = ( n1184 & n1968 ) | ( n1184 & ~n4890 ) | ( n1968 & ~n4890 ) ;
  assign n5395 = n2594 ^ n1901 ^ n1354 ;
  assign n5396 = n5394 | n5395 ;
  assign n5397 = x199 & ~n5396 ;
  assign n5399 = n5398 ^ n5397 ^ 1'b0 ;
  assign n5400 = ( x95 & n3126 ) | ( x95 & n4451 ) | ( n3126 & n4451 ) ;
  assign n5401 = n5400 ^ n2706 ^ 1'b0 ;
  assign n5402 = n1736 & ~n5401 ;
  assign n5403 = n5399 & n5402 ;
  assign n5406 = n2760 ^ x188 ^ x157 ;
  assign n5404 = ( ~n1832 & n3083 ) | ( ~n1832 & n5195 ) | ( n3083 & n5195 ) ;
  assign n5405 = x148 & n5404 ;
  assign n5407 = n5406 ^ n5405 ^ n310 ;
  assign n5408 = n2858 | n3408 ;
  assign n5409 = n5408 ^ n5147 ^ 1'b0 ;
  assign n5410 = n5409 ^ n1987 ^ x0 ;
  assign n5411 = ( n1225 & ~n4911 ) | ( n1225 & n5410 ) | ( ~n4911 & n5410 ) ;
  assign n5412 = ( n1780 & n3214 ) | ( n1780 & ~n5411 ) | ( n3214 & ~n5411 ) ;
  assign n5413 = n1308 & ~n2610 ;
  assign n5414 = ~n3717 & n5413 ;
  assign n5415 = n5237 ^ n4599 ^ n822 ;
  assign n5416 = n280 & ~n856 ;
  assign n5417 = n2996 ^ n2217 ^ x33 ;
  assign n5418 = ( n361 & ~n5416 ) | ( n361 & n5417 ) | ( ~n5416 & n5417 ) ;
  assign n5419 = n5418 ^ n953 ^ n843 ;
  assign n5420 = ( ~n1064 & n1091 ) | ( ~n1064 & n4697 ) | ( n1091 & n4697 ) ;
  assign n5421 = n5420 ^ n3535 ^ x149 ;
  assign n5422 = n931 & n5421 ;
  assign n5423 = n3943 & n5422 ;
  assign n5424 = n4049 ^ n3363 ^ n2247 ;
  assign n5425 = ~n1689 & n5424 ;
  assign n5426 = n5425 ^ n3085 ^ x68 ;
  assign n5427 = ~n484 & n5426 ;
  assign n5428 = ~n650 & n3213 ;
  assign n5429 = n2718 ^ n2081 ^ n763 ;
  assign n5430 = n5429 ^ n4342 ^ n3973 ;
  assign n5431 = n5430 ^ n4697 ^ n3387 ;
  assign n5432 = ( n2181 & n5428 ) | ( n2181 & ~n5431 ) | ( n5428 & ~n5431 ) ;
  assign n5433 = n5427 & ~n5432 ;
  assign n5434 = ( n1487 & n3879 ) | ( n1487 & n3895 ) | ( n3879 & n3895 ) ;
  assign n5438 = n4597 ^ n3437 ^ n2590 ;
  assign n5435 = n1377 ^ n817 ^ 1'b0 ;
  assign n5436 = n5435 ^ n3265 ^ 1'b0 ;
  assign n5437 = x181 & n5436 ;
  assign n5439 = n5438 ^ n5437 ^ n4120 ;
  assign n5440 = n5439 ^ n5323 ^ 1'b0 ;
  assign n5441 = n5434 & n5440 ;
  assign n5442 = ~n2259 & n5441 ;
  assign n5456 = n385 ^ n318 ^ x233 ;
  assign n5457 = n789 | n5456 ;
  assign n5455 = x202 & ~n1565 ;
  assign n5458 = n5457 ^ n5455 ^ 1'b0 ;
  assign n5451 = n2097 ^ n2085 ^ 1'b0 ;
  assign n5452 = n5451 ^ n2520 ^ n1143 ;
  assign n5453 = ( n513 & n664 ) | ( n513 & n5452 ) | ( n664 & n5452 ) ;
  assign n5450 = n4225 ^ n2302 ^ n1921 ;
  assign n5454 = n5453 ^ n5450 ^ n683 ;
  assign n5443 = n3247 ^ n2664 ^ n2318 ;
  assign n5444 = ( n905 & n4230 ) | ( n905 & ~n5443 ) | ( n4230 & ~n5443 ) ;
  assign n5445 = n1979 & ~n2184 ;
  assign n5446 = ( n1838 & n2222 ) | ( n1838 & ~n5445 ) | ( n2222 & ~n5445 ) ;
  assign n5447 = n5446 ^ n2210 ^ 1'b0 ;
  assign n5448 = n5447 ^ n1093 ^ 1'b0 ;
  assign n5449 = ( n2697 & n5444 ) | ( n2697 & ~n5448 ) | ( n5444 & ~n5448 ) ;
  assign n5459 = n5458 ^ n5454 ^ n5449 ;
  assign n5460 = n2081 ^ n1003 ^ 1'b0 ;
  assign n5461 = n522 & ~n5460 ;
  assign n5462 = ( n689 & n2449 ) | ( n689 & n3561 ) | ( n2449 & n3561 ) ;
  assign n5463 = ( n2523 & ~n5461 ) | ( n2523 & n5462 ) | ( ~n5461 & n5462 ) ;
  assign n5464 = n4853 ^ n4068 ^ n950 ;
  assign n5465 = n5464 ^ n3441 ^ n1629 ;
  assign n5466 = ( n2842 & ~n5463 ) | ( n2842 & n5465 ) | ( ~n5463 & n5465 ) ;
  assign n5467 = x72 & ~n452 ;
  assign n5468 = n5467 ^ n2839 ^ n425 ;
  assign n5469 = n5468 ^ n4172 ^ 1'b0 ;
  assign n5470 = ( n3054 & n5466 ) | ( n3054 & n5469 ) | ( n5466 & n5469 ) ;
  assign n5471 = n4987 ^ n4771 ^ x235 ;
  assign n5472 = n694 & ~n2539 ;
  assign n5473 = n5472 ^ n2701 ^ 1'b0 ;
  assign n5474 = n1897 & n5473 ;
  assign n5475 = n5471 & n5474 ;
  assign n5476 = n4164 & ~n5475 ;
  assign n5477 = n5476 ^ n2565 ^ 1'b0 ;
  assign n5478 = n5332 ^ n3596 ^ n442 ;
  assign n5479 = n1594 | n1890 ;
  assign n5480 = n5479 ^ n5471 ^ n2948 ;
  assign n5501 = ( x198 & n372 ) | ( x198 & n636 ) | ( n372 & n636 ) ;
  assign n5496 = n732 & ~n1272 ;
  assign n5497 = n3151 ^ n2737 ^ 1'b0 ;
  assign n5498 = ~n3873 & n5497 ;
  assign n5499 = n5496 & n5498 ;
  assign n5500 = n5499 ^ n1693 ^ 1'b0 ;
  assign n5492 = ( n430 & n1702 ) | ( n430 & n3099 ) | ( n1702 & n3099 ) ;
  assign n5493 = n1503 | n5492 ;
  assign n5494 = n5493 ^ n4724 ^ n2742 ;
  assign n5481 = n442 & n981 ;
  assign n5482 = ( ~n1952 & n4514 ) | ( ~n1952 & n5481 ) | ( n4514 & n5481 ) ;
  assign n5483 = n1972 ^ n345 ^ 1'b0 ;
  assign n5484 = ~n4305 & n5483 ;
  assign n5485 = n4295 & ~n5484 ;
  assign n5488 = ( n2655 & ~n3134 ) | ( n2655 & n4063 ) | ( ~n3134 & n4063 ) ;
  assign n5489 = n5488 ^ n2792 ^ 1'b0 ;
  assign n5486 = n3501 ^ n2024 ^ 1'b0 ;
  assign n5487 = n3942 & ~n5486 ;
  assign n5490 = n5489 ^ n5487 ^ n3854 ;
  assign n5491 = ( ~n5482 & n5485 ) | ( ~n5482 & n5490 ) | ( n5485 & n5490 ) ;
  assign n5495 = n5494 ^ n5491 ^ n3608 ;
  assign n5502 = n5501 ^ n5500 ^ n5495 ;
  assign n5503 = ( ~n3333 & n5480 ) | ( ~n3333 & n5502 ) | ( n5480 & n5502 ) ;
  assign n5504 = n4867 & n5503 ;
  assign n5505 = n3457 ^ n2161 ^ n1242 ;
  assign n5506 = n2508 & ~n5505 ;
  assign n5507 = n1198 & n2580 ;
  assign n5508 = n5507 ^ n311 ^ 1'b0 ;
  assign n5509 = ( n606 & ~n3871 ) | ( n606 & n5508 ) | ( ~n3871 & n5508 ) ;
  assign n5510 = n2364 & ~n5509 ;
  assign n5511 = n2760 & n5510 ;
  assign n5512 = ( n1131 & ~n2592 ) | ( n1131 & n4100 ) | ( ~n2592 & n4100 ) ;
  assign n5513 = ~n531 & n1758 ;
  assign n5514 = n5513 ^ n3557 ^ 1'b0 ;
  assign n5515 = n5514 ^ n3933 ^ n3024 ;
  assign n5516 = ( ~n2826 & n3449 ) | ( ~n2826 & n5515 ) | ( n3449 & n5515 ) ;
  assign n5517 = ( ~n5153 & n5512 ) | ( ~n5153 & n5516 ) | ( n5512 & n5516 ) ;
  assign n5518 = n711 & n2960 ;
  assign n5519 = n5518 ^ n4579 ^ 1'b0 ;
  assign n5520 = ( x49 & n1391 ) | ( x49 & n1783 ) | ( n1391 & n1783 ) ;
  assign n5521 = n5520 ^ n5492 ^ n1754 ;
  assign n5522 = n5519 & n5521 ;
  assign n5525 = ( n815 & n1032 ) | ( n815 & n1839 ) | ( n1032 & n1839 ) ;
  assign n5526 = ( n2461 & n5165 ) | ( n2461 & n5525 ) | ( n5165 & n5525 ) ;
  assign n5523 = ( n351 & ~n1006 ) | ( n351 & n2697 ) | ( ~n1006 & n2697 ) ;
  assign n5524 = n2660 & ~n5523 ;
  assign n5527 = n5526 ^ n5524 ^ n3729 ;
  assign n5528 = ~n2655 & n2836 ;
  assign n5529 = n2033 & n5528 ;
  assign n5530 = ( n1799 & n3175 ) | ( n1799 & ~n5529 ) | ( n3175 & ~n5529 ) ;
  assign n5531 = n5530 ^ n3213 ^ 1'b0 ;
  assign n5532 = ~n874 & n3211 ;
  assign n5533 = ( n1595 & ~n3002 ) | ( n1595 & n5532 ) | ( ~n3002 & n5532 ) ;
  assign n5534 = ( n3262 & ~n3758 ) | ( n3262 & n5533 ) | ( ~n3758 & n5533 ) ;
  assign n5535 = n5531 & n5534 ;
  assign n5536 = n1777 & n5535 ;
  assign n5537 = n271 & n2040 ;
  assign n5538 = n5537 ^ n2058 ^ 1'b0 ;
  assign n5539 = n5538 ^ n3263 ^ 1'b0 ;
  assign n5540 = ~n1254 & n5539 ;
  assign n5541 = n3472 ^ n1345 ^ 1'b0 ;
  assign n5542 = ~n431 & n5541 ;
  assign n5543 = n5542 ^ n3185 ^ n2660 ;
  assign n5544 = ( n2758 & n3541 ) | ( n2758 & ~n3887 ) | ( n3541 & ~n3887 ) ;
  assign n5545 = n2271 | n2929 ;
  assign n5546 = n5544 & ~n5545 ;
  assign n5547 = n4781 ^ n2509 ^ n2176 ;
  assign n5548 = ( n1651 & n2741 ) | ( n1651 & n4919 ) | ( n2741 & n4919 ) ;
  assign n5549 = n5548 ^ n3185 ^ 1'b0 ;
  assign n5550 = n1668 & ~n5549 ;
  assign n5551 = n5479 ^ n1361 ^ 1'b0 ;
  assign n5552 = n280 & n5551 ;
  assign n5553 = ( n3320 & n5550 ) | ( n3320 & ~n5552 ) | ( n5550 & ~n5552 ) ;
  assign n5554 = ( n997 & ~n2209 ) | ( n997 & n4852 ) | ( ~n2209 & n4852 ) ;
  assign n5555 = ( n1948 & n4080 ) | ( n1948 & n5554 ) | ( n4080 & n5554 ) ;
  assign n5556 = ( x134 & ~n3292 ) | ( x134 & n5555 ) | ( ~n3292 & n5555 ) ;
  assign n5557 = ~n528 & n2445 ;
  assign n5558 = n5557 ^ n3626 ^ 1'b0 ;
  assign n5559 = n5558 ^ n3102 ^ 1'b0 ;
  assign n5560 = n5556 & n5559 ;
  assign n5561 = n5560 ^ n1020 ^ 1'b0 ;
  assign n5562 = n5002 ^ n2894 ^ n1355 ;
  assign n5563 = ( ~n644 & n977 ) | ( ~n644 & n5562 ) | ( n977 & n5562 ) ;
  assign n5565 = n2591 ^ x233 ^ 1'b0 ;
  assign n5564 = ( ~n1290 & n1762 ) | ( ~n1290 & n2832 ) | ( n1762 & n2832 ) ;
  assign n5566 = n5565 ^ n5564 ^ 1'b0 ;
  assign n5567 = n5566 ^ n2553 ^ n462 ;
  assign n5568 = n1181 & ~n2318 ;
  assign n5569 = n369 & n5568 ;
  assign n5570 = n4990 ^ n3481 ^ n2435 ;
  assign n5571 = n374 & ~n890 ;
  assign n5572 = n5571 ^ n600 ^ n408 ;
  assign n5573 = ~n2039 & n5572 ;
  assign n5574 = n5573 ^ n3166 ^ 1'b0 ;
  assign n5575 = n755 ^ n740 ^ n325 ;
  assign n5576 = ( ~n1245 & n4381 ) | ( ~n1245 & n5575 ) | ( n4381 & n5575 ) ;
  assign n5577 = ( ~x157 & n932 ) | ( ~x157 & n1827 ) | ( n932 & n1827 ) ;
  assign n5578 = n5577 ^ n4841 ^ x212 ;
  assign n5579 = ( n5574 & ~n5576 ) | ( n5574 & n5578 ) | ( ~n5576 & n5578 ) ;
  assign n5580 = n4284 ^ n1775 ^ n1299 ;
  assign n5581 = n1257 ^ n549 ^ x154 ;
  assign n5582 = n5581 ^ n1003 ^ n887 ;
  assign n5583 = ~x72 & n2178 ;
  assign n5584 = n2412 | n5583 ;
  assign n5585 = n5584 ^ n587 ^ 1'b0 ;
  assign n5586 = n1240 | n5585 ;
  assign n5587 = n556 | n5586 ;
  assign n5588 = n261 & n5587 ;
  assign n5589 = n4275 ^ n3837 ^ 1'b0 ;
  assign n5591 = n4597 ^ n931 ^ n326 ;
  assign n5590 = n405 | n2066 ;
  assign n5592 = n5591 ^ n5590 ^ 1'b0 ;
  assign n5593 = n1425 | n3991 ;
  assign n5594 = n468 & n5593 ;
  assign n5595 = n5594 ^ n1529 ^ 1'b0 ;
  assign n5596 = ( n592 & n5592 ) | ( n592 & ~n5595 ) | ( n5592 & ~n5595 ) ;
  assign n5597 = ( n5588 & ~n5589 ) | ( n5588 & n5596 ) | ( ~n5589 & n5596 ) ;
  assign n5598 = n5496 ^ n2484 ^ n1168 ;
  assign n5599 = n2889 ^ n2132 ^ x187 ;
  assign n5600 = ( n807 & n5555 ) | ( n807 & n5599 ) | ( n5555 & n5599 ) ;
  assign n5601 = n4788 & ~n5600 ;
  assign n5602 = n5601 ^ n3713 ^ 1'b0 ;
  assign n5603 = ( n2699 & n4010 ) | ( n2699 & ~n5602 ) | ( n4010 & ~n5602 ) ;
  assign n5606 = n639 ^ n415 ^ 1'b0 ;
  assign n5607 = ~n1925 & n5606 ;
  assign n5604 = ( ~n1316 & n1858 ) | ( ~n1316 & n1955 ) | ( n1858 & n1955 ) ;
  assign n5605 = n1035 | n5604 ;
  assign n5608 = n5607 ^ n5605 ^ 1'b0 ;
  assign n5614 = n1475 & n3600 ;
  assign n5615 = n5614 ^ n4931 ^ 1'b0 ;
  assign n5616 = n4970 & n5615 ;
  assign n5610 = ~n576 & n754 ;
  assign n5611 = n5610 ^ n3262 ^ 1'b0 ;
  assign n5612 = ( x20 & n850 ) | ( x20 & ~n5611 ) | ( n850 & ~n5611 ) ;
  assign n5613 = ( n1287 & n2516 ) | ( n1287 & n5612 ) | ( n2516 & n5612 ) ;
  assign n5609 = n5493 ^ n2774 ^ 1'b0 ;
  assign n5617 = n5616 ^ n5613 ^ n5609 ;
  assign n5618 = ( n4902 & n5608 ) | ( n4902 & n5617 ) | ( n5608 & n5617 ) ;
  assign n5619 = ( n1308 & ~n3239 ) | ( n1308 & n5618 ) | ( ~n3239 & n5618 ) ;
  assign n5620 = ( ~n5598 & n5603 ) | ( ~n5598 & n5619 ) | ( n5603 & n5619 ) ;
  assign n5622 = n3217 ^ n1670 ^ 1'b0 ;
  assign n5623 = n5622 ^ n5335 ^ 1'b0 ;
  assign n5621 = n5409 ^ n2764 ^ 1'b0 ;
  assign n5624 = n5623 ^ n5621 ^ n1703 ;
  assign n5625 = n345 & n5624 ;
  assign n5626 = ~n2881 & n5625 ;
  assign n5627 = n2474 & n2884 ;
  assign n5630 = n5435 ^ n4248 ^ x171 ;
  assign n5628 = n3871 ^ n2397 ^ n1250 ;
  assign n5629 = ( n2070 & ~n2565 ) | ( n2070 & n5628 ) | ( ~n2565 & n5628 ) ;
  assign n5631 = n5630 ^ n5629 ^ 1'b0 ;
  assign n5632 = n566 | n5631 ;
  assign n5633 = ( n2303 & n4447 ) | ( n2303 & n5534 ) | ( n4447 & n5534 ) ;
  assign n5634 = ( n2471 & ~n5252 ) | ( n2471 & n5418 ) | ( ~n5252 & n5418 ) ;
  assign n5635 = n1095 ^ n1003 ^ x60 ;
  assign n5636 = ( n1091 & n3426 ) | ( n1091 & n3759 ) | ( n3426 & n3759 ) ;
  assign n5637 = n5636 ^ n1898 ^ n1236 ;
  assign n5638 = ( ~n3917 & n5635 ) | ( ~n3917 & n5637 ) | ( n5635 & n5637 ) ;
  assign n5639 = ( n2552 & n3377 ) | ( n2552 & n5638 ) | ( n3377 & n5638 ) ;
  assign n5640 = ~n689 & n2401 ;
  assign n5641 = n5640 ^ n1573 ^ n1535 ;
  assign n5642 = ( ~n3103 & n5320 ) | ( ~n3103 & n5641 ) | ( n5320 & n5641 ) ;
  assign n5643 = ( ~n1780 & n5639 ) | ( ~n1780 & n5642 ) | ( n5639 & n5642 ) ;
  assign n5644 = n1740 | n4784 ;
  assign n5645 = n2059 | n5644 ;
  assign n5647 = n3802 & ~n4407 ;
  assign n5648 = ~n427 & n5647 ;
  assign n5646 = n1862 & n2717 ;
  assign n5649 = n5648 ^ n5646 ^ 1'b0 ;
  assign n5650 = ~n628 & n1530 ;
  assign n5651 = n1122 & n5650 ;
  assign n5652 = n5651 ^ x44 ^ 1'b0 ;
  assign n5653 = x195 & ~n1710 ;
  assign n5654 = n5653 ^ n4841 ^ 1'b0 ;
  assign n5655 = x10 & n5654 ;
  assign n5656 = n5655 ^ n4285 ^ n2200 ;
  assign n5657 = ( n4917 & n5652 ) | ( n4917 & n5656 ) | ( n5652 & n5656 ) ;
  assign n5661 = n1632 & n3113 ;
  assign n5659 = n436 & ~n2636 ;
  assign n5660 = n5659 ^ n1070 ^ 1'b0 ;
  assign n5658 = ( n1467 & ~n2807 ) | ( n1467 & n3238 ) | ( ~n2807 & n3238 ) ;
  assign n5662 = n5661 ^ n5660 ^ n5658 ;
  assign n5663 = n1875 | n3083 ;
  assign n5664 = ( n3352 & n4182 ) | ( n3352 & n4969 ) | ( n4182 & n4969 ) ;
  assign n5665 = n5623 ^ n3649 ^ n870 ;
  assign n5666 = ( n371 & ~n975 ) | ( n371 & n1659 ) | ( ~n975 & n1659 ) ;
  assign n5667 = ~n796 & n3922 ;
  assign n5668 = ( n1296 & n5666 ) | ( n1296 & n5667 ) | ( n5666 & n5667 ) ;
  assign n5669 = n5668 ^ n2689 ^ n1113 ;
  assign n5670 = ( ~n720 & n2184 ) | ( ~n720 & n2620 ) | ( n2184 & n2620 ) ;
  assign n5671 = ( ~x187 & n1291 ) | ( ~x187 & n5305 ) | ( n1291 & n5305 ) ;
  assign n5672 = n5044 ^ n4971 ^ 1'b0 ;
  assign n5673 = n5274 ^ n2786 ^ n1595 ;
  assign n5677 = n1717 & n2923 ;
  assign n5678 = n2092 & n5677 ;
  assign n5679 = ~n939 & n5678 ;
  assign n5680 = n2170 & ~n5679 ;
  assign n5674 = n1196 ^ n934 ^ 1'b0 ;
  assign n5675 = ( ~n3008 & n5062 ) | ( ~n3008 & n5674 ) | ( n5062 & n5674 ) ;
  assign n5676 = n5675 ^ n3017 ^ n308 ;
  assign n5681 = n5680 ^ n5676 ^ n790 ;
  assign n5682 = ( n1146 & n2114 ) | ( n1146 & n3747 ) | ( n2114 & n3747 ) ;
  assign n5683 = n3163 ^ n1855 ^ 1'b0 ;
  assign n5684 = n5682 & ~n5683 ;
  assign n5685 = ( ~n1202 & n2474 ) | ( ~n1202 & n3381 ) | ( n2474 & n3381 ) ;
  assign n5686 = ( ~n736 & n1774 ) | ( ~n736 & n5685 ) | ( n1774 & n5685 ) ;
  assign n5687 = n2884 ^ n2179 ^ n347 ;
  assign n5688 = n5686 | n5687 ;
  assign n5689 = ( n3084 & n4177 ) | ( n3084 & ~n5688 ) | ( n4177 & ~n5688 ) ;
  assign n5690 = ( n5681 & n5684 ) | ( n5681 & n5689 ) | ( n5684 & n5689 ) ;
  assign n5691 = n5690 ^ n1581 ^ 1'b0 ;
  assign n5693 = ( n1534 & n2779 ) | ( n1534 & n4924 ) | ( n2779 & n4924 ) ;
  assign n5692 = n2286 | n2673 ;
  assign n5694 = n5693 ^ n5692 ^ 1'b0 ;
  assign n5695 = ( n1748 & n2517 ) | ( n1748 & n5366 ) | ( n2517 & n5366 ) ;
  assign n5696 = n3674 ^ n3305 ^ 1'b0 ;
  assign n5697 = x134 & n1840 ;
  assign n5698 = n5697 ^ n4379 ^ n1290 ;
  assign n5699 = n5696 & n5698 ;
  assign n5700 = n5699 ^ n2425 ^ 1'b0 ;
  assign n5701 = n5700 ^ n3848 ^ n1038 ;
  assign n5702 = n2077 & ~n2263 ;
  assign n5703 = n3401 & n5702 ;
  assign n5704 = n2586 | n4223 ;
  assign n5705 = n5704 ^ n2462 ^ n2426 ;
  assign n5706 = ( ~n4196 & n5703 ) | ( ~n4196 & n5705 ) | ( n5703 & n5705 ) ;
  assign n5707 = n5706 ^ n2631 ^ 1'b0 ;
  assign n5717 = n2850 ^ n2456 ^ 1'b0 ;
  assign n5714 = ( n2020 & ~n2315 ) | ( n2020 & n3415 ) | ( ~n2315 & n3415 ) ;
  assign n5713 = ( n1752 & ~n2042 ) | ( n1752 & n2605 ) | ( ~n2042 & n2605 ) ;
  assign n5715 = n5714 ^ n5713 ^ 1'b0 ;
  assign n5716 = n5574 | n5715 ;
  assign n5710 = ( ~n1967 & n2243 ) | ( ~n1967 & n2961 ) | ( n2243 & n2961 ) ;
  assign n5711 = ( ~n2427 & n4712 ) | ( ~n2427 & n5710 ) | ( n4712 & n5710 ) ;
  assign n5708 = n3710 ^ n1675 ^ 1'b0 ;
  assign n5709 = x168 & n5708 ;
  assign n5712 = n5711 ^ n5709 ^ n363 ;
  assign n5718 = n5717 ^ n5716 ^ n5712 ;
  assign n5719 = ( ~n525 & n1534 ) | ( ~n525 & n3397 ) | ( n1534 & n3397 ) ;
  assign n5720 = n5719 ^ n4122 ^ 1'b0 ;
  assign n5721 = n5720 ^ n4017 ^ n1914 ;
  assign n5727 = n951 | n2479 ;
  assign n5728 = n4841 & ~n5727 ;
  assign n5729 = ~n3710 & n5728 ;
  assign n5725 = n3515 ^ n1647 ^ n644 ;
  assign n5722 = ( n690 & n1980 ) | ( n690 & ~n2555 ) | ( n1980 & ~n2555 ) ;
  assign n5723 = n5722 ^ n722 ^ 1'b0 ;
  assign n5724 = ( n925 & n3272 ) | ( n925 & n5723 ) | ( n3272 & n5723 ) ;
  assign n5726 = n5725 ^ n5724 ^ n2827 ;
  assign n5730 = n5729 ^ n5726 ^ 1'b0 ;
  assign n5731 = ( n3309 & n3549 ) | ( n3309 & ~n4197 ) | ( n3549 & ~n4197 ) ;
  assign n5732 = ( n1242 & n1692 ) | ( n1242 & n5731 ) | ( n1692 & n5731 ) ;
  assign n5733 = n4180 ^ n1554 ^ n416 ;
  assign n5734 = n5733 ^ n3742 ^ 1'b0 ;
  assign n5735 = n5732 | n5734 ;
  assign n5736 = ( n4306 & n5196 ) | ( n4306 & ~n5735 ) | ( n5196 & ~n5735 ) ;
  assign n5737 = ( n1080 & n1185 ) | ( n1080 & n4937 ) | ( n1185 & n4937 ) ;
  assign n5738 = ( ~n657 & n750 ) | ( ~n657 & n1330 ) | ( n750 & n1330 ) ;
  assign n5739 = n5738 ^ n3355 ^ 1'b0 ;
  assign n5740 = n5739 ^ n1809 ^ 1'b0 ;
  assign n5741 = n5740 ^ n2254 ^ 1'b0 ;
  assign n5742 = n5737 & ~n5741 ;
  assign n5743 = n2321 ^ n301 ^ 1'b0 ;
  assign n5744 = ( ~n1979 & n3489 ) | ( ~n1979 & n3585 ) | ( n3489 & n3585 ) ;
  assign n5745 = n4363 ^ n2870 ^ n1453 ;
  assign n5746 = n3374 & n5745 ;
  assign n5747 = ( n5743 & ~n5744 ) | ( n5743 & n5746 ) | ( ~n5744 & n5746 ) ;
  assign n5748 = n3943 | n5747 ;
  assign n5749 = n5131 ^ n3318 ^ n2705 ;
  assign n5754 = n4180 ^ n1327 ^ n410 ;
  assign n5752 = n5679 ^ n1539 ^ 1'b0 ;
  assign n5753 = n4876 | n5752 ;
  assign n5750 = n5406 ^ x156 ^ x109 ;
  assign n5751 = n5750 ^ n4830 ^ n2576 ;
  assign n5755 = n5754 ^ n5753 ^ n5751 ;
  assign n5756 = ( ~n1325 & n3456 ) | ( ~n1325 & n5755 ) | ( n3456 & n5755 ) ;
  assign n5757 = ( n2827 & n5749 ) | ( n2827 & ~n5756 ) | ( n5749 & ~n5756 ) ;
  assign n5763 = n4052 ^ n1528 ^ 1'b0 ;
  assign n5764 = n5763 ^ n4937 ^ n1417 ;
  assign n5765 = n5764 ^ n3312 ^ x145 ;
  assign n5759 = n2168 ^ n288 ^ x220 ;
  assign n5760 = ( n856 & n1240 ) | ( n856 & ~n5759 ) | ( n1240 & ~n5759 ) ;
  assign n5761 = n5760 ^ n2189 ^ n401 ;
  assign n5762 = n5761 ^ n1957 ^ n707 ;
  assign n5758 = n4666 ^ n3073 ^ n495 ;
  assign n5766 = n5765 ^ n5762 ^ n5758 ;
  assign n5767 = n2438 ^ n2266 ^ n1061 ;
  assign n5768 = ~n3203 & n5403 ;
  assign n5769 = ~n5767 & n5768 ;
  assign n5770 = n1376 ^ n872 ^ 1'b0 ;
  assign n5771 = n2190 ^ n682 ^ 1'b0 ;
  assign n5772 = n5770 & ~n5771 ;
  assign n5773 = n4784 & n5772 ;
  assign n5774 = n2743 ^ n545 ^ x131 ;
  assign n5775 = n278 & ~n3928 ;
  assign n5776 = n5304 ^ n3323 ^ 1'b0 ;
  assign n5777 = n3840 ^ n3562 ^ n3212 ;
  assign n5778 = n5777 ^ n2635 ^ n1692 ;
  assign n5779 = n3978 ^ n732 ^ 1'b0 ;
  assign n5780 = n447 & n5779 ;
  assign n5781 = ~n1695 & n3493 ;
  assign n5782 = ~n2127 & n5781 ;
  assign n5783 = n5782 ^ n5190 ^ 1'b0 ;
  assign n5784 = n5780 & ~n5783 ;
  assign n5788 = n4225 ^ n3022 ^ 1'b0 ;
  assign n5789 = n614 | n5788 ;
  assign n5785 = ~n670 & n1460 ;
  assign n5786 = n299 & n5785 ;
  assign n5787 = n5786 ^ n2333 ^ n517 ;
  assign n5790 = n5789 ^ n5787 ^ n711 ;
  assign n5791 = n3077 & n5790 ;
  assign n5792 = n5791 ^ n970 ^ 1'b0 ;
  assign n5793 = n1349 | n3530 ;
  assign n5794 = n2078 | n5793 ;
  assign n5795 = ( n3948 & n5195 ) | ( n3948 & n5794 ) | ( n5195 & n5794 ) ;
  assign n5796 = n2806 ^ n524 ^ 1'b0 ;
  assign n5797 = n2089 ^ n920 ^ x91 ;
  assign n5798 = ( x188 & ~n947 ) | ( x188 & n5797 ) | ( ~n947 & n5797 ) ;
  assign n5799 = n5798 ^ n3958 ^ n3414 ;
  assign n5800 = n5799 ^ n4983 ^ n4481 ;
  assign n5801 = ( n711 & ~n1795 ) | ( n711 & n5800 ) | ( ~n1795 & n5800 ) ;
  assign n5802 = n3226 ^ n3141 ^ n2793 ;
  assign n5803 = n791 ^ x15 ^ 1'b0 ;
  assign n5804 = n2717 & ~n5803 ;
  assign n5805 = n1756 & n5804 ;
  assign n5806 = n4257 & n5805 ;
  assign n5807 = ~n1935 & n2885 ;
  assign n5808 = ~n749 & n5807 ;
  assign n5809 = n5808 ^ n2827 ^ n1851 ;
  assign n5810 = ( n4381 & ~n5806 ) | ( n4381 & n5809 ) | ( ~n5806 & n5809 ) ;
  assign n5811 = n3024 ^ n2099 ^ n916 ;
  assign n5812 = n5811 ^ n3296 ^ n1594 ;
  assign n5815 = n4969 ^ n4005 ^ x86 ;
  assign n5813 = n504 ^ x229 ^ 1'b0 ;
  assign n5814 = n1665 & ~n5813 ;
  assign n5816 = n5815 ^ n5814 ^ 1'b0 ;
  assign n5817 = n5812 & n5816 ;
  assign n5820 = n3902 ^ n2395 ^ n1436 ;
  assign n5821 = ( x29 & n614 ) | ( x29 & n2052 ) | ( n614 & n2052 ) ;
  assign n5822 = n1205 & n5821 ;
  assign n5823 = ~n5820 & n5822 ;
  assign n5818 = ~n1018 & n4131 ;
  assign n5819 = n5818 ^ n5608 ^ n653 ;
  assign n5824 = n5823 ^ n5819 ^ n3221 ;
  assign n5825 = n2455 ^ n771 ^ 1'b0 ;
  assign n5831 = ( n677 & ~n1012 ) | ( n677 & n2124 ) | ( ~n1012 & n2124 ) ;
  assign n5832 = ( n597 & n1200 ) | ( n597 & ~n5831 ) | ( n1200 & ~n5831 ) ;
  assign n5833 = ( x196 & ~n2549 ) | ( x196 & n5832 ) | ( ~n2549 & n5832 ) ;
  assign n5830 = n2899 ^ n523 ^ n463 ;
  assign n5826 = x134 & ~n680 ;
  assign n5827 = n5826 ^ n2164 ^ 1'b0 ;
  assign n5828 = n5827 ^ n3151 ^ x203 ;
  assign n5829 = ( n755 & n1708 ) | ( n755 & n5828 ) | ( n1708 & n5828 ) ;
  assign n5834 = n5833 ^ n5830 ^ n5829 ;
  assign n5837 = n735 & ~n3496 ;
  assign n5835 = n3355 | n3505 ;
  assign n5836 = n5835 ^ n5668 ^ 1'b0 ;
  assign n5838 = n5837 ^ n5836 ^ n467 ;
  assign n5839 = ( n5825 & n5834 ) | ( n5825 & n5838 ) | ( n5834 & n5838 ) ;
  assign n5840 = n5318 ^ n3096 ^ n2366 ;
  assign n5849 = ( n1006 & ~n2326 ) | ( n1006 & n2393 ) | ( ~n2326 & n2393 ) ;
  assign n5846 = n4005 ^ n956 ^ x204 ;
  assign n5841 = x250 & ~n1042 ;
  assign n5842 = ( n538 & ~n2397 ) | ( n538 & n5841 ) | ( ~n2397 & n5841 ) ;
  assign n5843 = n1090 ^ x137 ^ 1'b0 ;
  assign n5844 = ( ~n3812 & n5842 ) | ( ~n3812 & n5843 ) | ( n5842 & n5843 ) ;
  assign n5845 = n3695 & n5844 ;
  assign n5847 = n5846 ^ n5845 ^ 1'b0 ;
  assign n5848 = n5847 ^ n2871 ^ n2662 ;
  assign n5850 = n5849 ^ n5848 ^ n1889 ;
  assign n5851 = ( n755 & n1463 ) | ( n755 & ~n4493 ) | ( n1463 & ~n4493 ) ;
  assign n5855 = x9 & n1758 ;
  assign n5856 = ~x112 & n5855 ;
  assign n5857 = ( n504 & ~n606 ) | ( n504 & n5856 ) | ( ~n606 & n5856 ) ;
  assign n5852 = n3443 ^ n2842 ^ n273 ;
  assign n5853 = n1237 & n5852 ;
  assign n5854 = ~n2846 & n5853 ;
  assign n5858 = n5857 ^ n5854 ^ 1'b0 ;
  assign n5859 = ( n4130 & ~n4645 ) | ( n4130 & n5858 ) | ( ~n4645 & n5858 ) ;
  assign n5860 = ( n959 & n5851 ) | ( n959 & n5859 ) | ( n5851 & n5859 ) ;
  assign n5861 = ( ~n1650 & n3084 ) | ( ~n1650 & n3828 ) | ( n3084 & n3828 ) ;
  assign n5862 = n2124 & ~n5293 ;
  assign n5863 = n5862 ^ n5789 ^ 1'b0 ;
  assign n5864 = ~x41 & n594 ;
  assign n5865 = n5864 ^ n3963 ^ 1'b0 ;
  assign n5866 = n2101 & ~n5865 ;
  assign n5867 = n5863 & n5866 ;
  assign n5868 = ~n915 & n5562 ;
  assign n5869 = n5868 ^ n4023 ^ 1'b0 ;
  assign n5870 = n5869 ^ n2896 ^ n1678 ;
  assign n5871 = x35 & ~n3991 ;
  assign n5872 = n5871 ^ n4909 ^ n1774 ;
  assign n5874 = n2301 & ~n4894 ;
  assign n5873 = ( n2737 & n3752 ) | ( n2737 & ~n5205 ) | ( n3752 & ~n5205 ) ;
  assign n5875 = n5874 ^ n5873 ^ n2058 ;
  assign n5878 = n4248 ^ n1137 ^ 1'b0 ;
  assign n5876 = n5328 ^ n5118 ^ n1911 ;
  assign n5877 = n5876 ^ n1656 ^ 1'b0 ;
  assign n5879 = n5878 ^ n5877 ^ n2774 ;
  assign n5880 = ( n3228 & n5875 ) | ( n3228 & n5879 ) | ( n5875 & n5879 ) ;
  assign n5881 = ( n5870 & n5872 ) | ( n5870 & n5880 ) | ( n5872 & n5880 ) ;
  assign n5882 = n1295 ^ x253 ^ 1'b0 ;
  assign n5884 = ( n836 & n1048 ) | ( n836 & n2372 ) | ( n1048 & n2372 ) ;
  assign n5885 = n5884 ^ n3799 ^ 1'b0 ;
  assign n5886 = x241 & ~n5885 ;
  assign n5883 = n1391 | n1788 ;
  assign n5887 = n5886 ^ n5883 ^ n5503 ;
  assign n5888 = n5696 ^ n529 ^ n286 ;
  assign n5890 = n1225 ^ n683 ^ n299 ;
  assign n5891 = n1817 & n5890 ;
  assign n5892 = n270 & n5891 ;
  assign n5893 = ( ~n2364 & n2411 ) | ( ~n2364 & n2545 ) | ( n2411 & n2545 ) ;
  assign n5894 = n5893 ^ n3504 ^ n1241 ;
  assign n5895 = n1771 & ~n5894 ;
  assign n5896 = n5892 & n5895 ;
  assign n5889 = ~n4331 & n4410 ;
  assign n5897 = n5896 ^ n5889 ^ 1'b0 ;
  assign n5898 = ( ~n424 & n5447 ) | ( ~n424 & n5897 ) | ( n5447 & n5897 ) ;
  assign n5899 = n4361 ^ n2301 ^ 1'b0 ;
  assign n5906 = ( x91 & ~n739 ) | ( x91 & n3933 ) | ( ~n739 & n3933 ) ;
  assign n5907 = n5906 ^ n5118 ^ 1'b0 ;
  assign n5908 = ( n456 & ~n4353 ) | ( n456 & n5907 ) | ( ~n4353 & n5907 ) ;
  assign n5904 = n1564 ^ n1301 ^ x41 ;
  assign n5900 = n1330 ^ x146 ^ 1'b0 ;
  assign n5901 = n531 & ~n5900 ;
  assign n5902 = n5901 ^ n2394 ^ 1'b0 ;
  assign n5903 = n5902 ^ n2024 ^ n1736 ;
  assign n5905 = n5904 ^ n5903 ^ x219 ;
  assign n5909 = n5908 ^ n5905 ^ n4503 ;
  assign n5910 = n5015 ^ n3580 ^ n282 ;
  assign n5911 = n5910 ^ n3556 ^ 1'b0 ;
  assign n5915 = n2454 ^ x27 ^ 1'b0 ;
  assign n5914 = n758 | n3710 ;
  assign n5916 = n5915 ^ n5914 ^ 1'b0 ;
  assign n5912 = n4926 ^ n3035 ^ n858 ;
  assign n5913 = n5912 ^ n310 ^ 1'b0 ;
  assign n5917 = n5916 ^ n5913 ^ 1'b0 ;
  assign n5918 = ( n1392 & n1884 ) | ( n1392 & ~n3052 ) | ( n1884 & ~n3052 ) ;
  assign n5919 = n3981 ^ n1655 ^ n261 ;
  assign n5920 = ( ~n4293 & n5918 ) | ( ~n4293 & n5919 ) | ( n5918 & n5919 ) ;
  assign n5921 = ( n1898 & n5707 ) | ( n1898 & n5920 ) | ( n5707 & n5920 ) ;
  assign n5924 = ( n1365 & n2632 ) | ( n1365 & n3350 ) | ( n2632 & n3350 ) ;
  assign n5923 = n5173 ^ n3963 ^ n1197 ;
  assign n5922 = ~n4275 & n5682 ;
  assign n5925 = n5924 ^ n5923 ^ n5922 ;
  assign n5926 = ~n4865 & n5129 ;
  assign n5927 = n4406 ^ n1294 ^ 1'b0 ;
  assign n5928 = ~n2693 & n5927 ;
  assign n5929 = ~n5926 & n5928 ;
  assign n5930 = ( n2089 & n5925 ) | ( n2089 & n5929 ) | ( n5925 & n5929 ) ;
  assign n5931 = x42 & ~n1556 ;
  assign n5932 = n5931 ^ n3068 ^ n1896 ;
  assign n5933 = n5932 ^ n860 ^ 1'b0 ;
  assign n5934 = n5933 ^ n5033 ^ 1'b0 ;
  assign n5939 = n2527 ^ x13 ^ 1'b0 ;
  assign n5940 = x84 & n421 ;
  assign n5941 = n5940 ^ n4188 ^ 1'b0 ;
  assign n5942 = ( ~n1139 & n2849 ) | ( ~n1139 & n5941 ) | ( n2849 & n5941 ) ;
  assign n5943 = ( n2658 & n5939 ) | ( n2658 & ~n5942 ) | ( n5939 & ~n5942 ) ;
  assign n5935 = ~n2535 & n3414 ;
  assign n5936 = n5935 ^ n1936 ^ n1037 ;
  assign n5937 = ~n2133 & n2546 ;
  assign n5938 = ( n5690 & n5936 ) | ( n5690 & ~n5937 ) | ( n5936 & ~n5937 ) ;
  assign n5944 = n5943 ^ n5938 ^ n4895 ;
  assign n5945 = n4472 ^ n2819 ^ n1130 ;
  assign n5946 = x22 & n874 ;
  assign n5947 = ~n617 & n5946 ;
  assign n5948 = ( n1096 & n2143 ) | ( n1096 & ~n5947 ) | ( n2143 & ~n5947 ) ;
  assign n5952 = ~n1589 & n2111 ;
  assign n5949 = n2583 ^ n1650 ^ 1'b0 ;
  assign n5950 = ~n2824 & n5949 ;
  assign n5951 = ( n3208 & n5594 ) | ( n3208 & n5950 ) | ( n5594 & n5950 ) ;
  assign n5953 = n5952 ^ n5951 ^ n3690 ;
  assign n5954 = n5948 & n5953 ;
  assign n5955 = ~n5945 & n5954 ;
  assign n5956 = ( n1210 & n2528 ) | ( n1210 & n5400 ) | ( n2528 & n5400 ) ;
  assign n5957 = n1961 & ~n5956 ;
  assign n5958 = n2444 & ~n4475 ;
  assign n5960 = x50 & n1603 ;
  assign n5961 = ~n4780 & n5960 ;
  assign n5959 = ( n1110 & ~n3765 ) | ( n1110 & n4188 ) | ( ~n3765 & n4188 ) ;
  assign n5962 = n5961 ^ n5959 ^ n2193 ;
  assign n5963 = n5962 ^ n3609 ^ n1229 ;
  assign n5964 = n1271 & ~n1894 ;
  assign n5965 = ( ~x73 & n3048 ) | ( ~x73 & n5964 ) | ( n3048 & n5964 ) ;
  assign n5966 = n5965 ^ n634 ^ 1'b0 ;
  assign n5967 = n1276 & ~n1588 ;
  assign n5968 = n5967 ^ n2042 ^ n1619 ;
  assign n5969 = n5968 ^ x135 ^ 1'b0 ;
  assign n5970 = ( n2466 & ~n3040 ) | ( n2466 & n3117 ) | ( ~n3040 & n3117 ) ;
  assign n5971 = n5071 & n5970 ;
  assign n5972 = n5971 ^ n325 ^ 1'b0 ;
  assign n5977 = n883 & n2175 ;
  assign n5978 = ~n2927 & n5977 ;
  assign n5979 = ( n1577 & n5555 ) | ( n1577 & ~n5978 ) | ( n5555 & ~n5978 ) ;
  assign n5980 = ( ~x12 & n1480 ) | ( ~x12 & n2591 ) | ( n1480 & n2591 ) ;
  assign n5981 = ( ~x86 & n1142 ) | ( ~x86 & n5980 ) | ( n1142 & n5980 ) ;
  assign n5982 = n5981 ^ n2019 ^ 1'b0 ;
  assign n5983 = n5979 & n5982 ;
  assign n5973 = n5585 ^ n809 ^ 1'b0 ;
  assign n5974 = n4301 ^ n3528 ^ n1118 ;
  assign n5975 = n5974 ^ n2042 ^ n1099 ;
  assign n5976 = ( n583 & n5973 ) | ( n583 & ~n5975 ) | ( n5973 & ~n5975 ) ;
  assign n5984 = n5983 ^ n5976 ^ n921 ;
  assign n5985 = n5984 ^ n2686 ^ 1'b0 ;
  assign n5986 = ( ~x14 & n1056 ) | ( ~x14 & n2759 ) | ( n1056 & n2759 ) ;
  assign n5987 = n5986 ^ n2200 ^ n1210 ;
  assign n5988 = n2710 ^ x235 ^ x130 ;
  assign n5997 = n1707 | n3048 ;
  assign n5998 = n5142 ^ n3429 ^ x217 ;
  assign n5999 = ( ~n289 & n5997 ) | ( ~n289 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6000 = n5999 ^ n2583 ^ 1'b0 ;
  assign n6001 = ~n955 & n6000 ;
  assign n5989 = n3437 & ~n3520 ;
  assign n5990 = n5989 ^ n3193 ^ 1'b0 ;
  assign n5991 = n1052 ^ n1031 ^ n570 ;
  assign n5992 = n5523 | n5991 ;
  assign n5993 = n5992 ^ n3178 ^ 1'b0 ;
  assign n5994 = n557 & n5993 ;
  assign n5995 = n5994 ^ n2315 ^ 1'b0 ;
  assign n5996 = n5990 & n5995 ;
  assign n6002 = n6001 ^ n5996 ^ 1'b0 ;
  assign n6003 = ( n2740 & n5004 ) | ( n2740 & n5930 ) | ( n5004 & n5930 ) ;
  assign n6006 = ( x22 & n2264 ) | ( x22 & n4301 ) | ( n2264 & n4301 ) ;
  assign n6004 = ( n2973 & n3535 ) | ( n2973 & n4176 ) | ( n3535 & n4176 ) ;
  assign n6005 = n6004 ^ n5354 ^ n1541 ;
  assign n6007 = n6006 ^ n6005 ^ 1'b0 ;
  assign n6008 = ( n3030 & n3185 ) | ( n3030 & ~n6007 ) | ( n3185 & ~n6007 ) ;
  assign n6009 = ( n3694 & n3979 ) | ( n3694 & ~n6008 ) | ( n3979 & ~n6008 ) ;
  assign n6010 = ( n2548 & ~n2780 ) | ( n2548 & n2916 ) | ( ~n2780 & n2916 ) ;
  assign n6017 = n306 & ~n4962 ;
  assign n6018 = n6017 ^ n2566 ^ n1728 ;
  assign n6019 = ( n2658 & ~n5981 ) | ( n2658 & n6018 ) | ( ~n5981 & n6018 ) ;
  assign n6012 = ( ~n955 & n2108 ) | ( ~n955 & n3485 ) | ( n2108 & n3485 ) ;
  assign n6013 = n5464 ^ n777 ^ 1'b0 ;
  assign n6014 = n6012 & n6013 ;
  assign n6011 = ~n1947 & n2028 ;
  assign n6015 = n6014 ^ n6011 ^ 1'b0 ;
  assign n6016 = ~n1619 & n6015 ;
  assign n6020 = n6019 ^ n6016 ^ 1'b0 ;
  assign n6021 = n874 & ~n6020 ;
  assign n6028 = x134 & n442 ;
  assign n6027 = ( n845 & n1437 ) | ( n845 & ~n1575 ) | ( n1437 & ~n1575 ) ;
  assign n6022 = x62 & n4937 ;
  assign n6023 = ~n853 & n6022 ;
  assign n6024 = ( x12 & ~n1729 ) | ( x12 & n6023 ) | ( ~n1729 & n6023 ) ;
  assign n6025 = ( ~n3316 & n3833 ) | ( ~n3316 & n6024 ) | ( n3833 & n6024 ) ;
  assign n6026 = ( n3505 & ~n4420 ) | ( n3505 & n6025 ) | ( ~n4420 & n6025 ) ;
  assign n6029 = n6028 ^ n6027 ^ n6026 ;
  assign n6030 = n5572 ^ n3390 ^ n1620 ;
  assign n6031 = n5396 ^ n1797 ^ 1'b0 ;
  assign n6032 = n3494 | n6031 ;
  assign n6033 = n2224 & ~n6032 ;
  assign n6034 = ( x212 & n6030 ) | ( x212 & n6033 ) | ( n6030 & n6033 ) ;
  assign n6035 = n2913 ^ n2360 ^ 1'b0 ;
  assign n6036 = ( ~n834 & n5888 ) | ( ~n834 & n6035 ) | ( n5888 & n6035 ) ;
  assign n6037 = n3854 ^ x65 ^ 1'b0 ;
  assign n6038 = n6037 ^ x253 ^ x96 ;
  assign n6042 = ( ~n552 & n2003 ) | ( ~n552 & n2995 ) | ( n2003 & n2995 ) ;
  assign n6043 = n6042 ^ n4139 ^ n414 ;
  assign n6040 = n3855 ^ n3337 ^ n1085 ;
  assign n6039 = n2074 | n5363 ;
  assign n6041 = n6040 ^ n6039 ^ n4919 ;
  assign n6044 = n6043 ^ n6041 ^ 1'b0 ;
  assign n6045 = n6038 & n6044 ;
  assign n6046 = ( ~n2568 & n4150 ) | ( ~n2568 & n6045 ) | ( n4150 & n6045 ) ;
  assign n6047 = ( n476 & n1331 ) | ( n476 & n1442 ) | ( n1331 & n1442 ) ;
  assign n6048 = ( x224 & n2428 ) | ( x224 & ~n6047 ) | ( n2428 & ~n6047 ) ;
  assign n6049 = ( n421 & n1184 ) | ( n421 & n3502 ) | ( n1184 & n3502 ) ;
  assign n6050 = n6048 | n6049 ;
  assign n6064 = n1139 & ~n3336 ;
  assign n6051 = n5219 ^ n1645 ^ 1'b0 ;
  assign n6052 = n947 & ~n1377 ;
  assign n6053 = n6052 ^ n4205 ^ n3986 ;
  assign n6054 = n4641 ^ n4190 ^ n3225 ;
  assign n6055 = n6054 ^ n2254 ^ 1'b0 ;
  assign n6056 = ~n6053 & n6055 ;
  assign n6059 = n488 ^ x124 ^ 1'b0 ;
  assign n6057 = n5636 ^ n3184 ^ 1'b0 ;
  assign n6058 = ~n5205 & n6057 ;
  assign n6060 = n6059 ^ n6058 ^ n2208 ;
  assign n6061 = n6056 & ~n6060 ;
  assign n6062 = n6051 & n6061 ;
  assign n6063 = n6062 ^ n4271 ^ n1960 ;
  assign n6065 = n6064 ^ n6063 ^ n698 ;
  assign n6066 = n5236 & ~n6065 ;
  assign n6067 = n5339 & n6066 ;
  assign n6069 = ( n2668 & n3048 ) | ( n2668 & n3918 ) | ( n3048 & n3918 ) ;
  assign n6068 = ( n2995 & n3661 ) | ( n2995 & n4219 ) | ( n3661 & n4219 ) ;
  assign n6070 = n6069 ^ n6068 ^ 1'b0 ;
  assign n6071 = ~n6067 & n6070 ;
  assign n6072 = x14 & n1215 ;
  assign n6073 = n3250 & n6072 ;
  assign n6074 = n6073 ^ n5118 ^ 1'b0 ;
  assign n6078 = n1722 | n2823 ;
  assign n6079 = n6078 ^ n1246 ^ 1'b0 ;
  assign n6076 = n2449 ^ n2175 ^ n2160 ;
  assign n6075 = n5195 ^ n4838 ^ n2040 ;
  assign n6077 = n6076 ^ n6075 ^ 1'b0 ;
  assign n6080 = n6079 ^ n6077 ^ 1'b0 ;
  assign n6081 = ~n6074 & n6080 ;
  assign n6087 = ( ~n2474 & n3317 ) | ( ~n2474 & n4594 ) | ( n3317 & n4594 ) ;
  assign n6083 = ( n424 & n1486 ) | ( n424 & n2326 ) | ( n1486 & n2326 ) ;
  assign n6084 = n6083 ^ n2899 ^ 1'b0 ;
  assign n6085 = ~n352 & n6084 ;
  assign n6086 = n4342 & n6085 ;
  assign n6088 = n6087 ^ n6086 ^ 1'b0 ;
  assign n6082 = n1711 & n3727 ;
  assign n6089 = n6088 ^ n6082 ^ 1'b0 ;
  assign n6090 = ~n5213 & n6089 ;
  assign n6091 = n1032 | n2318 ;
  assign n6092 = n3810 ^ n2749 ^ n1476 ;
  assign n6093 = n6092 ^ n2206 ^ n1701 ;
  assign n6094 = n1278 & ~n2802 ;
  assign n6095 = n4239 ^ n1321 ^ 1'b0 ;
  assign n6096 = ~n3037 & n6095 ;
  assign n6097 = n6094 & n6096 ;
  assign n6098 = n5919 ^ n3025 ^ 1'b0 ;
  assign n6099 = n2033 | n6098 ;
  assign n6100 = n6097 | n6099 ;
  assign n6101 = n6093 & ~n6100 ;
  assign n6102 = ( x53 & n3489 ) | ( x53 & ~n6101 ) | ( n3489 & ~n6101 ) ;
  assign n6103 = n5843 ^ n3733 ^ n1082 ;
  assign n6104 = ( n1463 & ~n3207 ) | ( n1463 & n6103 ) | ( ~n3207 & n6103 ) ;
  assign n6105 = ( n2839 & ~n3279 ) | ( n2839 & n3658 ) | ( ~n3279 & n3658 ) ;
  assign n6106 = n3037 ^ n2688 ^ 1'b0 ;
  assign n6107 = ( n6104 & n6105 ) | ( n6104 & ~n6106 ) | ( n6105 & ~n6106 ) ;
  assign n6108 = n1789 | n2643 ;
  assign n6109 = n6108 ^ n5832 ^ 1'b0 ;
  assign n6110 = n6109 ^ n4623 ^ n1741 ;
  assign n6111 = n6110 ^ n3422 ^ n2550 ;
  assign n6112 = ~n2865 & n6111 ;
  assign n6113 = ( n861 & n3504 ) | ( n861 & ~n5846 ) | ( n3504 & ~n5846 ) ;
  assign n6114 = ( ~n1811 & n2994 ) | ( ~n1811 & n6113 ) | ( n2994 & n6113 ) ;
  assign n6118 = n3995 ^ n3139 ^ 1'b0 ;
  assign n6119 = ~n5825 & n6118 ;
  assign n6115 = n1928 & ~n3065 ;
  assign n6116 = n6115 ^ n2175 ^ 1'b0 ;
  assign n6117 = n6116 ^ n4641 ^ n3404 ;
  assign n6120 = n6119 ^ n6117 ^ n2949 ;
  assign n6121 = n6120 ^ n5451 ^ 1'b0 ;
  assign n6122 = n6114 & ~n6121 ;
  assign n6123 = ( n2707 & n5718 ) | ( n2707 & n5758 ) | ( n5718 & n5758 ) ;
  assign n6124 = n1726 | n4881 ;
  assign n6125 = n6124 ^ n3938 ^ n627 ;
  assign n6126 = ( ~n275 & n1256 ) | ( ~n275 & n1750 ) | ( n1256 & n1750 ) ;
  assign n6127 = n6126 ^ n5417 ^ n2103 ;
  assign n6128 = n6127 ^ n2654 ^ 1'b0 ;
  assign n6129 = n6125 | n6128 ;
  assign n6130 = n5998 ^ n2083 ^ 1'b0 ;
  assign n6131 = n3271 ^ n2393 ^ 1'b0 ;
  assign n6135 = n3638 ^ n3525 ^ n2841 ;
  assign n6132 = n2966 ^ n948 ^ x116 ;
  assign n6133 = ~n5381 & n6132 ;
  assign n6134 = n5252 & n6133 ;
  assign n6136 = n6135 ^ n6134 ^ n1830 ;
  assign n6137 = n3910 ^ n1906 ^ n1232 ;
  assign n6138 = n4384 & n6137 ;
  assign n6139 = ( n2129 & n4876 ) | ( n2129 & ~n5360 ) | ( n4876 & ~n5360 ) ;
  assign n6140 = n6139 ^ n2133 ^ 1'b0 ;
  assign n6141 = n1117 & n6140 ;
  assign n6145 = n478 ^ x218 ^ 1'b0 ;
  assign n6146 = n1497 | n6145 ;
  assign n6147 = n754 & ~n3185 ;
  assign n6148 = n6147 ^ n1349 ^ 1'b0 ;
  assign n6149 = ( ~n1122 & n6146 ) | ( ~n1122 & n6148 ) | ( n6146 & n6148 ) ;
  assign n6143 = ( n422 & ~n1151 ) | ( n422 & n1760 ) | ( ~n1151 & n1760 ) ;
  assign n6142 = ( n340 & ~n381 ) | ( n340 & n3937 ) | ( ~n381 & n3937 ) ;
  assign n6144 = n6143 ^ n6142 ^ n492 ;
  assign n6150 = n6149 ^ n6144 ^ n5034 ;
  assign n6151 = n2135 ^ n932 ^ n312 ;
  assign n6152 = n6151 ^ n6037 ^ 1'b0 ;
  assign n6153 = n427 & ~n6152 ;
  assign n6154 = x182 & ~n2408 ;
  assign n6155 = ~n1115 & n6154 ;
  assign n6156 = n555 & n4623 ;
  assign n6157 = ~n2280 & n6156 ;
  assign n6158 = n6157 ^ n5016 ^ n921 ;
  assign n6159 = ( n3881 & n6151 ) | ( n3881 & n6158 ) | ( n6151 & n6158 ) ;
  assign n6160 = ( n3795 & n6155 ) | ( n3795 & ~n6159 ) | ( n6155 & ~n6159 ) ;
  assign n6161 = n3606 ^ n1777 ^ n1201 ;
  assign n6162 = ( ~n2547 & n5697 ) | ( ~n2547 & n5892 ) | ( n5697 & n5892 ) ;
  assign n6163 = n6162 ^ n3241 ^ 1'b0 ;
  assign n6164 = n2367 & ~n6163 ;
  assign n6165 = ~n5710 & n6164 ;
  assign n6166 = ~n6161 & n6165 ;
  assign n6167 = n2913 ^ n1926 ^ n1140 ;
  assign n6168 = n6167 ^ n5373 ^ n787 ;
  assign n6171 = ( n768 & ~n907 ) | ( n768 & n3268 ) | ( ~n907 & n3268 ) ;
  assign n6172 = n6171 ^ n4181 ^ n2399 ;
  assign n6170 = n3795 ^ n1217 ^ n1079 ;
  assign n6169 = ( x149 & n969 ) | ( x149 & ~n2733 ) | ( n969 & ~n2733 ) ;
  assign n6173 = n6172 ^ n6170 ^ n6169 ;
  assign n6177 = n1224 ^ n423 ^ 1'b0 ;
  assign n6174 = n1729 ^ n658 ^ 1'b0 ;
  assign n6175 = n1768 | n6174 ;
  assign n6176 = n6175 ^ n2068 ^ n1589 ;
  assign n6178 = n6177 ^ n6176 ^ n6039 ;
  assign n6179 = n3381 ^ n2581 ^ n1481 ;
  assign n6180 = n5538 & n5924 ;
  assign n6181 = n6179 & n6180 ;
  assign n6184 = n3309 ^ n3018 ^ n484 ;
  assign n6182 = ( x145 & n849 ) | ( x145 & n1225 ) | ( n849 & n1225 ) ;
  assign n6183 = n284 & n6182 ;
  assign n6185 = n6184 ^ n6183 ^ 1'b0 ;
  assign n6187 = ( x11 & n2450 ) | ( x11 & n2553 ) | ( n2450 & n2553 ) ;
  assign n6188 = n6187 ^ n2860 ^ 1'b0 ;
  assign n6186 = ( ~n2006 & n5032 ) | ( ~n2006 & n5676 ) | ( n5032 & n5676 ) ;
  assign n6189 = n6188 ^ n6186 ^ 1'b0 ;
  assign n6191 = ( ~x67 & n2729 ) | ( ~x67 & n5843 ) | ( n2729 & n5843 ) ;
  assign n6192 = n6191 ^ n1652 ^ 1'b0 ;
  assign n6193 = ~n1175 & n6192 ;
  assign n6190 = n2224 ^ n1358 ^ 1'b0 ;
  assign n6194 = n6193 ^ n6190 ^ 1'b0 ;
  assign n6195 = n5635 & ~n6194 ;
  assign n6196 = n6195 ^ n5944 ^ 1'b0 ;
  assign n6197 = n4012 ^ x201 ^ 1'b0 ;
  assign n6205 = n4954 ^ n4022 ^ n2406 ;
  assign n6201 = n535 | n758 ;
  assign n6202 = n2033 & ~n6201 ;
  assign n6203 = n6202 ^ n4267 ^ 1'b0 ;
  assign n6204 = n4583 | n6203 ;
  assign n6198 = n2069 ^ n1738 ^ 1'b0 ;
  assign n6199 = n1555 & ~n6198 ;
  assign n6200 = ~n5051 & n6199 ;
  assign n6206 = n6205 ^ n6204 ^ n6200 ;
  assign n6207 = ~n6197 & n6206 ;
  assign n6208 = ( ~n744 & n1677 ) | ( ~n744 & n6207 ) | ( n1677 & n6207 ) ;
  assign n6209 = ( x98 & n1909 ) | ( x98 & ~n6208 ) | ( n1909 & ~n6208 ) ;
  assign n6210 = n2366 & n3547 ;
  assign n6211 = ( x48 & n2615 ) | ( x48 & n3330 ) | ( n2615 & n3330 ) ;
  assign n6212 = n6211 ^ n4510 ^ x50 ;
  assign n6213 = n6212 ^ n5444 ^ n2854 ;
  assign n6214 = ( n1414 & ~n4166 ) | ( n1414 & n6213 ) | ( ~n4166 & n6213 ) ;
  assign n6215 = n1771 & ~n5757 ;
  assign n6216 = n6214 & n6215 ;
  assign n6217 = ( ~n707 & n1655 ) | ( ~n707 & n1942 ) | ( n1655 & n1942 ) ;
  assign n6218 = n6217 ^ n1381 ^ 1'b0 ;
  assign n6219 = n5662 & n6218 ;
  assign n6220 = n6219 ^ n2456 ^ 1'b0 ;
  assign n6222 = n3253 ^ n1950 ^ x233 ;
  assign n6221 = ~n694 & n3945 ;
  assign n6223 = n6222 ^ n6221 ^ n5255 ;
  assign n6224 = x111 & n1085 ;
  assign n6225 = n6223 & ~n6224 ;
  assign n6226 = n6225 ^ n3909 ^ 1'b0 ;
  assign n6227 = n6226 ^ n536 ^ n289 ;
  assign n6228 = n1909 ^ n455 ^ 1'b0 ;
  assign n6229 = n719 & n6228 ;
  assign n6230 = n6229 ^ n935 ^ 1'b0 ;
  assign n6232 = ( n2072 & n4072 ) | ( n2072 & n5496 ) | ( n4072 & n5496 ) ;
  assign n6233 = ~n5525 & n6232 ;
  assign n6234 = ~n3525 & n6233 ;
  assign n6231 = n2899 ^ n2512 ^ n1761 ;
  assign n6235 = n6234 ^ n6231 ^ n2213 ;
  assign n6236 = ( n1090 & ~n1164 ) | ( n1090 & n6235 ) | ( ~n1164 & n6235 ) ;
  assign n6237 = n1463 & ~n2468 ;
  assign n6238 = n2558 & ~n4487 ;
  assign n6239 = n6238 ^ n1343 ^ x15 ;
  assign n6240 = ( n715 & n1632 ) | ( n715 & n4077 ) | ( n1632 & n4077 ) ;
  assign n6241 = ~n735 & n6240 ;
  assign n6242 = n5367 ^ n4787 ^ n3220 ;
  assign n6243 = n6241 | n6242 ;
  assign n6244 = n6243 ^ n3323 ^ 1'b0 ;
  assign n6245 = x24 & n3005 ;
  assign n6246 = ( n1309 & n2158 ) | ( n1309 & n6245 ) | ( n2158 & n6245 ) ;
  assign n6247 = n2188 & ~n3629 ;
  assign n6248 = ~x180 & n6247 ;
  assign n6249 = ( x35 & n3738 ) | ( x35 & n6248 ) | ( n3738 & n6248 ) ;
  assign n6250 = ( ~n298 & n6246 ) | ( ~n298 & n6249 ) | ( n6246 & n6249 ) ;
  assign n6251 = n4440 ^ n2427 ^ n1299 ;
  assign n6252 = n410 & n2122 ;
  assign n6253 = ~n3119 & n6252 ;
  assign n6254 = n6253 ^ n3251 ^ 1'b0 ;
  assign n6255 = ~n6251 & n6254 ;
  assign n6261 = n4983 ^ n3781 ^ n2076 ;
  assign n6259 = n2058 ^ x130 ^ 1'b0 ;
  assign n6256 = n3191 ^ n2142 ^ 1'b0 ;
  assign n6257 = n1480 & n6256 ;
  assign n6258 = ~n4693 & n6257 ;
  assign n6260 = n6259 ^ n6258 ^ 1'b0 ;
  assign n6262 = n6261 ^ n6260 ^ n3938 ;
  assign n6263 = ( x234 & n717 ) | ( x234 & n2736 ) | ( n717 & n2736 ) ;
  assign n6264 = n5947 & n6263 ;
  assign n6270 = ~n545 & n3326 ;
  assign n6271 = n6270 ^ n5051 ^ n2115 ;
  assign n6268 = n1677 ^ n1653 ^ n1487 ;
  assign n6269 = n6268 ^ n6257 ^ 1'b0 ;
  assign n6272 = n6271 ^ n6269 ^ n4859 ;
  assign n6265 = n1645 & n3244 ;
  assign n6266 = n6265 ^ n2292 ^ 1'b0 ;
  assign n6267 = n3384 | n6266 ;
  assign n6273 = n6272 ^ n6267 ^ n5071 ;
  assign n6274 = n6264 | n6273 ;
  assign n6275 = n6274 ^ n3487 ^ 1'b0 ;
  assign n6276 = n4876 | n6275 ;
  assign n6277 = n4790 | n6276 ;
  assign n6280 = n1980 ^ n1107 ^ 1'b0 ;
  assign n6278 = n4971 & ~n5066 ;
  assign n6279 = n6278 ^ n4623 ^ 1'b0 ;
  assign n6281 = n6280 ^ n6279 ^ n1405 ;
  assign n6282 = n6281 ^ n6028 ^ n5442 ;
  assign n6283 = n3885 & ~n6282 ;
  assign n6284 = ( x96 & ~n3550 ) | ( x96 & n4417 ) | ( ~n3550 & n4417 ) ;
  assign n6285 = n1225 | n4271 ;
  assign n6286 = n4197 & ~n6285 ;
  assign n6287 = ( n4750 & n6284 ) | ( n4750 & n6286 ) | ( n6284 & n6286 ) ;
  assign n6293 = ( x63 & ~x214 ) | ( x63 & n619 ) | ( ~x214 & n619 ) ;
  assign n6294 = ( n1536 & n3381 ) | ( n1536 & ~n6293 ) | ( n3381 & ~n6293 ) ;
  assign n6290 = ( n2339 & n2454 ) | ( n2339 & ~n3395 ) | ( n2454 & ~n3395 ) ;
  assign n6291 = n6290 ^ n2871 ^ 1'b0 ;
  assign n6292 = x11 & n6291 ;
  assign n6288 = n5144 ^ n2509 ^ 1'b0 ;
  assign n6289 = n4077 & ~n6288 ;
  assign n6295 = n6294 ^ n6292 ^ n6289 ;
  assign n6296 = n6295 ^ n1077 ^ x226 ;
  assign n6297 = ~n6287 & n6296 ;
  assign n6298 = n6297 ^ n5687 ^ 1'b0 ;
  assign n6299 = n5146 ^ n1565 ^ n482 ;
  assign n6300 = n6299 ^ n3351 ^ n2608 ;
  assign n6301 = n6300 ^ x49 ^ 1'b0 ;
  assign n6302 = n5742 ^ n2399 ^ n1477 ;
  assign n6303 = n1463 & n5857 ;
  assign n6304 = n6303 ^ n3399 ^ 1'b0 ;
  assign n6305 = n5825 ^ n321 ^ n288 ;
  assign n6308 = n2625 & n4180 ;
  assign n6309 = ~n2228 & n6308 ;
  assign n6306 = ( ~n1395 & n3385 ) | ( ~n1395 & n4022 ) | ( n3385 & n4022 ) ;
  assign n6307 = n6306 ^ n3068 ^ n2555 ;
  assign n6310 = n6309 ^ n6307 ^ n732 ;
  assign n6311 = ( ~n2691 & n6305 ) | ( ~n2691 & n6310 ) | ( n6305 & n6310 ) ;
  assign n6312 = n6311 ^ n3989 ^ n2729 ;
  assign n6318 = ( ~n452 & n802 ) | ( ~n452 & n1686 ) | ( n802 & n1686 ) ;
  assign n6319 = n3045 ^ n1650 ^ 1'b0 ;
  assign n6320 = n6318 | n6319 ;
  assign n6315 = n1475 & ~n2133 ;
  assign n6316 = ~x210 & n6315 ;
  assign n6313 = n5856 ^ n1713 ^ 1'b0 ;
  assign n6314 = n3061 | n6313 ;
  assign n6317 = n6316 ^ n6314 ^ n1948 ;
  assign n6321 = n6320 ^ n6317 ^ n2227 ;
  assign n6322 = n357 & n532 ;
  assign n6323 = n6322 ^ n917 ^ 1'b0 ;
  assign n6324 = n2214 & n5533 ;
  assign n6325 = n5144 ^ n2995 ^ 1'b0 ;
  assign n6326 = ( n6323 & ~n6324 ) | ( n6323 & n6325 ) | ( ~n6324 & n6325 ) ;
  assign n6327 = ( n1231 & n1602 ) | ( n1231 & n5110 ) | ( n1602 & n5110 ) ;
  assign n6328 = n2085 ^ n1743 ^ n1102 ;
  assign n6329 = n4441 ^ n1655 ^ x106 ;
  assign n6330 = n6329 ^ n852 ^ n326 ;
  assign n6331 = ( n930 & n1418 ) | ( n930 & n2842 ) | ( n1418 & n2842 ) ;
  assign n6332 = n1954 ^ n266 ^ 1'b0 ;
  assign n6333 = n3025 & ~n6332 ;
  assign n6334 = ( n2510 & ~n6331 ) | ( n2510 & n6333 ) | ( ~n6331 & n6333 ) ;
  assign n6335 = n5764 ^ n5212 ^ 1'b0 ;
  assign n6336 = n6334 & n6335 ;
  assign n6337 = ( n6328 & ~n6330 ) | ( n6328 & n6336 ) | ( ~n6330 & n6336 ) ;
  assign n6338 = n3266 ^ n3167 ^ n2774 ;
  assign n6339 = n6338 ^ n4817 ^ n2486 ;
  assign n6342 = n963 ^ n610 ^ 1'b0 ;
  assign n6340 = n3244 ^ n1527 ^ 1'b0 ;
  assign n6341 = n6340 ^ n913 ^ 1'b0 ;
  assign n6343 = n6342 ^ n6341 ^ n1452 ;
  assign n6344 = ( x85 & n1925 ) | ( x85 & n3528 ) | ( n1925 & n3528 ) ;
  assign n6345 = n6344 ^ n5941 ^ n4743 ;
  assign n6346 = n5815 ^ n4834 ^ n1637 ;
  assign n6347 = ( n1655 & n3415 ) | ( n1655 & n6346 ) | ( n3415 & n6346 ) ;
  assign n6348 = ( n1682 & ~n5726 ) | ( n1682 & n6132 ) | ( ~n5726 & n6132 ) ;
  assign n6349 = n5435 ^ n5253 ^ x62 ;
  assign n6350 = n6349 ^ n5307 ^ 1'b0 ;
  assign n6351 = n6348 & ~n6350 ;
  assign n6354 = x23 & ~n1783 ;
  assign n6355 = ~n1928 & n6354 ;
  assign n6352 = n3638 ^ n1958 ^ n1599 ;
  assign n6353 = ~n620 & n6352 ;
  assign n6356 = n6355 ^ n6353 ^ 1'b0 ;
  assign n6357 = n2244 | n6356 ;
  assign n6358 = n378 & ~n1906 ;
  assign n6359 = n6358 ^ n3247 ^ 1'b0 ;
  assign n6360 = n6359 ^ n3098 ^ 1'b0 ;
  assign n6361 = ~n5873 & n6360 ;
  assign n6362 = ~n289 & n1477 ;
  assign n6363 = ( x2 & ~n903 ) | ( x2 & n6362 ) | ( ~n903 & n6362 ) ;
  assign n6364 = n6363 ^ n1623 ^ n1595 ;
  assign n6365 = ( n2244 & n3053 ) | ( n2244 & ~n6364 ) | ( n3053 & ~n6364 ) ;
  assign n6366 = ( n2795 & n6361 ) | ( n2795 & n6365 ) | ( n6361 & n6365 ) ;
  assign n6367 = ~n2569 & n5997 ;
  assign n6368 = n2728 & n6367 ;
  assign n6369 = n1421 ^ n592 ^ 1'b0 ;
  assign n6370 = n1264 | n6369 ;
  assign n6371 = x220 & ~n6370 ;
  assign n6372 = n6368 & n6371 ;
  assign n6373 = n2550 & ~n6372 ;
  assign n6374 = n6200 & n6373 ;
  assign n6375 = n6374 ^ n484 ^ 1'b0 ;
  assign n6376 = n4603 ^ n2373 ^ n1394 ;
  assign n6377 = ( ~n4101 & n5289 ) | ( ~n4101 & n6376 ) | ( n5289 & n6376 ) ;
  assign n6378 = n6377 ^ n6116 ^ 1'b0 ;
  assign n6379 = n6378 ^ n4625 ^ n3733 ;
  assign n6380 = ( n783 & n2072 ) | ( n783 & n6112 ) | ( n2072 & n6112 ) ;
  assign n6381 = n1709 ^ n865 ^ 1'b0 ;
  assign n6382 = n3397 ^ n697 ^ 1'b0 ;
  assign n6383 = n856 & ~n6382 ;
  assign n6385 = n1636 & ~n2034 ;
  assign n6384 = n665 & n5603 ;
  assign n6386 = n6385 ^ n6384 ^ 1'b0 ;
  assign n6387 = ( n6381 & n6383 ) | ( n6381 & ~n6386 ) | ( n6383 & ~n6386 ) ;
  assign n6388 = ( x109 & n5343 ) | ( x109 & n6387 ) | ( n5343 & n6387 ) ;
  assign n6389 = n6135 ^ n5751 ^ 1'b0 ;
  assign n6390 = n5872 ^ n5255 ^ 1'b0 ;
  assign n6391 = ~n6389 & n6390 ;
  assign n6393 = n1131 ^ n799 ^ 1'b0 ;
  assign n6394 = ~n2875 & n6393 ;
  assign n6392 = ( n1188 & ~n1817 ) | ( n1188 & n2589 ) | ( ~n1817 & n2589 ) ;
  assign n6395 = n6394 ^ n6392 ^ n302 ;
  assign n6396 = ( n1938 & ~n3106 ) | ( n1938 & n6395 ) | ( ~n3106 & n6395 ) ;
  assign n6398 = n4955 ^ n3099 ^ n874 ;
  assign n6399 = n6398 ^ n5222 ^ n1360 ;
  assign n6397 = n1760 | n4042 ;
  assign n6400 = n6399 ^ n6397 ^ n5890 ;
  assign n6401 = ( ~x164 & n1151 ) | ( ~x164 & n1882 ) | ( n1151 & n1882 ) ;
  assign n6404 = n3959 ^ n2767 ^ n412 ;
  assign n6402 = ( ~x18 & x235 ) | ( ~x18 & n5196 ) | ( x235 & n5196 ) ;
  assign n6403 = n6402 ^ n3947 ^ n614 ;
  assign n6405 = n6404 ^ n6403 ^ n1561 ;
  assign n6406 = n6401 & ~n6405 ;
  assign n6407 = n6406 ^ n1904 ^ 1'b0 ;
  assign n6409 = ~n1433 & n3301 ;
  assign n6408 = ~n325 & n2815 ;
  assign n6410 = n6409 ^ n6408 ^ n342 ;
  assign n6411 = n6410 ^ n1949 ^ 1'b0 ;
  assign n6412 = n5890 ^ n2311 ^ 1'b0 ;
  assign n6413 = n2998 | n6412 ;
  assign n6414 = n6413 ^ n4003 ^ n733 ;
  assign n6415 = n6414 ^ n2952 ^ 1'b0 ;
  assign n6416 = n2126 & n3143 ;
  assign n6417 = n1223 & n6416 ;
  assign n6418 = n2066 ^ n1196 ^ 1'b0 ;
  assign n6419 = n2910 | n6418 ;
  assign n6420 = n843 | n2310 ;
  assign n6421 = n2389 | n6420 ;
  assign n6422 = n3463 & ~n6421 ;
  assign n6423 = n2754 | n6422 ;
  assign n6424 = ( n823 & n6419 ) | ( n823 & n6423 ) | ( n6419 & n6423 ) ;
  assign n6425 = ( n1440 & ~n6417 ) | ( n1440 & n6424 ) | ( ~n6417 & n6424 ) ;
  assign n6426 = n5393 ^ n1628 ^ 1'b0 ;
  assign n6427 = n3977 & ~n6426 ;
  assign n6428 = ( n2892 & n5665 ) | ( n2892 & n6232 ) | ( n5665 & n6232 ) ;
  assign n6429 = x221 & n2105 ;
  assign n6430 = n6429 ^ n2750 ^ n1609 ;
  assign n6431 = n6430 ^ n5339 ^ n735 ;
  assign n6432 = n2540 & ~n4291 ;
  assign n6433 = n1025 & n6432 ;
  assign n6434 = n6433 ^ n4942 ^ n398 ;
  assign n6435 = n4773 ^ n3038 ^ 1'b0 ;
  assign n6436 = ( n418 & ~n1080 ) | ( n418 & n2273 ) | ( ~n1080 & n2273 ) ;
  assign n6437 = n320 | n2051 ;
  assign n6438 = n6436 | n6437 ;
  assign n6439 = n2549 | n6438 ;
  assign n6440 = n6435 & n6439 ;
  assign n6441 = n6434 & n6440 ;
  assign n6442 = ( n1260 & n3866 ) | ( n1260 & n6027 ) | ( n3866 & n6027 ) ;
  assign n6443 = n6135 ^ n2367 ^ 1'b0 ;
  assign n6444 = n6442 | n6443 ;
  assign n6445 = ( ~n2360 & n3906 ) | ( ~n2360 & n6333 ) | ( n3906 & n6333 ) ;
  assign n6446 = n2154 ^ n1807 ^ 1'b0 ;
  assign n6447 = n5832 & ~n6446 ;
  assign n6448 = ( ~n683 & n2286 ) | ( ~n683 & n6447 ) | ( n2286 & n6447 ) ;
  assign n6449 = n6445 & ~n6448 ;
  assign n6450 = n6449 ^ n1019 ^ 1'b0 ;
  assign n6451 = n6444 & n6450 ;
  assign n6452 = n4507 ^ x105 ^ 1'b0 ;
  assign n6453 = n963 ^ n837 ^ 1'b0 ;
  assign n6454 = n2408 & n4205 ;
  assign n6455 = n6454 ^ n1775 ^ 1'b0 ;
  assign n6456 = ( n4538 & n6453 ) | ( n4538 & ~n6455 ) | ( n6453 & ~n6455 ) ;
  assign n6457 = n6026 ^ n5015 ^ n1486 ;
  assign n6458 = ( n504 & n775 ) | ( n504 & n5550 ) | ( n775 & n5550 ) ;
  assign n6459 = n1842 & ~n6458 ;
  assign n6465 = n4636 ^ n2677 ^ n1372 ;
  assign n6466 = ( n4247 & ~n5800 ) | ( n4247 & n6465 ) | ( ~n5800 & n6465 ) ;
  assign n6461 = ( x179 & n4096 ) | ( x179 & n6110 ) | ( n4096 & n6110 ) ;
  assign n6460 = x168 & n3313 ;
  assign n6462 = n6461 ^ n6460 ^ 1'b0 ;
  assign n6463 = n1091 & ~n6462 ;
  assign n6464 = n6463 ^ n925 ^ 1'b0 ;
  assign n6467 = n6466 ^ n6464 ^ n2949 ;
  assign n6468 = ( ~n1920 & n4572 ) | ( ~n1920 & n6323 ) | ( n4572 & n6323 ) ;
  assign n6469 = n4271 ^ x33 ^ 1'b0 ;
  assign n6470 = n4794 ^ n1682 ^ n1461 ;
  assign n6471 = n6469 | n6470 ;
  assign n6472 = n1479 | n6471 ;
  assign n6473 = n6472 ^ n1961 ^ n381 ;
  assign n6474 = n5662 ^ n552 ^ 1'b0 ;
  assign n6475 = n1020 & ~n6474 ;
  assign n6476 = n6475 ^ n3923 ^ n3502 ;
  assign n6477 = n6202 ^ n2540 ^ 1'b0 ;
  assign n6478 = ( n1405 & ~n3253 ) | ( n1405 & n6477 ) | ( ~n3253 & n6477 ) ;
  assign n6479 = n2770 | n3484 ;
  assign n6480 = ( n1448 & n2445 ) | ( n1448 & ~n2462 ) | ( n2445 & ~n2462 ) ;
  assign n6481 = n2174 ^ n1665 ^ x140 ;
  assign n6482 = ( n3938 & n6132 ) | ( n3938 & n6481 ) | ( n6132 & n6481 ) ;
  assign n6483 = n6021 & ~n6482 ;
  assign n6484 = n6480 & n6483 ;
  assign n6485 = n552 & ~n666 ;
  assign n6486 = n6485 ^ n1817 ^ 1'b0 ;
  assign n6487 = n2169 | n6486 ;
  assign n6488 = n978 | n6487 ;
  assign n6489 = ( n1578 & ~n2644 ) | ( n1578 & n6488 ) | ( ~n2644 & n6488 ) ;
  assign n6490 = ( ~n4952 & n6052 ) | ( ~n4952 & n6489 ) | ( n6052 & n6489 ) ;
  assign n6491 = ( x85 & x163 ) | ( x85 & ~n995 ) | ( x163 & ~n995 ) ;
  assign n6492 = n938 & ~n2309 ;
  assign n6493 = n6492 ^ x91 ^ 1'b0 ;
  assign n6494 = ( ~n6490 & n6491 ) | ( ~n6490 & n6493 ) | ( n6491 & n6493 ) ;
  assign n6495 = ( n1100 & ~n3693 ) | ( n1100 & n6494 ) | ( ~n3693 & n6494 ) ;
  assign n6496 = ( ~n1368 & n4657 ) | ( ~n1368 & n6495 ) | ( n4657 & n6495 ) ;
  assign n6497 = ( n3165 & ~n3892 ) | ( n3165 & n5500 ) | ( ~n3892 & n5500 ) ;
  assign n6498 = n6497 ^ n989 ^ 1'b0 ;
  assign n6499 = n6498 ^ n3288 ^ n2059 ;
  assign n6504 = x42 & n1001 ;
  assign n6505 = ~n1845 & n6504 ;
  assign n6507 = n4291 ^ n1417 ^ 1'b0 ;
  assign n6508 = n1695 & ~n6507 ;
  assign n6506 = n1510 & n3753 ;
  assign n6509 = n6508 ^ n6506 ^ 1'b0 ;
  assign n6510 = n508 ^ n431 ^ 1'b0 ;
  assign n6511 = n6509 & ~n6510 ;
  assign n6512 = ( n538 & ~n6505 ) | ( n538 & n6511 ) | ( ~n6505 & n6511 ) ;
  assign n6500 = n1655 ^ n683 ^ 1'b0 ;
  assign n6501 = n6500 ^ n693 ^ x113 ;
  assign n6502 = n4025 ^ n3911 ^ 1'b0 ;
  assign n6503 = ~n6501 & n6502 ;
  assign n6513 = n6512 ^ n6503 ^ 1'b0 ;
  assign n6519 = n3441 ^ n1394 ^ 1'b0 ;
  assign n6520 = ~n486 & n6519 ;
  assign n6521 = ( n405 & n5556 ) | ( n405 & n6520 ) | ( n5556 & n6520 ) ;
  assign n6514 = n821 | n4901 ;
  assign n6515 = n4000 | n6514 ;
  assign n6516 = n6515 ^ n4820 ^ n4054 ;
  assign n6517 = n6516 ^ n3445 ^ n2508 ;
  assign n6518 = ( n1954 & n2094 ) | ( n1954 & n6517 ) | ( n2094 & n6517 ) ;
  assign n6522 = n6521 ^ n6518 ^ 1'b0 ;
  assign n6523 = n3468 | n6522 ;
  assign n6524 = ( n275 & ~n3635 ) | ( n275 & n4033 ) | ( ~n3635 & n4033 ) ;
  assign n6525 = n6524 ^ n4420 ^ 1'b0 ;
  assign n6533 = ( n641 & n2124 ) | ( n641 & ~n4940 ) | ( n2124 & ~n4940 ) ;
  assign n6534 = n1020 & ~n2348 ;
  assign n6535 = n6533 & n6534 ;
  assign n6529 = ( n406 & ~n3303 ) | ( n406 & n4590 ) | ( ~n3303 & n4590 ) ;
  assign n6530 = n6529 ^ n2638 ^ 1'b0 ;
  assign n6531 = n1355 | n6530 ;
  assign n6526 = x228 & ~n1663 ;
  assign n6527 = n6526 ^ n1695 ^ 1'b0 ;
  assign n6528 = n6527 ^ n2849 ^ n2728 ;
  assign n6532 = n6531 ^ n6528 ^ n5571 ;
  assign n6536 = n6535 ^ n6532 ^ 1'b0 ;
  assign n6537 = n3213 & n6536 ;
  assign n6538 = n3835 ^ n547 ^ 1'b0 ;
  assign n6563 = n3463 ^ n1738 ^ 1'b0 ;
  assign n6564 = n5719 | n6563 ;
  assign n6550 = n1866 ^ n1819 ^ n1656 ;
  assign n6551 = n801 & ~n6550 ;
  assign n6552 = n6551 ^ n1074 ^ 1'b0 ;
  assign n6553 = n1770 & n6552 ;
  assign n6554 = n2388 & n6553 ;
  assign n6555 = n4291 ^ n1360 ^ 1'b0 ;
  assign n6556 = n2725 & ~n6555 ;
  assign n6557 = ( n765 & n1746 ) | ( n765 & ~n2539 ) | ( n1746 & ~n2539 ) ;
  assign n6558 = ( n458 & n1080 ) | ( n458 & ~n6557 ) | ( n1080 & ~n6557 ) ;
  assign n6559 = ~n799 & n5965 ;
  assign n6560 = n6558 & n6559 ;
  assign n6561 = ( n5292 & n6556 ) | ( n5292 & ~n6560 ) | ( n6556 & ~n6560 ) ;
  assign n6562 = ~n6554 & n6561 ;
  assign n6565 = n6564 ^ n6562 ^ 1'b0 ;
  assign n6539 = n522 & n2432 ;
  assign n6540 = ~n438 & n6539 ;
  assign n6541 = n6540 ^ n725 ^ n496 ;
  assign n6542 = n1863 & ~n3986 ;
  assign n6543 = n6542 ^ n1290 ^ 1'b0 ;
  assign n6544 = n1023 ^ n904 ^ 1'b0 ;
  assign n6545 = ( n6541 & ~n6543 ) | ( n6541 & n6544 ) | ( ~n6543 & n6544 ) ;
  assign n6546 = x234 & ~n2360 ;
  assign n6547 = n6546 ^ n4518 ^ n971 ;
  assign n6548 = n6547 ^ n4812 ^ n3963 ;
  assign n6549 = n6545 | n6548 ;
  assign n6566 = n6565 ^ n6549 ^ 1'b0 ;
  assign n6567 = n3146 & ~n6029 ;
  assign n6568 = ~n1588 & n6567 ;
  assign n6569 = n631 & n6568 ;
  assign n6570 = n418 & ~n6569 ;
  assign n6571 = ~n2360 & n6570 ;
  assign n6572 = ( n2160 & ~n2746 ) | ( n2160 & n6541 ) | ( ~n2746 & n6541 ) ;
  assign n6573 = n2615 & n5918 ;
  assign n6574 = n4196 ^ n1882 ^ 1'b0 ;
  assign n6575 = n4086 & n6574 ;
  assign n6576 = n6575 ^ n3780 ^ n2544 ;
  assign n6577 = ( ~n1663 & n2807 ) | ( ~n1663 & n4135 ) | ( n2807 & n4135 ) ;
  assign n6578 = n3196 ^ n1320 ^ x60 ;
  assign n6579 = ( n1295 & ~n1610 ) | ( n1295 & n6578 ) | ( ~n1610 & n6578 ) ;
  assign n6584 = ( ~n563 & n3061 ) | ( ~n563 & n3575 ) | ( n3061 & n3575 ) ;
  assign n6582 = ( ~n333 & n1238 ) | ( ~n333 & n3501 ) | ( n1238 & n3501 ) ;
  assign n6580 = n3134 ^ n787 ^ 1'b0 ;
  assign n6581 = n6408 & ~n6580 ;
  assign n6583 = n6582 ^ n6581 ^ n5046 ;
  assign n6585 = n6584 ^ n6583 ^ n2843 ;
  assign n6586 = ( n6577 & ~n6579 ) | ( n6577 & n6585 ) | ( ~n6579 & n6585 ) ;
  assign n6587 = ( n283 & ~n334 ) | ( n283 & n3599 ) | ( ~n334 & n3599 ) ;
  assign n6588 = n1147 & n3181 ;
  assign n6589 = n4341 & n6588 ;
  assign n6590 = n3336 ^ n470 ^ n356 ;
  assign n6591 = ( ~x88 & n1955 ) | ( ~x88 & n6052 ) | ( n1955 & n6052 ) ;
  assign n6592 = ( ~n4586 & n6590 ) | ( ~n4586 & n6591 ) | ( n6590 & n6591 ) ;
  assign n6593 = ( n1822 & n2410 ) | ( n1822 & ~n4340 ) | ( n2410 & ~n4340 ) ;
  assign n6594 = n1668 & ~n2471 ;
  assign n6595 = ( n4919 & n6593 ) | ( n4919 & ~n6594 ) | ( n6593 & ~n6594 ) ;
  assign n6596 = n3628 ^ x31 ^ 1'b0 ;
  assign n6597 = ~n3454 & n6596 ;
  assign n6598 = ~n3056 & n6597 ;
  assign n6599 = n2477 ^ n1518 ^ 1'b0 ;
  assign n6600 = ( ~n4397 & n5021 ) | ( ~n4397 & n6599 ) | ( n5021 & n6599 ) ;
  assign n6601 = ( n3304 & n4240 ) | ( n3304 & n4924 ) | ( n4240 & n4924 ) ;
  assign n6602 = ( n356 & n2105 ) | ( n356 & ~n2823 ) | ( n2105 & ~n2823 ) ;
  assign n6603 = ( n5991 & ~n6601 ) | ( n5991 & n6602 ) | ( ~n6601 & n6602 ) ;
  assign n6604 = n6603 ^ n5792 ^ n3862 ;
  assign n6613 = ( ~n633 & n1650 ) | ( ~n633 & n3414 ) | ( n1650 & n3414 ) ;
  assign n6612 = ( ~x91 & n378 ) | ( ~x91 & n905 ) | ( n378 & n905 ) ;
  assign n6614 = n6613 ^ n6612 ^ n672 ;
  assign n6605 = n2122 ^ n1828 ^ 1'b0 ;
  assign n6606 = ~n1927 & n6605 ;
  assign n6607 = n1675 & n6606 ;
  assign n6608 = n6607 ^ n5583 ^ 1'b0 ;
  assign n6609 = n4501 ^ n4012 ^ n3923 ;
  assign n6610 = ( n290 & n6608 ) | ( n290 & n6609 ) | ( n6608 & n6609 ) ;
  assign n6611 = n6610 ^ n4477 ^ 1'b0 ;
  assign n6615 = n6614 ^ n6611 ^ 1'b0 ;
  assign n6619 = ~n3236 & n3431 ;
  assign n6620 = ~n389 & n5941 ;
  assign n6621 = n6620 ^ n2526 ^ 1'b0 ;
  assign n6622 = ( n2846 & n6619 ) | ( n2846 & n6621 ) | ( n6619 & n6621 ) ;
  assign n6616 = n2676 & n4070 ;
  assign n6617 = n6616 ^ n5008 ^ n1154 ;
  assign n6618 = n6617 ^ n4529 ^ n3300 ;
  assign n6623 = n6622 ^ n6618 ^ n2428 ;
  assign n6624 = ( n620 & ~n6410 ) | ( n620 & n6623 ) | ( ~n6410 & n6623 ) ;
  assign n6625 = n657 & n852 ;
  assign n6626 = n2389 & n6625 ;
  assign n6627 = ( n1200 & n3332 ) | ( n1200 & ~n6626 ) | ( n3332 & ~n6626 ) ;
  assign n6628 = n6627 ^ n6362 ^ n3422 ;
  assign n6629 = n263 & ~n2388 ;
  assign n6630 = n6628 & n6629 ;
  assign n6631 = n5740 | n6630 ;
  assign n6632 = n3068 & ~n6631 ;
  assign n6633 = ( n3050 & ~n3828 ) | ( n3050 & n6632 ) | ( ~n3828 & n6632 ) ;
  assign n6640 = n4852 ^ n4010 ^ n3399 ;
  assign n6639 = n4609 ^ n4139 ^ n3525 ;
  assign n6641 = n6640 ^ n6639 ^ 1'b0 ;
  assign n6642 = n3291 | n6641 ;
  assign n6634 = ( n781 & n2144 ) | ( n781 & ~n4163 ) | ( n2144 & ~n4163 ) ;
  assign n6635 = n6041 & n6634 ;
  assign n6636 = ( n1304 & n4510 ) | ( n1304 & n5233 ) | ( n4510 & n5233 ) ;
  assign n6637 = n6636 ^ n2771 ^ n2118 ;
  assign n6638 = ( n3922 & ~n6635 ) | ( n3922 & n6637 ) | ( ~n6635 & n6637 ) ;
  assign n6643 = n6642 ^ n6638 ^ 1'b0 ;
  assign n6646 = n1068 & ~n5942 ;
  assign n6647 = ~n715 & n4885 ;
  assign n6648 = ~n883 & n6647 ;
  assign n6649 = ~n6646 & n6648 ;
  assign n6650 = n5042 | n6649 ;
  assign n6651 = ( n1161 & ~n1554 ) | ( n1161 & n6650 ) | ( ~n1554 & n6650 ) ;
  assign n6644 = n2865 ^ x24 ^ 1'b0 ;
  assign n6645 = ( n2217 & n3326 ) | ( n2217 & n6644 ) | ( n3326 & n6644 ) ;
  assign n6652 = n6651 ^ n6645 ^ n6046 ;
  assign n6662 = x192 & n1433 ;
  assign n6663 = n6662 ^ n3286 ^ 1'b0 ;
  assign n6653 = ( n598 & ~n1218 ) | ( n598 & n2591 ) | ( ~n1218 & n2591 ) ;
  assign n6654 = ~n1118 & n6653 ;
  assign n6655 = ( n1757 & n2793 ) | ( n1757 & n5611 ) | ( n2793 & n5611 ) ;
  assign n6656 = ~n1562 & n6655 ;
  assign n6657 = n6654 & n6656 ;
  assign n6658 = ( n282 & n434 ) | ( n282 & ~n3281 ) | ( n434 & ~n3281 ) ;
  assign n6659 = ( n2185 & ~n3671 ) | ( n2185 & n6658 ) | ( ~n3671 & n6658 ) ;
  assign n6660 = n6659 ^ n408 ^ 1'b0 ;
  assign n6661 = ~n6657 & n6660 ;
  assign n6664 = n6663 ^ n6661 ^ 1'b0 ;
  assign n6668 = ( n1503 & ~n2319 ) | ( n1503 & n2635 ) | ( ~n2319 & n2635 ) ;
  assign n6669 = n5363 ^ n530 ^ n278 ;
  assign n6670 = ( ~n5724 & n6668 ) | ( ~n5724 & n6669 ) | ( n6668 & n6669 ) ;
  assign n6666 = n2851 ^ n2064 ^ x193 ;
  assign n6665 = n1291 & n4541 ;
  assign n6667 = n6666 ^ n6665 ^ 1'b0 ;
  assign n6671 = n6670 ^ n6667 ^ n2377 ;
  assign n6672 = n4748 ^ n2932 ^ n2094 ;
  assign n6673 = ( n3664 & n6671 ) | ( n3664 & n6672 ) | ( n6671 & n6672 ) ;
  assign n6674 = n1794 & n3996 ;
  assign n6675 = n6674 ^ n2625 ^ 1'b0 ;
  assign n6676 = n4983 ^ n3015 ^ n881 ;
  assign n6677 = n6676 ^ n3427 ^ 1'b0 ;
  assign n6678 = ~x31 & n2075 ;
  assign n6679 = n1197 & ~n6678 ;
  assign n6680 = ~n2504 & n6679 ;
  assign n6681 = n286 & n6680 ;
  assign n6682 = n6681 ^ n3961 ^ 1'b0 ;
  assign n6683 = ( ~n857 & n1858 ) | ( ~n857 & n2684 ) | ( n1858 & n2684 ) ;
  assign n6686 = n2795 ^ n815 ^ 1'b0 ;
  assign n6687 = x118 & n6686 ;
  assign n6684 = n6655 ^ n1325 ^ n755 ;
  assign n6685 = n5736 & n6684 ;
  assign n6688 = n6687 ^ n6685 ^ 1'b0 ;
  assign n6689 = n5797 & n6688 ;
  assign n6691 = n3905 ^ n886 ^ x107 ;
  assign n6692 = ( n669 & n4408 ) | ( n669 & ~n6691 ) | ( n4408 & ~n6691 ) ;
  assign n6690 = n918 & ~n5164 ;
  assign n6693 = n6692 ^ n6690 ^ 1'b0 ;
  assign n6698 = n3641 ^ n929 ^ 1'b0 ;
  assign n6699 = n6698 ^ n1020 ^ 1'b0 ;
  assign n6697 = n3549 ^ n1997 ^ n1039 ;
  assign n6700 = n6699 ^ n6697 ^ n2031 ;
  assign n6694 = n5893 ^ n1830 ^ 1'b0 ;
  assign n6695 = n6463 ^ n5844 ^ 1'b0 ;
  assign n6696 = n6694 & ~n6695 ;
  assign n6701 = n6700 ^ n6696 ^ 1'b0 ;
  assign n6703 = n4487 ^ n3585 ^ n1558 ;
  assign n6702 = n1865 | n2018 ;
  assign n6704 = n6703 ^ n6702 ^ n3248 ;
  assign n6705 = n6704 ^ n4856 ^ n4011 ;
  assign n6706 = n6705 ^ n1940 ^ 1'b0 ;
  assign n6707 = n5236 ^ n4145 ^ n494 ;
  assign n6708 = n6368 | n6707 ;
  assign n6709 = n901 ^ n836 ^ n818 ;
  assign n6710 = ( n840 & n1848 ) | ( n840 & ~n4128 ) | ( n1848 & ~n4128 ) ;
  assign n6711 = ( n4644 & n6709 ) | ( n4644 & ~n6710 ) | ( n6709 & ~n6710 ) ;
  assign n6712 = ( n576 & n4000 ) | ( n576 & n6711 ) | ( n4000 & n6711 ) ;
  assign n6713 = ( n1835 & n3556 ) | ( n1835 & n4623 ) | ( n3556 & n4623 ) ;
  assign n6714 = ( ~n2025 & n6712 ) | ( ~n2025 & n6713 ) | ( n6712 & n6713 ) ;
  assign n6715 = n4472 ^ n3980 ^ 1'b0 ;
  assign n6716 = ( ~x82 & n1079 ) | ( ~x82 & n1465 ) | ( n1079 & n1465 ) ;
  assign n6717 = n1455 & n6716 ;
  assign n6718 = n6717 ^ n5983 ^ n399 ;
  assign n6721 = n4279 ^ n928 ^ 1'b0 ;
  assign n6722 = n1421 | n6721 ;
  assign n6719 = ( n637 & n1002 ) | ( n637 & ~n2603 ) | ( n1002 & ~n2603 ) ;
  assign n6720 = n2477 & n6719 ;
  assign n6723 = n6722 ^ n6720 ^ 1'b0 ;
  assign n6724 = n6723 ^ n5072 ^ n3583 ;
  assign n6725 = n356 & n6724 ;
  assign n6726 = ( n621 & n4342 ) | ( n621 & n6725 ) | ( n4342 & n6725 ) ;
  assign n6727 = n1005 & n6494 ;
  assign n6728 = n6727 ^ n1363 ^ 1'b0 ;
  assign n6729 = n3064 | n5599 ;
  assign n6730 = n6728 | n6729 ;
  assign n6731 = n6730 ^ n5762 ^ n4130 ;
  assign n6732 = n1155 & ~n2564 ;
  assign n6733 = ( n1852 & n2461 ) | ( n1852 & ~n3401 ) | ( n2461 & ~n3401 ) ;
  assign n6734 = ~n333 & n6733 ;
  assign n6735 = ~n3579 & n6734 ;
  assign n6736 = n6735 ^ n3143 ^ n547 ;
  assign n6737 = n3614 & n6736 ;
  assign n6738 = ( n886 & n2737 ) | ( n886 & ~n6737 ) | ( n2737 & ~n6737 ) ;
  assign n6739 = ( ~n2978 & n6732 ) | ( ~n2978 & n6738 ) | ( n6732 & n6738 ) ;
  assign n6740 = n6739 ^ n6430 ^ n3509 ;
  assign n6748 = n1758 & n3490 ;
  assign n6749 = n6748 ^ n3169 ^ 1'b0 ;
  assign n6741 = n575 | n3250 ;
  assign n6742 = x215 | n6741 ;
  assign n6743 = n6742 ^ n4512 ^ n628 ;
  assign n6744 = n6743 ^ n3063 ^ 1'b0 ;
  assign n6745 = n898 & n6744 ;
  assign n6746 = n1000 & n6745 ;
  assign n6747 = n6746 ^ n302 ^ 1'b0 ;
  assign n6750 = n6749 ^ n6747 ^ n5576 ;
  assign n6751 = n1154 | n5213 ;
  assign n6752 = n2289 & ~n6751 ;
  assign n6753 = n6752 ^ n1175 ^ 1'b0 ;
  assign n6754 = n6750 & n6753 ;
  assign n6755 = ( n1538 & ~n1555 ) | ( n1538 & n2679 ) | ( ~n1555 & n2679 ) ;
  assign n6756 = n3173 ^ n1320 ^ 1'b0 ;
  assign n6757 = n6755 | n6756 ;
  assign n6758 = n1260 ^ x98 ^ 1'b0 ;
  assign n6759 = n1327 & ~n6758 ;
  assign n6760 = ( n6478 & n6757 ) | ( n6478 & n6759 ) | ( n6757 & n6759 ) ;
  assign n6761 = ( n2485 & n6300 ) | ( n2485 & n6452 ) | ( n6300 & n6452 ) ;
  assign n6765 = n5220 ^ n873 ^ n872 ;
  assign n6762 = ~n1726 & n4796 ;
  assign n6763 = n5680 | n6762 ;
  assign n6764 = n6763 ^ n1417 ^ 1'b0 ;
  assign n6766 = n6765 ^ n6764 ^ n4368 ;
  assign n6767 = n3248 ^ n3109 ^ n846 ;
  assign n6768 = ( ~n5937 & n6766 ) | ( ~n5937 & n6767 ) | ( n6766 & n6767 ) ;
  assign n6769 = ( ~n2091 & n3000 ) | ( ~n2091 & n6768 ) | ( n3000 & n6768 ) ;
  assign n6770 = n4578 ^ n3612 ^ n337 ;
  assign n6771 = n1120 & n6770 ;
  assign n6772 = ( n530 & ~n6769 ) | ( n530 & n6771 ) | ( ~n6769 & n6771 ) ;
  assign n6774 = ( n657 & n4192 ) | ( n657 & n5484 ) | ( n4192 & n5484 ) ;
  assign n6773 = n3859 & ~n4935 ;
  assign n6775 = n6774 ^ n6773 ^ 1'b0 ;
  assign n6783 = n1405 | n2918 ;
  assign n6784 = n6783 ^ n6038 ^ n1287 ;
  assign n6780 = n4164 ^ n1376 ^ x90 ;
  assign n6781 = n6780 ^ n5462 ^ n298 ;
  assign n6782 = n2988 & ~n6781 ;
  assign n6785 = n6784 ^ n6782 ^ 1'b0 ;
  assign n6776 = n374 ^ n288 ^ 1'b0 ;
  assign n6777 = n733 & n4110 ;
  assign n6778 = n6776 & n6777 ;
  assign n6779 = n3933 & ~n6778 ;
  assign n6786 = n6785 ^ n6779 ^ 1'b0 ;
  assign n6787 = n2486 ^ x67 ^ 1'b0 ;
  assign n6788 = ~n6786 & n6787 ;
  assign n6789 = n4825 ^ n785 ^ x73 ;
  assign n6790 = n380 & n805 ;
  assign n6791 = n6790 ^ n4798 ^ 1'b0 ;
  assign n6792 = n6789 | n6791 ;
  assign n6793 = x1 & x93 ;
  assign n6794 = n6793 ^ n925 ^ 1'b0 ;
  assign n6795 = n6724 ^ n5054 ^ 1'b0 ;
  assign n6796 = n6794 | n6795 ;
  assign n6797 = n6796 ^ n5506 ^ 1'b0 ;
  assign n6798 = n5164 ^ n2980 ^ n1321 ;
  assign n6799 = ( n325 & n4436 ) | ( n325 & ~n6798 ) | ( n4436 & ~n6798 ) ;
  assign n6800 = n6511 & ~n6799 ;
  assign n6801 = ~n2087 & n6800 ;
  assign n6802 = n6124 ^ n2884 ^ n2694 ;
  assign n6803 = n5329 ^ n3583 ^ n3424 ;
  assign n6804 = ( n719 & ~n1703 ) | ( n719 & n2634 ) | ( ~n1703 & n2634 ) ;
  assign n6805 = n6803 | n6804 ;
  assign n6806 = n6805 ^ n1155 ^ 1'b0 ;
  assign n6813 = x26 | n495 ;
  assign n6809 = n5997 ^ n4734 ^ n2691 ;
  assign n6807 = x83 & n2765 ;
  assign n6808 = ~n6622 & n6807 ;
  assign n6810 = n6809 ^ n6808 ^ n2285 ;
  assign n6811 = ~n1200 & n3960 ;
  assign n6812 = ~n6810 & n6811 ;
  assign n6814 = n6813 ^ n6812 ^ n975 ;
  assign n6815 = ( ~n2047 & n6806 ) | ( ~n2047 & n6814 ) | ( n6806 & n6814 ) ;
  assign n6816 = n2622 ^ n1741 ^ 1'b0 ;
  assign n6817 = n5884 ^ n4070 ^ n2878 ;
  assign n6818 = n4533 ^ n4486 ^ 1'b0 ;
  assign n6819 = n6817 & n6818 ;
  assign n6823 = n2913 ^ n2216 ^ n492 ;
  assign n6822 = n5498 & ~n5501 ;
  assign n6824 = n6823 ^ n6822 ^ 1'b0 ;
  assign n6820 = n4841 ^ n4002 ^ 1'b0 ;
  assign n6821 = ( n1873 & ~n6088 ) | ( n1873 & n6820 ) | ( ~n6088 & n6820 ) ;
  assign n6825 = n6824 ^ n6821 ^ n2027 ;
  assign n6826 = n2426 | n3178 ;
  assign n6827 = n6826 ^ n1894 ^ 1'b0 ;
  assign n6828 = n6827 ^ n4518 ^ n2999 ;
  assign n6829 = n4670 & n6828 ;
  assign n6830 = x99 & n2886 ;
  assign n6831 = n1299 & n6830 ;
  assign n6832 = n641 | n6831 ;
  assign n6833 = n6829 & ~n6832 ;
  assign n6841 = n1287 ^ n1151 ^ 1'b0 ;
  assign n6842 = n2573 | n6841 ;
  assign n6840 = n6051 & ~n6465 ;
  assign n6837 = ~n908 & n4848 ;
  assign n6838 = ~n1616 & n6837 ;
  assign n6834 = ( n431 & n1168 ) | ( n431 & ~n2224 ) | ( n1168 & ~n2224 ) ;
  assign n6835 = n6834 ^ n2227 ^ 1'b0 ;
  assign n6836 = n1605 & ~n6835 ;
  assign n6839 = n6838 ^ n6836 ^ n2509 ;
  assign n6843 = n6842 ^ n6840 ^ n6839 ;
  assign n6844 = n481 & n6843 ;
  assign n6845 = n5777 ^ n1592 ^ x75 ;
  assign n6846 = n6067 ^ n4682 ^ n2053 ;
  assign n6847 = ( x140 & n3754 ) | ( x140 & ~n3803 ) | ( n3754 & ~n3803 ) ;
  assign n6848 = n4122 ^ n3349 ^ 1'b0 ;
  assign n6849 = n6847 & ~n6848 ;
  assign n6850 = n4750 ^ n2755 ^ n2298 ;
  assign n6851 = ( n5617 & n6849 ) | ( n5617 & ~n6850 ) | ( n6849 & ~n6850 ) ;
  assign n6852 = n6851 ^ n6368 ^ n3737 ;
  assign n6853 = x180 & n3084 ;
  assign n6854 = n6853 ^ n3323 ^ 1'b0 ;
  assign n6855 = n5328 ^ n2382 ^ n298 ;
  assign n6856 = n3460 ^ n348 ^ 1'b0 ;
  assign n6857 = n2214 & n6856 ;
  assign n6858 = n6855 & n6857 ;
  assign n6859 = n582 ^ x85 ^ 1'b0 ;
  assign n6860 = n4897 & n6859 ;
  assign n6861 = n2508 ^ n1863 ^ n364 ;
  assign n6862 = n6861 ^ n431 ^ 1'b0 ;
  assign n6863 = n6862 ^ n6444 ^ n589 ;
  assign n6864 = n1674 ^ n1567 ^ n1149 ;
  assign n6865 = n563 & ~n6864 ;
  assign n6866 = n6865 ^ n1117 ^ 1'b0 ;
  assign n6867 = ( n814 & n2050 ) | ( n814 & n3303 ) | ( n2050 & n3303 ) ;
  assign n6868 = n6824 ^ n5863 ^ n1195 ;
  assign n6869 = ( n4237 & n6867 ) | ( n4237 & ~n6868 ) | ( n6867 & ~n6868 ) ;
  assign n6870 = n6869 ^ n4254 ^ n3749 ;
  assign n6876 = n1972 | n3315 ;
  assign n6877 = n3948 | n6876 ;
  assign n6874 = n2998 ^ n2212 ^ n1982 ;
  assign n6875 = ( x83 & n1485 ) | ( x83 & n6874 ) | ( n1485 & n6874 ) ;
  assign n6872 = n385 & ~n478 ;
  assign n6871 = ( n1748 & ~n3185 ) | ( n1748 & n3787 ) | ( ~n3185 & n3787 ) ;
  assign n6873 = n6872 ^ n6871 ^ n6255 ;
  assign n6878 = n6877 ^ n6875 ^ n6873 ;
  assign n6879 = n1405 ^ x147 ^ 1'b0 ;
  assign n6880 = x99 & ~n6879 ;
  assign n6881 = n2935 & n6880 ;
  assign n6882 = n6881 ^ n720 ^ 1'b0 ;
  assign n6883 = n6882 ^ n4838 ^ x246 ;
  assign n6884 = n1951 | n4177 ;
  assign n6885 = n6884 ^ n5242 ^ 1'b0 ;
  assign n6886 = ( n1554 & ~n3904 ) | ( n1554 & n4963 ) | ( ~n3904 & n4963 ) ;
  assign n6887 = n4316 ^ n2918 ^ x131 ;
  assign n6888 = n6887 ^ n4952 ^ 1'b0 ;
  assign n6889 = ( n632 & n6886 ) | ( n632 & ~n6888 ) | ( n6886 & ~n6888 ) ;
  assign n6890 = n5798 ^ n3599 ^ n3304 ;
  assign n6891 = n6890 ^ n1976 ^ 1'b0 ;
  assign n6892 = n4394 ^ n1244 ^ n1050 ;
  assign n6893 = ~n3101 & n6892 ;
  assign n6894 = n2393 & n6893 ;
  assign n6895 = ( ~n1673 & n6891 ) | ( ~n1673 & n6894 ) | ( n6891 & n6894 ) ;
  assign n6896 = n1739 ^ n491 ^ 1'b0 ;
  assign n6897 = ~n1217 & n2722 ;
  assign n6898 = ~n853 & n6897 ;
  assign n6899 = n6898 ^ n6231 ^ n2158 ;
  assign n6900 = n6896 & ~n6899 ;
  assign n6910 = n3561 ^ n2401 ^ n1158 ;
  assign n6909 = x20 & ~n513 ;
  assign n6911 = n6910 ^ n6909 ^ 1'b0 ;
  assign n6908 = ( n896 & ~n5284 ) | ( n896 & n5635 ) | ( ~n5284 & n5635 ) ;
  assign n6904 = n1194 ^ n353 ^ 1'b0 ;
  assign n6905 = n1323 & ~n6904 ;
  assign n6903 = ( n375 & n1574 ) | ( n375 & n5216 ) | ( n1574 & n5216 ) ;
  assign n6906 = n6905 ^ n6903 ^ n2648 ;
  assign n6901 = n1911 ^ n813 ^ 1'b0 ;
  assign n6902 = n3097 & ~n6901 ;
  assign n6907 = n6906 ^ n6902 ^ 1'b0 ;
  assign n6912 = n6911 ^ n6908 ^ n6907 ;
  assign n6913 = n6912 ^ n4613 ^ n1369 ;
  assign n6918 = n6118 ^ n1875 ^ n733 ;
  assign n6914 = n1601 ^ n883 ^ n449 ;
  assign n6915 = ( n2629 & n4194 ) | ( n2629 & n6914 ) | ( n4194 & n6914 ) ;
  assign n6916 = n306 & n6915 ;
  assign n6917 = ~n2144 & n6916 ;
  assign n6919 = n6918 ^ n6917 ^ n1488 ;
  assign n6920 = ( ~n950 & n2950 ) | ( ~n950 & n6919 ) | ( n2950 & n6919 ) ;
  assign n6921 = ( ~n3857 & n5767 ) | ( ~n3857 & n6804 ) | ( n5767 & n6804 ) ;
  assign n6922 = ( n367 & n2091 ) | ( n367 & ~n6921 ) | ( n2091 & ~n6921 ) ;
  assign n6923 = n2463 & ~n6922 ;
  assign n6924 = n2905 & n6923 ;
  assign n6937 = n1479 ^ x244 ^ x123 ;
  assign n6938 = n6937 ^ n4135 ^ 1'b0 ;
  assign n6939 = n6938 ^ n828 ^ 1'b0 ;
  assign n6932 = n2506 ^ n557 ^ 1'b0 ;
  assign n6933 = n546 & ~n6932 ;
  assign n6934 = ~n3158 & n6933 ;
  assign n6935 = ~n1459 & n6934 ;
  assign n6926 = ( n765 & n2792 ) | ( n765 & ~n3368 ) | ( n2792 & ~n3368 ) ;
  assign n6925 = n2143 & n3679 ;
  assign n6927 = n6926 ^ n6925 ^ n379 ;
  assign n6928 = n6927 ^ n1276 ^ 1'b0 ;
  assign n6929 = x104 & n563 ;
  assign n6930 = ~n5495 & n6929 ;
  assign n6931 = n6928 & ~n6930 ;
  assign n6936 = n6935 ^ n6931 ^ 1'b0 ;
  assign n6940 = n6939 ^ n6936 ^ n5637 ;
  assign n6955 = n6231 ^ n1422 ^ x116 ;
  assign n6956 = n6955 ^ x184 ^ 1'b0 ;
  assign n6953 = n6527 ^ x213 ^ 1'b0 ;
  assign n6954 = x53 & n6953 ;
  assign n6943 = ( ~x112 & n360 ) | ( ~x112 & n2076 ) | ( n360 & n2076 ) ;
  assign n6944 = n6943 ^ n3693 ^ 1'b0 ;
  assign n6941 = n2570 ^ x23 ^ 1'b0 ;
  assign n6942 = n3840 & n6941 ;
  assign n6945 = n6944 ^ n6942 ^ n2317 ;
  assign n6946 = ~n854 & n2809 ;
  assign n6947 = n6946 ^ n5733 ^ 1'b0 ;
  assign n6948 = n749 & n6947 ;
  assign n6949 = ~x197 & n6948 ;
  assign n6950 = n6949 ^ n1407 ^ 1'b0 ;
  assign n6951 = n6945 | n6950 ;
  assign n6952 = n6951 ^ n4904 ^ n4014 ;
  assign n6957 = n6956 ^ n6954 ^ n6952 ;
  assign n6958 = n2043 | n6142 ;
  assign n6959 = n6958 ^ n765 ^ 1'b0 ;
  assign n6960 = n3599 ^ n1965 ^ n1945 ;
  assign n6961 = ( n376 & n6959 ) | ( n376 & ~n6960 ) | ( n6959 & ~n6960 ) ;
  assign n6962 = n5163 & ~n6666 ;
  assign n6963 = n1627 & n6962 ;
  assign n6964 = ( n1457 & ~n3813 ) | ( n1457 & n6963 ) | ( ~n3813 & n6963 ) ;
  assign n6965 = n4856 ^ n4665 ^ n2129 ;
  assign n6973 = n3299 ^ n2062 ^ x116 ;
  assign n6969 = ~n997 & n1220 ;
  assign n6970 = ~n1880 & n6969 ;
  assign n6971 = n6970 ^ n4689 ^ n1475 ;
  assign n6966 = ( ~n1293 & n2124 ) | ( ~n1293 & n6755 ) | ( n2124 & n6755 ) ;
  assign n6967 = n6966 ^ n6890 ^ n610 ;
  assign n6968 = ( n4319 & n4863 ) | ( n4319 & n6967 ) | ( n4863 & n6967 ) ;
  assign n6972 = n6971 ^ n6968 ^ n5786 ;
  assign n6974 = n6973 ^ n6972 ^ n6053 ;
  assign n6975 = ( n2328 & ~n5334 ) | ( n2328 & n6337 ) | ( ~n5334 & n6337 ) ;
  assign n6976 = n4735 | n5585 ;
  assign n6977 = ( n1457 & n2652 ) | ( n1457 & ~n4070 ) | ( n2652 & ~n4070 ) ;
  assign n6978 = ( ~n2443 & n6970 ) | ( ~n2443 & n6977 ) | ( n6970 & n6977 ) ;
  assign n6983 = ( n528 & n1113 ) | ( n528 & ~n2506 ) | ( n1113 & ~n2506 ) ;
  assign n6979 = n3474 ^ n1896 ^ 1'b0 ;
  assign n6980 = ( n2255 & ~n3010 ) | ( n2255 & n3953 ) | ( ~n3010 & n3953 ) ;
  assign n6981 = ~n5978 & n6980 ;
  assign n6982 = ( ~n5720 & n6979 ) | ( ~n5720 & n6981 ) | ( n6979 & n6981 ) ;
  assign n6984 = n6983 ^ n6982 ^ n3716 ;
  assign n6987 = ( n359 & ~n1807 ) | ( n359 & n1960 ) | ( ~n1807 & n1960 ) ;
  assign n6988 = n1607 ^ n1087 ^ n838 ;
  assign n6989 = ~n393 & n6988 ;
  assign n6990 = ~n2960 & n6989 ;
  assign n6991 = ~n6987 & n6990 ;
  assign n6985 = ( n616 & n868 ) | ( n616 & n3872 ) | ( n868 & n3872 ) ;
  assign n6986 = ( n2610 & n5886 ) | ( n2610 & n6985 ) | ( n5886 & n6985 ) ;
  assign n6992 = n6991 ^ n6986 ^ 1'b0 ;
  assign n6993 = ( ~x67 & n4853 ) | ( ~x67 & n6992 ) | ( n4853 & n6992 ) ;
  assign n6994 = ( x89 & n3813 ) | ( x89 & ~n5740 ) | ( n3813 & ~n5740 ) ;
  assign n6995 = n6994 ^ n6511 ^ n4122 ;
  assign n6996 = ( n1465 & n3811 ) | ( n1465 & n4139 ) | ( n3811 & n4139 ) ;
  assign n6997 = n4288 ^ n2695 ^ n950 ;
  assign n6998 = n3372 & n6997 ;
  assign n6999 = n6998 ^ n5753 ^ n2450 ;
  assign n7000 = n3241 ^ n899 ^ 1'b0 ;
  assign n7001 = ( n6224 & n6999 ) | ( n6224 & ~n7000 ) | ( n6999 & ~n7000 ) ;
  assign n7004 = n5595 ^ n3017 ^ n1665 ;
  assign n7002 = n6915 ^ n3325 ^ n3305 ;
  assign n7003 = n1962 | n7002 ;
  assign n7005 = n7004 ^ n7003 ^ 1'b0 ;
  assign n7014 = n4883 ^ n1349 ^ 1'b0 ;
  assign n7015 = ~n835 & n7014 ;
  assign n7013 = n1899 | n2494 ;
  assign n7016 = n7015 ^ n7013 ^ 1'b0 ;
  assign n7017 = x250 & n7016 ;
  assign n7012 = ( n597 & ~n4128 ) | ( n597 & n5429 ) | ( ~n4128 & n5429 ) ;
  assign n7006 = n1127 | n1968 ;
  assign n7018 = n7017 ^ n7012 ^ n7006 ;
  assign n7019 = n2847 | n7018 ;
  assign n7020 = n4297 | n7019 ;
  assign n7021 = n7020 ^ n4389 ^ n585 ;
  assign n7009 = n971 & n4734 ;
  assign n7007 = n2662 ^ n2311 ^ n755 ;
  assign n7008 = n3097 & ~n7007 ;
  assign n7010 = n7009 ^ n7008 ^ 1'b0 ;
  assign n7011 = n7006 | n7010 ;
  assign n7022 = n7021 ^ n7011 ^ 1'b0 ;
  assign n7023 = ( n969 & n7005 ) | ( n969 & n7022 ) | ( n7005 & n7022 ) ;
  assign n7024 = n7023 ^ n1709 ^ 1'b0 ;
  assign n7025 = n6949 ^ n6794 ^ n4817 ;
  assign n7026 = ( n1112 & n2820 ) | ( n1112 & ~n7025 ) | ( n2820 & ~n7025 ) ;
  assign n7037 = n6377 ^ n3583 ^ n3175 ;
  assign n7035 = ( ~n2826 & n3596 ) | ( ~n2826 & n3962 ) | ( n3596 & n3962 ) ;
  assign n7028 = ( ~n3841 & n4976 ) | ( ~n3841 & n5724 ) | ( n4976 & n5724 ) ;
  assign n7029 = n2376 ^ n498 ^ x225 ;
  assign n7030 = ( n1278 & n1298 ) | ( n1278 & n6042 ) | ( n1298 & n6042 ) ;
  assign n7031 = ( n6381 & n7029 ) | ( n6381 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7032 = ( n407 & n6234 ) | ( n407 & n7031 ) | ( n6234 & n7031 ) ;
  assign n7033 = n7032 ^ n2166 ^ 1'b0 ;
  assign n7034 = n7028 & ~n7033 ;
  assign n7027 = n6774 ^ n2867 ^ 1'b0 ;
  assign n7036 = n7035 ^ n7034 ^ n7027 ;
  assign n7038 = n7037 ^ n7036 ^ 1'b0 ;
  assign n7039 = n2309 | n2553 ;
  assign n7040 = n5275 | n7039 ;
  assign n7041 = x241 | n7040 ;
  assign n7042 = n3592 ^ n2548 ^ n2481 ;
  assign n7043 = n3872 ^ n1844 ^ n1638 ;
  assign n7044 = n1967 ^ n1579 ^ n600 ;
  assign n7045 = ( n1142 & ~n2538 ) | ( n1142 & n3639 ) | ( ~n2538 & n3639 ) ;
  assign n7046 = ( ~n1556 & n7044 ) | ( ~n1556 & n7045 ) | ( n7044 & n7045 ) ;
  assign n7047 = n6653 ^ n1410 ^ n1344 ;
  assign n7048 = n7047 ^ x60 ^ 1'b0 ;
  assign n7049 = ~n5352 & n7048 ;
  assign n7050 = n7049 ^ n2290 ^ n1146 ;
  assign n7051 = ( ~n7043 & n7046 ) | ( ~n7043 & n7050 ) | ( n7046 & n7050 ) ;
  assign n7052 = n5069 & ~n7051 ;
  assign n7053 = ~n7042 & n7052 ;
  assign n7055 = n4240 ^ n2228 ^ 1'b0 ;
  assign n7056 = n1397 & ~n7055 ;
  assign n7057 = n7056 ^ n4449 ^ n3799 ;
  assign n7054 = ( n4541 & ~n6148 ) | ( n4541 & n6955 ) | ( ~n6148 & n6955 ) ;
  assign n7058 = n7057 ^ n7054 ^ n3280 ;
  assign n7059 = n7058 ^ n920 ^ 1'b0 ;
  assign n7060 = n7053 | n7059 ;
  assign n7061 = n6236 ^ n4169 ^ n903 ;
  assign n7062 = ( n988 & n5131 ) | ( n988 & ~n5789 ) | ( n5131 & ~n5789 ) ;
  assign n7063 = n7062 ^ n2053 ^ n486 ;
  assign n7064 = n2818 ^ n1918 ^ 1'b0 ;
  assign n7065 = n1827 & ~n7064 ;
  assign n7066 = n6293 ^ n1392 ^ 1'b0 ;
  assign n7067 = n4139 | n7066 ;
  assign n7068 = n7067 ^ n6892 ^ n2171 ;
  assign n7069 = ( n5829 & ~n7065 ) | ( n5829 & n7068 ) | ( ~n7065 & n7068 ) ;
  assign n7070 = ( n2935 & ~n7063 ) | ( n2935 & n7069 ) | ( ~n7063 & n7069 ) ;
  assign n7071 = ~n3593 & n7070 ;
  assign n7072 = ( n5089 & ~n6561 ) | ( n5089 & n7071 ) | ( ~n6561 & n7071 ) ;
  assign n7079 = ( x163 & ~n1565 ) | ( x163 & n4539 ) | ( ~n1565 & n4539 ) ;
  assign n7076 = n1959 & n2011 ;
  assign n7077 = n7076 ^ n402 ^ 1'b0 ;
  assign n7074 = n5376 ^ n3976 ^ n2456 ;
  assign n7073 = n3454 ^ n2981 ^ n2678 ;
  assign n7075 = n7074 ^ n7073 ^ n3736 ;
  assign n7078 = n7077 ^ n7075 ^ n1979 ;
  assign n7080 = n7079 ^ n7078 ^ n6600 ;
  assign n7081 = n895 & ~n1378 ;
  assign n7082 = n7081 ^ n6560 ^ 1'b0 ;
  assign n7083 = ( ~n912 & n2066 ) | ( ~n912 & n7082 ) | ( n2066 & n7082 ) ;
  assign n7084 = n4145 ^ n271 ^ 1'b0 ;
  assign n7088 = ( n1495 & n3293 ) | ( n1495 & n5242 ) | ( n3293 & n5242 ) ;
  assign n7089 = n7088 ^ n5662 ^ n2683 ;
  assign n7085 = n4070 ^ n1301 ^ n988 ;
  assign n7086 = n7085 ^ n459 ^ 1'b0 ;
  assign n7087 = n6454 & n7086 ;
  assign n7090 = n7089 ^ n7087 ^ 1'b0 ;
  assign n7091 = ( n1821 & ~n2134 ) | ( n1821 & n3343 ) | ( ~n2134 & n3343 ) ;
  assign n7092 = ( n2585 & ~n3511 ) | ( n2585 & n7091 ) | ( ~n3511 & n7091 ) ;
  assign n7093 = ~n5661 & n7092 ;
  assign n7094 = n7093 ^ n3076 ^ n1706 ;
  assign n7095 = n7094 ^ n259 ^ 1'b0 ;
  assign n7096 = n4549 & n5886 ;
  assign n7097 = n7096 ^ n5021 ^ 1'b0 ;
  assign n7098 = n7097 ^ n2852 ^ 1'b0 ;
  assign n7099 = n2432 ^ n1714 ^ n728 ;
  assign n7100 = n1347 & n2531 ;
  assign n7101 = n2240 ^ n1972 ^ 1'b0 ;
  assign n7102 = n4444 ^ n2257 ^ n288 ;
  assign n7103 = n7102 ^ n911 ^ 1'b0 ;
  assign n7104 = n2750 & ~n7103 ;
  assign n7105 = n7104 ^ n3536 ^ x172 ;
  assign n7106 = n478 ^ x29 ^ 1'b0 ;
  assign n7107 = ( n7101 & n7105 ) | ( n7101 & n7106 ) | ( n7105 & n7106 ) ;
  assign n7108 = ( n7099 & ~n7100 ) | ( n7099 & n7107 ) | ( ~n7100 & n7107 ) ;
  assign n7109 = n4268 ^ n3716 ^ 1'b0 ;
  assign n7110 = n3433 ^ n474 ^ 1'b0 ;
  assign n7111 = n7110 ^ n5111 ^ n1949 ;
  assign n7112 = n3247 ^ n2965 ^ 1'b0 ;
  assign n7113 = n7112 ^ n3967 ^ n2055 ;
  assign n7114 = ( ~n1590 & n3814 ) | ( ~n1590 & n6355 ) | ( n3814 & n6355 ) ;
  assign n7115 = ( n1860 & n3136 ) | ( n1860 & n4147 ) | ( n3136 & n4147 ) ;
  assign n7116 = n5890 ^ n2221 ^ x143 ;
  assign n7117 = n7115 & ~n7116 ;
  assign n7118 = ~n7114 & n7117 ;
  assign n7119 = n7118 ^ n6605 ^ 1'b0 ;
  assign n7120 = n6132 & ~n7119 ;
  assign n7121 = ( n523 & n6801 ) | ( n523 & n7120 ) | ( n6801 & n7120 ) ;
  assign n7122 = n4890 | n5508 ;
  assign n7128 = n1362 | n2514 ;
  assign n7123 = n2566 & ~n2809 ;
  assign n7124 = ~n5300 & n7123 ;
  assign n7125 = n7124 ^ n1291 ^ 1'b0 ;
  assign n7126 = n7125 ^ n2328 ^ 1'b0 ;
  assign n7127 = n749 & n7126 ;
  assign n7129 = n7128 ^ n7127 ^ n1015 ;
  assign n7134 = ~n1224 & n5611 ;
  assign n7133 = n4309 ^ n1553 ^ n834 ;
  assign n7130 = n6110 ^ n1705 ^ x239 ;
  assign n7131 = n4496 & ~n7130 ;
  assign n7132 = n843 & n7131 ;
  assign n7135 = n7134 ^ n7133 ^ n7132 ;
  assign n7136 = ( x105 & n2905 ) | ( x105 & ~n7135 ) | ( n2905 & ~n7135 ) ;
  assign n7137 = n7136 ^ n4238 ^ 1'b0 ;
  assign n7138 = n5777 ^ n2028 ^ 1'b0 ;
  assign n7139 = n2962 & n7138 ;
  assign n7140 = ( n928 & ~n1954 ) | ( n928 & n7139 ) | ( ~n1954 & n7139 ) ;
  assign n7141 = ( ~n5352 & n6863 ) | ( ~n5352 & n7140 ) | ( n6863 & n7140 ) ;
  assign n7142 = n3463 ^ n1601 ^ n1152 ;
  assign n7143 = n415 & ~n7142 ;
  assign n7144 = ~n1594 & n4526 ;
  assign n7145 = ( n4899 & ~n5394 ) | ( n4899 & n7144 ) | ( ~n5394 & n7144 ) ;
  assign n7148 = n5398 ^ n4767 ^ n2185 ;
  assign n7146 = n561 | n5294 ;
  assign n7147 = n1231 & ~n7146 ;
  assign n7149 = n7148 ^ n7147 ^ n4271 ;
  assign n7153 = ( n522 & n798 ) | ( n522 & ~n1433 ) | ( n798 & ~n1433 ) ;
  assign n7150 = ( ~x43 & n1088 ) | ( ~x43 & n2570 ) | ( n1088 & n2570 ) ;
  assign n7151 = n7150 ^ n2867 ^ n1943 ;
  assign n7152 = n7151 ^ n1716 ^ 1'b0 ;
  assign n7154 = n7153 ^ n7152 ^ n2256 ;
  assign n7155 = n2923 ^ n1384 ^ n1170 ;
  assign n7156 = n6769 & n7155 ;
  assign n7157 = n911 & ~n7156 ;
  assign n7158 = ~x226 & n7157 ;
  assign n7159 = n7158 ^ n5258 ^ n4225 ;
  assign n7160 = ( x233 & n2684 ) | ( x233 & n7159 ) | ( n2684 & n7159 ) ;
  assign n7183 = n683 ^ n277 ^ n274 ;
  assign n7184 = n7183 ^ n1670 ^ n1485 ;
  assign n7185 = n7184 ^ n2456 ^ n1507 ;
  assign n7169 = n5253 ^ n1142 ^ n784 ;
  assign n7170 = n2300 | n4946 ;
  assign n7171 = n7170 ^ n4534 ^ 1'b0 ;
  assign n7174 = n2605 ^ n2076 ^ n1340 ;
  assign n7175 = n1678 & ~n7174 ;
  assign n7176 = n7175 ^ n1168 ^ 1'b0 ;
  assign n7177 = ( x62 & n1175 ) | ( x62 & n7176 ) | ( n1175 & n7176 ) ;
  assign n7178 = n2139 | n6184 ;
  assign n7179 = n7177 & n7178 ;
  assign n7180 = n6599 & n7179 ;
  assign n7172 = ( ~n1295 & n4309 ) | ( ~n1295 & n5022 ) | ( n4309 & n5022 ) ;
  assign n7173 = n7172 ^ n3386 ^ n2997 ;
  assign n7181 = n7180 ^ n7173 ^ 1'b0 ;
  assign n7182 = ( n7169 & n7171 ) | ( n7169 & n7181 ) | ( n7171 & n7181 ) ;
  assign n7186 = n7185 ^ n7182 ^ n5320 ;
  assign n7161 = n1694 ^ n869 ^ 1'b0 ;
  assign n7162 = n5234 & n7161 ;
  assign n7163 = n7162 ^ n5302 ^ n1491 ;
  assign n7164 = n647 | n2329 ;
  assign n7165 = n7164 ^ n1238 ^ 1'b0 ;
  assign n7166 = n6824 | n7165 ;
  assign n7167 = n6659 ^ n476 ^ 1'b0 ;
  assign n7168 = ( n7163 & n7166 ) | ( n7163 & n7167 ) | ( n7166 & n7167 ) ;
  assign n7187 = n7186 ^ n7168 ^ n5376 ;
  assign n7188 = n5118 ^ n2199 ^ n1719 ;
  assign n7189 = n7188 ^ n573 ^ 1'b0 ;
  assign n7190 = ( n3566 & n6839 ) | ( n3566 & ~n7189 ) | ( n6839 & ~n7189 ) ;
  assign n7201 = n2436 & ~n6030 ;
  assign n7202 = ~n398 & n7201 ;
  assign n7203 = n7012 | n7202 ;
  assign n7204 = n7203 ^ n916 ^ 1'b0 ;
  assign n7191 = n2705 ^ n2609 ^ n298 ;
  assign n7192 = n4257 ^ n3158 ^ x97 ;
  assign n7193 = n2213 ^ n765 ^ 1'b0 ;
  assign n7194 = n7193 ^ n2183 ^ 1'b0 ;
  assign n7195 = n7192 | n7194 ;
  assign n7198 = ( ~n267 & n800 ) | ( ~n267 & n2711 ) | ( n800 & n2711 ) ;
  assign n7196 = n849 & n2657 ;
  assign n7197 = ( n1144 & n3638 ) | ( n1144 & n7196 ) | ( n3638 & n7196 ) ;
  assign n7199 = n7198 ^ n7197 ^ 1'b0 ;
  assign n7200 = ( ~n7191 & n7195 ) | ( ~n7191 & n7199 ) | ( n7195 & n7199 ) ;
  assign n7205 = n7204 ^ n7200 ^ 1'b0 ;
  assign n7206 = n4164 & n7205 ;
  assign n7207 = n6733 & ~n7206 ;
  assign n7208 = n5374 ^ n1943 ^ 1'b0 ;
  assign n7209 = n5886 ^ n1898 ^ n909 ;
  assign n7210 = n987 | n7209 ;
  assign n7211 = n7210 ^ n2115 ^ 1'b0 ;
  assign n7212 = n1308 & ~n6135 ;
  assign n7213 = n7212 ^ n1428 ^ 1'b0 ;
  assign n7214 = ( n5817 & ~n6604 ) | ( n5817 & n7213 ) | ( ~n6604 & n7213 ) ;
  assign n7215 = n2024 ^ n2002 ^ 1'b0 ;
  assign n7216 = n1668 & ~n7215 ;
  assign n7217 = ( n5247 & n7027 ) | ( n5247 & n7216 ) | ( n7027 & n7216 ) ;
  assign n7218 = ( n2323 & ~n2542 ) | ( n2323 & n5530 ) | ( ~n2542 & n5530 ) ;
  assign n7219 = n5194 ^ n3539 ^ x84 ;
  assign n7220 = n7218 & n7219 ;
  assign n7221 = n6235 & ~n7220 ;
  assign n7227 = n2631 ^ n1894 ^ n1032 ;
  assign n7228 = ( ~n3372 & n5074 ) | ( ~n3372 & n7227 ) | ( n5074 & n7227 ) ;
  assign n7222 = n4471 ^ n1122 ^ n379 ;
  assign n7223 = n2072 ^ n1913 ^ n1200 ;
  assign n7224 = n7223 ^ x115 ^ 1'b0 ;
  assign n7225 = n7224 ^ n3330 ^ n1801 ;
  assign n7226 = ( n1155 & ~n7222 ) | ( n1155 & n7225 ) | ( ~n7222 & n7225 ) ;
  assign n7229 = n7228 ^ n7226 ^ 1'b0 ;
  assign n7232 = n1863 & n3769 ;
  assign n7233 = n7232 ^ n1550 ^ 1'b0 ;
  assign n7234 = n7233 ^ n1449 ^ 1'b0 ;
  assign n7230 = n4228 ^ n4022 ^ 1'b0 ;
  assign n7231 = ( x57 & n3214 ) | ( x57 & n7230 ) | ( n3214 & n7230 ) ;
  assign n7235 = n7234 ^ n7231 ^ n1231 ;
  assign n7236 = n300 ^ x204 ^ x41 ;
  assign n7237 = n7236 ^ n6603 ^ 1'b0 ;
  assign n7243 = n3641 ^ n1674 ^ 1'b0 ;
  assign n7244 = n1110 & ~n7243 ;
  assign n7238 = n5165 ^ n1357 ^ n688 ;
  assign n7239 = n7238 ^ n4165 ^ 1'b0 ;
  assign n7240 = n4923 & n7239 ;
  assign n7241 = n7240 ^ n7114 ^ 1'b0 ;
  assign n7242 = n7241 ^ n2747 ^ 1'b0 ;
  assign n7245 = n7244 ^ n7242 ^ n6417 ;
  assign n7254 = n1503 & n5864 ;
  assign n7246 = n2389 | n2983 ;
  assign n7250 = ( n1101 & ~n1110 ) | ( n1101 & n2016 ) | ( ~n1110 & n2016 ) ;
  assign n7251 = n2994 | n7250 ;
  assign n7247 = ( ~n1044 & n5724 ) | ( ~n1044 & n6054 ) | ( n5724 & n6054 ) ;
  assign n7248 = n5965 & n7247 ;
  assign n7249 = ~n1071 & n7248 ;
  assign n7252 = n7251 ^ n7249 ^ n4998 ;
  assign n7253 = ( n5608 & n7246 ) | ( n5608 & n7252 ) | ( n7246 & n7252 ) ;
  assign n7255 = n7254 ^ n7253 ^ n7015 ;
  assign n7256 = n3704 ^ x122 ^ 1'b0 ;
  assign n7258 = n2139 & n3747 ;
  assign n7259 = n7258 ^ n2452 ^ 1'b0 ;
  assign n7257 = n6111 ^ n962 ^ n864 ;
  assign n7260 = n7259 ^ n7257 ^ n1974 ;
  assign n7261 = n6246 ^ n6244 ^ n1727 ;
  assign n7262 = n1590 ^ n271 ^ 1'b0 ;
  assign n7263 = n3016 & ~n7262 ;
  assign n7268 = ( n529 & n1315 ) | ( n529 & ~n1412 ) | ( n1315 & ~n1412 ) ;
  assign n7269 = n3514 ^ n3262 ^ 1'b0 ;
  assign n7270 = n7268 | n7269 ;
  assign n7266 = ~n1505 & n2525 ;
  assign n7267 = n7266 ^ x147 ^ 1'b0 ;
  assign n7264 = n296 | n5067 ;
  assign n7265 = n7264 ^ n1565 ^ n1055 ;
  assign n7271 = n7270 ^ n7267 ^ n7265 ;
  assign n7272 = n7271 ^ n4676 ^ 1'b0 ;
  assign n7273 = n6887 ^ n1027 ^ n415 ;
  assign n7274 = n6299 & n7273 ;
  assign n7275 = n7274 ^ n2479 ^ 1'b0 ;
  assign n7276 = n6042 ^ n3962 ^ 1'b0 ;
  assign n7277 = n5903 ^ n3782 ^ n1245 ;
  assign n7278 = ( n4175 & n4704 ) | ( n4175 & ~n7277 ) | ( n4704 & ~n7277 ) ;
  assign n7279 = ( n2216 & ~n5498 ) | ( n2216 & n5658 ) | ( ~n5498 & n5658 ) ;
  assign n7280 = ( n3401 & n4925 ) | ( n3401 & ~n7279 ) | ( n4925 & ~n7279 ) ;
  assign n7281 = ( n6528 & n7278 ) | ( n6528 & n7280 ) | ( n7278 & n7280 ) ;
  assign n7282 = ( n547 & n1996 ) | ( n547 & ~n2531 ) | ( n1996 & ~n2531 ) ;
  assign n7283 = ( ~n764 & n4221 ) | ( ~n764 & n7282 ) | ( n4221 & n7282 ) ;
  assign n7285 = ( n500 & n2840 ) | ( n500 & n5242 ) | ( n2840 & n5242 ) ;
  assign n7286 = ( n1806 & n2827 ) | ( n1806 & n7285 ) | ( n2827 & n7285 ) ;
  assign n7287 = n7286 ^ n6229 ^ n895 ;
  assign n7284 = ( x248 & n5380 ) | ( x248 & n5491 ) | ( n5380 & n5491 ) ;
  assign n7288 = n7287 ^ n7284 ^ n2876 ;
  assign n7289 = ( n3208 & n7283 ) | ( n3208 & ~n7288 ) | ( n7283 & ~n7288 ) ;
  assign n7290 = n3754 ^ n3399 ^ 1'b0 ;
  assign n7291 = n7290 ^ n5818 ^ n1385 ;
  assign n7294 = n6238 ^ n3185 ^ n836 ;
  assign n7292 = ( x41 & ~n610 ) | ( x41 & n2348 ) | ( ~n610 & n2348 ) ;
  assign n7293 = ( n4581 & n5760 ) | ( n4581 & ~n7292 ) | ( n5760 & ~n7292 ) ;
  assign n7295 = n7294 ^ n7293 ^ n5720 ;
  assign n7296 = ( n1315 & ~n2288 ) | ( n1315 & n2928 ) | ( ~n2288 & n2928 ) ;
  assign n7297 = n7296 ^ n4462 ^ x105 ;
  assign n7298 = n7297 ^ n5514 ^ n5479 ;
  assign n7299 = ( ~n6076 & n6865 ) | ( ~n6076 & n7298 ) | ( n6865 & n7298 ) ;
  assign n7300 = ( n2150 & ~n6719 ) | ( n2150 & n7299 ) | ( ~n6719 & n7299 ) ;
  assign n7304 = ( ~x239 & n909 ) | ( ~x239 & n2948 ) | ( n909 & n2948 ) ;
  assign n7303 = n6025 ^ n4255 ^ n1319 ;
  assign n7301 = n1273 | n3518 ;
  assign n7302 = n7301 ^ n5437 ^ n4940 ;
  assign n7305 = n7304 ^ n7303 ^ n7302 ;
  assign n7306 = ( n3630 & ~n5842 ) | ( n3630 & n6613 ) | ( ~n5842 & n6613 ) ;
  assign n7307 = n7306 ^ n3323 ^ n3002 ;
  assign n7308 = n7307 ^ n7264 ^ n1938 ;
  assign n7314 = n6395 ^ n6012 ^ 1'b0 ;
  assign n7309 = n3242 ^ n2199 ^ n1305 ;
  assign n7310 = ~n3631 & n4216 ;
  assign n7311 = n3303 | n7310 ;
  assign n7312 = ( n1705 & n7309 ) | ( n1705 & ~n7311 ) | ( n7309 & ~n7311 ) ;
  assign n7313 = ( n3452 & n5587 ) | ( n3452 & ~n7312 ) | ( n5587 & ~n7312 ) ;
  assign n7315 = n7314 ^ n7313 ^ 1'b0 ;
  assign n7317 = ( ~n418 & n2779 ) | ( ~n418 & n5280 ) | ( n2779 & n5280 ) ;
  assign n7316 = ( n2124 & n4291 ) | ( n2124 & n5875 ) | ( n4291 & n5875 ) ;
  assign n7318 = n7317 ^ n7316 ^ n4496 ;
  assign n7319 = n3146 & n7318 ;
  assign n7321 = n5932 ^ n1156 ^ x122 ;
  assign n7322 = ( n1241 & n4888 ) | ( n1241 & n7321 ) | ( n4888 & n7321 ) ;
  assign n7323 = n6529 & n7322 ;
  assign n7324 = ~x56 & n7323 ;
  assign n7320 = n4449 & n6342 ;
  assign n7325 = n7324 ^ n7320 ^ 1'b0 ;
  assign n7326 = ( x220 & ~n2945 ) | ( x220 & n5352 ) | ( ~n2945 & n5352 ) ;
  assign n7327 = n5893 & n6069 ;
  assign n7328 = ( n3474 & ~n7326 ) | ( n3474 & n7327 ) | ( ~n7326 & n7327 ) ;
  assign n7329 = ( n1209 & n1665 ) | ( n1209 & ~n7328 ) | ( n1665 & ~n7328 ) ;
  assign n7330 = ( n6312 & ~n7315 ) | ( n6312 & n7329 ) | ( ~n7315 & n7329 ) ;
  assign n7331 = x67 & ~n1504 ;
  assign n7332 = ( ~n5108 & n5383 ) | ( ~n5108 & n7331 ) | ( n5383 & n7331 ) ;
  assign n7342 = ( n1558 & n2745 ) | ( n1558 & n3303 ) | ( n2745 & n3303 ) ;
  assign n7343 = ( x207 & ~n5904 ) | ( x207 & n7342 ) | ( ~n5904 & n7342 ) ;
  assign n7333 = n5202 & ~n5808 ;
  assign n7334 = n945 | n1920 ;
  assign n7335 = n7334 ^ n1250 ^ 1'b0 ;
  assign n7336 = n1340 & ~n5328 ;
  assign n7337 = n7336 ^ n7250 ^ 1'b0 ;
  assign n7338 = ~n3265 & n7337 ;
  assign n7339 = ( ~n482 & n7335 ) | ( ~n482 & n7338 ) | ( n7335 & n7338 ) ;
  assign n7340 = ( n501 & n1820 ) | ( n501 & ~n7339 ) | ( n1820 & ~n7339 ) ;
  assign n7341 = ( n1967 & n7333 ) | ( n1967 & n7340 ) | ( n7333 & n7340 ) ;
  assign n7344 = n7343 ^ n7341 ^ 1'b0 ;
  assign n7345 = n2562 & ~n5024 ;
  assign n7346 = n7345 ^ n600 ^ 1'b0 ;
  assign n7347 = n4875 ^ n3173 ^ 1'b0 ;
  assign n7348 = n6861 ^ n4682 ^ n3393 ;
  assign n7349 = n6028 | n7348 ;
  assign n7350 = n1433 & ~n7349 ;
  assign n7351 = n7347 & n7350 ;
  assign n7352 = n7351 ^ n4418 ^ n1519 ;
  assign n7353 = n2389 ^ n648 ^ 1'b0 ;
  assign n7354 = ~n1127 & n5600 ;
  assign n7355 = n5294 ^ n1549 ^ n345 ;
  assign n7356 = n7354 | n7355 ;
  assign n7357 = n7353 | n7356 ;
  assign n7358 = n7357 ^ n2661 ^ n346 ;
  assign n7361 = n2277 ^ n2202 ^ n600 ;
  assign n7362 = n854 & n7361 ;
  assign n7359 = n6372 ^ n4815 ^ n3881 ;
  assign n7360 = n7359 ^ n5998 ^ 1'b0 ;
  assign n7363 = n7362 ^ n7360 ^ n2046 ;
  assign n7369 = ( n1046 & n2635 ) | ( n1046 & n3151 ) | ( n2635 & n3151 ) ;
  assign n7364 = ( n1218 & ~n5154 ) | ( n1218 & n5302 ) | ( ~n5154 & n5302 ) ;
  assign n7365 = n4164 & n7364 ;
  assign n7366 = n2272 ^ n993 ^ n522 ;
  assign n7367 = n7366 ^ n5182 ^ 1'b0 ;
  assign n7368 = ( n1856 & n7365 ) | ( n1856 & n7367 ) | ( n7365 & n7367 ) ;
  assign n7370 = n7369 ^ n7368 ^ 1'b0 ;
  assign n7371 = n3578 | n7370 ;
  assign n7372 = n7363 & ~n7371 ;
  assign n7373 = ( n1973 & n5442 ) | ( n1973 & n5996 ) | ( n5442 & n5996 ) ;
  assign n7374 = n872 | n5825 ;
  assign n7375 = n5367 ^ n2993 ^ 1'b0 ;
  assign n7376 = n7375 ^ n2610 ^ 1'b0 ;
  assign n7377 = n7376 ^ n864 ^ 1'b0 ;
  assign n7381 = n2684 ^ n1733 ^ 1'b0 ;
  assign n7382 = n1280 | n7381 ;
  assign n7383 = n6991 ^ n5608 ^ 1'b0 ;
  assign n7384 = n7382 | n7383 ;
  assign n7378 = ( n4554 & ~n6914 ) | ( n4554 & n7176 ) | ( ~n6914 & n7176 ) ;
  assign n7379 = n7378 ^ n7318 ^ n5143 ;
  assign n7380 = x48 & n7379 ;
  assign n7385 = n7384 ^ n7380 ^ 1'b0 ;
  assign n7386 = n2286 ^ n1416 ^ n754 ;
  assign n7387 = ( n6306 & n6611 ) | ( n6306 & ~n7386 ) | ( n6611 & ~n7386 ) ;
  assign n7388 = ( n2712 & ~n3181 ) | ( n2712 & n3598 ) | ( ~n3181 & n3598 ) ;
  assign n7389 = n7388 ^ n3748 ^ n1047 ;
  assign n7390 = n5760 ^ n4444 ^ n1510 ;
  assign n7391 = n3653 & ~n7390 ;
  assign n7392 = n788 & n7391 ;
  assign n7393 = ( ~n704 & n2510 ) | ( ~n704 & n2617 ) | ( n2510 & n2617 ) ;
  assign n7394 = n2989 ^ n2413 ^ 1'b0 ;
  assign n7395 = n3725 & ~n7394 ;
  assign n7396 = ~n2305 & n3212 ;
  assign n7397 = n3538 & n7396 ;
  assign n7398 = ( x10 & n2694 ) | ( x10 & n7397 ) | ( n2694 & n7397 ) ;
  assign n7399 = n7395 & n7398 ;
  assign n7400 = n7198 & n7399 ;
  assign n7401 = n3043 ^ n2031 ^ n1497 ;
  assign n7402 = ( n2501 & n2641 ) | ( n2501 & n6880 ) | ( n2641 & n6880 ) ;
  assign n7403 = ( ~n1926 & n5178 ) | ( ~n1926 & n7402 ) | ( n5178 & n7402 ) ;
  assign n7404 = n3476 & n7403 ;
  assign n7405 = ( n4166 & n7401 ) | ( n4166 & n7404 ) | ( n7401 & n7404 ) ;
  assign n7406 = ~n7400 & n7405 ;
  assign n7407 = n7406 ^ x141 ^ 1'b0 ;
  assign n7408 = n7393 & ~n7407 ;
  assign n7409 = n7392 & n7408 ;
  assign n7410 = n4282 ^ x140 ^ 1'b0 ;
  assign n7411 = ~n1546 & n7410 ;
  assign n7412 = n7411 ^ n4527 ^ n925 ;
  assign n7413 = ~n5623 & n7412 ;
  assign n7414 = n7085 ^ n6646 ^ n3915 ;
  assign n7415 = n7414 ^ n3234 ^ n2697 ;
  assign n7416 = ( ~n478 & n5884 ) | ( ~n478 & n6234 ) | ( n5884 & n6234 ) ;
  assign n7417 = ( n2046 & n3250 ) | ( n2046 & n5743 ) | ( n3250 & n5743 ) ;
  assign n7418 = n7417 ^ n5141 ^ n4685 ;
  assign n7419 = ( n3132 & n7416 ) | ( n3132 & ~n7418 ) | ( n7416 & ~n7418 ) ;
  assign n7420 = n7419 ^ n7135 ^ 1'b0 ;
  assign n7421 = ~n705 & n7420 ;
  assign n7422 = n4198 ^ n2079 ^ 1'b0 ;
  assign n7423 = n5458 | n7422 ;
  assign n7424 = ( n7222 & n7421 ) | ( n7222 & ~n7423 ) | ( n7421 & ~n7423 ) ;
  assign n7433 = x75 & ~n1240 ;
  assign n7434 = n1527 & n7433 ;
  assign n7431 = n5722 ^ n339 ^ 1'b0 ;
  assign n7432 = n312 & n7431 ;
  assign n7435 = n7434 ^ n7432 ^ n4318 ;
  assign n7425 = ( n2996 & n3363 ) | ( n2996 & ~n4548 ) | ( n3363 & ~n4548 ) ;
  assign n7426 = n4795 | n7425 ;
  assign n7427 = x166 & ~n2272 ;
  assign n7428 = ~n2257 & n7427 ;
  assign n7429 = n7428 ^ n3974 ^ n3912 ;
  assign n7430 = ( n3004 & n7426 ) | ( n3004 & ~n7429 ) | ( n7426 & ~n7429 ) ;
  assign n7436 = n7435 ^ n7430 ^ n6752 ;
  assign n7437 = n2189 ^ n597 ^ n459 ;
  assign n7438 = n7437 ^ n3911 ^ n1880 ;
  assign n7452 = n537 ^ x230 ^ x73 ;
  assign n7453 = n7452 ^ n3157 ^ 1'b0 ;
  assign n7454 = x254 & ~n7453 ;
  assign n7449 = ~n1101 & n2260 ;
  assign n7439 = n3248 ^ n2516 ^ n502 ;
  assign n7440 = ( n1325 & ~n2707 ) | ( n1325 & n7439 ) | ( ~n2707 & n7439 ) ;
  assign n7441 = ( ~n4002 & n4175 ) | ( ~n4002 & n6535 ) | ( n4175 & n6535 ) ;
  assign n7442 = ( n883 & n2453 ) | ( n883 & n7441 ) | ( n2453 & n7441 ) ;
  assign n7443 = x239 & ~n1642 ;
  assign n7444 = ( n6520 & n7442 ) | ( n6520 & n7443 ) | ( n7442 & n7443 ) ;
  assign n7446 = n3887 | n5216 ;
  assign n7445 = ~n302 & n3695 ;
  assign n7447 = n7446 ^ n7445 ^ n6025 ;
  assign n7448 = ( ~n7440 & n7444 ) | ( ~n7440 & n7447 ) | ( n7444 & n7447 ) ;
  assign n7450 = n7449 ^ n7448 ^ 1'b0 ;
  assign n7451 = n7450 ^ n2305 ^ n835 ;
  assign n7455 = n7454 ^ n7451 ^ n4062 ;
  assign n7465 = ~n3918 & n4757 ;
  assign n7456 = ~n3852 & n4754 ;
  assign n7459 = n2743 | n3804 ;
  assign n7460 = n7459 ^ n3042 ^ 1'b0 ;
  assign n7461 = ( n1320 & n3484 ) | ( n1320 & ~n7460 ) | ( n3484 & ~n7460 ) ;
  assign n7462 = ( n2465 & n4303 ) | ( n2465 & ~n7461 ) | ( n4303 & ~n7461 ) ;
  assign n7457 = n4931 ^ n2895 ^ n534 ;
  assign n7458 = n7457 ^ n7379 ^ n5480 ;
  assign n7463 = n7462 ^ n7458 ^ n4417 ;
  assign n7464 = ( ~x181 & n7456 ) | ( ~x181 & n7463 ) | ( n7456 & n7463 ) ;
  assign n7466 = n7465 ^ n7464 ^ n914 ;
  assign n7467 = ( n1724 & ~n2362 ) | ( n1724 & n7015 ) | ( ~n2362 & n7015 ) ;
  assign n7468 = ( n1954 & n5230 ) | ( n1954 & n7467 ) | ( n5230 & n7467 ) ;
  assign n7469 = n4715 ^ n1578 ^ 1'b0 ;
  assign n7470 = n7469 ^ n1307 ^ 1'b0 ;
  assign n7471 = n7468 & n7470 ;
  assign n7472 = n1729 & n4865 ;
  assign n7473 = n1280 & n7472 ;
  assign n7474 = n6489 ^ n853 ^ 1'b0 ;
  assign n7475 = ~n7473 & n7474 ;
  assign n7476 = ( n2296 & n2356 ) | ( n2296 & n7475 ) | ( n2356 & n7475 ) ;
  assign n7477 = n5800 ^ n908 ^ 1'b0 ;
  assign n7478 = n7476 & n7477 ;
  assign n7479 = n7478 ^ n5756 ^ n2040 ;
  assign n7480 = n5659 ^ n2223 ^ n1565 ;
  assign n7481 = n7480 ^ n7273 ^ 1'b0 ;
  assign n7482 = n5882 | n7481 ;
  assign n7487 = n3525 ^ n1793 ^ n1232 ;
  assign n7483 = ( n2377 & ~n3368 ) | ( n2377 & n4744 ) | ( ~n3368 & n4744 ) ;
  assign n7484 = ~n3735 & n7483 ;
  assign n7485 = ~n1209 & n7484 ;
  assign n7486 = n7485 ^ n5609 ^ n1925 ;
  assign n7488 = n7487 ^ n7486 ^ n6232 ;
  assign n7489 = n904 ^ n863 ^ 1'b0 ;
  assign n7490 = ( n2914 & n3606 ) | ( n2914 & n7489 ) | ( n3606 & n7489 ) ;
  assign n7491 = ( n2627 & n5589 ) | ( n2627 & n7490 ) | ( n5589 & n7490 ) ;
  assign n7502 = n2120 ^ n1688 ^ 1'b0 ;
  assign n7503 = n2635 & n7502 ;
  assign n7501 = n2006 | n2557 ;
  assign n7504 = n7503 ^ n7501 ^ 1'b0 ;
  assign n7494 = n7191 ^ n5488 ^ 1'b0 ;
  assign n7492 = ( ~n1101 & n1229 ) | ( ~n1101 & n1510 ) | ( n1229 & n1510 ) ;
  assign n7493 = ( ~n777 & n3598 ) | ( ~n777 & n7492 ) | ( n3598 & n7492 ) ;
  assign n7495 = n7494 ^ n7493 ^ n1003 ;
  assign n7496 = n4489 ^ n4449 ^ 1'b0 ;
  assign n7497 = n2090 & n7496 ;
  assign n7498 = n7497 ^ n6547 ^ 1'b0 ;
  assign n7499 = n1120 | n7498 ;
  assign n7500 = n7495 | n7499 ;
  assign n7505 = n7504 ^ n7500 ^ n3630 ;
  assign n7509 = ~n1801 & n4697 ;
  assign n7506 = n684 | n2923 ;
  assign n7507 = n6048 & ~n7506 ;
  assign n7508 = n7507 ^ n1464 ^ 1'b0 ;
  assign n7510 = n7509 ^ n7508 ^ 1'b0 ;
  assign n7511 = n4904 & ~n5488 ;
  assign n7512 = n7511 ^ n1297 ^ 1'b0 ;
  assign n7513 = n7512 ^ n6362 ^ 1'b0 ;
  assign n7514 = n7513 ^ n1505 ^ x158 ;
  assign n7515 = n7063 ^ n4434 ^ n4143 ;
  assign n7516 = ( n5658 & n6202 ) | ( n5658 & ~n7515 ) | ( n6202 & ~n7515 ) ;
  assign n7517 = ( n1970 & n7514 ) | ( n1970 & n7516 ) | ( n7514 & n7516 ) ;
  assign n7518 = n7510 | n7517 ;
  assign n7519 = n7518 ^ n7069 ^ 1'b0 ;
  assign n7520 = n4331 ^ n4029 ^ 1'b0 ;
  assign n7521 = ( n2479 & n7009 ) | ( n2479 & n7520 ) | ( n7009 & n7520 ) ;
  assign n7522 = ( n546 & n6722 ) | ( n546 & ~n7521 ) | ( n6722 & ~n7521 ) ;
  assign n7523 = n2105 ^ n1426 ^ n687 ;
  assign n7524 = n6461 & ~n7523 ;
  assign n7525 = n7524 ^ n798 ^ 1'b0 ;
  assign n7526 = n7525 ^ n4404 ^ x71 ;
  assign n7527 = ( n2015 & n2811 ) | ( n2015 & ~n5083 ) | ( n2811 & ~n5083 ) ;
  assign n7528 = n548 & ~n7527 ;
  assign n7529 = ~n7526 & n7528 ;
  assign n7530 = n266 & n1666 ;
  assign n7531 = ( ~n1233 & n4906 ) | ( ~n1233 & n5384 ) | ( n4906 & n5384 ) ;
  assign n7532 = ( n3841 & n5898 ) | ( n3841 & ~n7531 ) | ( n5898 & ~n7531 ) ;
  assign n7533 = x37 & n3561 ;
  assign n7534 = n7533 ^ n3173 ^ 1'b0 ;
  assign n7535 = ( n296 & ~n6344 ) | ( n296 & n7534 ) | ( ~n6344 & n7534 ) ;
  assign n7536 = n6917 ^ n2130 ^ n1846 ;
  assign n7537 = n7536 ^ n3439 ^ 1'b0 ;
  assign n7538 = ~n3351 & n4312 ;
  assign n7539 = n4673 & n7538 ;
  assign n7540 = n3971 ^ n3218 ^ n1737 ;
  assign n7541 = n3130 ^ x229 ^ 1'b0 ;
  assign n7542 = n3026 | n7541 ;
  assign n7543 = n7542 ^ n605 ^ 1'b0 ;
  assign n7544 = n7540 & ~n7543 ;
  assign n7545 = ( ~n1151 & n7539 ) | ( ~n1151 & n7544 ) | ( n7539 & n7544 ) ;
  assign n7546 = ( n4091 & n7537 ) | ( n4091 & ~n7545 ) | ( n7537 & ~n7545 ) ;
  assign n7547 = ~n7535 & n7546 ;
  assign n7548 = n2706 | n6554 ;
  assign n7549 = n7548 ^ n4623 ^ 1'b0 ;
  assign n7550 = ( ~n1997 & n3487 ) | ( ~n1997 & n7549 ) | ( n3487 & n7549 ) ;
  assign n7551 = ( ~x179 & n2036 ) | ( ~x179 & n7176 ) | ( n2036 & n7176 ) ;
  assign n7552 = ~n1891 & n2519 ;
  assign n7553 = ~n4626 & n7552 ;
  assign n7554 = ( n5749 & n7551 ) | ( n5749 & n7553 ) | ( n7551 & n7553 ) ;
  assign n7566 = n6817 ^ n829 ^ n304 ;
  assign n7556 = ( x119 & ~n5697 ) | ( x119 & n6783 ) | ( ~n5697 & n6783 ) ;
  assign n7557 = x159 & ~n4069 ;
  assign n7558 = ~n2546 & n7557 ;
  assign n7559 = n7558 ^ x227 ^ 1'b0 ;
  assign n7560 = ~n7556 & n7559 ;
  assign n7561 = n3039 & n7100 ;
  assign n7562 = n7561 ^ n3230 ^ 1'b0 ;
  assign n7563 = ( ~n4603 & n7100 ) | ( ~n4603 & n7562 ) | ( n7100 & n7562 ) ;
  assign n7564 = n7563 ^ n4630 ^ 1'b0 ;
  assign n7565 = n7560 & n7564 ;
  assign n7567 = n7566 ^ n7565 ^ 1'b0 ;
  assign n7555 = x1 & n931 ;
  assign n7568 = n7567 ^ n7555 ^ 1'b0 ;
  assign n7572 = n7259 ^ n6776 ^ n1327 ;
  assign n7569 = ( n423 & ~n1420 ) | ( n423 & n2233 ) | ( ~n1420 & n2233 ) ;
  assign n7570 = n1616 & ~n7569 ;
  assign n7571 = x234 & n7570 ;
  assign n7573 = n7572 ^ n7571 ^ n7054 ;
  assign n7578 = n2459 | n4944 ;
  assign n7574 = ( x208 & n2786 ) | ( x208 & n3021 ) | ( n2786 & n3021 ) ;
  assign n7575 = n7574 ^ n6409 ^ n1063 ;
  assign n7576 = n7575 ^ n2652 ^ 1'b0 ;
  assign n7577 = x179 & n7576 ;
  assign n7579 = n7578 ^ n7577 ^ n2918 ;
  assign n7580 = ( ~x187 & x188 ) | ( ~x187 & n1425 ) | ( x188 & n1425 ) ;
  assign n7581 = n7580 ^ n3737 ^ n1710 ;
  assign n7582 = ( n2127 & n3291 ) | ( n2127 & n4651 ) | ( n3291 & n4651 ) ;
  assign n7583 = n5833 & n7582 ;
  assign n7584 = n7581 & n7583 ;
  assign n7585 = n2752 ^ n790 ^ n438 ;
  assign n7586 = ( ~x111 & n2564 ) | ( ~x111 & n7585 ) | ( n2564 & n7585 ) ;
  assign n7587 = n7586 ^ n699 ^ 1'b0 ;
  assign n7588 = n2045 & n7587 ;
  assign n7589 = ( x161 & n1764 ) | ( x161 & n7588 ) | ( n1764 & n7588 ) ;
  assign n7590 = n7589 ^ n6954 ^ n1428 ;
  assign n7592 = n4426 ^ n3649 ^ n909 ;
  assign n7591 = n7082 ^ n4152 ^ 1'b0 ;
  assign n7593 = n7592 ^ n7591 ^ n617 ;
  assign n7594 = ( n542 & ~n2156 ) | ( n542 & n5725 ) | ( ~n2156 & n5725 ) ;
  assign n7595 = n7594 ^ n3129 ^ 1'b0 ;
  assign n7596 = n3450 | n7595 ;
  assign n7597 = ~n7593 & n7596 ;
  assign n7598 = n7597 ^ n3191 ^ 1'b0 ;
  assign n7599 = n4326 ^ n1299 ^ 1'b0 ;
  assign n7600 = n2523 ^ n1014 ^ 1'b0 ;
  assign n7601 = ( n1476 & ~n2213 ) | ( n1476 & n2470 ) | ( ~n2213 & n2470 ) ;
  assign n7602 = n7601 ^ n4776 ^ 1'b0 ;
  assign n7603 = n7600 | n7602 ;
  assign n7604 = ~n919 & n5318 ;
  assign n7605 = n7603 & n7604 ;
  assign n7606 = n7605 ^ x173 ^ 1'b0 ;
  assign n7607 = n2028 & n7606 ;
  assign n7608 = ( n2345 & ~n5852 ) | ( n2345 & n6132 ) | ( ~n5852 & n6132 ) ;
  assign n7609 = n5192 | n7608 ;
  assign n7610 = x39 & n5080 ;
  assign n7611 = n7610 ^ n7192 ^ 1'b0 ;
  assign n7612 = n7611 ^ n3427 ^ 1'b0 ;
  assign n7613 = n7609 | n7612 ;
  assign n7614 = ~n2210 & n5481 ;
  assign n7615 = n7613 & n7614 ;
  assign n7616 = n4365 ^ n2443 ^ 1'b0 ;
  assign n7617 = n2618 & ~n7616 ;
  assign n7618 = n7617 ^ n6097 ^ n2270 ;
  assign n7619 = ~n4875 & n7618 ;
  assign n7620 = n7615 & n7619 ;
  assign n7621 = n874 & n2630 ;
  assign n7622 = n7621 ^ n6866 ^ 1'b0 ;
  assign n7623 = n4634 ^ n4250 ^ n2090 ;
  assign n7624 = n7623 ^ n2263 ^ x46 ;
  assign n7626 = x215 & ~n2971 ;
  assign n7627 = ~n5557 & n7626 ;
  assign n7625 = ( x114 & n398 ) | ( x114 & n1709 ) | ( n398 & n1709 ) ;
  assign n7628 = n7627 ^ n7625 ^ n4100 ;
  assign n7629 = n2878 ^ n2426 ^ 1'b0 ;
  assign n7630 = ( n688 & n720 ) | ( n688 & ~n3897 ) | ( n720 & ~n3897 ) ;
  assign n7631 = x107 & ~n7630 ;
  assign n7632 = ~n7629 & n7631 ;
  assign n7633 = n3447 ^ x106 ^ 1'b0 ;
  assign n7634 = ( n4774 & n6146 ) | ( n4774 & ~n7633 ) | ( n6146 & ~n7633 ) ;
  assign n7635 = n1536 ^ n953 ^ 1'b0 ;
  assign n7636 = n7635 ^ n6113 ^ n3408 ;
  assign n7637 = n2811 ^ n475 ^ 1'b0 ;
  assign n7638 = ~n1588 & n4541 ;
  assign n7639 = n7638 ^ n853 ^ 1'b0 ;
  assign n7640 = ( n1067 & n6359 ) | ( n1067 & ~n6687 ) | ( n6359 & ~n6687 ) ;
  assign n7645 = ( n2150 & n2412 ) | ( n2150 & n2670 ) | ( n2412 & n2670 ) ;
  assign n7646 = n974 & ~n7645 ;
  assign n7647 = ~n3285 & n7646 ;
  assign n7648 = n7647 ^ n295 ^ 1'b0 ;
  assign n7649 = n5172 & n7648 ;
  assign n7644 = ( n1695 & n2067 ) | ( n1695 & n2175 ) | ( n2067 & n2175 ) ;
  assign n7641 = ( x168 & n1412 ) | ( x168 & n5133 ) | ( n1412 & n5133 ) ;
  assign n7642 = x244 & n7641 ;
  assign n7643 = n7642 ^ n5599 ^ n374 ;
  assign n7650 = n7649 ^ n7644 ^ n7643 ;
  assign n7651 = ~n983 & n993 ;
  assign n7652 = ( x106 & ~n2086 ) | ( x106 & n7651 ) | ( ~n2086 & n7651 ) ;
  assign n7653 = n7652 ^ n1399 ^ n885 ;
  assign n7654 = ( n5711 & n7062 ) | ( n5711 & ~n7653 ) | ( n7062 & ~n7653 ) ;
  assign n7655 = ( n1703 & n4555 ) | ( n1703 & ~n5910 ) | ( n4555 & ~n5910 ) ;
  assign n7656 = n7302 ^ n7102 ^ n2088 ;
  assign n7657 = n7656 ^ n1464 ^ 1'b0 ;
  assign n7658 = n2482 & ~n7657 ;
  assign n7659 = ~n7655 & n7658 ;
  assign n7669 = n4348 & ~n5383 ;
  assign n7670 = n7669 ^ n4234 ^ 1'b0 ;
  assign n7671 = n7670 ^ n1492 ^ x176 ;
  assign n7667 = ( n1242 & ~n1720 ) | ( n1242 & n2193 ) | ( ~n1720 & n2193 ) ;
  assign n7666 = n3469 ^ n3363 ^ n1806 ;
  assign n7668 = n7667 ^ n7666 ^ n2399 ;
  assign n7662 = n1709 | n3820 ;
  assign n7660 = n6454 & n7264 ;
  assign n7661 = n7660 ^ n7176 ^ 1'b0 ;
  assign n7663 = n7662 ^ n7661 ^ n6915 ;
  assign n7664 = ( x111 & n2598 ) | ( x111 & n3287 ) | ( n2598 & n3287 ) ;
  assign n7665 = ( ~n1868 & n7663 ) | ( ~n1868 & n7664 ) | ( n7663 & n7664 ) ;
  assign n7672 = n7671 ^ n7668 ^ n7665 ;
  assign n7673 = ( ~n2166 & n5991 ) | ( ~n2166 & n7509 ) | ( n5991 & n7509 ) ;
  assign n7674 = n7673 ^ n4255 ^ 1'b0 ;
  assign n7680 = x135 & ~n1099 ;
  assign n7681 = n7680 ^ n880 ^ 1'b0 ;
  assign n7682 = ( n1416 & n6450 ) | ( n1416 & ~n7681 ) | ( n6450 & ~n7681 ) ;
  assign n7683 = n6144 & n7682 ;
  assign n7684 = n2098 & n7683 ;
  assign n7675 = n2659 ^ n1738 ^ n1492 ;
  assign n7676 = n4333 & n7675 ;
  assign n7677 = n1290 | n7676 ;
  assign n7678 = n5329 | n7677 ;
  assign n7679 = ( n4001 & n4694 ) | ( n4001 & n7678 ) | ( n4694 & n7678 ) ;
  assign n7685 = n7684 ^ n7679 ^ n1438 ;
  assign n7686 = n6340 ^ n2408 ^ 1'b0 ;
  assign n7687 = n7686 ^ n5952 ^ 1'b0 ;
  assign n7688 = n6169 & ~n6302 ;
  assign n7689 = ( ~n407 & n7687 ) | ( ~n407 & n7688 ) | ( n7687 & n7688 ) ;
  assign n7690 = ( n378 & n2802 ) | ( n378 & ~n3490 ) | ( n2802 & ~n3490 ) ;
  assign n7691 = n7690 ^ n2377 ^ n891 ;
  assign n7692 = ( n3211 & n4168 ) | ( n3211 & ~n7691 ) | ( n4168 & ~n7691 ) ;
  assign n7693 = n3030 ^ n1419 ^ 1'b0 ;
  assign n7694 = ( ~n3758 & n6527 ) | ( ~n3758 & n7693 ) | ( n6527 & n7693 ) ;
  assign n7695 = n4795 ^ n3429 ^ 1'b0 ;
  assign n7696 = n3393 & n7695 ;
  assign n7697 = n7696 ^ n5607 ^ 1'b0 ;
  assign n7703 = ( x92 & n1668 ) | ( x92 & n2005 ) | ( n1668 & n2005 ) ;
  assign n7698 = n5237 ^ n1292 ^ 1'b0 ;
  assign n7699 = ( n4507 & n6933 ) | ( n4507 & n7698 ) | ( n6933 & n7698 ) ;
  assign n7700 = n7699 ^ n748 ^ x19 ;
  assign n7701 = n7188 & n7700 ;
  assign n7702 = n7701 ^ n481 ^ 1'b0 ;
  assign n7704 = n7703 ^ n7702 ^ 1'b0 ;
  assign n7705 = n574 & ~n7704 ;
  assign n7706 = n3015 ^ n1204 ^ n674 ;
  assign n7707 = n7706 ^ n7448 ^ n3959 ;
  assign n7708 = n1836 & ~n7150 ;
  assign n7709 = ( x125 & ~n922 ) | ( x125 & n4972 ) | ( ~n922 & n4972 ) ;
  assign n7710 = n7709 ^ n956 ^ 1'b0 ;
  assign n7711 = n7708 & n7710 ;
  assign n7712 = ( n3147 & n5164 ) | ( n3147 & ~n7711 ) | ( n5164 & ~n7711 ) ;
  assign n7715 = n2903 ^ n461 ^ 1'b0 ;
  assign n7713 = ( n1058 & n2667 ) | ( n1058 & n2735 ) | ( n2667 & n2735 ) ;
  assign n7714 = n7713 ^ n6952 ^ 1'b0 ;
  assign n7716 = n7715 ^ n7714 ^ 1'b0 ;
  assign n7717 = ~n528 & n7716 ;
  assign n7719 = n1442 ^ n489 ^ 1'b0 ;
  assign n7720 = n913 & n7719 ;
  assign n7718 = n1678 & ~n5604 ;
  assign n7721 = n7720 ^ n7718 ^ 1'b0 ;
  assign n7722 = n7721 ^ x42 ^ 1'b0 ;
  assign n7723 = ( ~n2559 & n3280 ) | ( ~n2559 & n5974 ) | ( n3280 & n5974 ) ;
  assign n7724 = n4372 ^ n3097 ^ n1009 ;
  assign n7725 = n7724 ^ n6626 ^ 1'b0 ;
  assign n7726 = n7723 & n7725 ;
  assign n7727 = ~n7643 & n7726 ;
  assign n7735 = n3235 ^ n1759 ^ n1242 ;
  assign n7729 = n621 & ~n1516 ;
  assign n7730 = ( ~n1463 & n2171 ) | ( ~n1463 & n7729 ) | ( n2171 & n7729 ) ;
  assign n7731 = n817 & ~n7730 ;
  assign n7732 = n7731 ^ n1645 ^ 1'b0 ;
  assign n7728 = x1 | n3399 ;
  assign n7733 = n7732 ^ n7728 ^ n5659 ;
  assign n7734 = ~n5394 & n7733 ;
  assign n7736 = n7735 ^ n7734 ^ 1'b0 ;
  assign n7737 = n3829 | n7736 ;
  assign n7738 = n7327 & ~n7737 ;
  assign n7740 = n2668 ^ n871 ^ x163 ;
  assign n7739 = ( n838 & ~n3117 ) | ( n838 & n4168 ) | ( ~n3117 & n4168 ) ;
  assign n7741 = n7740 ^ n7739 ^ 1'b0 ;
  assign n7742 = n7741 ^ n787 ^ 1'b0 ;
  assign n7743 = n7742 ^ n1251 ^ 1'b0 ;
  assign n7744 = n7743 ^ n5546 ^ 1'b0 ;
  assign n7745 = n7738 | n7744 ;
  assign n7746 = n6352 ^ n4566 ^ 1'b0 ;
  assign n7747 = n6104 ^ n5519 ^ n4781 ;
  assign n7748 = n7746 & ~n7747 ;
  assign n7749 = ( ~n2687 & n2710 ) | ( ~n2687 & n7257 ) | ( n2710 & n7257 ) ;
  assign n7750 = n2950 & ~n3472 ;
  assign n7751 = n7123 & n7750 ;
  assign n7752 = n7751 ^ n7208 ^ 1'b0 ;
  assign n7753 = ~n7749 & n7752 ;
  assign n7754 = n2005 ^ x239 ^ 1'b0 ;
  assign n7755 = n7754 ^ n5580 ^ n277 ;
  assign n7756 = n7421 ^ n2202 ^ n890 ;
  assign n7757 = n3041 & n3624 ;
  assign n7758 = n2141 ^ n973 ^ n665 ;
  assign n7759 = ( ~n2163 & n4705 ) | ( ~n2163 & n5651 ) | ( n4705 & n5651 ) ;
  assign n7760 = ( n5172 & n7758 ) | ( n5172 & n7759 ) | ( n7758 & n7759 ) ;
  assign n7764 = n1668 & n3210 ;
  assign n7761 = n6187 ^ n4955 ^ n4800 ;
  assign n7762 = n5595 & ~n7761 ;
  assign n7763 = n773 & n7762 ;
  assign n7765 = n7764 ^ n7763 ^ n7005 ;
  assign n7766 = n4342 ^ n1939 ^ n1788 ;
  assign n7767 = n529 ^ x197 ^ 1'b0 ;
  assign n7768 = n5206 & n7767 ;
  assign n7769 = ( ~n670 & n2848 ) | ( ~n670 & n7768 ) | ( n2848 & n7768 ) ;
  assign n7770 = ~n7766 & n7769 ;
  assign n7771 = n7770 ^ n5315 ^ 1'b0 ;
  assign n7772 = n4923 & ~n7771 ;
  assign n7778 = ~x145 & n1538 ;
  assign n7779 = n7778 ^ n2002 ^ n912 ;
  assign n7780 = n7779 ^ n7577 ^ n1297 ;
  assign n7773 = x227 & n1672 ;
  assign n7774 = ~n1466 & n7773 ;
  assign n7775 = n7774 ^ n3463 ^ n527 ;
  assign n7776 = ~n5372 & n7775 ;
  assign n7777 = ~n4365 & n7776 ;
  assign n7781 = n7780 ^ n7777 ^ 1'b0 ;
  assign n7782 = n5418 ^ n3407 ^ 1'b0 ;
  assign n7783 = ( n5780 & ~n7781 ) | ( n5780 & n7782 ) | ( ~n7781 & n7782 ) ;
  assign n7784 = ( n2585 & ~n3071 ) | ( n2585 & n6232 ) | ( ~n3071 & n6232 ) ;
  assign n7785 = n979 & n7784 ;
  assign n7786 = ( n974 & ~n6933 ) | ( n974 & n7785 ) | ( ~n6933 & n7785 ) ;
  assign n7787 = n7786 ^ n1707 ^ 1'b0 ;
  assign n7788 = n5579 & n7787 ;
  assign n7789 = ( n3074 & n4156 ) | ( n3074 & ~n6774 ) | ( n4156 & ~n6774 ) ;
  assign n7790 = ~n380 & n4192 ;
  assign n7791 = ( n2176 & ~n2370 ) | ( n2176 & n7461 ) | ( ~n2370 & n7461 ) ;
  assign n7792 = x207 & n1564 ;
  assign n7793 = n4311 ^ n3399 ^ 1'b0 ;
  assign n7794 = n7793 ^ n7230 ^ n3630 ;
  assign n7795 = n7794 ^ n4610 ^ n2565 ;
  assign n7796 = n726 & ~n7795 ;
  assign n7797 = n7796 ^ n7387 ^ 1'b0 ;
  assign n7798 = ( n1153 & ~n2394 ) | ( n1153 & n6177 ) | ( ~n2394 & n6177 ) ;
  assign n7799 = n7798 ^ n4099 ^ n3592 ;
  assign n7800 = n7799 ^ n6550 ^ n2346 ;
  assign n7801 = ( n1735 & n2242 ) | ( n1735 & ~n3184 ) | ( n2242 & ~n3184 ) ;
  assign n7802 = n7801 ^ n3757 ^ n2565 ;
  assign n7803 = n7802 ^ n3817 ^ 1'b0 ;
  assign n7804 = n6190 ^ n5479 ^ n4470 ;
  assign n7805 = n7804 ^ n3023 ^ 1'b0 ;
  assign n7806 = n4685 ^ n4673 ^ 1'b0 ;
  assign n7807 = n5832 & n7806 ;
  assign n7808 = x66 & x103 ;
  assign n7809 = ( n570 & n2730 ) | ( n570 & ~n7808 ) | ( n2730 & ~n7808 ) ;
  assign n7810 = n7809 ^ n3759 ^ n2470 ;
  assign n7811 = n7807 & n7810 ;
  assign n7812 = n7811 ^ n927 ^ 1'b0 ;
  assign n7813 = n3043 ^ n2660 ^ n1113 ;
  assign n7814 = ( ~n3467 & n3853 ) | ( ~n3467 & n7813 ) | ( n3853 & n7813 ) ;
  assign n7815 = n7814 ^ n6630 ^ n4136 ;
  assign n7816 = x42 & ~n716 ;
  assign n7817 = n7816 ^ n1813 ^ 1'b0 ;
  assign n7818 = ( x163 & n496 ) | ( x163 & n686 ) | ( n496 & n686 ) ;
  assign n7819 = ( ~n6691 & n7817 ) | ( ~n6691 & n7818 ) | ( n7817 & n7818 ) ;
  assign n7820 = ( n5587 & ~n7815 ) | ( n5587 & n7819 ) | ( ~n7815 & n7819 ) ;
  assign n7826 = ( n3292 & n5733 ) | ( n3292 & ~n6293 ) | ( n5733 & ~n6293 ) ;
  assign n7824 = n7625 ^ n1062 ^ x206 ;
  assign n7825 = ~n2964 & n7824 ;
  assign n7827 = n7826 ^ n7825 ^ n6505 ;
  assign n7828 = n7827 ^ n4168 ^ n1368 ;
  assign n7821 = n4250 ^ n2586 ^ n598 ;
  assign n7822 = n7821 ^ n2589 ^ 1'b0 ;
  assign n7823 = ( n3917 & n5190 ) | ( n3917 & ~n7822 ) | ( n5190 & ~n7822 ) ;
  assign n7829 = n7828 ^ n7823 ^ x70 ;
  assign n7830 = ( n948 & ~n1661 ) | ( n948 & n2055 ) | ( ~n1661 & n2055 ) ;
  assign n7831 = n2577 ^ n793 ^ 1'b0 ;
  assign n7832 = n7830 & ~n7831 ;
  assign n7836 = n3029 ^ x91 ^ 1'b0 ;
  assign n7837 = ~n5398 & n7836 ;
  assign n7834 = ( n1601 & n1606 ) | ( n1601 & n5398 ) | ( n1606 & n5398 ) ;
  assign n7835 = n7834 ^ n1916 ^ n594 ;
  assign n7838 = n7837 ^ n7835 ^ 1'b0 ;
  assign n7839 = n6087 & n7838 ;
  assign n7833 = ~n5259 & n6132 ;
  assign n7840 = n7839 ^ n7833 ^ 1'b0 ;
  assign n7841 = n7832 & ~n7840 ;
  assign n7842 = n3130 & n7841 ;
  assign n7843 = n7022 ^ n5693 ^ n4391 ;
  assign n7844 = n5086 ^ n2088 ^ n1763 ;
  assign n7845 = n7844 ^ n7571 ^ 1'b0 ;
  assign n7846 = ~n2678 & n4380 ;
  assign n7847 = n6589 & n7846 ;
  assign n7848 = n3519 ^ n3325 ^ 1'b0 ;
  assign n7849 = ( n2866 & n6604 ) | ( n2866 & n7848 ) | ( n6604 & n7848 ) ;
  assign n7858 = n7093 ^ n3410 ^ 1'b0 ;
  assign n7855 = ( x173 & ~n1155 ) | ( x173 & n2632 ) | ( ~n1155 & n2632 ) ;
  assign n7856 = n7855 ^ n4835 ^ 1'b0 ;
  assign n7853 = n5269 ^ n2927 ^ 1'b0 ;
  assign n7850 = n3352 & ~n5479 ;
  assign n7851 = n2950 & n7850 ;
  assign n7852 = n7851 ^ n3116 ^ 1'b0 ;
  assign n7854 = n7853 ^ n7852 ^ n2054 ;
  assign n7857 = n7856 ^ n7854 ^ n5941 ;
  assign n7859 = n7858 ^ n7857 ^ 1'b0 ;
  assign n7860 = n4027 ^ n3896 ^ n1292 ;
  assign n7861 = n6828 ^ n5922 ^ x96 ;
  assign n7862 = n7861 ^ n4437 ^ n555 ;
  assign n7864 = ( n1524 & n2948 ) | ( n1524 & ~n5496 ) | ( n2948 & ~n5496 ) ;
  assign n7865 = n7864 ^ n3276 ^ n2224 ;
  assign n7866 = n7865 ^ n7353 ^ n1683 ;
  assign n7863 = ( n2448 & n3595 ) | ( n2448 & n6529 ) | ( n3595 & n6529 ) ;
  assign n7867 = n7866 ^ n7863 ^ n1222 ;
  assign n7868 = ( n498 & n1437 ) | ( n498 & ~n1643 ) | ( n1437 & ~n1643 ) ;
  assign n7869 = n495 | n3534 ;
  assign n7870 = ( n4933 & n7868 ) | ( n4933 & n7869 ) | ( n7868 & n7869 ) ;
  assign n7871 = ( ~n371 & n5704 ) | ( ~n371 & n7809 ) | ( n5704 & n7809 ) ;
  assign n7872 = ~n4586 & n6075 ;
  assign n7873 = ~n7871 & n7872 ;
  assign n7874 = n7069 ^ n2612 ^ 1'b0 ;
  assign n7875 = ~n7873 & n7874 ;
  assign n7876 = n7641 ^ n1384 ^ n496 ;
  assign n7877 = n1093 & ~n4347 ;
  assign n7878 = n4350 & n7877 ;
  assign n7879 = ( n3814 & n4942 ) | ( n3814 & n7878 ) | ( n4942 & n7878 ) ;
  assign n7880 = ( n1414 & ~n2166 ) | ( n1414 & n7664 ) | ( ~n2166 & n7664 ) ;
  assign n7881 = ( n764 & n1774 ) | ( n764 & ~n2558 ) | ( n1774 & ~n2558 ) ;
  assign n7882 = n4224 | n7881 ;
  assign n7883 = n6212 ^ n2499 ^ n2301 ;
  assign n7884 = n7883 ^ n2516 ^ x158 ;
  assign n7885 = n7884 ^ n7837 ^ n2365 ;
  assign n7886 = n7885 ^ n7027 ^ n3323 ;
  assign n7887 = n5303 ^ n4509 ^ 1'b0 ;
  assign n7888 = ~n2668 & n7887 ;
  assign n7890 = n5622 ^ n5352 ^ n2711 ;
  assign n7889 = n3376 ^ n2857 ^ n2313 ;
  assign n7891 = n7890 ^ n7889 ^ n4840 ;
  assign n7892 = ( ~n280 & n7888 ) | ( ~n280 & n7891 ) | ( n7888 & n7891 ) ;
  assign n7893 = n6690 ^ n1027 ^ 1'b0 ;
  assign n7894 = ~n1568 & n7893 ;
  assign n7895 = ~n2633 & n5373 ;
  assign n7896 = n6265 | n7895 ;
  assign n7898 = n7588 ^ n3919 ^ n1553 ;
  assign n7897 = ( n892 & n2308 ) | ( n892 & n5997 ) | ( n2308 & n5997 ) ;
  assign n7899 = n7898 ^ n7897 ^ 1'b0 ;
  assign n7900 = n383 & ~n7899 ;
  assign n7901 = ( n595 & ~n1890 ) | ( n595 & n7900 ) | ( ~n1890 & n7900 ) ;
  assign n7902 = n5594 & n7901 ;
  assign n7903 = n7902 ^ n1222 ^ 1'b0 ;
  assign n7904 = ( n1113 & ~n4472 ) | ( n1113 & n7903 ) | ( ~n4472 & n7903 ) ;
  assign n7906 = ( n3107 & n3472 ) | ( n3107 & n5931 ) | ( n3472 & n5931 ) ;
  assign n7907 = n7906 ^ n3859 ^ n2514 ;
  assign n7905 = ( ~n1046 & n3703 ) | ( ~n1046 & n5014 ) | ( n3703 & n5014 ) ;
  assign n7908 = n7907 ^ n7905 ^ 1'b0 ;
  assign n7909 = n880 ^ x80 ^ 1'b0 ;
  assign n7910 = n3142 ^ n836 ^ 1'b0 ;
  assign n7911 = ( n4851 & n7909 ) | ( n4851 & ~n7910 ) | ( n7909 & ~n7910 ) ;
  assign n7912 = n6586 & n7911 ;
  assign n7913 = n5572 ^ n3694 ^ 1'b0 ;
  assign n7914 = n4694 ^ x248 ^ 1'b0 ;
  assign n7915 = ( x23 & ~n7313 ) | ( x23 & n7914 ) | ( ~n7313 & n7914 ) ;
  assign n7916 = n4134 ^ n3227 ^ 1'b0 ;
  assign n7917 = n2085 | n7916 ;
  assign n7923 = n3081 ^ x42 ^ 1'b0 ;
  assign n7924 = ~n901 & n7923 ;
  assign n7922 = n4048 ^ n2234 ^ n765 ;
  assign n7925 = n7924 ^ n7922 ^ n4067 ;
  assign n7918 = n3525 ^ n2066 ^ 1'b0 ;
  assign n7919 = n1868 | n7918 ;
  assign n7920 = n910 & ~n7919 ;
  assign n7921 = n2017 & n7920 ;
  assign n7926 = n7925 ^ n7921 ^ 1'b0 ;
  assign n7927 = ( n2610 & n4451 ) | ( n2610 & n7926 ) | ( n4451 & n7926 ) ;
  assign n7936 = n5074 | n5485 ;
  assign n7937 = n7936 ^ n1416 ^ 1'b0 ;
  assign n7928 = ( n1434 & ~n2074 ) | ( n1434 & n2342 ) | ( ~n2074 & n2342 ) ;
  assign n7929 = n3061 | n5849 ;
  assign n7930 = n7928 & ~n7929 ;
  assign n7931 = ~n1016 & n2010 ;
  assign n7932 = n2643 & n7931 ;
  assign n7933 = n7930 | n7932 ;
  assign n7934 = n7933 ^ n6210 ^ 1'b0 ;
  assign n7935 = n3989 & ~n7934 ;
  assign n7938 = n7937 ^ n7935 ^ 1'b0 ;
  assign n7939 = n5991 ^ n3332 ^ n2510 ;
  assign n7940 = ( n1173 & n7572 ) | ( n1173 & ~n7939 ) | ( n7572 & ~n7939 ) ;
  assign n7941 = n3471 & ~n7940 ;
  assign n7948 = ( n1482 & n1668 ) | ( n1482 & ~n3158 ) | ( n1668 & ~n3158 ) ;
  assign n7945 = ~n3060 & n5194 ;
  assign n7946 = n3193 & n7945 ;
  assign n7947 = ( n2365 & ~n3184 ) | ( n2365 & n7946 ) | ( ~n3184 & n7946 ) ;
  assign n7943 = ( n277 & ~n394 ) | ( n277 & n1788 ) | ( ~n394 & n1788 ) ;
  assign n7942 = ( n615 & n3045 ) | ( n615 & n6612 ) | ( n3045 & n6612 ) ;
  assign n7944 = n7943 ^ n7942 ^ n3922 ;
  assign n7949 = n7948 ^ n7947 ^ n7944 ;
  assign n7952 = n2224 ^ n935 ^ x157 ;
  assign n7953 = n4924 ^ n2273 ^ 1'b0 ;
  assign n7954 = n7952 & ~n7953 ;
  assign n7955 = n7954 ^ n5411 ^ n4243 ;
  assign n7950 = ( n707 & n1184 ) | ( n707 & ~n2096 ) | ( n1184 & ~n2096 ) ;
  assign n7951 = n1082 | n7950 ;
  assign n7956 = n7955 ^ n7951 ^ 1'b0 ;
  assign n7957 = ~n973 & n5736 ;
  assign n7958 = n1386 | n3313 ;
  assign n7959 = n7115 | n7958 ;
  assign n7960 = n7959 ^ n3401 ^ 1'b0 ;
  assign n7961 = n4001 | n7960 ;
  assign n7962 = ( n1805 & ~n2011 ) | ( n1805 & n4172 ) | ( ~n2011 & n4172 ) ;
  assign n7963 = ( ~n416 & n4984 ) | ( ~n416 & n5462 ) | ( n4984 & n5462 ) ;
  assign n7964 = ~n2186 & n5763 ;
  assign n7965 = n7964 ^ n3432 ^ 1'b0 ;
  assign n7966 = ~n3210 & n6988 ;
  assign n7967 = n7965 & n7966 ;
  assign n7968 = ( x99 & n2007 ) | ( x99 & n7967 ) | ( n2007 & n7967 ) ;
  assign n7970 = n3431 ^ n2801 ^ x44 ;
  assign n7971 = n2998 ^ n2778 ^ x72 ;
  assign n7972 = ( x126 & n7428 ) | ( x126 & ~n7971 ) | ( n7428 & ~n7971 ) ;
  assign n7973 = ( n5828 & n7970 ) | ( n5828 & n7972 ) | ( n7970 & n7972 ) ;
  assign n7969 = ~n3355 & n4475 ;
  assign n7974 = n7973 ^ n7969 ^ 1'b0 ;
  assign n7975 = n3631 ^ n3530 ^ n488 ;
  assign n7976 = n7975 ^ n1298 ^ 1'b0 ;
  assign n7977 = x38 & ~n7976 ;
  assign n7978 = n1202 | n7366 ;
  assign n7979 = n7978 ^ n5883 ^ 1'b0 ;
  assign n7980 = ( x119 & ~n7977 ) | ( x119 & n7979 ) | ( ~n7977 & n7979 ) ;
  assign n7981 = n5852 ^ n3771 ^ n2378 ;
  assign n7982 = ( ~n3795 & n4746 ) | ( ~n3795 & n7981 ) | ( n4746 & n7981 ) ;
  assign n7983 = n7982 ^ n5425 ^ n2404 ;
  assign n7984 = n5500 ^ n4050 ^ n3074 ;
  assign n7985 = n3649 ^ n1805 ^ 1'b0 ;
  assign n7986 = ( n275 & n7984 ) | ( n275 & n7985 ) | ( n7984 & n7985 ) ;
  assign n7987 = n1995 ^ n1967 ^ n1023 ;
  assign n7988 = ( n5458 & n7147 ) | ( n5458 & ~n7987 ) | ( n7147 & ~n7987 ) ;
  assign n7989 = ( n2444 & ~n2976 ) | ( n2444 & n6434 ) | ( ~n2976 & n6434 ) ;
  assign n7990 = n1272 ^ n664 ^ 1'b0 ;
  assign n7991 = n7990 ^ n1949 ^ n643 ;
  assign n7995 = n2019 ^ n1634 ^ n367 ;
  assign n7992 = n1307 ^ n970 ^ n644 ;
  assign n7993 = n2775 & n7992 ;
  assign n7994 = ~n5481 & n7993 ;
  assign n7996 = n7995 ^ n7994 ^ n2311 ;
  assign n7997 = n7996 ^ n2122 ^ 1'b0 ;
  assign n7998 = n1507 | n2827 ;
  assign n7999 = n3207 | n7998 ;
  assign n8000 = ( ~n5773 & n6318 ) | ( ~n5773 & n7999 ) | ( n6318 & n7999 ) ;
  assign n8001 = n3383 ^ n1616 ^ n1508 ;
  assign n8002 = n2456 ^ n2403 ^ x122 ;
  assign n8003 = n8001 & ~n8002 ;
  assign n8004 = ~n5878 & n8003 ;
  assign n8005 = n5442 | n8004 ;
  assign n8006 = n4539 & ~n8005 ;
  assign n8007 = n2830 | n6392 ;
  assign n8008 = n4312 | n8007 ;
  assign n8009 = ( x110 & n6394 ) | ( x110 & n7188 ) | ( n6394 & n7188 ) ;
  assign n8010 = ( n6143 & n8008 ) | ( n6143 & ~n8009 ) | ( n8008 & ~n8009 ) ;
  assign n8011 = n431 | n6894 ;
  assign n8012 = ( n4563 & n8010 ) | ( n4563 & n8011 ) | ( n8010 & n8011 ) ;
  assign n8013 = ( n2679 & n6918 ) | ( n2679 & ~n8012 ) | ( n6918 & ~n8012 ) ;
  assign n8014 = n5852 ^ n2026 ^ n2006 ;
  assign n8015 = n3723 ^ n3351 ^ n988 ;
  assign n8016 = ( ~n282 & n2662 ) | ( ~n282 & n6560 ) | ( n2662 & n6560 ) ;
  assign n8017 = ( n8014 & n8015 ) | ( n8014 & ~n8016 ) | ( n8015 & ~n8016 ) ;
  assign n8018 = n8017 ^ n4631 ^ n961 ;
  assign n8020 = ( ~n1711 & n3493 ) | ( ~n1711 & n6053 ) | ( n3493 & n6053 ) ;
  assign n8019 = n3732 ^ n2300 ^ n1404 ;
  assign n8021 = n8020 ^ n8019 ^ n1339 ;
  assign n8022 = ( n5731 & n7401 ) | ( n5731 & n8021 ) | ( n7401 & n8021 ) ;
  assign n8023 = ( n1813 & n3780 ) | ( n1813 & ~n6997 ) | ( n3780 & ~n6997 ) ;
  assign n8024 = n7629 ^ n3221 ^ 1'b0 ;
  assign n8025 = n8023 & ~n8024 ;
  assign n8026 = n1858 & n8025 ;
  assign n8027 = ( n3022 & n8022 ) | ( n3022 & n8026 ) | ( n8022 & n8026 ) ;
  assign n8028 = n3184 ^ n2629 ^ n644 ;
  assign n8029 = ~n642 & n1784 ;
  assign n8030 = ~n702 & n8029 ;
  assign n8031 = n8030 ^ n2630 ^ 1'b0 ;
  assign n8032 = n2961 & n5467 ;
  assign n8033 = ~n723 & n8032 ;
  assign n8034 = n7943 ^ n4550 ^ n1759 ;
  assign n8035 = ( n1095 & n3547 ) | ( n1095 & n6712 ) | ( n3547 & n6712 ) ;
  assign n8036 = ( n8033 & n8034 ) | ( n8033 & n8035 ) | ( n8034 & n8035 ) ;
  assign n8037 = n5313 ^ n4465 ^ n1599 ;
  assign n8038 = n1590 | n2100 ;
  assign n8039 = n8037 & n8038 ;
  assign n8040 = n2663 & n2775 ;
  assign n8041 = n8040 ^ n7174 ^ 1'b0 ;
  assign n8042 = n6189 & n8041 ;
  assign n8043 = n3727 ^ n1264 ^ 1'b0 ;
  assign n8044 = n8043 ^ n4077 ^ 1'b0 ;
  assign n8045 = x92 & ~n3311 ;
  assign n8046 = ( n3600 & n8044 ) | ( n3600 & n8045 ) | ( n8044 & n8045 ) ;
  assign n8047 = n1332 ^ n336 ^ 1'b0 ;
  assign n8048 = n8047 ^ n763 ^ x212 ;
  assign n8049 = n606 | n6666 ;
  assign n8050 = n8049 ^ n4627 ^ 1'b0 ;
  assign n8051 = ( ~n4269 & n8048 ) | ( ~n4269 & n8050 ) | ( n8048 & n8050 ) ;
  assign n8052 = n4954 ^ n2365 ^ x150 ;
  assign n8053 = ( n306 & n5565 ) | ( n306 & n6595 ) | ( n5565 & n6595 ) ;
  assign n8060 = n3062 ^ n1109 ^ 1'b0 ;
  assign n8061 = n4147 | n8060 ;
  assign n8062 = n8061 ^ n5581 ^ n2179 ;
  assign n8063 = n2977 & n8062 ;
  assign n8064 = ( ~n1568 & n3761 ) | ( ~n1568 & n8063 ) | ( n3761 & n8063 ) ;
  assign n8056 = n1898 ^ n1655 ^ 1'b0 ;
  assign n8057 = n3973 | n8056 ;
  assign n8058 = n8057 ^ n1223 ^ 1'b0 ;
  assign n8054 = n321 | n430 ;
  assign n8055 = n8054 ^ n7185 ^ n2015 ;
  assign n8059 = n8058 ^ n8055 ^ n2433 ;
  assign n8065 = n8064 ^ n8059 ^ 1'b0 ;
  assign n8066 = n5243 ^ n2107 ^ x32 ;
  assign n8067 = ( n981 & n1780 ) | ( n981 & n4132 ) | ( n1780 & n4132 ) ;
  assign n8068 = ( ~n1755 & n4081 ) | ( ~n1755 & n8067 ) | ( n4081 & n8067 ) ;
  assign n8069 = ~n4234 & n8068 ;
  assign n8070 = n5364 & ~n7166 ;
  assign n8071 = n6771 & n8070 ;
  assign n8072 = n8069 | n8071 ;
  assign n8073 = ~x225 & n2833 ;
  assign n8074 = n8073 ^ n4870 ^ n823 ;
  assign n8075 = ( n2326 & n5264 ) | ( n2326 & n6783 ) | ( n5264 & n6783 ) ;
  assign n8076 = n8075 ^ n6408 ^ 1'b0 ;
  assign n8077 = n3242 ^ n2581 ^ n725 ;
  assign n8078 = ~n3221 & n8077 ;
  assign n8079 = n4705 | n8078 ;
  assign n8080 = n3765 & ~n6824 ;
  assign n8081 = n3525 ^ n2526 ^ n2389 ;
  assign n8082 = n8081 ^ n4922 ^ n2648 ;
  assign n8092 = n5249 ^ n5187 ^ n4470 ;
  assign n8083 = n4466 ^ n487 ^ 1'b0 ;
  assign n8084 = n1809 | n3303 ;
  assign n8085 = n8084 ^ x189 ^ 1'b0 ;
  assign n8086 = n8085 ^ n7729 ^ n6712 ;
  assign n8087 = n8086 ^ n2083 ^ n578 ;
  assign n8088 = n8087 ^ n6217 ^ 1'b0 ;
  assign n8089 = n8088 ^ n6447 ^ n4824 ;
  assign n8090 = ( n1789 & ~n8083 ) | ( n1789 & n8089 ) | ( ~n8083 & n8089 ) ;
  assign n8091 = n5725 & ~n8090 ;
  assign n8093 = n8092 ^ n8091 ^ 1'b0 ;
  assign n8094 = ( ~x7 & n2650 ) | ( ~x7 & n3074 ) | ( n2650 & n3074 ) ;
  assign n8095 = n8094 ^ n5203 ^ n2612 ;
  assign n8096 = n1372 & ~n2704 ;
  assign n8097 = ~n3877 & n8096 ;
  assign n8098 = ( n1590 & n8095 ) | ( n1590 & n8097 ) | ( n8095 & n8097 ) ;
  assign n8101 = n7728 ^ n3858 ^ 1'b0 ;
  assign n8102 = n3517 & ~n8101 ;
  assign n8103 = n4579 & n8102 ;
  assign n8104 = n8103 ^ n5149 ^ 1'b0 ;
  assign n8099 = n6042 ^ n4787 ^ n286 ;
  assign n8100 = n8099 ^ n7629 ^ 1'b0 ;
  assign n8105 = n8104 ^ n8100 ^ 1'b0 ;
  assign n8106 = n4131 & ~n8105 ;
  assign n8107 = n4311 ^ n2561 ^ 1'b0 ;
  assign n8108 = ( n573 & n2008 ) | ( n573 & ~n3487 ) | ( n2008 & ~n3487 ) ;
  assign n8109 = ( n7234 & n8107 ) | ( n7234 & ~n8108 ) | ( n8107 & ~n8108 ) ;
  assign n8110 = ( ~n2846 & n7028 ) | ( ~n2846 & n8109 ) | ( n7028 & n8109 ) ;
  assign n8111 = ~x44 & n1247 ;
  assign n8112 = n4092 & n6745 ;
  assign n8113 = n7850 & n8112 ;
  assign n8114 = n3094 & n8113 ;
  assign n8115 = n6491 & n8114 ;
  assign n8118 = n2047 & n2059 ;
  assign n8119 = n8118 ^ n1377 ^ 1'b0 ;
  assign n8116 = ( x118 & n1514 ) | ( x118 & ~n6359 ) | ( n1514 & ~n6359 ) ;
  assign n8117 = ( n4859 & ~n5498 ) | ( n4859 & n8116 ) | ( ~n5498 & n8116 ) ;
  assign n8120 = n8119 ^ n8117 ^ n3033 ;
  assign n8121 = ( ~n8111 & n8115 ) | ( ~n8111 & n8120 ) | ( n8115 & n8120 ) ;
  assign n8123 = n5607 ^ n1407 ^ 1'b0 ;
  assign n8122 = n6430 ^ n5724 ^ n2559 ;
  assign n8124 = n8123 ^ n8122 ^ n5817 ;
  assign n8125 = ( n1972 & ~n6301 ) | ( n1972 & n8124 ) | ( ~n6301 & n8124 ) ;
  assign n8128 = n1232 ^ n1215 ^ n470 ;
  assign n8129 = n846 & ~n8128 ;
  assign n8130 = n8129 ^ n1500 ^ 1'b0 ;
  assign n8126 = n5991 ^ n856 ^ 1'b0 ;
  assign n8127 = n8126 ^ n4265 ^ n2199 ;
  assign n8131 = n8130 ^ n8127 ^ 1'b0 ;
  assign n8132 = n619 | n8131 ;
  assign n8135 = x142 & n1087 ;
  assign n8136 = n8135 ^ n2084 ^ n1058 ;
  assign n8133 = n2931 ^ n1586 ^ n1224 ;
  assign n8134 = n8133 ^ n3078 ^ 1'b0 ;
  assign n8137 = n8136 ^ n8134 ^ n5948 ;
  assign n8138 = n2960 ^ n1763 ^ n1035 ;
  assign n8139 = n8138 ^ n7209 ^ 1'b0 ;
  assign n8140 = n3067 ^ n1884 ^ 1'b0 ;
  assign n8141 = n4533 | n8140 ;
  assign n8142 = n301 | n8141 ;
  assign n8143 = ( n3538 & ~n8139 ) | ( n3538 & n8142 ) | ( ~n8139 & n8142 ) ;
  assign n8144 = n6364 ^ n5672 ^ 1'b0 ;
  assign n8145 = n7809 ^ n5557 ^ 1'b0 ;
  assign n8146 = ( x42 & n3334 ) | ( x42 & ~n8145 ) | ( n3334 & ~n8145 ) ;
  assign n8148 = ~n5458 & n5886 ;
  assign n8149 = n2519 ^ n698 ^ 1'b0 ;
  assign n8150 = ~n2606 & n8149 ;
  assign n8151 = ~n5952 & n8150 ;
  assign n8152 = ~n8148 & n8151 ;
  assign n8147 = ( n1830 & n2538 ) | ( n1830 & ~n7506 ) | ( n2538 & ~n7506 ) ;
  assign n8153 = n8152 ^ n8147 ^ n5076 ;
  assign n8154 = n8153 ^ n6874 ^ n6454 ;
  assign n8164 = ( n427 & ~n3965 ) | ( n427 & n7589 ) | ( ~n3965 & n7589 ) ;
  assign n8155 = n2345 ^ n2162 ^ 1'b0 ;
  assign n8156 = n8155 ^ n6037 ^ n2737 ;
  assign n8157 = n8156 ^ n2953 ^ n2491 ;
  assign n8158 = ( n1194 & n6926 ) | ( n1194 & ~n8157 ) | ( n6926 & ~n8157 ) ;
  assign n8159 = n2813 ^ n2658 ^ n1167 ;
  assign n8160 = x96 & n8159 ;
  assign n8161 = n8160 ^ n6590 ^ n1657 ;
  assign n8162 = n8158 | n8161 ;
  assign n8163 = n6804 & ~n8162 ;
  assign n8165 = n8164 ^ n8163 ^ n7020 ;
  assign n8169 = ( ~n2017 & n4086 ) | ( ~n2017 & n4566 ) | ( n4086 & n4566 ) ;
  assign n8170 = n8169 ^ n487 ^ 1'b0 ;
  assign n8167 = x128 & ~n2865 ;
  assign n8166 = ~n3948 & n7864 ;
  assign n8168 = n8167 ^ n8166 ^ n4935 ;
  assign n8171 = n8170 ^ n8168 ^ n7071 ;
  assign n8172 = ~x108 & x167 ;
  assign n8173 = ( n1431 & ~n4258 ) | ( n1431 & n8172 ) | ( ~n4258 & n8172 ) ;
  assign n8174 = n8173 ^ n2408 ^ n270 ;
  assign n8175 = n5282 ^ n4223 ^ n1420 ;
  assign n8187 = n4744 ^ n2527 ^ n1539 ;
  assign n8177 = n429 & ~n1459 ;
  assign n8178 = n920 | n1729 ;
  assign n8179 = n1768 | n2599 ;
  assign n8180 = n8178 & ~n8179 ;
  assign n8181 = n6490 ^ n2979 ^ 1'b0 ;
  assign n8182 = n4460 | n8181 ;
  assign n8183 = n8180 | n8182 ;
  assign n8184 = n8177 & ~n8183 ;
  assign n8185 = n3945 ^ n1022 ^ 1'b0 ;
  assign n8186 = n8184 | n8185 ;
  assign n8188 = n8187 ^ n8186 ^ 1'b0 ;
  assign n8176 = n4160 & ~n7596 ;
  assign n8189 = n8188 ^ n8176 ^ 1'b0 ;
  assign n8190 = n5924 ^ n4013 ^ x74 ;
  assign n8191 = ( n2634 & n2984 ) | ( n2634 & ~n8190 ) | ( n2984 & ~n8190 ) ;
  assign n8192 = ~n566 & n8191 ;
  assign n8193 = ~x49 & n8192 ;
  assign n8194 = n8193 ^ n6667 ^ n2701 ;
  assign n8195 = ( n8175 & n8189 ) | ( n8175 & ~n8194 ) | ( n8189 & ~n8194 ) ;
  assign n8197 = ( ~x56 & n3143 ) | ( ~x56 & n4548 ) | ( n3143 & n4548 ) ;
  assign n8196 = n1853 & ~n6210 ;
  assign n8198 = n8197 ^ n8196 ^ n6985 ;
  assign n8199 = n6252 ^ n3213 ^ n1952 ;
  assign n8200 = ( n2139 & ~n2684 ) | ( n2139 & n2818 ) | ( ~n2684 & n2818 ) ;
  assign n8201 = ( n1078 & n2474 ) | ( n1078 & ~n2480 ) | ( n2474 & ~n2480 ) ;
  assign n8202 = n5396 ^ n2895 ^ 1'b0 ;
  assign n8203 = ( n4482 & n8201 ) | ( n4482 & ~n8202 ) | ( n8201 & ~n8202 ) ;
  assign n8204 = n1820 ^ n600 ^ 1'b0 ;
  assign n8205 = n394 & n8204 ;
  assign n8206 = ( ~n2875 & n4225 ) | ( ~n2875 & n4597 ) | ( n4225 & n4597 ) ;
  assign n8207 = n8206 ^ n2766 ^ 1'b0 ;
  assign n8208 = n8205 & n8207 ;
  assign n8209 = ( n2858 & n5478 ) | ( n2858 & n8208 ) | ( n5478 & n8208 ) ;
  assign n8210 = ( n8200 & n8203 ) | ( n8200 & n8209 ) | ( n8203 & n8209 ) ;
  assign n8218 = n3236 ^ n2630 ^ n2057 ;
  assign n8211 = n3742 ^ n1257 ^ x158 ;
  assign n8212 = n5979 ^ n4026 ^ n1399 ;
  assign n8213 = ( n4043 & ~n8211 ) | ( n4043 & n8212 ) | ( ~n8211 & n8212 ) ;
  assign n8214 = n5444 ^ n373 ^ x158 ;
  assign n8215 = n8214 ^ n7885 ^ 1'b0 ;
  assign n8216 = n2644 & n8215 ;
  assign n8217 = n8213 & n8216 ;
  assign n8219 = n8218 ^ n8217 ^ 1'b0 ;
  assign n8220 = ( ~n798 & n2170 ) | ( ~n798 & n2800 ) | ( n2170 & n2800 ) ;
  assign n8221 = n8220 ^ n3282 ^ 1'b0 ;
  assign n8222 = n2521 | n8221 ;
  assign n8223 = ( n2956 & ~n3605 ) | ( n2956 & n6480 ) | ( ~n3605 & n6480 ) ;
  assign n8224 = ~n8222 & n8223 ;
  assign n8225 = n4397 ^ n4297 ^ n3956 ;
  assign n8226 = n5843 ^ n3253 ^ n2926 ;
  assign n8227 = n410 & n1475 ;
  assign n8228 = n8227 ^ x163 ^ 1'b0 ;
  assign n8229 = n4265 ^ n2878 ^ n835 ;
  assign n8230 = ( n531 & n1295 ) | ( n531 & n8229 ) | ( n1295 & n8229 ) ;
  assign n8231 = ( ~n7050 & n8228 ) | ( ~n7050 & n8230 ) | ( n8228 & n8230 ) ;
  assign n8232 = n8226 & n8231 ;
  assign n8233 = n8232 ^ n7286 ^ n2630 ;
  assign n8234 = ( ~n2550 & n6058 ) | ( ~n2550 & n8233 ) | ( n6058 & n8233 ) ;
  assign n8235 = ~n2004 & n8234 ;
  assign n8236 = n3539 & ~n5359 ;
  assign n8237 = n2715 ^ n1982 ^ x158 ;
  assign n8238 = ( ~n3468 & n4326 ) | ( ~n3468 & n8237 ) | ( n4326 & n8237 ) ;
  assign n8239 = n2995 & n3332 ;
  assign n8240 = ( ~n4190 & n8238 ) | ( ~n4190 & n8239 ) | ( n8238 & n8239 ) ;
  assign n8254 = n5843 ^ n2858 ^ n1903 ;
  assign n8255 = n8254 ^ n2277 ^ n1191 ;
  assign n8256 = n1727 & n8255 ;
  assign n8257 = n8256 ^ n2495 ^ 1'b0 ;
  assign n8249 = n5581 ^ n1950 ^ 1'b0 ;
  assign n8250 = n3802 & ~n8249 ;
  assign n8251 = n1680 & n8250 ;
  assign n8252 = ~n1248 & n8251 ;
  assign n8247 = n5526 ^ n5378 ^ 1'b0 ;
  assign n8248 = ( n2208 & ~n6450 ) | ( n2208 & n8247 ) | ( ~n6450 & n8247 ) ;
  assign n8253 = n8252 ^ n8248 ^ 1'b0 ;
  assign n8241 = n2576 ^ n2055 ^ n1312 ;
  assign n8242 = ( n3484 & ~n3797 ) | ( n3484 & n8241 ) | ( ~n3797 & n8241 ) ;
  assign n8243 = n2255 | n8242 ;
  assign n8244 = n2507 & ~n8243 ;
  assign n8245 = n6264 ^ n5349 ^ x190 ;
  assign n8246 = n8244 & ~n8245 ;
  assign n8258 = n8257 ^ n8253 ^ n8246 ;
  assign n8259 = n1607 & n3408 ;
  assign n8260 = n7093 & ~n8259 ;
  assign n8261 = ~n3150 & n8260 ;
  assign n8262 = n8261 ^ n6270 ^ n3588 ;
  assign n8263 = ( x231 & ~n489 ) | ( x231 & n8262 ) | ( ~n489 & n8262 ) ;
  assign n8264 = ( n1152 & ~n1246 ) | ( n1152 & n8001 ) | ( ~n1246 & n8001 ) ;
  assign n8265 = n8264 ^ n5844 ^ n4030 ;
  assign n8266 = n6875 & n7504 ;
  assign n8267 = ~n4122 & n8266 ;
  assign n8268 = ( ~n598 & n3928 ) | ( ~n598 & n6051 ) | ( n3928 & n6051 ) ;
  assign n8269 = ( n2370 & n5490 ) | ( n2370 & ~n8268 ) | ( n5490 & ~n8268 ) ;
  assign n8270 = ( n8265 & n8267 ) | ( n8265 & ~n8269 ) | ( n8267 & ~n8269 ) ;
  assign n8271 = n7344 | n8270 ;
  assign n8272 = n4877 & ~n8271 ;
  assign n8275 = n3309 ^ n751 ^ 1'b0 ;
  assign n8273 = ( n283 & ~n785 ) | ( n283 & n1151 ) | ( ~n785 & n1151 ) ;
  assign n8274 = n8273 ^ n6963 ^ n5108 ;
  assign n8276 = n8275 ^ n8274 ^ n2506 ;
  assign n8285 = x56 & n1332 ;
  assign n8286 = n8285 ^ n4033 ^ n2473 ;
  assign n8287 = n1666 & n8286 ;
  assign n8288 = n8287 ^ n1889 ^ 1'b0 ;
  assign n8281 = ~n1231 & n4800 ;
  assign n8282 = n8281 ^ n2717 ^ 1'b0 ;
  assign n8283 = n8282 ^ n1600 ^ 1'b0 ;
  assign n8277 = ( ~n4341 & n7013 ) | ( ~n4341 & n7174 ) | ( n7013 & n7174 ) ;
  assign n8278 = x140 & ~n2914 ;
  assign n8279 = n8278 ^ n6619 ^ 1'b0 ;
  assign n8280 = n8277 & ~n8279 ;
  assign n8284 = n8283 ^ n8280 ^ 1'b0 ;
  assign n8289 = n8288 ^ n8284 ^ n7930 ;
  assign n8290 = n3986 ^ n2585 ^ n2160 ;
  assign n8291 = n903 & ~n2169 ;
  assign n8292 = n8290 & n8291 ;
  assign n8293 = n7512 ^ n3349 ^ 1'b0 ;
  assign n8294 = n6921 ^ n1129 ^ 1'b0 ;
  assign n8295 = x22 | n7759 ;
  assign n8296 = n8294 & n8295 ;
  assign n8297 = ~n8293 & n8296 ;
  assign n8299 = x12 & ~n1262 ;
  assign n8300 = n3526 & n8299 ;
  assign n8298 = n3126 ^ n2125 ^ n1380 ;
  assign n8301 = n8300 ^ n8298 ^ n3347 ;
  assign n8302 = n8301 ^ n3272 ^ n1672 ;
  assign n8303 = ( n853 & n2947 ) | ( n853 & ~n4499 ) | ( n2947 & ~n4499 ) ;
  assign n8304 = n8303 ^ n5135 ^ n3943 ;
  assign n8305 = n8304 ^ n1787 ^ 1'b0 ;
  assign n8306 = ( n431 & n2626 ) | ( n431 & ~n6143 ) | ( n2626 & ~n6143 ) ;
  assign n8310 = ( ~n775 & n1320 ) | ( ~n775 & n2042 ) | ( n1320 & n2042 ) ;
  assign n8307 = ( n2568 & ~n3029 ) | ( n2568 & n5727 ) | ( ~n3029 & n5727 ) ;
  assign n8308 = n8307 ^ n3811 ^ n2615 ;
  assign n8309 = n7110 & n8308 ;
  assign n8311 = n8310 ^ n8309 ^ 1'b0 ;
  assign n8312 = n8306 | n8311 ;
  assign n8313 = n8312 ^ n6967 ^ 1'b0 ;
  assign n8314 = ~n892 & n8313 ;
  assign n8315 = n8160 & n8314 ;
  assign n8316 = ( n308 & ~n687 ) | ( n308 & n983 ) | ( ~n687 & n983 ) ;
  assign n8317 = n5335 | n5555 ;
  assign n8318 = n8317 ^ n833 ^ 1'b0 ;
  assign n8319 = ( n6757 & ~n8316 ) | ( n6757 & n8318 ) | ( ~n8316 & n8318 ) ;
  assign n8323 = ( n3208 & ~n3265 ) | ( n3208 & n4894 ) | ( ~n3265 & n4894 ) ;
  assign n8322 = n1748 ^ n1589 ^ n1583 ;
  assign n8320 = n3645 & n6349 ;
  assign n8321 = n8320 ^ n7785 ^ 1'b0 ;
  assign n8324 = n8323 ^ n8322 ^ n8321 ;
  assign n8325 = n8324 ^ n7676 ^ n7084 ;
  assign n8326 = n5953 ^ x76 ^ 1'b0 ;
  assign n8327 = ( n4351 & n4363 ) | ( n4351 & n8326 ) | ( n4363 & n8326 ) ;
  assign n8328 = x198 | n8327 ;
  assign n8329 = n8328 ^ n4613 ^ n1265 ;
  assign n8330 = n3691 ^ n2718 ^ 1'b0 ;
  assign n8337 = ( n1371 & ~n2376 ) | ( n1371 & n3399 ) | ( ~n2376 & n3399 ) ;
  assign n8334 = n3542 ^ n1252 ^ 1'b0 ;
  assign n8335 = n6463 & n8334 ;
  assign n8336 = ~n3262 & n8335 ;
  assign n8338 = n8337 ^ n8336 ^ n7101 ;
  assign n8331 = n3540 | n5188 ;
  assign n8332 = n7636 | n8331 ;
  assign n8333 = ~n1999 & n8332 ;
  assign n8339 = n8338 ^ n8333 ^ 1'b0 ;
  assign n8340 = n5171 ^ n3214 ^ n2432 ;
  assign n8345 = ( n1436 & n4735 ) | ( n1436 & n7580 ) | ( n4735 & n7580 ) ;
  assign n8346 = n8345 ^ n2174 ^ 1'b0 ;
  assign n8341 = x186 & n1232 ;
  assign n8342 = ~n4498 & n8341 ;
  assign n8343 = n4049 & n8342 ;
  assign n8344 = n6980 & n8343 ;
  assign n8347 = n8346 ^ n8344 ^ n3043 ;
  assign n8348 = n5425 ^ n4523 ^ 1'b0 ;
  assign n8349 = n6841 ^ n4348 ^ n1953 ;
  assign n8350 = ~n4284 & n5141 ;
  assign n8351 = ~n7799 & n8350 ;
  assign n8352 = ( n8348 & n8349 ) | ( n8348 & ~n8351 ) | ( n8349 & ~n8351 ) ;
  assign n8353 = n4591 & n8352 ;
  assign n8354 = n8353 ^ n4585 ^ 1'b0 ;
  assign n8355 = n6282 ^ n4957 ^ 1'b0 ;
  assign n8356 = n2100 & n2300 ;
  assign n8357 = ( n1805 & ~n6488 ) | ( n1805 & n8356 ) | ( ~n6488 & n8356 ) ;
  assign n8358 = n7920 & ~n8357 ;
  assign n8359 = ~n2394 & n8358 ;
  assign n8360 = n5932 ^ n1459 ^ 1'b0 ;
  assign n8361 = n3764 & n8360 ;
  assign n8362 = n3916 & n8361 ;
  assign n8363 = ~x209 & n1949 ;
  assign n8364 = n8363 ^ n6531 ^ n1508 ;
  assign n8365 = n2818 ^ n1714 ^ n820 ;
  assign n8366 = n570 ^ x212 ^ 1'b0 ;
  assign n8367 = n2069 | n8366 ;
  assign n8369 = ( x152 & n5462 ) | ( x152 & n6074 ) | ( n5462 & n6074 ) ;
  assign n8368 = n595 | n5789 ;
  assign n8370 = n8369 ^ n8368 ^ 1'b0 ;
  assign n8371 = n5271 ^ n681 ^ n538 ;
  assign n8372 = n5674 ^ n3530 ^ n2592 ;
  assign n8373 = n4575 & n8372 ;
  assign n8374 = ( n1998 & n8371 ) | ( n1998 & ~n8373 ) | ( n8371 & ~n8373 ) ;
  assign n8375 = ( n8367 & ~n8370 ) | ( n8367 & n8374 ) | ( ~n8370 & n8374 ) ;
  assign n8376 = ( n1716 & n8365 ) | ( n1716 & n8375 ) | ( n8365 & n8375 ) ;
  assign n8377 = n5196 ^ n3067 ^ n1496 ;
  assign n8378 = n1274 & ~n4094 ;
  assign n8379 = ( n728 & n1870 ) | ( n728 & ~n8378 ) | ( n1870 & ~n8378 ) ;
  assign n8380 = n1650 | n8379 ;
  assign n8381 = n8377 | n8380 ;
  assign n8383 = ( n2288 & ~n2683 ) | ( n2288 & n8273 ) | ( ~n2683 & n8273 ) ;
  assign n8382 = n2319 & ~n6513 ;
  assign n8384 = n8383 ^ n8382 ^ 1'b0 ;
  assign n8385 = n6599 ^ n1052 ^ 1'b0 ;
  assign n8386 = ~n8384 & n8385 ;
  assign n8387 = ( n311 & n5069 ) | ( n311 & n7574 ) | ( n5069 & n7574 ) ;
  assign n8388 = n2324 ^ n1433 ^ 1'b0 ;
  assign n8389 = x124 | n3530 ;
  assign n8390 = n4048 ^ x227 ^ 1'b0 ;
  assign n8391 = ( n1707 & n8389 ) | ( n1707 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8392 = n8391 ^ n4496 ^ n866 ;
  assign n8393 = ~n4621 & n8390 ;
  assign n8394 = n3839 & ~n4574 ;
  assign n8395 = n8394 ^ n3165 ^ 1'b0 ;
  assign n8396 = ~n5488 & n8395 ;
  assign n8397 = n3921 & n8396 ;
  assign n8398 = ( ~n2579 & n3025 ) | ( ~n2579 & n8397 ) | ( n3025 & n8397 ) ;
  assign n8400 = ~n2753 & n3506 ;
  assign n8399 = ( n2767 & ~n7128 ) | ( n2767 & n7193 ) | ( ~n7128 & n7193 ) ;
  assign n8401 = n8400 ^ n8399 ^ n2905 ;
  assign n8402 = ( x47 & n2050 ) | ( x47 & n3448 ) | ( n2050 & n3448 ) ;
  assign n8403 = ( n1339 & n4730 ) | ( n1339 & ~n5248 ) | ( n4730 & ~n5248 ) ;
  assign n8404 = n8402 & n8403 ;
  assign n8405 = ~n8401 & n8404 ;
  assign n8406 = ( ~n8175 & n8398 ) | ( ~n8175 & n8405 ) | ( n8398 & n8405 ) ;
  assign n8407 = n8406 ^ n4538 ^ 1'b0 ;
  assign n8408 = n7849 | n8407 ;
  assign n8409 = ( n760 & n8393 ) | ( n760 & ~n8408 ) | ( n8393 & ~n8408 ) ;
  assign n8412 = ~n732 & n1380 ;
  assign n8410 = n7290 ^ n2045 ^ n1469 ;
  assign n8411 = n8410 ^ n5124 ^ n1490 ;
  assign n8413 = n8412 ^ n8411 ^ n7684 ;
  assign n8417 = ( n1601 & ~n2631 ) | ( n1601 & n3502 ) | ( ~n2631 & n3502 ) ;
  assign n8418 = n8417 ^ n2759 ^ 1'b0 ;
  assign n8414 = ~n3315 & n4576 ;
  assign n8415 = n7506 | n8414 ;
  assign n8416 = n3681 & n8415 ;
  assign n8419 = n8418 ^ n8416 ^ 1'b0 ;
  assign n8420 = n3963 & ~n7763 ;
  assign n8421 = n7240 ^ n5043 ^ 1'b0 ;
  assign n8422 = n8421 ^ n7713 ^ n4022 ;
  assign n8423 = n1351 ^ n1251 ^ n536 ;
  assign n8424 = ( x97 & n5130 ) | ( x97 & ~n8423 ) | ( n5130 & ~n8423 ) ;
  assign n8425 = ( n452 & n2303 ) | ( n452 & n8424 ) | ( n2303 & n8424 ) ;
  assign n8429 = n2241 ^ n750 ^ x81 ;
  assign n8426 = n1155 | n3117 ;
  assign n8427 = ( n519 & n2957 ) | ( n519 & n7017 ) | ( n2957 & n7017 ) ;
  assign n8428 = ( ~n2277 & n8426 ) | ( ~n2277 & n8427 ) | ( n8426 & n8427 ) ;
  assign n8430 = n8429 ^ n8428 ^ 1'b0 ;
  assign n8436 = n5716 ^ n3853 ^ x182 ;
  assign n8437 = ~n5458 & n5739 ;
  assign n8438 = ~n8436 & n8437 ;
  assign n8431 = ( n283 & n2930 ) | ( n283 & n4080 ) | ( n2930 & n4080 ) ;
  assign n8432 = n2342 & n8431 ;
  assign n8433 = n8432 ^ n6040 ^ 1'b0 ;
  assign n8434 = n5564 | n8433 ;
  assign n8435 = ( n1827 & ~n3518 ) | ( n1827 & n8434 ) | ( ~n3518 & n8434 ) ;
  assign n8439 = n8438 ^ n8435 ^ n938 ;
  assign n8440 = n5451 ^ n1628 ^ 1'b0 ;
  assign n8441 = n1080 | n8440 ;
  assign n8442 = n1966 ^ n914 ^ 1'b0 ;
  assign n8443 = n8441 | n8442 ;
  assign n8444 = n8443 ^ n1048 ^ 1'b0 ;
  assign n8445 = n6712 ^ n6207 ^ n3483 ;
  assign n8446 = n8445 ^ n5913 ^ n3029 ;
  assign n8447 = ( ~n1195 & n2382 ) | ( ~n1195 & n7563 ) | ( n2382 & n7563 ) ;
  assign n8448 = ( n1485 & n4638 ) | ( n1485 & ~n8447 ) | ( n4638 & ~n8447 ) ;
  assign n8449 = n8448 ^ n4789 ^ 1'b0 ;
  assign n8450 = n8446 & n8449 ;
  assign n8451 = ( ~n4585 & n5152 ) | ( ~n4585 & n7300 ) | ( n5152 & n7300 ) ;
  assign n8452 = n7315 ^ n6216 ^ 1'b0 ;
  assign n8453 = ~n8451 & n8452 ;
  assign n8454 = ( n341 & ~n2143 ) | ( n341 & n3438 ) | ( ~n2143 & n3438 ) ;
  assign n8455 = n2438 ^ n461 ^ 1'b0 ;
  assign n8456 = n6933 ^ n3685 ^ n555 ;
  assign n8457 = n8455 & n8456 ;
  assign n8458 = ~n8075 & n8457 ;
  assign n8459 = ~n4687 & n8458 ;
  assign n8460 = n8454 | n8459 ;
  assign n8461 = n7333 & ~n8460 ;
  assign n8462 = ( n2317 & n3915 ) | ( n2317 & ~n4368 ) | ( n3915 & ~n4368 ) ;
  assign n8463 = n8456 ^ n8336 ^ n2802 ;
  assign n8464 = n8463 ^ n6752 ^ n6612 ;
  assign n8465 = ( n6119 & n8462 ) | ( n6119 & ~n8464 ) | ( n8462 & ~n8464 ) ;
  assign n8471 = n5117 & ~n6970 ;
  assign n8472 = n8471 ^ n1323 ^ 1'b0 ;
  assign n8473 = n5980 ^ n931 ^ 1'b0 ;
  assign n8474 = n8472 | n8473 ;
  assign n8466 = n7047 ^ n2862 ^ n624 ;
  assign n8467 = ~n2184 & n2363 ;
  assign n8468 = n8467 ^ n3019 ^ 1'b0 ;
  assign n8469 = n8468 ^ n4072 ^ x35 ;
  assign n8470 = ( n5748 & n8466 ) | ( n5748 & ~n8469 ) | ( n8466 & ~n8469 ) ;
  assign n8475 = n8474 ^ n8470 ^ 1'b0 ;
  assign n8476 = n1755 & ~n8475 ;
  assign n8477 = n6546 & n8476 ;
  assign n8478 = n721 & n722 ;
  assign n8479 = ( ~n1635 & n4608 ) | ( ~n1635 & n8478 ) | ( n4608 & n8478 ) ;
  assign n8480 = n3727 ^ n3688 ^ n1337 ;
  assign n8481 = ( ~n3281 & n4626 ) | ( ~n3281 & n8480 ) | ( n4626 & n8480 ) ;
  assign n8482 = n4459 | n7826 ;
  assign n8483 = n8481 & ~n8482 ;
  assign n8484 = n8479 & n8483 ;
  assign n8485 = n2680 & n6634 ;
  assign n8486 = n8484 & n8485 ;
  assign n8488 = n4997 ^ n3915 ^ n3838 ;
  assign n8489 = n3577 & n8488 ;
  assign n8490 = n8489 ^ n6554 ^ 1'b0 ;
  assign n8487 = ( ~n409 & n1701 ) | ( ~n409 & n8031 ) | ( n1701 & n8031 ) ;
  assign n8491 = n8490 ^ n8487 ^ n4512 ;
  assign n8492 = n6139 ^ n1429 ^ n889 ;
  assign n8493 = ( n3275 & ~n3328 ) | ( n3275 & n8492 ) | ( ~n3328 & n8492 ) ;
  assign n8494 = n1406 & ~n1690 ;
  assign n8495 = ( n749 & ~n6841 ) | ( n749 & n8494 ) | ( ~n6841 & n8494 ) ;
  assign n8496 = n3006 & n8315 ;
  assign n8497 = n2309 | n7517 ;
  assign n8498 = n8497 ^ n5481 ^ 1'b0 ;
  assign n8499 = n4293 ^ n2197 ^ n1126 ;
  assign n8500 = n5157 | n5800 ;
  assign n8501 = n8500 ^ n1330 ^ 1'b0 ;
  assign n8502 = n8501 ^ n1446 ^ n566 ;
  assign n8503 = ( n6585 & n8499 ) | ( n6585 & ~n8502 ) | ( n8499 & ~n8502 ) ;
  assign n8504 = ~n694 & n1384 ;
  assign n8505 = ( n2395 & n3002 ) | ( n2395 & ~n5612 ) | ( n3002 & ~n5612 ) ;
  assign n8506 = n8504 & ~n8505 ;
  assign n8507 = n2006 | n8506 ;
  assign n8508 = n8507 ^ n5123 ^ 1'b0 ;
  assign n8509 = n6760 ^ n6324 ^ n2115 ;
  assign n8513 = n2213 ^ n1505 ^ x154 ;
  assign n8512 = ( n928 & ~n1577 ) | ( n928 & n3926 ) | ( ~n1577 & n3926 ) ;
  assign n8510 = ( x173 & ~n1201 ) | ( x173 & n2194 ) | ( ~n1201 & n2194 ) ;
  assign n8511 = ( n649 & ~n5151 ) | ( n649 & n8510 ) | ( ~n5151 & n8510 ) ;
  assign n8514 = n8513 ^ n8512 ^ n8511 ;
  assign n8515 = n7834 ^ n4026 ^ 1'b0 ;
  assign n8516 = ( ~n1887 & n5771 ) | ( ~n1887 & n8515 ) | ( n5771 & n8515 ) ;
  assign n8517 = ( ~n1775 & n7722 ) | ( ~n1775 & n8516 ) | ( n7722 & n8516 ) ;
  assign n8518 = n1213 & ~n3299 ;
  assign n8519 = n3920 & n8518 ;
  assign n8520 = n5612 | n8519 ;
  assign n8521 = ( n2194 & n3523 ) | ( n2194 & n6557 ) | ( n3523 & n6557 ) ;
  assign n8522 = n2271 ^ n528 ^ n458 ;
  assign n8523 = n8521 & ~n8522 ;
  assign n8524 = ( ~n2599 & n8520 ) | ( ~n2599 & n8523 ) | ( n8520 & n8523 ) ;
  assign n8528 = n3673 ^ n1269 ^ x133 ;
  assign n8529 = n2489 | n8528 ;
  assign n8526 = n2679 ^ n2518 ^ n1789 ;
  assign n8525 = n4760 ^ n4015 ^ n916 ;
  assign n8527 = n8526 ^ n8525 ^ n5243 ;
  assign n8530 = n8529 ^ n8527 ^ n7043 ;
  assign n8531 = n2549 & n8530 ;
  assign n8532 = ~n8436 & n8531 ;
  assign n8533 = n1675 ^ n716 ^ 1'b0 ;
  assign n8534 = x36 & n8533 ;
  assign n8535 = n8534 ^ n2544 ^ 1'b0 ;
  assign n8536 = n8535 ^ n3574 ^ n1793 ;
  assign n8537 = n6789 ^ n676 ^ 1'b0 ;
  assign n8538 = n5926 & n8537 ;
  assign n8539 = n8173 ^ n4450 ^ n383 ;
  assign n8540 = ( n4788 & n5830 ) | ( n4788 & n8539 ) | ( n5830 & n8539 ) ;
  assign n8542 = n4665 ^ n4518 ^ n1451 ;
  assign n8543 = n8542 ^ n5732 ^ n1794 ;
  assign n8541 = n2585 ^ n2319 ^ 1'b0 ;
  assign n8544 = n8543 ^ n8541 ^ 1'b0 ;
  assign n8545 = ( ~x152 & n3355 ) | ( ~x152 & n7573 ) | ( n3355 & n7573 ) ;
  assign n8548 = ( n586 & n1736 ) | ( n586 & n3319 ) | ( n1736 & n3319 ) ;
  assign n8549 = n8548 ^ n2837 ^ n2752 ;
  assign n8550 = n8549 ^ n6711 ^ n3056 ;
  assign n8551 = ( n271 & ~n4706 ) | ( n271 & n8550 ) | ( ~n4706 & n8550 ) ;
  assign n8546 = n3416 & n5366 ;
  assign n8547 = n6930 & n8546 ;
  assign n8552 = n8551 ^ n8547 ^ n369 ;
  assign n8553 = n8552 ^ n1680 ^ 1'b0 ;
  assign n8554 = n6700 & ~n8553 ;
  assign n8558 = ~n3492 & n4693 ;
  assign n8557 = ( n1449 & ~n6960 ) | ( n1449 & n8277 ) | ( ~n6960 & n8277 ) ;
  assign n8555 = n4564 | n8402 ;
  assign n8556 = n8555 ^ n8504 ^ n3638 ;
  assign n8559 = n8558 ^ n8557 ^ n8556 ;
  assign n8560 = n8559 ^ n8551 ^ n6564 ;
  assign n8561 = n331 | n5300 ;
  assign n8562 = ( n1987 & n3351 ) | ( n1987 & n8561 ) | ( n3351 & n8561 ) ;
  assign n8563 = ~n8175 & n8562 ;
  assign n8564 = ~n6503 & n8563 ;
  assign n8565 = n8564 ^ n412 ^ 1'b0 ;
  assign n8566 = ( ~n615 & n8560 ) | ( ~n615 & n8565 ) | ( n8560 & n8565 ) ;
  assign n8567 = n7910 ^ n5130 ^ n501 ;
  assign n8568 = n1698 | n8567 ;
  assign n8569 = n8568 ^ n5952 ^ 1'b0 ;
  assign n8570 = n8569 ^ n6348 ^ n5113 ;
  assign n8575 = n8102 ^ n6221 ^ n3184 ;
  assign n8571 = n3551 & ~n4555 ;
  assign n8572 = n2331 | n8571 ;
  assign n8573 = n5129 | n8572 ;
  assign n8574 = ( n5402 & ~n5844 ) | ( n5402 & n8573 ) | ( ~n5844 & n8573 ) ;
  assign n8576 = n8575 ^ n8574 ^ 1'b0 ;
  assign n8577 = ( n1306 & ~n3630 ) | ( n1306 & n8576 ) | ( ~n3630 & n8576 ) ;
  assign n8578 = ( n932 & n8570 ) | ( n932 & n8577 ) | ( n8570 & n8577 ) ;
  assign n8582 = ( x42 & n789 ) | ( x42 & n2827 ) | ( n789 & n2827 ) ;
  assign n8580 = n4145 ^ n2676 ^ n275 ;
  assign n8579 = ~n3651 & n4475 ;
  assign n8581 = n8580 ^ n8579 ^ 1'b0 ;
  assign n8583 = n8582 ^ n8581 ^ 1'b0 ;
  assign n8584 = n3041 ^ n2777 ^ 1'b0 ;
  assign n8585 = n7603 ^ n2843 ^ 1'b0 ;
  assign n8586 = n8585 ^ n3713 ^ n3044 ;
  assign n8587 = n8586 ^ n1072 ^ 1'b0 ;
  assign n8588 = n1072 & ~n8587 ;
  assign n8589 = n5621 & n8588 ;
  assign n8590 = ~n8584 & n8589 ;
  assign n8591 = n8590 ^ n5516 ^ n1957 ;
  assign n8592 = ~n5501 & n6284 ;
  assign n8593 = n8592 ^ n4192 ^ 1'b0 ;
  assign n8597 = n5233 ^ n491 ^ 1'b0 ;
  assign n8598 = ~n6363 & n8597 ;
  assign n8594 = n4180 & ~n4306 ;
  assign n8595 = n8594 ^ n2492 ^ 1'b0 ;
  assign n8596 = ~n2816 & n8595 ;
  assign n8599 = n8598 ^ n8596 ^ 1'b0 ;
  assign n8600 = n1974 | n8599 ;
  assign n8601 = n2947 | n8600 ;
  assign n8602 = n2189 ^ n2160 ^ 1'b0 ;
  assign n8603 = n8602 ^ n5981 ^ n1196 ;
  assign n8604 = n1516 ^ n1304 ^ 1'b0 ;
  assign n8605 = n8603 | n8604 ;
  assign n8606 = ( n4697 & n5654 ) | ( n4697 & n8605 ) | ( n5654 & n8605 ) ;
  assign n8607 = ( n866 & n5613 ) | ( n866 & ~n8606 ) | ( n5613 & ~n8606 ) ;
  assign n8609 = n3286 ^ n1331 ^ x212 ;
  assign n8610 = n1316 & ~n6294 ;
  assign n8611 = ( n407 & ~n1806 ) | ( n407 & n5475 ) | ( ~n1806 & n5475 ) ;
  assign n8612 = ( ~n8609 & n8610 ) | ( ~n8609 & n8611 ) | ( n8610 & n8611 ) ;
  assign n8608 = n2367 & n7912 ;
  assign n8613 = n8612 ^ n8608 ^ 1'b0 ;
  assign n8614 = n4388 ^ n2001 ^ 1'b0 ;
  assign n8615 = ( n2941 & n5348 ) | ( n2941 & n8614 ) | ( n5348 & n8614 ) ;
  assign n8616 = ( n4630 & ~n5040 ) | ( n4630 & n8615 ) | ( ~n5040 & n8615 ) ;
  assign n8617 = n6730 ^ n5230 ^ n536 ;
  assign n8624 = n4123 ^ n1269 ^ 1'b0 ;
  assign n8625 = n1194 | n8624 ;
  assign n8618 = n5165 ^ n4194 ^ n4139 ;
  assign n8620 = n6470 ^ n2255 ^ 1'b0 ;
  assign n8619 = n3371 & ~n7698 ;
  assign n8621 = n8620 ^ n8619 ^ 1'b0 ;
  assign n8622 = n8621 ^ n2506 ^ 1'b0 ;
  assign n8623 = ~n8618 & n8622 ;
  assign n8626 = n8625 ^ n8623 ^ n5289 ;
  assign n8627 = n8617 & n8626 ;
  assign n8635 = n3728 ^ n3453 ^ n2964 ;
  assign n8628 = n5941 ^ n3216 ^ n321 ;
  assign n8629 = ~n3125 & n3424 ;
  assign n8630 = ~n8628 & n8629 ;
  assign n8631 = n1732 | n8630 ;
  assign n8632 = n8631 ^ n6997 ^ 1'b0 ;
  assign n8633 = n8632 ^ n3035 ^ 1'b0 ;
  assign n8634 = ~n6311 & n8633 ;
  assign n8636 = n8635 ^ n8634 ^ n5132 ;
  assign n8637 = n8636 ^ n8626 ^ n7253 ;
  assign n8638 = ( n2580 & n3710 ) | ( n2580 & n6157 ) | ( n3710 & n6157 ) ;
  assign n8639 = ( n3976 & n4576 ) | ( n3976 & ~n6116 ) | ( n4576 & ~n6116 ) ;
  assign n8640 = n2381 ^ n2010 ^ 1'b0 ;
  assign n8641 = ( x65 & n2470 ) | ( x65 & ~n8640 ) | ( n2470 & ~n8640 ) ;
  assign n8642 = n8639 & ~n8641 ;
  assign n8643 = ~n8638 & n8642 ;
  assign n8644 = ( n860 & ~n1949 ) | ( n860 & n6654 ) | ( ~n1949 & n6654 ) ;
  assign n8645 = n3158 ^ n1722 ^ n1589 ;
  assign n8646 = n7075 & ~n8645 ;
  assign n8647 = ( ~n7514 & n8644 ) | ( ~n7514 & n8646 ) | ( n8644 & n8646 ) ;
  assign n8648 = n8647 ^ n4257 ^ n3116 ;
  assign n8655 = ~n3163 & n3619 ;
  assign n8656 = n8655 ^ n749 ^ 1'b0 ;
  assign n8654 = ( n295 & ~n2801 ) | ( n295 & n4196 ) | ( ~n2801 & n4196 ) ;
  assign n8649 = n2792 ^ x114 ^ 1'b0 ;
  assign n8650 = n1407 & ~n4926 ;
  assign n8651 = n8650 ^ n7123 ^ 1'b0 ;
  assign n8652 = ( ~n2158 & n4549 ) | ( ~n2158 & n8651 ) | ( n4549 & n8651 ) ;
  assign n8653 = ( ~n5972 & n8649 ) | ( ~n5972 & n8652 ) | ( n8649 & n8652 ) ;
  assign n8657 = n8656 ^ n8654 ^ n8653 ;
  assign n8658 = n257 ^ x160 ^ 1'b0 ;
  assign n8659 = x56 & n8658 ;
  assign n8660 = ( n3833 & ~n8228 ) | ( n3833 & n8659 ) | ( ~n8228 & n8659 ) ;
  assign n8661 = ( n430 & ~n4910 ) | ( n430 & n8660 ) | ( ~n4910 & n8660 ) ;
  assign n8662 = ( ~n556 & n1794 ) | ( ~n556 & n8505 ) | ( n1794 & n8505 ) ;
  assign n8663 = n8662 ^ n7530 ^ n4682 ;
  assign n8664 = ( n3858 & ~n8269 ) | ( n3858 & n8345 ) | ( ~n8269 & n8345 ) ;
  assign n8665 = n5656 & n7999 ;
  assign n8666 = ~n7483 & n8665 ;
  assign n8670 = ( ~n1977 & n5256 ) | ( ~n1977 & n8335 ) | ( n5256 & n8335 ) ;
  assign n8667 = n4383 & n7074 ;
  assign n8668 = ~n4239 & n8667 ;
  assign n8669 = n8668 ^ n6523 ^ n1807 ;
  assign n8671 = n8670 ^ n8669 ^ n7525 ;
  assign n8672 = ~n6249 & n8529 ;
  assign n8673 = ( n987 & n1636 ) | ( n987 & ~n4260 ) | ( n1636 & ~n4260 ) ;
  assign n8674 = n8673 ^ n5207 ^ n1784 ;
  assign n8675 = ( n2781 & ~n3469 ) | ( n2781 & n8674 ) | ( ~n3469 & n8674 ) ;
  assign n8676 = n1835 ^ n1011 ^ n602 ;
  assign n8677 = n8273 ^ n1852 ^ n1850 ;
  assign n8678 = ~n2557 & n8677 ;
  assign n8679 = ~n8676 & n8678 ;
  assign n8680 = n8679 ^ n4285 ^ 1'b0 ;
  assign n8681 = ( x68 & x172 ) | ( x68 & n2174 ) | ( x172 & n2174 ) ;
  assign n8682 = n8681 ^ n2548 ^ n2142 ;
  assign n8683 = ( n2813 & ~n8680 ) | ( n2813 & n8682 ) | ( ~n8680 & n8682 ) ;
  assign n8684 = n4457 & ~n8550 ;
  assign n8685 = n340 ^ x208 ^ 1'b0 ;
  assign n8686 = ( ~n3415 & n6524 ) | ( ~n3415 & n8685 ) | ( n6524 & n8685 ) ;
  assign n8698 = n1433 ^ n829 ^ 1'b0 ;
  assign n8699 = x62 & ~n8698 ;
  assign n8697 = ( ~n1179 & n3573 ) | ( ~n1179 & n6423 ) | ( n3573 & n6423 ) ;
  assign n8690 = ( n1048 & n2164 ) | ( n1048 & ~n4724 ) | ( n2164 & ~n4724 ) ;
  assign n8691 = n5179 ^ n2559 ^ n1097 ;
  assign n8692 = n5682 ^ n2336 ^ n1921 ;
  assign n8693 = n8692 ^ n3377 ^ 1'b0 ;
  assign n8694 = ~n8691 & n8693 ;
  assign n8695 = n8694 ^ n1031 ^ 1'b0 ;
  assign n8696 = ~n8690 & n8695 ;
  assign n8700 = n8699 ^ n8697 ^ n8696 ;
  assign n8687 = ( n418 & n958 ) | ( n418 & n1824 ) | ( n958 & n1824 ) ;
  assign n8688 = ( ~n407 & n3960 ) | ( ~n407 & n8687 ) | ( n3960 & n8687 ) ;
  assign n8689 = n1596 | n8688 ;
  assign n8701 = n8700 ^ n8689 ^ 1'b0 ;
  assign n8702 = ( n8684 & n8686 ) | ( n8684 & n8701 ) | ( n8686 & n8701 ) ;
  assign n8703 = n5251 ^ n3062 ^ n726 ;
  assign n8704 = ~n3734 & n8703 ;
  assign n8705 = n6535 & n8704 ;
  assign n8706 = n823 & n1688 ;
  assign n8707 = n3800 & n8706 ;
  assign n8708 = n8705 | n8707 ;
  assign n8709 = n8708 ^ n1007 ^ 1'b0 ;
  assign n8711 = ( n831 & n7120 ) | ( n831 & n7990 ) | ( n7120 & n7990 ) ;
  assign n8710 = n6520 ^ n3794 ^ x227 ;
  assign n8712 = n8711 ^ n8710 ^ n3942 ;
  assign n8713 = n5635 ^ n2827 ^ 1'b0 ;
  assign n8714 = n1390 | n8713 ;
  assign n8715 = ~n3643 & n4285 ;
  assign n8716 = n8714 & n8715 ;
  assign n8717 = n603 ^ n329 ^ 1'b0 ;
  assign n8718 = n6383 ^ n1514 ^ n1379 ;
  assign n8719 = n5484 & n8718 ;
  assign n8720 = n3290 & n8719 ;
  assign n8721 = n3405 ^ n1510 ^ 1'b0 ;
  assign n8722 = ~n8720 & n8721 ;
  assign n8725 = ~n2965 & n6823 ;
  assign n8726 = n8725 ^ n4735 ^ 1'b0 ;
  assign n8723 = n2615 | n3841 ;
  assign n8724 = ( ~n4629 & n6681 ) | ( ~n4629 & n8723 ) | ( n6681 & n8723 ) ;
  assign n8727 = n8726 ^ n8724 ^ n2113 ;
  assign n8728 = n8722 | n8727 ;
  assign n8729 = n8728 ^ n6279 ^ 1'b0 ;
  assign n8730 = n8729 ^ n2303 ^ 1'b0 ;
  assign n8731 = ( x174 & ~n644 ) | ( x174 & n2318 ) | ( ~n644 & n2318 ) ;
  assign n8732 = n8731 ^ n376 ^ x157 ;
  assign n8733 = ( ~n902 & n2332 ) | ( ~n902 & n3031 ) | ( n2332 & n3031 ) ;
  assign n8734 = n8732 | n8733 ;
  assign n8735 = n3254 ^ x99 ^ 1'b0 ;
  assign n8736 = ~n1971 & n8735 ;
  assign n8737 = n3991 ^ n2803 ^ 1'b0 ;
  assign n8738 = ~n3115 & n8737 ;
  assign n8739 = ( n962 & n1330 ) | ( n962 & ~n8738 ) | ( n1330 & ~n8738 ) ;
  assign n8740 = ( n4487 & n5821 ) | ( n4487 & ~n8739 ) | ( n5821 & ~n8739 ) ;
  assign n8741 = ~n6762 & n8740 ;
  assign n8742 = ~n8736 & n8741 ;
  assign n8743 = ( n3959 & ~n6905 ) | ( n3959 & n7189 ) | ( ~n6905 & n7189 ) ;
  assign n8744 = ( n5181 & ~n8742 ) | ( n5181 & n8743 ) | ( ~n8742 & n8743 ) ;
  assign n8745 = n1985 & ~n8744 ;
  assign n8748 = n697 ^ n491 ^ 1'b0 ;
  assign n8749 = n5304 & ~n8748 ;
  assign n8750 = n8749 ^ n5282 ^ 1'b0 ;
  assign n8746 = n3088 & ~n7417 ;
  assign n8747 = n7994 & n8746 ;
  assign n8751 = n8750 ^ n8747 ^ n4169 ;
  assign n8752 = n3958 ^ x52 ^ 1'b0 ;
  assign n8753 = n8752 ^ n6123 ^ 1'b0 ;
  assign n8754 = n6277 & ~n8753 ;
  assign n8755 = n1293 | n6749 ;
  assign n8756 = ( ~n8751 & n8754 ) | ( ~n8751 & n8755 ) | ( n8754 & n8755 ) ;
  assign n8757 = n8756 ^ n8592 ^ n1254 ;
  assign n8758 = ~n4204 & n5521 ;
  assign n8759 = ( n1237 & ~n4139 ) | ( n1237 & n8363 ) | ( ~n4139 & n8363 ) ;
  assign n8760 = n8759 ^ n4986 ^ n3657 ;
  assign n8761 = n640 & n2795 ;
  assign n8762 = ~n1146 & n8761 ;
  assign n8763 = x13 & n4983 ;
  assign n8764 = n8762 & n8763 ;
  assign n8765 = n8760 | n8764 ;
  assign n8766 = n5141 & ~n8429 ;
  assign n8767 = n2999 & n7306 ;
  assign n8768 = n8766 & n8767 ;
  assign n8770 = n4525 ^ n3452 ^ n2390 ;
  assign n8771 = n8770 ^ n7414 ^ n4060 ;
  assign n8769 = n1867 & ~n6992 ;
  assign n8772 = n8771 ^ n8769 ^ n4045 ;
  assign n8773 = n3488 | n4625 ;
  assign n8774 = n5178 & ~n8773 ;
  assign n8775 = n7183 ^ n4850 ^ 1'b0 ;
  assign n8776 = ( n2068 & n8774 ) | ( n2068 & ~n8775 ) | ( n8774 & ~n8775 ) ;
  assign n8777 = ( ~n3851 & n6329 ) | ( ~n3851 & n8549 ) | ( n6329 & n8549 ) ;
  assign n8778 = n2105 | n2217 ;
  assign n8779 = n8777 | n8778 ;
  assign n8780 = n5549 ^ n301 ^ 1'b0 ;
  assign n8781 = n8780 ^ n1491 ^ 1'b0 ;
  assign n8782 = ( n1899 & n4788 ) | ( n1899 & ~n8781 ) | ( n4788 & ~n8781 ) ;
  assign n8783 = ( n6470 & n8779 ) | ( n6470 & ~n8782 ) | ( n8779 & ~n8782 ) ;
  assign n8784 = ( n286 & ~n803 ) | ( n286 & n1433 ) | ( ~n803 & n1433 ) ;
  assign n8785 = n8784 ^ x68 ^ 1'b0 ;
  assign n8786 = n8783 & ~n8785 ;
  assign n8792 = n1422 ^ n501 ^ n485 ;
  assign n8793 = ( n6361 & ~n6839 ) | ( n6361 & n8792 ) | ( ~n6839 & n8792 ) ;
  assign n8789 = n5767 ^ n5716 ^ n2343 ;
  assign n8788 = n2923 & n2962 ;
  assign n8790 = n8789 ^ n8788 ^ 1'b0 ;
  assign n8787 = n3998 | n7361 ;
  assign n8791 = n8790 ^ n8787 ^ 1'b0 ;
  assign n8794 = n8793 ^ n8791 ^ n3130 ;
  assign n8795 = n7015 & n7419 ;
  assign n8796 = n459 & n8795 ;
  assign n8797 = n4015 | n8796 ;
  assign n8798 = n8797 ^ n3653 ^ 1'b0 ;
  assign n8799 = n4679 ^ n1924 ^ n393 ;
  assign n8802 = n324 & ~n815 ;
  assign n8803 = n8802 ^ n5896 ^ n4100 ;
  assign n8800 = ( n2686 & n6439 ) | ( n2686 & ~n7403 ) | ( n6439 & ~n7403 ) ;
  assign n8801 = ~n5358 & n8800 ;
  assign n8804 = n8803 ^ n8801 ^ 1'b0 ;
  assign n8805 = ( n5423 & n8799 ) | ( n5423 & n8804 ) | ( n8799 & n8804 ) ;
  assign n8806 = n6024 ^ n5723 ^ n1119 ;
  assign n8807 = n3258 ^ n765 ^ 1'b0 ;
  assign n8808 = n5434 & ~n8807 ;
  assign n8809 = n1520 & n3678 ;
  assign n8810 = ( ~n1778 & n1835 ) | ( ~n1778 & n3377 ) | ( n1835 & n3377 ) ;
  assign n8811 = n5599 | n8810 ;
  assign n8812 = n1706 | n2053 ;
  assign n8813 = n936 | n8812 ;
  assign n8814 = n8231 ^ n4830 ^ n669 ;
  assign n8815 = n8813 & n8814 ;
  assign n8816 = n2362 & n8815 ;
  assign n8817 = n8816 ^ n7301 ^ 1'b0 ;
  assign n8828 = ( ~x205 & n2135 ) | ( ~x205 & n2189 ) | ( n2135 & n2189 ) ;
  assign n8829 = x171 | n8828 ;
  assign n8821 = n1101 & n3332 ;
  assign n8822 = n8821 ^ n1544 ^ 1'b0 ;
  assign n8823 = ~n1735 & n8822 ;
  assign n8824 = n7673 & n8823 ;
  assign n8825 = ( n823 & ~n2614 ) | ( n823 & n8824 ) | ( ~n2614 & n8824 ) ;
  assign n8826 = n8825 ^ n2506 ^ 1'b0 ;
  assign n8818 = n6087 ^ n4517 ^ n1248 ;
  assign n8819 = ( n1225 & n3976 ) | ( n1225 & ~n8818 ) | ( n3976 & ~n8818 ) ;
  assign n8820 = ( n424 & ~n7029 ) | ( n424 & n8819 ) | ( ~n7029 & n8819 ) ;
  assign n8827 = n8826 ^ n8820 ^ n3808 ;
  assign n8830 = n8829 ^ n8827 ^ n5021 ;
  assign n8831 = ( ~n4729 & n5648 ) | ( ~n4729 & n8677 ) | ( n5648 & n8677 ) ;
  assign n8832 = n3301 | n5464 ;
  assign n8833 = n2810 & ~n8832 ;
  assign n8834 = ( ~n2976 & n3767 ) | ( ~n2976 & n8833 ) | ( n3767 & n8833 ) ;
  assign n8835 = ( n390 & ~n6037 ) | ( n390 & n8834 ) | ( ~n6037 & n8834 ) ;
  assign n8836 = ~n891 & n2735 ;
  assign n8837 = n8836 ^ x207 ^ 1'b0 ;
  assign n8838 = n8835 & ~n8837 ;
  assign n8839 = n3866 ^ n3524 ^ n525 ;
  assign n8840 = n8839 ^ n4636 ^ n1418 ;
  assign n8841 = ( n278 & n3956 ) | ( n278 & n8840 ) | ( n3956 & n8840 ) ;
  assign n8842 = n8841 ^ n2290 ^ n1938 ;
  assign n8843 = n763 & ~n8842 ;
  assign n8844 = n3319 ^ n3188 ^ n1490 ;
  assign n8845 = n8844 ^ n6967 ^ 1'b0 ;
  assign n8846 = n8845 ^ n8208 ^ n6838 ;
  assign n8847 = ( n1244 & n4156 ) | ( n1244 & ~n8846 ) | ( n4156 & ~n8846 ) ;
  assign n8848 = n8400 ^ n4327 ^ 1'b0 ;
  assign n8849 = n5371 & n6081 ;
  assign n8850 = n2244 & n8849 ;
  assign n8851 = n8850 ^ n4772 ^ 1'b0 ;
  assign n8852 = n5286 ^ n4694 ^ n4486 ;
  assign n8853 = n2509 | n4945 ;
  assign n8854 = n8853 ^ n2688 ^ 1'b0 ;
  assign n8855 = n8854 ^ n6654 ^ n1635 ;
  assign n8856 = n8855 ^ n6029 ^ 1'b0 ;
  assign n8866 = ( x75 & n633 ) | ( x75 & ~n698 ) | ( n633 & ~n698 ) ;
  assign n8867 = n8866 ^ n3235 ^ 1'b0 ;
  assign n8861 = ( x90 & n283 ) | ( x90 & n3922 ) | ( n283 & n3922 ) ;
  assign n8862 = n7740 ^ n3862 ^ n1562 ;
  assign n8863 = n8862 ^ n5912 ^ 1'b0 ;
  assign n8864 = n8861 | n8863 ;
  assign n8858 = x32 & ~n2740 ;
  assign n8859 = n6053 & n8858 ;
  assign n8857 = x70 & n6270 ;
  assign n8860 = n8859 ^ n8857 ^ 1'b0 ;
  assign n8865 = n8864 ^ n8860 ^ x73 ;
  assign n8868 = n8867 ^ n8865 ^ n3397 ;
  assign n8869 = n2183 ^ n1219 ^ n1054 ;
  assign n8870 = n8869 ^ n1517 ^ n918 ;
  assign n8871 = ( ~n892 & n3002 ) | ( ~n892 & n8870 ) | ( n3002 & n8870 ) ;
  assign n8872 = ( n1254 & n2369 ) | ( n1254 & ~n2964 ) | ( n2369 & ~n2964 ) ;
  assign n8873 = ( n4736 & n5103 ) | ( n4736 & ~n8872 ) | ( n5103 & ~n8872 ) ;
  assign n8874 = n6684 ^ n5224 ^ n750 ;
  assign n8875 = n6750 ^ n5596 ^ n2728 ;
  assign n8876 = ~n8874 & n8875 ;
  assign n8877 = n8876 ^ n6111 ^ 1'b0 ;
  assign n8878 = ( n8871 & ~n8873 ) | ( n8871 & n8877 ) | ( ~n8873 & n8877 ) ;
  assign n8879 = n8878 ^ n3949 ^ 1'b0 ;
  assign n8880 = n928 & n8879 ;
  assign n8881 = n4342 & ~n8182 ;
  assign n8882 = n8881 ^ n3455 ^ n627 ;
  assign n8883 = ~n334 & n1327 ;
  assign n8884 = n8883 ^ n2797 ^ 1'b0 ;
  assign n8885 = ~n3306 & n8884 ;
  assign n8886 = ( ~n1175 & n7943 ) | ( ~n1175 & n8885 ) | ( n7943 & n8885 ) ;
  assign n8887 = n8886 ^ n7250 ^ n1261 ;
  assign n8888 = ~n8882 & n8887 ;
  assign n8889 = n8888 ^ n6043 ^ 1'b0 ;
  assign n8890 = n312 & ~n8889 ;
  assign n8891 = n8890 ^ n440 ^ 1'b0 ;
  assign n8892 = n8891 ^ n8651 ^ n7675 ;
  assign n8893 = n5651 ^ n4603 ^ n3661 ;
  assign n8894 = n5348 ^ n4404 ^ 1'b0 ;
  assign n8895 = n8893 & n8894 ;
  assign n8896 = ( n372 & n4310 ) | ( n372 & n8895 ) | ( n4310 & n8895 ) ;
  assign n8897 = ( n2717 & n8072 ) | ( n2717 & n8464 ) | ( n8072 & n8464 ) ;
  assign n8898 = n6285 ^ n1655 ^ 1'b0 ;
  assign n8899 = ( n970 & n1893 ) | ( n970 & n2835 ) | ( n1893 & n2835 ) ;
  assign n8900 = n414 & ~n8899 ;
  assign n8901 = ~n3338 & n8900 ;
  assign n8902 = n8901 ^ n2717 ^ n504 ;
  assign n8903 = n3349 ^ n3178 ^ n2005 ;
  assign n8904 = ( n3940 & n7615 ) | ( n3940 & n8903 ) | ( n7615 & n8903 ) ;
  assign n8905 = ( n2370 & n8902 ) | ( n2370 & n8904 ) | ( n8902 & n8904 ) ;
  assign n8906 = n6110 ^ n4139 ^ 1'b0 ;
  assign n8907 = n7328 ^ n4271 ^ n4072 ;
  assign n8908 = ( n4368 & ~n8906 ) | ( n4368 & n8907 ) | ( ~n8906 & n8907 ) ;
  assign n8909 = n3134 ^ n1169 ^ n473 ;
  assign n8910 = n8909 ^ n6489 ^ 1'b0 ;
  assign n8911 = n2833 ^ n2736 ^ n1126 ;
  assign n8912 = ( n2974 & n6270 ) | ( n2974 & n8911 ) | ( n6270 & n8911 ) ;
  assign n8913 = ~n7137 & n8912 ;
  assign n8914 = n7807 ^ n5901 ^ 1'b0 ;
  assign n8918 = ( n752 & n2415 ) | ( n752 & ~n6436 ) | ( n2415 & ~n6436 ) ;
  assign n8917 = n5252 ^ n491 ^ 1'b0 ;
  assign n8915 = ( n4685 & n6164 ) | ( n4685 & n7515 ) | ( n6164 & n7515 ) ;
  assign n8916 = n1574 & ~n8915 ;
  assign n8919 = n8918 ^ n8917 ^ n8916 ;
  assign n8920 = n4707 | n8919 ;
  assign n8921 = n8914 & ~n8920 ;
  assign n8922 = n3802 ^ n3411 ^ n1706 ;
  assign n8923 = n8922 ^ n8456 ^ 1'b0 ;
  assign n8930 = n4851 ^ n2569 ^ n1927 ;
  assign n8926 = n6905 ^ n4320 ^ n902 ;
  assign n8927 = ( ~n3555 & n6202 ) | ( ~n3555 & n8926 ) | ( n6202 & n8926 ) ;
  assign n8924 = n4012 ^ n917 ^ 1'b0 ;
  assign n8925 = ( ~n3857 & n6735 ) | ( ~n3857 & n8924 ) | ( n6735 & n8924 ) ;
  assign n8928 = n8927 ^ n8925 ^ n906 ;
  assign n8929 = n8928 ^ n8307 ^ n6765 ;
  assign n8931 = n8930 ^ n8929 ^ 1'b0 ;
  assign n8933 = n5918 ^ n3376 ^ n2703 ;
  assign n8932 = n6158 ^ n3668 ^ n605 ;
  assign n8934 = n8933 ^ n8932 ^ n5737 ;
  assign n8935 = n7041 & ~n8934 ;
  assign n8936 = ~n7086 & n8935 ;
  assign n8937 = n5335 ^ n3498 ^ 1'b0 ;
  assign n8938 = n3161 | n8937 ;
  assign n8939 = n1844 ^ n823 ^ 1'b0 ;
  assign n8940 = n4294 ^ n3430 ^ n1602 ;
  assign n8941 = ~n8939 & n8940 ;
  assign n8942 = ~n8938 & n8941 ;
  assign n8943 = ~n3971 & n8942 ;
  assign n8944 = ~n3481 & n5353 ;
  assign n8945 = n8944 ^ n8097 ^ 1'b0 ;
  assign n8946 = ~n608 & n8945 ;
  assign n8948 = ( n3933 & n4008 ) | ( n3933 & n5456 ) | ( n4008 & n5456 ) ;
  assign n8949 = n8948 ^ n1797 ^ n1577 ;
  assign n8947 = n2704 & ~n5491 ;
  assign n8950 = n8949 ^ n8947 ^ n7804 ;
  assign n8951 = ( x77 & n442 ) | ( x77 & n1739 ) | ( n442 & n1739 ) ;
  assign n8952 = n5418 & n8951 ;
  assign n8953 = n8950 & n8952 ;
  assign n8954 = n2240 ^ n2066 ^ n1752 ;
  assign n8955 = ( ~n2719 & n3416 ) | ( ~n2719 & n8954 ) | ( n3416 & n8954 ) ;
  assign n8956 = n2929 & ~n8955 ;
  assign n8957 = n6613 ^ n1889 ^ 1'b0 ;
  assign n8958 = n8956 | n8957 ;
  assign n8960 = n7030 ^ n3071 ^ 1'b0 ;
  assign n8961 = n1248 & ~n8960 ;
  assign n8959 = ~n3979 & n8902 ;
  assign n8962 = n8961 ^ n8959 ^ 1'b0 ;
  assign n8963 = n6523 | n8962 ;
  assign n8968 = ( ~n3681 & n5842 ) | ( ~n3681 & n7365 ) | ( n5842 & n7365 ) ;
  assign n8964 = ( n692 & n4976 ) | ( n692 & ~n5262 ) | ( n4976 & ~n5262 ) ;
  assign n8965 = n1404 & n8964 ;
  assign n8966 = n8965 ^ n3809 ^ n1657 ;
  assign n8967 = ( n3962 & n4855 ) | ( n3962 & n8966 ) | ( n4855 & n8966 ) ;
  assign n8969 = n8968 ^ n8967 ^ n6234 ;
  assign n8971 = n4630 ^ n3858 ^ n3030 ;
  assign n8970 = ( n3101 & ~n5832 ) | ( n3101 & n7015 ) | ( ~n5832 & n7015 ) ;
  assign n8972 = n8971 ^ n8970 ^ 1'b0 ;
  assign n8973 = x18 & ~n8972 ;
  assign n8974 = n6662 & ~n8973 ;
  assign n8975 = n1358 & n7252 ;
  assign n8976 = ~n8974 & n8975 ;
  assign n8977 = n617 & n1917 ;
  assign n8978 = n8456 ^ n4444 ^ n1338 ;
  assign n8979 = n8978 ^ n2722 ^ n1256 ;
  assign n8980 = n8977 & n8979 ;
  assign n8981 = ( n5508 & ~n8569 ) | ( n5508 & n8649 ) | ( ~n8569 & n8649 ) ;
  assign n8982 = ( n1068 & n3103 ) | ( n1068 & n8150 ) | ( n3103 & n8150 ) ;
  assign n8983 = x78 & n278 ;
  assign n8984 = n8983 ^ n1016 ^ 1'b0 ;
  assign n8985 = ( n1439 & n8982 ) | ( n1439 & ~n8984 ) | ( n8982 & ~n8984 ) ;
  assign n8986 = n2363 | n6442 ;
  assign n8987 = n8878 & n8986 ;
  assign n8988 = ~n8985 & n8987 ;
  assign n8990 = ~n3379 & n4947 ;
  assign n8989 = n3263 & n5476 ;
  assign n8991 = n8990 ^ n8989 ^ 1'b0 ;
  assign n8992 = n2224 | n8991 ;
  assign n8993 = ~n6804 & n8992 ;
  assign n8997 = x139 & n2148 ;
  assign n8998 = n8997 ^ n1636 ^ 1'b0 ;
  assign n8994 = ( ~n1838 & n4791 ) | ( ~n1838 & n6666 ) | ( n4791 & n6666 ) ;
  assign n8995 = n6842 ^ x205 ^ 1'b0 ;
  assign n8996 = n8994 & n8995 ;
  assign n8999 = n8998 ^ n8996 ^ n313 ;
  assign n9000 = ( n1304 & n4649 ) | ( n1304 & ~n6167 ) | ( n4649 & ~n6167 ) ;
  assign n9001 = ( n3287 & n3809 ) | ( n3287 & n9000 ) | ( n3809 & n9000 ) ;
  assign n9002 = n3646 ^ n2415 ^ n1060 ;
  assign n9003 = n8255 ^ n1099 ^ 1'b0 ;
  assign n9004 = n6323 ^ n2635 ^ 1'b0 ;
  assign n9005 = ( n4208 & ~n9003 ) | ( n4208 & n9004 ) | ( ~n9003 & n9004 ) ;
  assign n9006 = ~n400 & n3814 ;
  assign n9007 = n9006 ^ n5038 ^ 1'b0 ;
  assign n9008 = ~n4873 & n9007 ;
  assign n9009 = ( n1822 & n2286 ) | ( n1822 & n4993 ) | ( n2286 & n4993 ) ;
  assign n9010 = n9009 ^ n1980 ^ 1'b0 ;
  assign n9011 = ~n8390 & n9010 ;
  assign n9012 = ( n3963 & n5553 ) | ( n3963 & ~n9011 ) | ( n5553 & ~n9011 ) ;
  assign n9013 = n892 | n9012 ;
  assign n9014 = n9013 ^ n8677 ^ 1'b0 ;
  assign n9016 = n2294 & n7135 ;
  assign n9015 = n4057 | n8338 ;
  assign n9017 = n9016 ^ n9015 ^ 1'b0 ;
  assign n9018 = ( n5235 & ~n6531 ) | ( n5235 & n9017 ) | ( ~n6531 & n9017 ) ;
  assign n9019 = n8030 ^ n1493 ^ 1'b0 ;
  assign n9020 = n1429 & ~n9019 ;
  assign n9021 = n5189 ^ n1134 ^ 1'b0 ;
  assign n9022 = n3910 & ~n9021 ;
  assign n9023 = n9022 ^ x112 ^ 1'b0 ;
  assign n9024 = n869 | n9023 ;
  assign n9025 = n9024 ^ n1795 ^ 1'b0 ;
  assign n9027 = n6719 ^ n6294 ^ 1'b0 ;
  assign n9026 = n5363 | n6927 ;
  assign n9028 = n9027 ^ n9026 ^ 1'b0 ;
  assign n9029 = n9028 ^ n6693 ^ n1994 ;
  assign n9030 = n3014 ^ n2981 ^ n318 ;
  assign n9031 = n9030 ^ n3973 ^ 1'b0 ;
  assign n9032 = n4787 | n9031 ;
  assign n9033 = ( n1304 & n5526 ) | ( n1304 & ~n8781 ) | ( n5526 & ~n8781 ) ;
  assign n9034 = n2017 ^ x131 ^ 1'b0 ;
  assign n9035 = n6028 ^ n5394 ^ n1464 ;
  assign n9036 = n364 & n8328 ;
  assign n9037 = n2967 & n9036 ;
  assign n9039 = x33 & ~n1327 ;
  assign n9040 = n9039 ^ n5764 ^ n1410 ;
  assign n9038 = n5437 & ~n8745 ;
  assign n9041 = n9040 ^ n9038 ^ 1'b0 ;
  assign n9042 = ( ~x56 & n271 ) | ( ~x56 & n6453 ) | ( n271 & n6453 ) ;
  assign n9043 = n4885 & ~n7509 ;
  assign n9044 = n9043 ^ n7363 ^ 1'b0 ;
  assign n9045 = ( n3609 & n9042 ) | ( n3609 & ~n9044 ) | ( n9042 & ~n9044 ) ;
  assign n9046 = ( ~x19 & n1365 ) | ( ~x19 & n8247 ) | ( n1365 & n8247 ) ;
  assign n9047 = n4158 ^ n2974 ^ n982 ;
  assign n9048 = n7085 ^ n2905 ^ n1336 ;
  assign n9049 = ( n4599 & n9047 ) | ( n4599 & n9048 ) | ( n9047 & n9048 ) ;
  assign n9050 = n7192 ^ n3668 ^ n1639 ;
  assign n9051 = n9050 ^ n6572 ^ 1'b0 ;
  assign n9052 = n3899 & ~n9051 ;
  assign n9053 = n3910 & n7262 ;
  assign n9054 = n9053 ^ n2271 ^ 1'b0 ;
  assign n9055 = ~n4547 & n9054 ;
  assign n9056 = n9055 ^ n358 ^ 1'b0 ;
  assign n9057 = n9056 ^ n3366 ^ n3015 ;
  assign n9058 = n5155 ^ n5153 ^ 1'b0 ;
  assign n9066 = n2751 ^ n1832 ^ 1'b0 ;
  assign n9067 = ( n819 & ~n8075 ) | ( n819 & n9066 ) | ( ~n8075 & n9066 ) ;
  assign n9064 = n447 & n2836 ;
  assign n9065 = ~n3879 & n9064 ;
  assign n9061 = n6058 & n8542 ;
  assign n9062 = n9061 ^ n1323 ^ n598 ;
  assign n9059 = n328 & ~n2823 ;
  assign n9060 = ~n7245 & n9059 ;
  assign n9063 = n9062 ^ n9060 ^ n6667 ;
  assign n9068 = n9067 ^ n9065 ^ n9063 ;
  assign n9069 = n4846 ^ n4334 ^ n2412 ;
  assign n9070 = ~n5289 & n9069 ;
  assign n9071 = n9070 ^ n1380 ^ 1'b0 ;
  assign n9072 = n9071 ^ n2175 ^ n627 ;
  assign n9073 = ( n3018 & n5403 ) | ( n3018 & ~n9072 ) | ( n5403 & ~n9072 ) ;
  assign n9074 = ( n3120 & n7039 ) | ( n3120 & n9073 ) | ( n7039 & n9073 ) ;
  assign n9075 = ~x49 & n4379 ;
  assign n9077 = ~n4487 & n6043 ;
  assign n9076 = n2015 ^ n1285 ^ 1'b0 ;
  assign n9078 = n9077 ^ n9076 ^ n7416 ;
  assign n9079 = n9078 ^ n2168 ^ 1'b0 ;
  assign n9080 = ( n2720 & n4261 ) | ( n2720 & ~n7839 ) | ( n4261 & ~n7839 ) ;
  assign n9081 = ( n6672 & n9079 ) | ( n6672 & ~n9080 ) | ( n9079 & ~n9080 ) ;
  assign n9082 = n9081 ^ n8419 ^ n6396 ;
  assign n9083 = n3078 & ~n6831 ;
  assign n9084 = ~n1763 & n9083 ;
  assign n9085 = ( ~n4480 & n5260 ) | ( ~n4480 & n8814 ) | ( n5260 & n8814 ) ;
  assign n9086 = ( ~n3414 & n3641 ) | ( ~n3414 & n7367 ) | ( n3641 & n7367 ) ;
  assign n9087 = ( n6657 & ~n9085 ) | ( n6657 & n9086 ) | ( ~n9085 & n9086 ) ;
  assign n9088 = n8979 ^ n4373 ^ 1'b0 ;
  assign n9089 = n9088 ^ n5858 ^ x175 ;
  assign n9090 = n3207 ^ n3084 ^ 1'b0 ;
  assign n9091 = ~n887 & n8557 ;
  assign n9092 = n8061 & n9091 ;
  assign n9093 = n3165 | n9092 ;
  assign n9094 = ~n1204 & n9093 ;
  assign n9095 = n667 | n5014 ;
  assign n9096 = n5387 & ~n9095 ;
  assign n9097 = n9096 ^ n4301 ^ 1'b0 ;
  assign n9098 = ( x41 & ~n6293 ) | ( x41 & n7512 ) | ( ~n6293 & n7512 ) ;
  assign n9099 = ~n1679 & n7077 ;
  assign n9100 = ( n1544 & n2745 ) | ( n1544 & n6179 ) | ( n2745 & n6179 ) ;
  assign n9101 = ( n7416 & ~n9099 ) | ( n7416 & n9100 ) | ( ~n9099 & n9100 ) ;
  assign n9103 = ~n1423 & n3922 ;
  assign n9102 = ( n895 & n1693 ) | ( n895 & n5458 ) | ( n1693 & n5458 ) ;
  assign n9104 = n9103 ^ n9102 ^ n2435 ;
  assign n9105 = ( n831 & n1279 ) | ( n831 & n1371 ) | ( n1279 & n1371 ) ;
  assign n9106 = n789 ^ n764 ^ 1'b0 ;
  assign n9107 = n4551 & n9106 ;
  assign n9108 = ~n2457 & n4325 ;
  assign n9109 = ~n690 & n9108 ;
  assign n9110 = n9107 | n9109 ;
  assign n9111 = n7292 | n9110 ;
  assign n9122 = ( ~n1316 & n4902 ) | ( ~n1316 & n4940 ) | ( n4902 & n4940 ) ;
  assign n9112 = n5786 ^ n3668 ^ n1248 ;
  assign n9113 = ( n2539 & n5679 ) | ( n2539 & n9112 ) | ( n5679 & n9112 ) ;
  assign n9114 = n2681 | n5492 ;
  assign n9115 = ( ~x1 & n2318 ) | ( ~x1 & n4383 ) | ( n2318 & n4383 ) ;
  assign n9116 = n5448 & ~n9115 ;
  assign n9117 = n9116 ^ n8277 ^ 1'b0 ;
  assign n9118 = ( n3472 & n5164 ) | ( n3472 & n9117 ) | ( n5164 & n9117 ) ;
  assign n9119 = n9114 | n9118 ;
  assign n9120 = n3551 & ~n9119 ;
  assign n9121 = n9113 | n9120 ;
  assign n9123 = n9122 ^ n9121 ^ 1'b0 ;
  assign n9124 = n9111 & ~n9123 ;
  assign n9125 = ( n9104 & n9105 ) | ( n9104 & n9124 ) | ( n9105 & n9124 ) ;
  assign n9126 = n1938 ^ n313 ^ 1'b0 ;
  assign n9127 = n3103 | n9126 ;
  assign n9128 = n9127 ^ n7720 ^ n2590 ;
  assign n9129 = ~n3267 & n5749 ;
  assign n9130 = ~n7231 & n9129 ;
  assign n9131 = ( ~x43 & n9128 ) | ( ~x43 & n9130 ) | ( n9128 & n9130 ) ;
  assign n9132 = n9131 ^ n7026 ^ n463 ;
  assign n9133 = ~n1119 & n2550 ;
  assign n9134 = n9133 ^ n8901 ^ 1'b0 ;
  assign n9135 = ~n2590 & n9134 ;
  assign n9136 = ( n6585 & n7756 ) | ( n6585 & ~n9135 ) | ( n7756 & ~n9135 ) ;
  assign n9137 = n5011 | n7675 ;
  assign n9138 = ( n1805 & n5359 ) | ( n1805 & n8335 ) | ( n5359 & n8335 ) ;
  assign n9139 = n1688 & ~n9138 ;
  assign n9142 = n955 ^ n898 ^ 1'b0 ;
  assign n9141 = n9040 ^ n1320 ^ n455 ;
  assign n9140 = n7247 ^ n6429 ^ n532 ;
  assign n9143 = n9142 ^ n9141 ^ n9140 ;
  assign n9144 = n4951 ^ n2998 ^ n997 ;
  assign n9145 = n3319 ^ n2218 ^ n516 ;
  assign n9146 = n9145 ^ n3287 ^ 1'b0 ;
  assign n9147 = n8456 & n8977 ;
  assign n9148 = n364 & n9147 ;
  assign n9149 = ( n9144 & n9146 ) | ( n9144 & n9148 ) | ( n9146 & n9148 ) ;
  assign n9150 = n5312 ^ n3230 ^ n2352 ;
  assign n9151 = ( n2271 & n3685 ) | ( n2271 & n9150 ) | ( n3685 & n9150 ) ;
  assign n9152 = n4322 ^ n3441 ^ 1'b0 ;
  assign n9153 = ( n2508 & n9151 ) | ( n2508 & ~n9152 ) | ( n9151 & ~n9152 ) ;
  assign n9154 = ~n8041 & n8649 ;
  assign n9155 = n2342 | n9154 ;
  assign n9156 = n3959 | n9155 ;
  assign n9157 = ( ~n4721 & n5701 ) | ( ~n4721 & n6501 ) | ( n5701 & n6501 ) ;
  assign n9158 = n5172 & n5942 ;
  assign n9159 = n9158 ^ n4560 ^ 1'b0 ;
  assign n9160 = ( n1040 & n2955 ) | ( n1040 & ~n6328 ) | ( n2955 & ~n6328 ) ;
  assign n9161 = ( n8881 & n9159 ) | ( n8881 & ~n9160 ) | ( n9159 & ~n9160 ) ;
  assign n9162 = ( n5155 & n6074 ) | ( n5155 & n7603 ) | ( n6074 & n7603 ) ;
  assign n9163 = x83 | n9162 ;
  assign n9164 = n2857 ^ n1459 ^ 1'b0 ;
  assign n9165 = n9164 ^ n3931 ^ n2656 ;
  assign n9166 = n9165 ^ n374 ^ 1'b0 ;
  assign n9169 = n4605 ^ n3852 ^ n1711 ;
  assign n9167 = ( n1586 & ~n2057 ) | ( n1586 & n2555 ) | ( ~n2057 & n2555 ) ;
  assign n9168 = n9167 ^ n8252 ^ n1466 ;
  assign n9170 = n9169 ^ n9168 ^ n6287 ;
  assign n9171 = n1713 & n9170 ;
  assign n9172 = n9171 ^ n6138 ^ 1'b0 ;
  assign n9173 = n9166 & ~n9172 ;
  assign n9174 = n4152 ^ n818 ^ 1'b0 ;
  assign n9175 = n9174 ^ n7202 ^ n3874 ;
  assign n9176 = n5695 ^ n4437 ^ 1'b0 ;
  assign n9177 = n3365 | n4197 ;
  assign n9178 = n9177 ^ n8628 ^ n4372 ;
  assign n9179 = ( ~n956 & n3526 ) | ( ~n956 & n5621 ) | ( n3526 & n5621 ) ;
  assign n9180 = ( ~n1567 & n4597 ) | ( ~n1567 & n9179 ) | ( n4597 & n9179 ) ;
  assign n9181 = ~n1599 & n9180 ;
  assign n9182 = n3412 & n9181 ;
  assign n9183 = ~n1623 & n9182 ;
  assign n9186 = ( n545 & n1129 ) | ( n545 & n7367 ) | ( n1129 & n7367 ) ;
  assign n9184 = x82 & n5236 ;
  assign n9185 = ~n509 & n9184 ;
  assign n9187 = n9186 ^ n9185 ^ n2011 ;
  assign n9188 = n9187 ^ n7204 ^ n3949 ;
  assign n9189 = n9188 ^ n6362 ^ 1'b0 ;
  assign n9190 = n1472 ^ n1042 ^ 1'b0 ;
  assign n9191 = n1849 & n9190 ;
  assign n9192 = n9191 ^ n1029 ^ 1'b0 ;
  assign n9193 = ~n7774 & n9192 ;
  assign n9194 = n5764 | n9193 ;
  assign n9195 = n2462 & ~n4291 ;
  assign n9196 = ~n6500 & n9195 ;
  assign n9197 = n9196 ^ n1523 ^ 1'b0 ;
  assign n9198 = ( x8 & ~n1382 ) | ( x8 & n2166 ) | ( ~n1382 & n2166 ) ;
  assign n9204 = n4449 ^ n1439 ^ 1'b0 ;
  assign n9205 = n8310 & n9204 ;
  assign n9199 = n6946 ^ n1087 ^ 1'b0 ;
  assign n9200 = n6901 ^ n1278 ^ x23 ;
  assign n9201 = n9200 ^ n8767 ^ 1'b0 ;
  assign n9202 = n9199 & ~n9201 ;
  assign n9203 = ~n283 & n9202 ;
  assign n9206 = n9205 ^ n9203 ^ 1'b0 ;
  assign n9207 = n9198 | n9206 ;
  assign n9208 = n9207 ^ n3510 ^ 1'b0 ;
  assign n9209 = n5204 ^ n1717 ^ n766 ;
  assign n9210 = ( n9197 & n9208 ) | ( n9197 & n9209 ) | ( n9208 & n9209 ) ;
  assign n9216 = n6362 ^ n4601 ^ n2524 ;
  assign n9217 = ( ~n6890 & n6928 ) | ( ~n6890 & n9216 ) | ( n6928 & n9216 ) ;
  assign n9211 = n4502 ^ n2832 ^ x30 ;
  assign n9212 = n9211 ^ n9066 ^ n4396 ;
  assign n9213 = n9212 ^ n3849 ^ 1'b0 ;
  assign n9214 = n8377 & n9213 ;
  assign n9215 = n6705 & n9214 ;
  assign n9218 = n9217 ^ n9215 ^ 1'b0 ;
  assign n9219 = ( x92 & ~x93 ) | ( x92 & n4101 ) | ( ~x93 & n4101 ) ;
  assign n9220 = ( n4514 & n6005 ) | ( n4514 & ~n9219 ) | ( n6005 & ~n9219 ) ;
  assign n9221 = n5959 | n8961 ;
  assign n9222 = n1679 ^ n1025 ^ 1'b0 ;
  assign n9223 = n2213 ^ n1205 ^ x226 ;
  assign n9224 = n9223 ^ n6810 ^ n4225 ;
  assign n9225 = n9222 & ~n9224 ;
  assign n9232 = n6062 & n8205 ;
  assign n9226 = ( n382 & n677 ) | ( n382 & ~n7608 ) | ( n677 & ~n7608 ) ;
  assign n9227 = n2867 ^ n772 ^ n359 ;
  assign n9228 = n9227 ^ n1740 ^ n614 ;
  assign n9229 = n1219 & ~n2255 ;
  assign n9230 = ~n9228 & n9229 ;
  assign n9231 = n9226 | n9230 ;
  assign n9233 = n9232 ^ n9231 ^ 1'b0 ;
  assign n9234 = n9225 | n9233 ;
  assign n9235 = n9221 | n9234 ;
  assign n9236 = ~n2564 & n5444 ;
  assign n9237 = n1355 & n9236 ;
  assign n9238 = n3508 ^ n3308 ^ n3031 ;
  assign n9239 = ( n3745 & n9237 ) | ( n3745 & n9238 ) | ( n9237 & n9238 ) ;
  assign n9240 = n9239 ^ n5879 ^ n1694 ;
  assign n9241 = ( ~n3909 & n4921 ) | ( ~n3909 & n5494 ) | ( n4921 & n5494 ) ;
  assign n9242 = n2017 & n6284 ;
  assign n9243 = ~n856 & n9242 ;
  assign n9244 = n2125 & ~n8311 ;
  assign n9245 = ( ~n9241 & n9243 ) | ( ~n9241 & n9244 ) | ( n9243 & n9244 ) ;
  assign n9246 = ( ~n4221 & n5887 ) | ( ~n4221 & n6321 ) | ( n5887 & n6321 ) ;
  assign n9247 = ( n3309 & n9245 ) | ( n3309 & ~n9246 ) | ( n9245 & ~n9246 ) ;
  assign n9251 = n6033 ^ n4289 ^ n3131 ;
  assign n9248 = ( n642 & ~n845 ) | ( n642 & n1823 ) | ( ~n845 & n1823 ) ;
  assign n9249 = n9248 ^ n733 ^ 1'b0 ;
  assign n9250 = n5428 & ~n9249 ;
  assign n9252 = n9251 ^ n9250 ^ n1695 ;
  assign n9253 = n9177 ^ n5376 ^ n3038 ;
  assign n9254 = n9253 ^ n332 ^ x163 ;
  assign n9255 = n9254 ^ n5196 ^ n4019 ;
  assign n9256 = ( n2125 & n9252 ) | ( n2125 & ~n9255 ) | ( n9252 & ~n9255 ) ;
  assign n9257 = n9247 & n9256 ;
  assign n9261 = ( n1746 & n3645 ) | ( n1746 & ~n5811 ) | ( n3645 & ~n5811 ) ;
  assign n9258 = n3633 ^ n2385 ^ n1587 ;
  assign n9259 = ~x67 & n387 ;
  assign n9260 = ~n9258 & n9259 ;
  assign n9262 = n9261 ^ n9260 ^ n474 ;
  assign n9263 = n304 | n364 ;
  assign n9264 = n9263 ^ n1002 ^ 1'b0 ;
  assign n9265 = n9264 ^ n6289 ^ n3943 ;
  assign n9266 = n5579 & n7101 ;
  assign n9267 = ~n9265 & n9266 ;
  assign n9268 = ( n5871 & n6906 ) | ( n5871 & n9267 ) | ( n6906 & n9267 ) ;
  assign n9273 = n2085 ^ n1632 ^ 1'b0 ;
  assign n9274 = n9273 ^ n1712 ^ 1'b0 ;
  assign n9270 = ( x6 & n3519 ) | ( x6 & n6453 ) | ( n3519 & n6453 ) ;
  assign n9269 = ( ~n3146 & n5425 ) | ( ~n3146 & n6764 ) | ( n5425 & n6764 ) ;
  assign n9271 = n9270 ^ n9269 ^ n1992 ;
  assign n9272 = ~n4669 & n9271 ;
  assign n9275 = n9274 ^ n9272 ^ n9003 ;
  assign n9280 = n5131 | n7647 ;
  assign n9281 = n1367 | n9280 ;
  assign n9279 = n7844 ^ n3598 ^ n1102 ;
  assign n9276 = n6552 ^ n2494 ^ n1188 ;
  assign n9277 = n9276 ^ n8308 ^ n361 ;
  assign n9278 = n9277 ^ n8762 ^ n5882 ;
  assign n9282 = n9281 ^ n9279 ^ n9278 ;
  assign n9283 = n382 ^ n302 ^ 1'b0 ;
  assign n9284 = ~n3282 & n4634 ;
  assign n9285 = ~n9283 & n9284 ;
  assign n9286 = n7681 ^ n977 ^ 1'b0 ;
  assign n9287 = n508 & ~n9286 ;
  assign n9288 = n9287 ^ n6921 ^ n2244 ;
  assign n9289 = ( n4945 & n9285 ) | ( n4945 & n9288 ) | ( n9285 & n9288 ) ;
  assign n9290 = n4355 ^ n3906 ^ 1'b0 ;
  assign n9291 = n3061 | n9290 ;
  assign n9294 = ( ~n430 & n713 ) | ( ~n430 & n1609 ) | ( n713 & n1609 ) ;
  assign n9295 = n9294 ^ n4960 ^ n3888 ;
  assign n9292 = ( ~n470 & n1638 ) | ( ~n470 & n2325 ) | ( n1638 & n2325 ) ;
  assign n9293 = n9292 ^ n9130 ^ n434 ;
  assign n9296 = n9295 ^ n9293 ^ n2009 ;
  assign n9297 = ( ~n2413 & n3102 ) | ( ~n2413 & n3249 ) | ( n3102 & n3249 ) ;
  assign n9298 = n3268 & ~n9297 ;
  assign n9299 = n1223 ^ n1066 ^ 1'b0 ;
  assign n9300 = n9299 ^ n1040 ^ n664 ;
  assign n9301 = n1116 ^ n572 ^ 1'b0 ;
  assign n9302 = n9301 ^ n5820 ^ n2044 ;
  assign n9303 = ( ~n777 & n864 ) | ( ~n777 & n6864 ) | ( n864 & n6864 ) ;
  assign n9304 = n9303 ^ n9123 ^ n5698 ;
  assign n9305 = n3280 ^ n299 ^ 1'b0 ;
  assign n9306 = ( n606 & ~n3304 ) | ( n606 & n4448 ) | ( ~n3304 & n4448 ) ;
  assign n9307 = n9306 ^ n1959 ^ 1'b0 ;
  assign n9308 = n9305 & ~n9307 ;
  assign n9309 = ( n3841 & n7505 ) | ( n3841 & ~n9308 ) | ( n7505 & ~n9308 ) ;
  assign n9310 = ( x25 & n3548 ) | ( x25 & ~n4260 ) | ( n3548 & ~n4260 ) ;
  assign n9311 = n3898 | n6552 ;
  assign n9312 = ( n4493 & n5617 ) | ( n4493 & ~n9311 ) | ( n5617 & ~n9311 ) ;
  assign n9313 = ( ~n2428 & n9310 ) | ( ~n2428 & n9312 ) | ( n9310 & n9312 ) ;
  assign n9314 = n3226 ^ n1637 ^ n1297 ;
  assign n9315 = n9314 ^ n5641 ^ n1577 ;
  assign n9316 = n2185 ^ n1724 ^ x108 ;
  assign n9317 = ( x163 & n4152 ) | ( x163 & n4841 ) | ( n4152 & n4841 ) ;
  assign n9318 = n9317 ^ x191 ^ x32 ;
  assign n9319 = ~n7366 & n9318 ;
  assign n9320 = ~n9316 & n9319 ;
  assign n9321 = ~n9315 & n9320 ;
  assign n9322 = n4186 | n9321 ;
  assign n9323 = n9313 | n9322 ;
  assign n9324 = ( x159 & n7100 ) | ( x159 & ~n7460 ) | ( n7100 & ~n7460 ) ;
  assign n9325 = n3332 & ~n7053 ;
  assign n9326 = n7730 & n9325 ;
  assign n9327 = n5267 ^ n4501 ^ 1'b0 ;
  assign n9328 = n9327 ^ n5689 ^ n3879 ;
  assign n9329 = n5864 ^ n3191 ^ 1'b0 ;
  assign n9330 = n7903 & ~n9329 ;
  assign n9331 = ( n3022 & n5652 ) | ( n3022 & n9330 ) | ( n5652 & n9330 ) ;
  assign n9332 = n9331 ^ n7575 ^ n4509 ;
  assign n9333 = ( n3117 & ~n3777 ) | ( n3117 & n4273 ) | ( ~n3777 & n4273 ) ;
  assign n9334 = ( n1151 & ~n2026 ) | ( n1151 & n5613 ) | ( ~n2026 & n5613 ) ;
  assign n9335 = n9334 ^ n7283 ^ n2094 ;
  assign n9336 = n9335 ^ n3445 ^ n268 ;
  assign n9337 = ( n4909 & n9333 ) | ( n4909 & ~n9336 ) | ( n9333 & ~n9336 ) ;
  assign n9338 = n9337 ^ x216 ^ 1'b0 ;
  assign n9339 = n6668 ^ n3223 ^ n3010 ;
  assign n9340 = n9339 ^ n5335 ^ 1'b0 ;
  assign n9341 = ( n497 & n5913 ) | ( n497 & n9340 ) | ( n5913 & n9340 ) ;
  assign n9342 = ( ~n870 & n7585 ) | ( ~n870 & n9341 ) | ( n7585 & n9341 ) ;
  assign n9347 = n8784 ^ n7233 ^ n5214 ;
  assign n9344 = n3165 ^ n2166 ^ n1775 ;
  assign n9343 = ( n841 & ~n1838 ) | ( n841 & n4694 ) | ( ~n1838 & n4694 ) ;
  assign n9345 = n9344 ^ n9343 ^ 1'b0 ;
  assign n9346 = ( x227 & ~n8835 ) | ( x227 & n9345 ) | ( ~n8835 & n9345 ) ;
  assign n9348 = n9347 ^ n9346 ^ n3747 ;
  assign n9349 = x227 | n6608 ;
  assign n9350 = n9349 ^ n3347 ^ n693 ;
  assign n9351 = ( n2438 & ~n6450 ) | ( n2438 & n9350 ) | ( ~n6450 & n9350 ) ;
  assign n9352 = n4541 ^ n3933 ^ 1'b0 ;
  assign n9353 = ( ~n5903 & n9351 ) | ( ~n5903 & n9352 ) | ( n9351 & n9352 ) ;
  assign n9354 = n9353 ^ n2875 ^ 1'b0 ;
  assign n9355 = n717 & ~n9354 ;
  assign n9356 = ~n5719 & n9355 ;
  assign n9357 = ( ~n789 & n2427 ) | ( ~n789 & n7478 ) | ( n2427 & n7478 ) ;
  assign n9358 = n4842 ^ n2385 ^ n2382 ;
  assign n9359 = ( ~n8304 & n9357 ) | ( ~n8304 & n9358 ) | ( n9357 & n9358 ) ;
  assign n9360 = ( n6051 & ~n9294 ) | ( n6051 & n9359 ) | ( ~n9294 & n9359 ) ;
  assign n9361 = ( n593 & n2905 ) | ( n593 & ~n3881 ) | ( n2905 & ~n3881 ) ;
  assign n9362 = n9361 ^ n6682 ^ 1'b0 ;
  assign n9363 = n4787 & n9362 ;
  assign n9364 = ( ~n692 & n1122 ) | ( ~n692 & n1250 ) | ( n1122 & n1250 ) ;
  assign n9365 = n9364 ^ n5874 ^ 1'b0 ;
  assign n9366 = n7017 & n9365 ;
  assign n9367 = ~n5013 & n9366 ;
  assign n9368 = n9367 ^ n8714 ^ 1'b0 ;
  assign n9369 = ( n2258 & ~n5511 ) | ( n2258 & n6030 ) | ( ~n5511 & n6030 ) ;
  assign n9370 = n9369 ^ n8182 ^ n3598 ;
  assign n9372 = ( n4281 & n6768 ) | ( n4281 & n8205 ) | ( n6768 & n8205 ) ;
  assign n9371 = ( n534 & ~n1791 ) | ( n534 & n4484 ) | ( ~n1791 & n4484 ) ;
  assign n9373 = n9372 ^ n9371 ^ n5468 ;
  assign n9374 = ( n1110 & n2146 ) | ( n1110 & ~n3541 ) | ( n2146 & ~n3541 ) ;
  assign n9375 = n664 ^ n505 ^ 1'b0 ;
  assign n9376 = n1992 & ~n9375 ;
  assign n9377 = n9376 ^ n9064 ^ 1'b0 ;
  assign n9378 = ~n1404 & n9377 ;
  assign n9379 = ( n1198 & ~n1761 ) | ( n1198 & n5640 ) | ( ~n1761 & n5640 ) ;
  assign n9380 = n9379 ^ n3520 ^ n1646 ;
  assign n9381 = n4734 & ~n9380 ;
  assign n9382 = n9381 ^ n2969 ^ 1'b0 ;
  assign n9383 = n9382 ^ n1232 ^ n952 ;
  assign n9384 = n2491 ^ n2038 ^ 1'b0 ;
  assign n9385 = n7540 & n9384 ;
  assign n9393 = ( n1298 & n3840 ) | ( n1298 & n8688 ) | ( n3840 & n8688 ) ;
  assign n9394 = ( n7596 & n7724 ) | ( n7596 & n9393 ) | ( n7724 & n9393 ) ;
  assign n9391 = n1389 | n3192 ;
  assign n9392 = ~n7825 & n9391 ;
  assign n9395 = n9394 ^ n9392 ^ n7865 ;
  assign n9386 = n2432 & n8431 ;
  assign n9387 = n1694 & n9386 ;
  assign n9388 = n1292 | n8371 ;
  assign n9389 = n9388 ^ n3331 ^ 1'b0 ;
  assign n9390 = ( n1527 & ~n9387 ) | ( n1527 & n9389 ) | ( ~n9387 & n9389 ) ;
  assign n9396 = n9395 ^ n9390 ^ n7574 ;
  assign n9397 = n9396 ^ n5000 ^ 1'b0 ;
  assign n9398 = n9385 & ~n9397 ;
  assign n9399 = ( ~x130 & n9383 ) | ( ~x130 & n9398 ) | ( n9383 & n9398 ) ;
  assign n9411 = n2846 & n3164 ;
  assign n9400 = n3239 & ~n4888 ;
  assign n9401 = n6465 ^ n2741 ^ 1'b0 ;
  assign n9402 = n3643 | n9401 ;
  assign n9403 = n9402 ^ n829 ^ 1'b0 ;
  assign n9404 = n2560 ^ n1858 ^ 1'b0 ;
  assign n9405 = n9403 & n9404 ;
  assign n9407 = n7901 ^ n1685 ^ 1'b0 ;
  assign n9408 = n2528 | n9407 ;
  assign n9406 = ( n366 & n854 ) | ( n366 & n5307 ) | ( n854 & n5307 ) ;
  assign n9409 = n9408 ^ n9406 ^ 1'b0 ;
  assign n9410 = ( n9400 & n9405 ) | ( n9400 & ~n9409 ) | ( n9405 & ~n9409 ) ;
  assign n9412 = n9411 ^ n9410 ^ n340 ;
  assign n9413 = ( n5304 & n8575 ) | ( n5304 & n9306 ) | ( n8575 & n9306 ) ;
  assign n9414 = n9413 ^ n5976 ^ 1'b0 ;
  assign n9415 = n6281 & ~n9414 ;
  assign n9430 = n3094 & n4123 ;
  assign n9431 = n9430 ^ n6723 ^ 1'b0 ;
  assign n9432 = ( n775 & n6272 ) | ( n775 & ~n9431 ) | ( n6272 & ~n9431 ) ;
  assign n9433 = ( x87 & ~n4350 ) | ( x87 & n9432 ) | ( ~n4350 & n9432 ) ;
  assign n9417 = n5142 ^ n1559 ^ 1'b0 ;
  assign n9418 = ~n4822 & n9417 ;
  assign n9419 = n1153 & n9418 ;
  assign n9420 = n9419 ^ n5732 ^ 1'b0 ;
  assign n9421 = n9420 ^ n4359 ^ n2390 ;
  assign n9416 = n7070 ^ n5725 ^ n1467 ;
  assign n9422 = n9421 ^ n9416 ^ 1'b0 ;
  assign n9423 = ( ~n266 & n1394 ) | ( ~n266 & n4408 ) | ( n1394 & n4408 ) ;
  assign n9424 = ( n5521 & ~n8071 ) | ( n5521 & n9423 ) | ( ~n8071 & n9423 ) ;
  assign n9425 = n1235 ^ n468 ^ 1'b0 ;
  assign n9426 = n1892 & ~n9425 ;
  assign n9427 = n9424 & ~n9426 ;
  assign n9428 = n2564 & n9427 ;
  assign n9429 = ( n5205 & n9422 ) | ( n5205 & ~n9428 ) | ( n9422 & ~n9428 ) ;
  assign n9434 = n9433 ^ n9429 ^ 1'b0 ;
  assign n9435 = n347 & n9434 ;
  assign n9436 = n4733 ^ x58 ^ 1'b0 ;
  assign n9437 = n5143 | n5343 ;
  assign n9438 = x103 & n5090 ;
  assign n9439 = ( n3414 & n6486 ) | ( n3414 & ~n9438 ) | ( n6486 & ~n9438 ) ;
  assign n9440 = n293 | n1610 ;
  assign n9441 = n9439 | n9440 ;
  assign n9442 = n9441 ^ n7253 ^ n6943 ;
  assign n9443 = n1793 ^ n1758 ^ x12 ;
  assign n9444 = n9443 ^ n8193 ^ n3185 ;
  assign n9445 = n9444 ^ n7467 ^ n6527 ;
  assign n9447 = ( n1548 & n1746 ) | ( n1548 & n1927 ) | ( n1746 & n1927 ) ;
  assign n9448 = n2453 | n9447 ;
  assign n9449 = n9448 ^ n6803 ^ 1'b0 ;
  assign n9450 = ( ~n1131 & n5827 ) | ( ~n1131 & n9449 ) | ( n5827 & n9449 ) ;
  assign n9446 = n7440 ^ n6557 ^ 1'b0 ;
  assign n9451 = n9450 ^ n9446 ^ n4578 ;
  assign n9452 = n1070 ^ x182 ^ 1'b0 ;
  assign n9453 = ~n729 & n1340 ;
  assign n9454 = n9453 ^ x248 ^ 1'b0 ;
  assign n9455 = ( n431 & n9452 ) | ( n431 & ~n9454 ) | ( n9452 & ~n9454 ) ;
  assign n9456 = ( n3292 & ~n5039 ) | ( n3292 & n9455 ) | ( ~n5039 & n9455 ) ;
  assign n9457 = n9451 & ~n9456 ;
  assign n9458 = ~n7505 & n9457 ;
  assign n9459 = n1151 & n1368 ;
  assign n9460 = n9459 ^ n892 ^ 1'b0 ;
  assign n9461 = ~n1354 & n9460 ;
  assign n9462 = n9461 ^ n2022 ^ 1'b0 ;
  assign n9463 = n9462 ^ n5404 ^ n4563 ;
  assign n9464 = n2341 & ~n9463 ;
  assign n9466 = n5915 ^ n748 ^ 1'b0 ;
  assign n9465 = n7774 ^ n1856 ^ 1'b0 ;
  assign n9467 = n9466 ^ n9465 ^ 1'b0 ;
  assign n9468 = n9467 ^ n1738 ^ 1'b0 ;
  assign n9469 = n9468 ^ n6537 ^ n2598 ;
  assign n9470 = x69 & ~n5092 ;
  assign n9471 = n9470 ^ x227 ^ 1'b0 ;
  assign n9472 = ( ~n1977 & n3369 ) | ( ~n1977 & n6810 ) | ( n3369 & n6810 ) ;
  assign n9473 = n6132 ^ n2494 ^ n1508 ;
  assign n9474 = ( n4336 & n6799 ) | ( n4336 & ~n9473 ) | ( n6799 & ~n9473 ) ;
  assign n9475 = ( ~n2158 & n9472 ) | ( ~n2158 & n9474 ) | ( n9472 & n9474 ) ;
  assign n9477 = ( n458 & n2079 ) | ( n458 & n2515 ) | ( n2079 & n2515 ) ;
  assign n9476 = n4042 & ~n8861 ;
  assign n9478 = n9477 ^ n9476 ^ n3765 ;
  assign n9479 = ( ~n2957 & n4040 ) | ( ~n2957 & n4486 ) | ( n4040 & n4486 ) ;
  assign n9480 = n9479 ^ n5462 ^ n4415 ;
  assign n9481 = n9480 ^ n8013 ^ n1067 ;
  assign n9482 = ( n1304 & n4588 ) | ( n1304 & ~n7732 ) | ( n4588 & ~n7732 ) ;
  assign n9483 = ( x134 & n1420 ) | ( x134 & n2931 ) | ( n1420 & n2931 ) ;
  assign n9484 = n3453 & n9483 ;
  assign n9485 = n9484 ^ n3332 ^ x64 ;
  assign n9486 = ( n4554 & ~n9482 ) | ( n4554 & n9485 ) | ( ~n9482 & n9485 ) ;
  assign n9487 = n9486 ^ n4741 ^ n1345 ;
  assign n9488 = n9487 ^ n5980 ^ n5632 ;
  assign n9490 = n5713 ^ n2974 ^ n1708 ;
  assign n9489 = ( n571 & n5275 ) | ( n571 & n6605 ) | ( n5275 & n6605 ) ;
  assign n9491 = n9490 ^ n9489 ^ n8370 ;
  assign n9492 = n8512 ^ n5207 ^ 1'b0 ;
  assign n9493 = ~n2005 & n3743 ;
  assign n9494 = n4506 ^ n3751 ^ n1325 ;
  assign n9495 = n5367 ^ n4294 ^ 1'b0 ;
  assign n9496 = ~n1386 & n9495 ;
  assign n9497 = n582 & n9496 ;
  assign n9498 = n9497 ^ n8218 ^ 1'b0 ;
  assign n9499 = ( n4442 & n7002 ) | ( n4442 & n7355 ) | ( n7002 & n7355 ) ;
  assign n9500 = n9498 & ~n9499 ;
  assign n9501 = n9500 ^ n2087 ^ 1'b0 ;
  assign n9502 = ( ~n8759 & n9494 ) | ( ~n8759 & n9501 ) | ( n9494 & n9501 ) ;
  assign n9503 = n7512 ^ n6164 ^ 1'b0 ;
  assign n9504 = n8627 | n9503 ;
  assign n9505 = n9504 ^ n7208 ^ 1'b0 ;
  assign n9506 = ( n566 & n9502 ) | ( n566 & ~n9505 ) | ( n9502 & ~n9505 ) ;
  assign n9507 = n4536 ^ x225 ^ 1'b0 ;
  assign n9508 = ~n1646 & n9507 ;
  assign n9509 = ~n4578 & n9508 ;
  assign n9510 = n5576 ^ n1916 ^ n1457 ;
  assign n9511 = n5564 | n8711 ;
  assign n9512 = n5698 | n9511 ;
  assign n9513 = n8525 ^ n296 ^ 1'b0 ;
  assign n9514 = n8699 & n9513 ;
  assign n9515 = n9514 ^ n1567 ^ 1'b0 ;
  assign n9516 = ( ~n5577 & n9512 ) | ( ~n5577 & n9515 ) | ( n9512 & n9515 ) ;
  assign n9517 = ~n8657 & n9516 ;
  assign n9518 = ~n9510 & n9517 ;
  assign n9519 = ( n7023 & ~n8825 ) | ( n7023 & n9518 ) | ( ~n8825 & n9518 ) ;
  assign n9520 = n6342 ^ n5395 ^ 1'b0 ;
  assign n9521 = n8699 & n9520 ;
  assign n9522 = n9521 ^ n3067 ^ n277 ;
  assign n9523 = n9522 ^ n8896 ^ n2803 ;
  assign n9525 = n4691 ^ n404 ^ 1'b0 ;
  assign n9524 = n4653 ^ n3804 ^ n2987 ;
  assign n9526 = n9525 ^ n9524 ^ n5182 ;
  assign n9527 = n3386 & ~n9343 ;
  assign n9528 = n9527 ^ n4673 ^ 1'b0 ;
  assign n9537 = n1511 & n6944 ;
  assign n9538 = ~n1530 & n9537 ;
  assign n9539 = x253 & ~n9538 ;
  assign n9540 = n6381 & n9539 ;
  assign n9541 = n9540 ^ n7834 ^ 1'b0 ;
  assign n9542 = n7850 & ~n9541 ;
  assign n9535 = ( x168 & ~n2750 ) | ( x168 & n8676 ) | ( ~n2750 & n8676 ) ;
  assign n9531 = ( n1449 & n2489 ) | ( n1449 & ~n5026 ) | ( n2489 & ~n5026 ) ;
  assign n9532 = n2025 & n9531 ;
  assign n9533 = ~n2364 & n9532 ;
  assign n9534 = ( n2454 & n4093 ) | ( n2454 & n9533 ) | ( n4093 & n9533 ) ;
  assign n9529 = n2977 ^ n2108 ^ 1'b0 ;
  assign n9530 = n9529 ^ n6361 ^ n5543 ;
  assign n9536 = n9535 ^ n9534 ^ n9530 ;
  assign n9543 = n9542 ^ n9536 ^ 1'b0 ;
  assign n9544 = n9528 & ~n9543 ;
  assign n9545 = n574 & n3963 ;
  assign n9546 = ~n5419 & n9545 ;
  assign n9547 = ( n787 & n2424 ) | ( n787 & ~n9546 ) | ( n2424 & ~n9546 ) ;
  assign n9548 = n2778 & n9283 ;
  assign n9549 = n2810 & n9548 ;
  assign n9550 = ( n1518 & n4089 ) | ( n1518 & ~n9549 ) | ( n4089 & ~n9549 ) ;
  assign n9552 = ( n1931 & ~n2092 ) | ( n1931 & n3967 ) | ( ~n2092 & n3967 ) ;
  assign n9553 = n5490 | n9552 ;
  assign n9551 = n324 & ~n4586 ;
  assign n9554 = n9553 ^ n9551 ^ 1'b0 ;
  assign n9555 = n9554 ^ n7121 ^ n1149 ;
  assign n9556 = n9550 & n9555 ;
  assign n9557 = n7234 ^ n5398 ^ n3160 ;
  assign n9558 = n6827 ^ n2586 ^ x19 ;
  assign n9559 = n4179 & n9558 ;
  assign n9560 = ~n9557 & n9559 ;
  assign n9561 = n9560 ^ n1093 ^ 1'b0 ;
  assign n9562 = n1505 | n9561 ;
  assign n9564 = ~n5051 & n6705 ;
  assign n9565 = ~n7398 & n9564 ;
  assign n9563 = ( n453 & n2329 ) | ( n453 & ~n6778 ) | ( n2329 & ~n6778 ) ;
  assign n9566 = n9565 ^ n9563 ^ 1'b0 ;
  assign n9567 = n2939 & ~n6243 ;
  assign n9568 = n9567 ^ n2443 ^ 1'b0 ;
  assign n9569 = n4591 & ~n9568 ;
  assign n9570 = n2199 ^ n418 ^ 1'b0 ;
  assign n9571 = ( x4 & n8423 ) | ( x4 & ~n9570 ) | ( n8423 & ~n9570 ) ;
  assign n9572 = ~n1264 & n9571 ;
  assign n9573 = n4707 & n9572 ;
  assign n9574 = ( ~n1657 & n9535 ) | ( ~n1657 & n9573 ) | ( n9535 & n9573 ) ;
  assign n9581 = n8844 ^ n6874 ^ 1'b0 ;
  assign n9582 = n4243 & ~n9581 ;
  assign n9583 = n9582 ^ n1154 ^ n562 ;
  assign n9577 = n4949 ^ n1304 ^ x66 ;
  assign n9578 = n9577 ^ n5253 ^ 1'b0 ;
  assign n9579 = x58 & n9578 ;
  assign n9575 = n8229 ^ n2526 ^ 1'b0 ;
  assign n9576 = n9575 ^ n5929 ^ x186 ;
  assign n9580 = n9579 ^ n9576 ^ n7057 ;
  assign n9584 = n9583 ^ n9580 ^ n2884 ;
  assign n9585 = n2725 & ~n4283 ;
  assign n9586 = n9585 ^ n7698 ^ 1'b0 ;
  assign n9587 = ~n3998 & n9586 ;
  assign n9601 = ~n1054 & n2404 ;
  assign n9602 = ( n628 & n3402 ) | ( n628 & n9601 ) | ( n3402 & n9601 ) ;
  assign n9603 = n5638 ^ n313 ^ x221 ;
  assign n9604 = ~n9602 & n9603 ;
  assign n9605 = n9604 ^ n1633 ^ 1'b0 ;
  assign n9595 = n924 & ~n3368 ;
  assign n9596 = n4550 & n9595 ;
  assign n9593 = ( n831 & n2325 ) | ( n831 & ~n2444 ) | ( n2325 & ~n2444 ) ;
  assign n9591 = ( n1805 & ~n3906 ) | ( n1805 & n3974 ) | ( ~n3906 & n3974 ) ;
  assign n9592 = n1467 | n9591 ;
  assign n9594 = n9593 ^ n9592 ^ x62 ;
  assign n9597 = n9596 ^ n9594 ^ n2334 ;
  assign n9598 = n6385 ^ n6307 ^ n1743 ;
  assign n9599 = ~n9597 & n9598 ;
  assign n9600 = n2535 & n9599 ;
  assign n9588 = ~n1646 & n2754 ;
  assign n9589 = n9588 ^ n2181 ^ 1'b0 ;
  assign n9590 = n9589 ^ n8068 ^ n962 ;
  assign n9606 = n9605 ^ n9600 ^ n9590 ;
  assign n9610 = ( n519 & n3973 ) | ( n519 & ~n5074 ) | ( n3973 & ~n5074 ) ;
  assign n9607 = ( n673 & n1449 ) | ( n673 & n5467 ) | ( n1449 & n5467 ) ;
  assign n9608 = n9607 ^ n4599 ^ n2634 ;
  assign n9609 = n9608 ^ n3092 ^ n1379 ;
  assign n9611 = n9610 ^ n9609 ^ n8178 ;
  assign n9612 = n9611 ^ n7155 ^ n607 ;
  assign n9613 = n1367 ^ n993 ^ n586 ;
  assign n9614 = n750 ^ n602 ^ 1'b0 ;
  assign n9615 = n9614 ^ n4583 ^ 1'b0 ;
  assign n9616 = n9613 | n9615 ;
  assign n9617 = n2106 | n2378 ;
  assign n9618 = n9616 & ~n9617 ;
  assign n9619 = n1602 | n6614 ;
  assign n9624 = n7172 ^ n5117 ^ n2243 ;
  assign n9625 = ( n3429 & n6212 ) | ( n3429 & n6377 ) | ( n6212 & n6377 ) ;
  assign n9626 = ( n4694 & n9624 ) | ( n4694 & ~n9625 ) | ( n9624 & ~n9625 ) ;
  assign n9620 = ~n1433 & n6361 ;
  assign n9621 = n9620 ^ n5607 ^ 1'b0 ;
  assign n9622 = n6182 & ~n6241 ;
  assign n9623 = n9621 & n9622 ;
  assign n9627 = n9626 ^ n9623 ^ n1752 ;
  assign n9632 = n5798 ^ n4931 ^ n979 ;
  assign n9633 = n7017 ^ n1143 ^ 1'b0 ;
  assign n9634 = n1313 | n9633 ;
  assign n9639 = ( x97 & n470 ) | ( x97 & n982 ) | ( n470 & n982 ) ;
  assign n9635 = ( n995 & n1689 ) | ( n995 & ~n1902 ) | ( n1689 & ~n1902 ) ;
  assign n9636 = n5194 & n9197 ;
  assign n9637 = n9635 & n9636 ;
  assign n9638 = ( n2598 & ~n2832 ) | ( n2598 & n9637 ) | ( ~n2832 & n9637 ) ;
  assign n9640 = n9639 ^ n9638 ^ n7398 ;
  assign n9641 = ( n9632 & n9634 ) | ( n9632 & n9640 ) | ( n9634 & n9640 ) ;
  assign n9628 = n1642 & n8584 ;
  assign n9629 = n9628 ^ n3484 ^ 1'b0 ;
  assign n9630 = n2044 | n9629 ;
  assign n9631 = n9630 ^ n5705 ^ 1'b0 ;
  assign n9642 = n9641 ^ n9631 ^ n5522 ;
  assign n9648 = n5774 ^ n3154 ^ n1737 ;
  assign n9643 = ( x100 & ~n4371 ) | ( x100 & n4928 ) | ( ~n4371 & n4928 ) ;
  assign n9644 = n9643 ^ n4341 ^ n266 ;
  assign n9645 = n4464 ^ n3596 ^ 1'b0 ;
  assign n9646 = n9644 & n9645 ;
  assign n9647 = ~n284 & n9646 ;
  assign n9649 = n9648 ^ n9647 ^ 1'b0 ;
  assign n9650 = n9460 ^ n4557 ^ n1378 ;
  assign n9651 = n8535 ^ n7768 ^ n366 ;
  assign n9652 = x97 & ~n9651 ;
  assign n9653 = n9652 ^ n6867 ^ 1'b0 ;
  assign n9654 = n2135 ^ n1496 ^ 1'b0 ;
  assign n9655 = n4431 & n9654 ;
  assign n9656 = ( n9650 & ~n9653 ) | ( n9650 & n9655 ) | ( ~n9653 & n9655 ) ;
  assign n9657 = n942 & n4428 ;
  assign n9658 = n7636 ^ n306 ^ 1'b0 ;
  assign n9659 = n7609 ^ n6754 ^ 1'b0 ;
  assign n9660 = n3802 ^ n1896 ^ 1'b0 ;
  assign n9661 = n8228 & ~n9660 ;
  assign n9662 = ( n704 & ~n1991 ) | ( n704 & n8673 ) | ( ~n1991 & n8673 ) ;
  assign n9663 = ( n6271 & n6776 ) | ( n6271 & ~n9662 ) | ( n6776 & ~n9662 ) ;
  assign n9664 = n9663 ^ n8871 ^ n5689 ;
  assign n9665 = n8705 ^ n3399 ^ 1'b0 ;
  assign n9666 = ~n6211 & n9665 ;
  assign n9667 = ( ~n3949 & n6170 ) | ( ~n3949 & n9666 ) | ( n6170 & n9666 ) ;
  assign n9668 = n9667 ^ n4440 ^ 1'b0 ;
  assign n9675 = ( n2094 & n2161 ) | ( n2094 & ~n3593 ) | ( n2161 & ~n3593 ) ;
  assign n9669 = ( n866 & n2791 ) | ( n866 & n4493 ) | ( n2791 & n4493 ) ;
  assign n9670 = n9669 ^ n2686 ^ n382 ;
  assign n9671 = n6039 ^ n3857 ^ n2880 ;
  assign n9672 = n4197 | n9671 ;
  assign n9673 = n9672 ^ n5261 ^ 1'b0 ;
  assign n9674 = ( ~n4623 & n9670 ) | ( ~n4623 & n9673 ) | ( n9670 & n9673 ) ;
  assign n9676 = n9675 ^ n9674 ^ n7961 ;
  assign n9677 = n3500 ^ n2579 ^ 1'b0 ;
  assign n9678 = n9677 ^ n300 ^ 1'b0 ;
  assign n9679 = n4079 ^ n2722 ^ n461 ;
  assign n9680 = n6175 | n7268 ;
  assign n9681 = n9679 | n9680 ;
  assign n9682 = n4277 ^ n3806 ^ 1'b0 ;
  assign n9683 = ~n2492 & n9682 ;
  assign n9684 = n9683 ^ n5829 ^ n1085 ;
  assign n9686 = ( n1565 & n4363 ) | ( n1565 & ~n4447 ) | ( n4363 & ~n4447 ) ;
  assign n9685 = x109 & n3310 ;
  assign n9687 = n9686 ^ n9685 ^ 1'b0 ;
  assign n9688 = ( n3165 & n7162 ) | ( n3165 & ~n9687 ) | ( n7162 & ~n9687 ) ;
  assign n9689 = ( ~n3858 & n9684 ) | ( ~n3858 & n9688 ) | ( n9684 & n9688 ) ;
  assign n9690 = n3039 & n5997 ;
  assign n9691 = n8855 ^ n8647 ^ n2705 ;
  assign n9692 = ( n552 & n2283 ) | ( n552 & ~n2950 ) | ( n2283 & ~n2950 ) ;
  assign n9694 = n3623 ^ n2161 ^ 1'b0 ;
  assign n9693 = ~n4181 & n5095 ;
  assign n9695 = n9694 ^ n9693 ^ 1'b0 ;
  assign n9696 = n7251 ^ n4017 ^ 1'b0 ;
  assign n9697 = n9695 | n9696 ;
  assign n9698 = x102 & n9697 ;
  assign n9699 = ~n1137 & n9698 ;
  assign n9700 = ~n3915 & n9699 ;
  assign n9701 = n1042 ^ x215 ^ 1'b0 ;
  assign n9702 = n9282 ^ n7000 ^ 1'b0 ;
  assign n9703 = n9701 | n9702 ;
  assign n9704 = ( n2885 & ~n3416 ) | ( n2885 & n9316 ) | ( ~n3416 & n9316 ) ;
  assign n9705 = n9704 ^ n8142 ^ n3803 ;
  assign n9706 = n1753 ^ n649 ^ x190 ;
  assign n9707 = n9706 ^ n6933 ^ n2125 ;
  assign n9708 = n9707 ^ n5291 ^ 1'b0 ;
  assign n9709 = n7335 & n9708 ;
  assign n9710 = ~n6776 & n9709 ;
  assign n9711 = ~n4723 & n9710 ;
  assign n9712 = n2055 | n2658 ;
  assign n9713 = n9712 ^ n7093 ^ 1'b0 ;
  assign n9714 = ~n9711 & n9713 ;
  assign n9715 = n9714 ^ n6954 ^ 1'b0 ;
  assign n9716 = ~n2515 & n9715 ;
  assign n9717 = n9716 ^ n4296 ^ 1'b0 ;
  assign n9718 = ( ~n2318 & n2352 ) | ( ~n2318 & n4069 ) | ( n2352 & n4069 ) ;
  assign n9719 = n2194 & n9718 ;
  assign n9720 = n6012 & n6317 ;
  assign n9721 = n9719 & n9720 ;
  assign n9722 = ( n7060 & n9717 ) | ( n7060 & ~n9721 ) | ( n9717 & ~n9721 ) ;
  assign n9723 = n9722 ^ n4465 ^ n2510 ;
  assign n9725 = ~n334 & n4154 ;
  assign n9726 = n3446 & n9725 ;
  assign n9727 = n1890 & n9726 ;
  assign n9724 = n5212 | n5588 ;
  assign n9728 = n9727 ^ n9724 ^ 1'b0 ;
  assign n9729 = ( ~n5838 & n8264 ) | ( ~n5838 & n9728 ) | ( n8264 & n9728 ) ;
  assign n9730 = ~n6798 & n8630 ;
  assign n9731 = n9730 ^ n8829 ^ n5952 ;
  assign n9732 = n2927 & n6957 ;
  assign n9733 = n9732 ^ n3258 ^ 1'b0 ;
  assign n9735 = n9589 ^ n6608 ^ n6242 ;
  assign n9736 = n9735 ^ n5415 ^ n2886 ;
  assign n9734 = x157 & n2452 ;
  assign n9737 = n9736 ^ n9734 ^ 1'b0 ;
  assign n9738 = ( n4066 & n6520 ) | ( n4066 & n9737 ) | ( n6520 & n9737 ) ;
  assign n9739 = ( n849 & n1904 ) | ( n849 & n9738 ) | ( n1904 & n9738 ) ;
  assign n9740 = n9733 | n9739 ;
  assign n9741 = n7967 ^ n2937 ^ n1052 ;
  assign n9743 = n2967 ^ n933 ^ 1'b0 ;
  assign n9744 = x136 & n9743 ;
  assign n9745 = n9744 ^ n5418 ^ n1735 ;
  assign n9746 = n9745 ^ n6813 ^ 1'b0 ;
  assign n9747 = n3593 ^ n2453 ^ 1'b0 ;
  assign n9748 = n7661 ^ n3745 ^ n615 ;
  assign n9749 = ( n9179 & n9747 ) | ( n9179 & ~n9748 ) | ( n9747 & ~n9748 ) ;
  assign n9750 = ( n4418 & n9746 ) | ( n4418 & n9749 ) | ( n9746 & n9749 ) ;
  assign n9742 = n7128 ^ n4991 ^ n3082 ;
  assign n9751 = n9750 ^ n9742 ^ n1120 ;
  assign n9753 = n7909 ^ n2688 ^ n2086 ;
  assign n9752 = n5381 | n5834 ;
  assign n9754 = n9753 ^ n9752 ^ 1'b0 ;
  assign n9755 = ( x26 & n1930 ) | ( x26 & n3111 ) | ( n1930 & n3111 ) ;
  assign n9756 = n9755 ^ n6054 ^ 1'b0 ;
  assign n9757 = ~n9754 & n9756 ;
  assign n9758 = n3342 ^ n1295 ^ n516 ;
  assign n9759 = ~n8145 & n9758 ;
  assign n9760 = ~n1511 & n9759 ;
  assign n9761 = n8090 ^ n2479 ^ 1'b0 ;
  assign n9762 = ~n4414 & n9761 ;
  assign n9763 = ( x243 & ~n585 ) | ( x243 & n5424 ) | ( ~n585 & n5424 ) ;
  assign n9764 = n5875 & ~n9763 ;
  assign n9765 = n9764 ^ n5790 ^ 1'b0 ;
  assign n9766 = ( n1341 & n2206 ) | ( n1341 & ~n9765 ) | ( n2206 & ~n9765 ) ;
  assign n9772 = n2591 ^ n2548 ^ n788 ;
  assign n9770 = n3906 ^ n1099 ^ 1'b0 ;
  assign n9771 = n340 & ~n9770 ;
  assign n9767 = n8770 & n9450 ;
  assign n9768 = n2826 ^ n2630 ^ 1'b0 ;
  assign n9769 = n9767 & ~n9768 ;
  assign n9773 = n9772 ^ n9771 ^ n9769 ;
  assign n9774 = ( n2764 & n3255 ) | ( n2764 & ~n7807 ) | ( n3255 & ~n7807 ) ;
  assign n9775 = ( ~n1736 & n2547 ) | ( ~n1736 & n9774 ) | ( n2547 & n9774 ) ;
  assign n9776 = ( ~n2489 & n3190 ) | ( ~n2489 & n9775 ) | ( n3190 & n9775 ) ;
  assign n9783 = n9283 ^ n8771 ^ n3651 ;
  assign n9778 = n8177 ^ n6149 ^ n536 ;
  assign n9779 = n1616 ^ n582 ^ 1'b0 ;
  assign n9780 = n8187 & n9779 ;
  assign n9781 = ( n1869 & n4406 ) | ( n1869 & n7490 ) | ( n4406 & n7490 ) ;
  assign n9782 = ( ~n9778 & n9780 ) | ( ~n9778 & n9781 ) | ( n9780 & n9781 ) ;
  assign n9777 = ( x245 & ~n2035 ) | ( x245 & n9624 ) | ( ~n2035 & n9624 ) ;
  assign n9784 = n9783 ^ n9782 ^ n9777 ;
  assign n9785 = n3528 & n7386 ;
  assign n9786 = n9785 ^ n5733 ^ 1'b0 ;
  assign n9787 = n7995 | n9786 ;
  assign n9788 = n3824 & n9787 ;
  assign n9789 = n3377 | n9788 ;
  assign n9790 = ( n2714 & n6117 ) | ( n2714 & n9789 ) | ( n6117 & n9789 ) ;
  assign n9791 = n3038 & n9790 ;
  assign n9792 = ~n4294 & n6402 ;
  assign n9806 = n9317 ^ n5638 ^ 1'b0 ;
  assign n9807 = n3695 & n9806 ;
  assign n9793 = n4092 ^ n2557 ^ n2342 ;
  assign n9794 = n4260 ^ n3166 ^ n1120 ;
  assign n9795 = n9794 ^ n6623 ^ n3326 ;
  assign n9797 = n3188 & ~n3222 ;
  assign n9798 = n7227 & ~n8630 ;
  assign n9799 = n9797 & n9798 ;
  assign n9800 = n9799 ^ n1845 ^ x70 ;
  assign n9796 = n2586 ^ x149 ^ 1'b0 ;
  assign n9801 = n9800 ^ n9796 ^ 1'b0 ;
  assign n9802 = n1206 & n9801 ;
  assign n9803 = n1344 & n9802 ;
  assign n9804 = n9803 ^ n9248 ^ 1'b0 ;
  assign n9805 = ( n9793 & ~n9795 ) | ( n9793 & n9804 ) | ( ~n9795 & n9804 ) ;
  assign n9808 = n9807 ^ n9805 ^ n4675 ;
  assign n9810 = n1883 | n7965 ;
  assign n9811 = n8609 ^ n1244 ^ n288 ;
  assign n9812 = n1943 | n9811 ;
  assign n9813 = ( n6862 & ~n9810 ) | ( n6862 & n9812 ) | ( ~n9810 & n9812 ) ;
  assign n9809 = n898 & n6933 ;
  assign n9814 = n9813 ^ n9809 ^ 1'b0 ;
  assign n9815 = ( n356 & ~n6709 ) | ( n356 & n6925 ) | ( ~n6709 & n6925 ) ;
  assign n9816 = n9815 ^ n5594 ^ n2729 ;
  assign n9817 = n1159 & ~n4149 ;
  assign n9818 = n7443 & n9817 ;
  assign n9819 = ~n2098 & n7275 ;
  assign n9820 = n9818 & n9819 ;
  assign n9821 = n2519 & ~n2809 ;
  assign n9822 = n9821 ^ n4437 ^ 1'b0 ;
  assign n9823 = n6875 & ~n9822 ;
  assign n9824 = n2715 ^ n2701 ^ 1'b0 ;
  assign n9825 = n3039 & n9824 ;
  assign n9826 = n7878 ^ x64 ^ 1'b0 ;
  assign n9827 = n9825 & ~n9826 ;
  assign n9828 = n6527 ^ n3429 ^ n1485 ;
  assign n9829 = n9828 ^ n3824 ^ n2043 ;
  assign n9830 = ( n3104 & ~n6917 ) | ( n3104 & n8402 ) | ( ~n6917 & n8402 ) ;
  assign n9831 = ( n2895 & n6378 ) | ( n2895 & n9830 ) | ( n6378 & n9830 ) ;
  assign n9832 = ~n798 & n9831 ;
  assign n9833 = ~n9829 & n9832 ;
  assign n9834 = n4564 ^ n3971 ^ 1'b0 ;
  assign n9835 = n4685 | n9834 ;
  assign n9836 = n9835 ^ n1868 ^ n1650 ;
  assign n9838 = n4894 ^ n2862 ^ n1317 ;
  assign n9837 = n1358 & ~n4191 ;
  assign n9839 = n9838 ^ n9837 ^ 1'b0 ;
  assign n9840 = ( ~x97 & x112 ) | ( ~x97 & n9839 ) | ( x112 & n9839 ) ;
  assign n9841 = n5658 ^ n541 ^ 1'b0 ;
  assign n9842 = n433 & n9841 ;
  assign n9843 = ( x100 & n9840 ) | ( x100 & n9842 ) | ( n9840 & n9842 ) ;
  assign n9844 = ( n5546 & n6660 ) | ( n5546 & n9843 ) | ( n6660 & n9843 ) ;
  assign n9845 = n5588 | n7661 ;
  assign n9846 = n9845 ^ n7022 ^ 1'b0 ;
  assign n9848 = n5080 ^ n360 ^ 1'b0 ;
  assign n9847 = n7544 ^ n6300 ^ n3012 ;
  assign n9849 = n9848 ^ n9847 ^ 1'b0 ;
  assign n9850 = n7779 | n9849 ;
  assign n9851 = ~n4503 & n5457 ;
  assign n9852 = ( ~n6430 & n9165 ) | ( ~n6430 & n9851 ) | ( n9165 & n9851 ) ;
  assign n9853 = ( ~n1265 & n1729 ) | ( ~n1265 & n2350 ) | ( n1729 & n2350 ) ;
  assign n9854 = n5751 & ~n9853 ;
  assign n9855 = ~n3268 & n3441 ;
  assign n9859 = ( n1185 & n3379 ) | ( n1185 & n4879 ) | ( n3379 & n4879 ) ;
  assign n9856 = n2429 & ~n5685 ;
  assign n9857 = n9856 ^ n5725 ^ 1'b0 ;
  assign n9858 = n1574 | n9857 ;
  assign n9860 = n9859 ^ n9858 ^ 1'b0 ;
  assign n9861 = n3833 & ~n9860 ;
  assign n9865 = ~n2018 & n7735 ;
  assign n9866 = n9865 ^ n6489 ^ 1'b0 ;
  assign n9863 = n4614 ^ n4211 ^ n1702 ;
  assign n9862 = ~n2865 & n4752 ;
  assign n9864 = n9863 ^ n9862 ^ 1'b0 ;
  assign n9867 = n9866 ^ n9864 ^ n1355 ;
  assign n9868 = ( n8771 & n9861 ) | ( n8771 & ~n9867 ) | ( n9861 & ~n9867 ) ;
  assign n9872 = n3417 ^ n1550 ^ n1093 ;
  assign n9871 = n3684 ^ n1950 ^ 1'b0 ;
  assign n9869 = n6420 ^ n2175 ^ 1'b0 ;
  assign n9870 = ( n4417 & n6590 ) | ( n4417 & ~n9869 ) | ( n6590 & ~n9869 ) ;
  assign n9873 = n9872 ^ n9871 ^ n9870 ;
  assign n9883 = n7230 ^ n2678 ^ 1'b0 ;
  assign n9882 = n3365 | n4101 ;
  assign n9884 = n9883 ^ n9882 ^ 1'b0 ;
  assign n9877 = n8389 ^ n5858 ^ n4284 ;
  assign n9876 = ~n901 & n5234 ;
  assign n9878 = n9877 ^ n9876 ^ 1'b0 ;
  assign n9879 = ( n2496 & n9193 ) | ( n2496 & n9878 ) | ( n9193 & n9878 ) ;
  assign n9880 = n9879 ^ n4405 ^ n288 ;
  assign n9874 = ( n1492 & ~n1773 ) | ( n1492 & n3958 ) | ( ~n1773 & n3958 ) ;
  assign n9875 = n9863 & ~n9874 ;
  assign n9881 = n9880 ^ n9875 ^ 1'b0 ;
  assign n9885 = n9884 ^ n9881 ^ n9562 ;
  assign n9886 = n2958 ^ n2895 ^ n1801 ;
  assign n9887 = ~n1622 & n5023 ;
  assign n9888 = ~n1326 & n9887 ;
  assign n9890 = ( n1355 & n1618 ) | ( n1355 & n6894 ) | ( n1618 & n6894 ) ;
  assign n9889 = n1210 | n5383 ;
  assign n9891 = n9890 ^ n9889 ^ 1'b0 ;
  assign n9892 = ( n9886 & ~n9888 ) | ( n9886 & n9891 ) | ( ~n9888 & n9891 ) ;
  assign n9893 = n8201 ^ n349 ^ 1'b0 ;
  assign n9894 = n9892 & ~n9893 ;
  assign n9895 = n7868 ^ n5194 ^ n1162 ;
  assign n9896 = n994 | n9895 ;
  assign n9897 = ( n2019 & ~n7035 ) | ( n2019 & n9896 ) | ( ~n7035 & n9896 ) ;
  assign n9898 = n2620 ^ n1266 ^ x77 ;
  assign n9899 = n9898 ^ n8775 ^ n2853 ;
  assign n9904 = n2055 | n2989 ;
  assign n9905 = n9904 ^ n7591 ^ 1'b0 ;
  assign n9901 = n6116 ^ n3227 ^ n2047 ;
  assign n9902 = n9901 ^ n5858 ^ n4063 ;
  assign n9903 = n9902 ^ n4983 ^ n3546 ;
  assign n9900 = ( n3214 & n5257 ) | ( n3214 & ~n6674 ) | ( n5257 & ~n6674 ) ;
  assign n9906 = n9905 ^ n9903 ^ n9900 ;
  assign n9907 = n7395 ^ n7233 ^ 1'b0 ;
  assign n9908 = ~n5386 & n9907 ;
  assign n9910 = n2347 ^ n1041 ^ 1'b0 ;
  assign n9909 = x28 & n9228 ;
  assign n9911 = n9910 ^ n9909 ^ 1'b0 ;
  assign n9912 = n9908 | n9911 ;
  assign n9913 = x91 | n620 ;
  assign n9914 = n9913 ^ n2640 ^ n2146 ;
  assign n9915 = n9914 ^ n2029 ^ n452 ;
  assign n9919 = n4644 ^ n1935 ^ x212 ;
  assign n9917 = ( n459 & ~n2645 ) | ( n459 & n3189 ) | ( ~n2645 & n3189 ) ;
  assign n9918 = n9917 ^ n4822 ^ n1852 ;
  assign n9920 = n9919 ^ n9918 ^ n2399 ;
  assign n9916 = n2694 & ~n4917 ;
  assign n9921 = n9920 ^ n9916 ^ 1'b0 ;
  assign n9922 = n4423 | n9921 ;
  assign n9923 = n7736 | n9922 ;
  assign n9924 = ( n2904 & n3622 ) | ( n2904 & n4640 ) | ( n3622 & n4640 ) ;
  assign n9925 = n500 & n9924 ;
  assign n9926 = ~n8513 & n9925 ;
  assign n9927 = ( n2901 & n4955 ) | ( n2901 & ~n7049 ) | ( n4955 & ~n7049 ) ;
  assign n9928 = n5968 | n9927 ;
  assign n9929 = n8300 & ~n9928 ;
  assign n9930 = n1793 | n9929 ;
  assign n9931 = ( ~n344 & n1487 ) | ( ~n344 & n4817 ) | ( n1487 & n4817 ) ;
  assign n9932 = ( n3624 & n4862 ) | ( n3624 & n9931 ) | ( n4862 & n9931 ) ;
  assign n9933 = n8020 | n9932 ;
  assign n9934 = n9930 | n9933 ;
  assign n9935 = ~n9926 & n9934 ;
  assign n9936 = ~n9923 & n9935 ;
  assign n9937 = n8611 ^ n6621 ^ n5062 ;
  assign n9938 = n6961 ^ n3255 ^ n1200 ;
  assign n9944 = n5764 ^ n2237 ^ 1'b0 ;
  assign n9939 = n8252 ^ n1599 ^ 1'b0 ;
  assign n9940 = ~n5750 & n9939 ;
  assign n9941 = ( n1738 & n4718 ) | ( n1738 & ~n9940 ) | ( n4718 & ~n9940 ) ;
  assign n9942 = n3742 ^ n3249 ^ 1'b0 ;
  assign n9943 = n9941 | n9942 ;
  assign n9945 = n9944 ^ n9943 ^ n1120 ;
  assign n9949 = n1290 | n3617 ;
  assign n9946 = n3447 ^ n1024 ^ n758 ;
  assign n9947 = ( ~n4581 & n7150 ) | ( ~n4581 & n9946 ) | ( n7150 & n9946 ) ;
  assign n9948 = n9313 & ~n9947 ;
  assign n9950 = n9949 ^ n9948 ^ 1'b0 ;
  assign n9951 = n3056 & ~n9950 ;
  assign n9952 = n849 & n4870 ;
  assign n9953 = n7885 | n9952 ;
  assign n9954 = ( n984 & n9951 ) | ( n984 & n9953 ) | ( n9951 & n9953 ) ;
  assign n9955 = n2295 ^ n563 ^ x45 ;
  assign n9956 = n9955 ^ n2516 ^ n2036 ;
  assign n9957 = n7125 ^ n3812 ^ 1'b0 ;
  assign n9958 = ( n9678 & n9956 ) | ( n9678 & n9957 ) | ( n9956 & n9957 ) ;
  assign n9959 = ( ~n755 & n3303 ) | ( ~n755 & n5129 ) | ( n3303 & n5129 ) ;
  assign n9960 = n6117 & n9959 ;
  assign n9961 = n7178 ^ n1402 ^ 1'b0 ;
  assign n9962 = n8270 ^ n3792 ^ x193 ;
  assign n9963 = n5383 ^ n3078 ^ 1'b0 ;
  assign n9964 = ( n4397 & n6468 ) | ( n4397 & n9963 ) | ( n6468 & n9963 ) ;
  assign n9965 = n1070 & n5477 ;
  assign n9966 = n9965 ^ n4743 ^ n3383 ;
  assign n9967 = ( n5109 & n7632 ) | ( n5109 & n9878 ) | ( n7632 & n9878 ) ;
  assign n9971 = n9269 ^ n6591 ^ 1'b0 ;
  assign n9972 = ( n4787 & n6880 ) | ( n4787 & n9064 ) | ( n6880 & n9064 ) ;
  assign n9973 = n9972 ^ n2932 ^ 1'b0 ;
  assign n9974 = x245 & ~n9973 ;
  assign n9975 = n4611 & n9974 ;
  assign n9976 = n9971 & n9975 ;
  assign n9968 = n6240 & n7848 ;
  assign n9969 = n9968 ^ n4295 ^ 1'b0 ;
  assign n9970 = n3108 | n9969 ;
  assign n9977 = n9976 ^ n9970 ^ 1'b0 ;
  assign n9983 = ( n668 & n762 ) | ( n668 & n1981 ) | ( n762 & n1981 ) ;
  assign n9979 = ~n659 & n1976 ;
  assign n9978 = n1376 & ~n5716 ;
  assign n9980 = n9979 ^ n9978 ^ 1'b0 ;
  assign n9981 = n9828 & n9980 ;
  assign n9982 = n9981 ^ n9955 ^ 1'b0 ;
  assign n9984 = n9983 ^ n9982 ^ 1'b0 ;
  assign n9985 = n1820 & n9984 ;
  assign n9986 = ( ~x58 & n4180 ) | ( ~x58 & n7362 ) | ( n4180 & n7362 ) ;
  assign n9987 = n9985 & n9986 ;
  assign n9988 = ~n3614 & n9987 ;
  assign n9989 = n1515 & ~n9988 ;
  assign n9990 = ~n7317 & n9989 ;
  assign n9991 = n2549 | n3872 ;
  assign n9992 = n9991 ^ n494 ^ 1'b0 ;
  assign n9993 = n9992 ^ n4368 ^ 1'b0 ;
  assign n9994 = ( x199 & ~n4134 ) | ( x199 & n9993 ) | ( ~n4134 & n9993 ) ;
  assign n9995 = n310 | n4807 ;
  assign n9996 = n9995 ^ n3129 ^ n2275 ;
  assign n10003 = ~n5287 & n6340 ;
  assign n10004 = ~n9716 & n10003 ;
  assign n10001 = ( ~n3208 & n6299 ) | ( ~n3208 & n7645 ) | ( n6299 & n7645 ) ;
  assign n9997 = ( ~n1188 & n2415 ) | ( ~n1188 & n3811 ) | ( n2415 & n3811 ) ;
  assign n9998 = n9997 ^ n7506 ^ n1473 ;
  assign n9999 = n7095 ^ n6346 ^ n2170 ;
  assign n10000 = n9998 & n9999 ;
  assign n10002 = n10001 ^ n10000 ^ 1'b0 ;
  assign n10005 = n10004 ^ n10002 ^ n5629 ;
  assign n10006 = ~n7102 & n10005 ;
  assign n10007 = n3707 ^ n3358 ^ n2969 ;
  assign n10008 = n10007 ^ n289 ^ 1'b0 ;
  assign n10009 = n7603 ^ n4501 ^ 1'b0 ;
  assign n10010 = n5740 | n10009 ;
  assign n10011 = ( n431 & n812 ) | ( n431 & ~n10010 ) | ( n812 & ~n10010 ) ;
  assign n10012 = n3606 ^ n333 ^ 1'b0 ;
  assign n10013 = ( ~n9014 & n10011 ) | ( ~n9014 & n10012 ) | ( n10011 & n10012 ) ;
  assign n10014 = n828 ^ n488 ^ 1'b0 ;
  assign n10015 = n3462 & ~n4440 ;
  assign n10016 = n10015 ^ n6754 ^ 1'b0 ;
  assign n10017 = ( ~n4635 & n10014 ) | ( ~n4635 & n10016 ) | ( n10014 & n10016 ) ;
  assign n10021 = n6330 ^ n4441 ^ n3856 ;
  assign n10022 = n10021 ^ n6383 ^ n3611 ;
  assign n10018 = n4717 | n8438 ;
  assign n10019 = n10018 ^ n1897 ^ 1'b0 ;
  assign n10020 = n10019 ^ n6270 ^ n3884 ;
  assign n10023 = n10022 ^ n10020 ^ 1'b0 ;
  assign n10024 = ( n5831 & n7944 ) | ( n5831 & ~n8258 ) | ( n7944 & ~n8258 ) ;
  assign n10025 = n6768 ^ n4404 ^ n3932 ;
  assign n10026 = n6849 ^ n471 ^ 1'b0 ;
  assign n10027 = ( n5812 & n8567 ) | ( n5812 & ~n10026 ) | ( n8567 & ~n10026 ) ;
  assign n10028 = n8311 ^ n4389 ^ 1'b0 ;
  assign n10029 = n1306 | n2205 ;
  assign n10030 = n3917 | n10029 ;
  assign n10031 = ( n2157 & n3420 ) | ( n2157 & n10030 ) | ( n3420 & n10030 ) ;
  assign n10032 = ( n8297 & ~n10028 ) | ( n8297 & n10031 ) | ( ~n10028 & n10031 ) ;
  assign n10037 = ( x15 & ~n2139 ) | ( x15 & n4064 ) | ( ~n2139 & n4064 ) ;
  assign n10033 = n6191 ^ n3391 ^ n1473 ;
  assign n10034 = n10033 ^ n4414 ^ n3793 ;
  assign n10035 = n3141 & ~n10034 ;
  assign n10036 = n4388 & n10035 ;
  assign n10038 = n10037 ^ n10036 ^ n8694 ;
  assign n10039 = n9570 ^ n2699 ^ 1'b0 ;
  assign n10040 = n468 & ~n10039 ;
  assign n10041 = n10040 ^ n6005 ^ 1'b0 ;
  assign n10042 = n4429 & n6376 ;
  assign n10043 = n10042 ^ n2311 ^ 1'b0 ;
  assign n10044 = n3802 & n10043 ;
  assign n10045 = n8720 & n10044 ;
  assign n10046 = n387 & ~n10045 ;
  assign n10047 = n10046 ^ n3721 ^ 1'b0 ;
  assign n10048 = n1570 | n2519 ;
  assign n10049 = n3379 & n10048 ;
  assign n10050 = n10049 ^ n3988 ^ n1995 ;
  assign n10051 = ( n4935 & n4991 ) | ( n4935 & ~n10050 ) | ( n4991 & ~n10050 ) ;
  assign n10052 = ( n3435 & ~n4925 ) | ( n3435 & n10051 ) | ( ~n4925 & n10051 ) ;
  assign n10053 = n3090 & n5353 ;
  assign n10054 = n8517 ^ n4780 ^ 1'b0 ;
  assign n10055 = x232 ^ x134 ^ 1'b0 ;
  assign n10056 = ~n7925 & n10055 ;
  assign n10057 = n10056 ^ n4006 ^ 1'b0 ;
  assign n10058 = n9226 ^ n4235 ^ n2712 ;
  assign n10059 = ( n1113 & n1384 ) | ( n1113 & ~n6041 ) | ( n1384 & ~n6041 ) ;
  assign n10060 = ( n4267 & n4460 ) | ( n4267 & n10059 ) | ( n4460 & n10059 ) ;
  assign n10061 = n10060 ^ n1431 ^ n598 ;
  assign n10062 = ~n10058 & n10061 ;
  assign n10063 = n4820 | n5753 ;
  assign n10064 = n2866 & ~n10063 ;
  assign n10067 = n8548 ^ n4487 ^ n471 ;
  assign n10068 = n10067 ^ n7627 ^ n1106 ;
  assign n10065 = ( n501 & ~n1574 ) | ( n501 & n2389 ) | ( ~n1574 & n2389 ) ;
  assign n10066 = n10065 ^ n4794 ^ x131 ;
  assign n10069 = n10068 ^ n10066 ^ 1'b0 ;
  assign n10070 = n2028 & ~n10069 ;
  assign n10078 = n1983 & n4476 ;
  assign n10079 = ~n8520 & n10078 ;
  assign n10073 = n1251 | n2877 ;
  assign n10074 = n10073 ^ n2798 ^ 1'b0 ;
  assign n10075 = n10074 ^ n5398 ^ n2256 ;
  assign n10071 = n728 & ~n1251 ;
  assign n10072 = n1732 & n10071 ;
  assign n10076 = n10075 ^ n10072 ^ 1'b0 ;
  assign n10077 = ~n4808 & n10076 ;
  assign n10080 = n10079 ^ n10077 ^ 1'b0 ;
  assign n10082 = ( n796 & ~n885 ) | ( n796 & n2382 ) | ( ~n885 & n2382 ) ;
  assign n10081 = n1555 | n3581 ;
  assign n10083 = n10082 ^ n10081 ^ n4903 ;
  assign n10084 = n10083 ^ n7099 ^ 1'b0 ;
  assign n10085 = ( n1219 & ~n3580 ) | ( n1219 & n10084 ) | ( ~n3580 & n10084 ) ;
  assign n10087 = n4937 ^ x218 ^ 1'b0 ;
  assign n10088 = n10087 ^ n9274 ^ n6709 ;
  assign n10086 = n8161 ^ n7429 ^ n1519 ;
  assign n10089 = n10088 ^ n10086 ^ n3525 ;
  assign n10095 = n3178 ^ n1296 ^ n956 ;
  assign n10093 = n7907 ^ n2526 ^ n783 ;
  assign n10094 = n10093 ^ n662 ^ 1'b0 ;
  assign n10091 = x68 & ~n920 ;
  assign n10090 = n3374 ^ n2470 ^ n1498 ;
  assign n10092 = n10091 ^ n10090 ^ 1'b0 ;
  assign n10096 = n10095 ^ n10094 ^ n10092 ;
  assign n10106 = n6397 ^ x73 ^ 1'b0 ;
  assign n10099 = n2319 & n3377 ;
  assign n10100 = ~n4919 & n10099 ;
  assign n10101 = n9317 ^ n6217 ^ n5022 ;
  assign n10102 = n10100 | n10101 ;
  assign n10103 = n6334 | n10102 ;
  assign n10104 = n10103 ^ n7866 ^ 1'b0 ;
  assign n10105 = n2353 | n10104 ;
  assign n10097 = n436 & ~n7174 ;
  assign n10098 = ~n7999 & n10097 ;
  assign n10107 = n10106 ^ n10105 ^ n10098 ;
  assign n10108 = ~n1152 & n8720 ;
  assign n10109 = n10108 ^ n5696 ^ n1959 ;
  assign n10114 = n6172 ^ n3036 ^ 1'b0 ;
  assign n10115 = n10114 ^ n4792 ^ n2889 ;
  assign n10116 = n6396 & ~n10115 ;
  assign n10117 = n10116 ^ n2454 ^ 1'b0 ;
  assign n10110 = n5581 ^ n4241 ^ 1'b0 ;
  assign n10111 = n4004 & n10110 ;
  assign n10112 = n2233 & ~n10111 ;
  assign n10113 = n6246 & ~n10112 ;
  assign n10118 = n10117 ^ n10113 ^ 1'b0 ;
  assign n10119 = ( n2795 & n10109 ) | ( n2795 & n10118 ) | ( n10109 & n10118 ) ;
  assign n10120 = n6489 & ~n9772 ;
  assign n10121 = n10120 ^ n1060 ^ 1'b0 ;
  assign n10122 = x53 & n10121 ;
  assign n10123 = ~x229 & n10122 ;
  assign n10124 = n8742 & ~n10123 ;
  assign n10125 = n10124 ^ n3152 ^ n1659 ;
  assign n10126 = n10125 ^ n4118 ^ 1'b0 ;
  assign n10127 = n3978 & ~n10126 ;
  assign n10128 = ( n2774 & n3084 ) | ( n2774 & n10127 ) | ( n3084 & n10127 ) ;
  assign n10138 = ~n666 & n3736 ;
  assign n10139 = n2827 & n10138 ;
  assign n10140 = n10139 ^ n3150 ^ n2106 ;
  assign n10136 = ~n430 & n6877 ;
  assign n10137 = ~n1745 & n10136 ;
  assign n10141 = n10140 ^ n10137 ^ 1'b0 ;
  assign n10142 = ~n5115 & n10141 ;
  assign n10143 = ~n624 & n10142 ;
  assign n10144 = n10143 ^ n3854 ^ 1'b0 ;
  assign n10129 = n10072 ^ n2617 ^ x67 ;
  assign n10130 = ( n3368 & ~n3777 ) | ( n3368 & n10129 ) | ( ~n3777 & n10129 ) ;
  assign n10131 = n744 & ~n10130 ;
  assign n10132 = n10131 ^ n5211 ^ 1'b0 ;
  assign n10133 = ( n2127 & n8994 ) | ( n2127 & n10132 ) | ( n8994 & n10132 ) ;
  assign n10134 = ( n1832 & n5787 ) | ( n1832 & n10133 ) | ( n5787 & n10133 ) ;
  assign n10135 = n10134 ^ n1818 ^ 1'b0 ;
  assign n10145 = n10144 ^ n10135 ^ 1'b0 ;
  assign n10146 = n6992 & ~n10145 ;
  assign n10149 = n1516 | n1926 ;
  assign n10150 = n10149 ^ n4110 ^ 1'b0 ;
  assign n10147 = n7984 ^ n4507 ^ 1'b0 ;
  assign n10148 = n433 & n10147 ;
  assign n10151 = n10150 ^ n10148 ^ n5461 ;
  assign n10152 = ( n548 & n4578 ) | ( n548 & n7123 ) | ( n4578 & n7123 ) ;
  assign n10153 = n3837 & n10152 ;
  assign n10154 = n10153 ^ n4962 ^ 1'b0 ;
  assign n10155 = n7343 ^ n5329 ^ n4190 ;
  assign n10156 = n10155 ^ n5008 ^ n4581 ;
  assign n10157 = n10156 ^ n3904 ^ n3731 ;
  assign n10158 = n10154 | n10157 ;
  assign n10159 = n8566 & ~n10158 ;
  assign n10160 = n6613 ^ n645 ^ 1'b0 ;
  assign n10161 = n3086 & n10160 ;
  assign n10162 = n10161 ^ n1596 ^ x206 ;
  assign n10163 = n6481 ^ n5592 ^ n2252 ;
  assign n10164 = n6292 ^ n5955 ^ n2905 ;
  assign n10165 = ( n5056 & ~n10163 ) | ( n5056 & n10164 ) | ( ~n10163 & n10164 ) ;
  assign n10166 = n6241 ^ n3841 ^ 1'b0 ;
  assign n10167 = ~n3268 & n10166 ;
  assign n10168 = n9639 ^ n2843 ^ 1'b0 ;
  assign n10169 = n5804 & n10168 ;
  assign n10170 = n10169 ^ n8701 ^ 1'b0 ;
  assign n10171 = ( n1267 & n10167 ) | ( n1267 & ~n10170 ) | ( n10167 & ~n10170 ) ;
  assign n10172 = ~n894 & n9185 ;
  assign n10173 = x96 & ~n5370 ;
  assign n10174 = ( ~n631 & n4507 ) | ( ~n631 & n6935 ) | ( n4507 & n6935 ) ;
  assign n10175 = n10174 ^ n6097 ^ n5008 ;
  assign n10176 = n10089 ^ n9763 ^ 1'b0 ;
  assign n10177 = ~n2043 & n6143 ;
  assign n10178 = n4331 & n10177 ;
  assign n10179 = n3812 ^ n1918 ^ 1'b0 ;
  assign n10180 = n10179 ^ n5387 ^ 1'b0 ;
  assign n10181 = n10180 ^ n9298 ^ 1'b0 ;
  assign n10182 = n10178 | n10181 ;
  assign n10183 = n987 | n5424 ;
  assign n10184 = n10183 ^ n4475 ^ 1'b0 ;
  assign n10185 = n5242 ^ n4654 ^ n3495 ;
  assign n10186 = ( n2476 & n6937 ) | ( n2476 & ~n10185 ) | ( n6937 & ~n10185 ) ;
  assign n10187 = ( ~n3868 & n10184 ) | ( ~n3868 & n10186 ) | ( n10184 & n10186 ) ;
  assign n10188 = n10187 ^ n1296 ^ 1'b0 ;
  assign n10189 = ( ~n8922 & n8947 ) | ( ~n8922 & n10040 ) | ( n8947 & n10040 ) ;
  assign n10190 = n3299 | n8705 ;
  assign n10191 = n10190 ^ n2662 ^ 1'b0 ;
  assign n10192 = n7650 ^ n755 ^ 1'b0 ;
  assign n10197 = n9069 ^ n6867 ^ x7 ;
  assign n10198 = n4664 | n10197 ;
  assign n10199 = n10198 ^ n1256 ^ 1'b0 ;
  assign n10193 = ~n2243 & n4049 ;
  assign n10194 = n10193 ^ n6657 ^ 1'b0 ;
  assign n10195 = ~n8833 & n10194 ;
  assign n10196 = n368 & n10195 ;
  assign n10200 = n10199 ^ n10196 ^ 1'b0 ;
  assign n10201 = n2395 & n6601 ;
  assign n10202 = n10201 ^ n9238 ^ n8160 ;
  assign n10203 = n10202 ^ n7301 ^ 1'b0 ;
  assign n10204 = n7834 & ~n10203 ;
  assign n10210 = ~n2545 & n2793 ;
  assign n10211 = ~n1029 & n10210 ;
  assign n10212 = n10211 ^ n2137 ^ n604 ;
  assign n10213 = n2815 & n9294 ;
  assign n10214 = n5874 ^ n1960 ^ 1'b0 ;
  assign n10215 = n10213 & n10214 ;
  assign n10216 = ( n6470 & ~n10212 ) | ( n6470 & n10215 ) | ( ~n10212 & n10215 ) ;
  assign n10217 = ~n4012 & n10216 ;
  assign n10218 = n7225 & ~n10217 ;
  assign n10219 = n7321 ^ n494 ^ n289 ;
  assign n10220 = n5686 & n10219 ;
  assign n10221 = n6877 ^ n3260 ^ 1'b0 ;
  assign n10222 = ~n10220 & n10221 ;
  assign n10223 = n10222 ^ n5016 ^ n1848 ;
  assign n10224 = ( n9651 & n10218 ) | ( n9651 & n10223 ) | ( n10218 & n10223 ) ;
  assign n10205 = n3144 & n4679 ;
  assign n10206 = n10205 ^ n4166 ^ 1'b0 ;
  assign n10207 = x191 & x218 ;
  assign n10208 = n10207 ^ n8747 ^ 1'b0 ;
  assign n10209 = ~n10206 & n10208 ;
  assign n10225 = n10224 ^ n10209 ^ 1'b0 ;
  assign n10228 = n5398 ^ n3216 ^ n2465 ;
  assign n10226 = n8014 ^ n4224 ^ n1467 ;
  assign n10227 = n10226 ^ n1947 ^ n1433 ;
  assign n10229 = n10228 ^ n10227 ^ n444 ;
  assign n10230 = n10229 ^ n7330 ^ n2758 ;
  assign n10231 = ( ~n3754 & n9608 ) | ( ~n3754 & n10230 ) | ( n9608 & n10230 ) ;
  assign n10232 = n9321 ^ n8067 ^ n5525 ;
  assign n10233 = n10232 ^ n7903 ^ n5467 ;
  assign n10234 = ( n3490 & ~n4067 ) | ( n3490 & n6092 ) | ( ~n4067 & n6092 ) ;
  assign n10241 = ( n2006 & n2643 ) | ( n2006 & ~n2905 ) | ( n2643 & ~n2905 ) ;
  assign n10236 = n897 ^ n575 ^ x15 ;
  assign n10237 = n3780 & n10236 ;
  assign n10238 = ~n3600 & n10237 ;
  assign n10239 = ( ~n2216 & n6037 ) | ( ~n2216 & n10238 ) | ( n6037 & n10238 ) ;
  assign n10235 = n942 | n1421 ;
  assign n10240 = n10239 ^ n10235 ^ n866 ;
  assign n10242 = n10241 ^ n10240 ^ n9473 ;
  assign n10243 = n10242 ^ n8557 ^ 1'b0 ;
  assign n10244 = n8571 ^ n295 ^ 1'b0 ;
  assign n10245 = n10243 & n10244 ;
  assign n10246 = n10245 ^ n3311 ^ 1'b0 ;
  assign n10249 = ( n1998 & n4531 ) | ( n1998 & ~n5242 ) | ( n4531 & ~n5242 ) ;
  assign n10250 = n4179 & ~n10249 ;
  assign n10247 = ( n1455 & n6409 ) | ( n1455 & n7437 ) | ( n6409 & n7437 ) ;
  assign n10248 = ( ~n6413 & n8961 ) | ( ~n6413 & n10247 ) | ( n8961 & n10247 ) ;
  assign n10251 = n10250 ^ n10248 ^ n863 ;
  assign n10254 = n9589 ^ n2676 ^ 1'b0 ;
  assign n10255 = n473 | n10254 ;
  assign n10252 = n8692 ^ n5928 ^ 1'b0 ;
  assign n10253 = ~n3591 & n10252 ;
  assign n10256 = n10255 ^ n10253 ^ n874 ;
  assign n10257 = n9237 ^ n6069 ^ 1'b0 ;
  assign n10258 = n3720 | n7987 ;
  assign n10259 = n10258 ^ n5619 ^ 1'b0 ;
  assign n10260 = n10259 ^ n8915 ^ n5843 ;
  assign n10261 = n2247 & ~n10260 ;
  assign n10262 = n10257 & n10261 ;
  assign n10264 = ( x107 & n3438 ) | ( x107 & n7062 ) | ( n3438 & n7062 ) ;
  assign n10265 = ~n8994 & n10264 ;
  assign n10263 = ( n1914 & n2034 ) | ( n1914 & n6164 ) | ( n2034 & n6164 ) ;
  assign n10266 = n10265 ^ n10263 ^ n4514 ;
  assign n10267 = n311 | n6781 ;
  assign n10268 = ( n3676 & n9346 ) | ( n3676 & ~n10267 ) | ( n9346 & ~n10267 ) ;
  assign n10269 = n10084 ^ n3629 ^ 1'b0 ;
  assign n10270 = ~n10268 & n10269 ;
  assign n10271 = n4701 & n5565 ;
  assign n10272 = n8115 ^ n6869 ^ n5709 ;
  assign n10273 = n4101 | n7251 ;
  assign n10274 = n10273 ^ n2308 ^ 1'b0 ;
  assign n10275 = n9390 ^ n9226 ^ 1'b0 ;
  assign n10276 = n10274 | n10275 ;
  assign n10277 = n9747 | n10276 ;
  assign n10278 = n3018 | n4925 ;
  assign n10279 = n10278 ^ n687 ^ 1'b0 ;
  assign n10280 = n10279 ^ n7784 ^ n1408 ;
  assign n10281 = n7905 & ~n10280 ;
  assign n10282 = ~n433 & n10281 ;
  assign n10283 = n10282 ^ n7652 ^ n4899 ;
  assign n10284 = n1700 ^ n1526 ^ 1'b0 ;
  assign n10285 = n3154 | n10284 ;
  assign n10286 = n353 & n938 ;
  assign n10287 = n10286 ^ n3787 ^ 1'b0 ;
  assign n10288 = n8641 | n10287 ;
  assign n10289 = n10288 ^ n4264 ^ 1'b0 ;
  assign n10290 = x189 & n10289 ;
  assign n10291 = ~n2089 & n10290 ;
  assign n10292 = n5018 ^ n2292 ^ n1475 ;
  assign n10293 = n10291 | n10292 ;
  assign n10294 = n5129 ^ n2800 ^ 1'b0 ;
  assign n10295 = n732 & ~n8714 ;
  assign n10296 = n10294 & n10295 ;
  assign n10297 = n4363 ^ x212 ^ 1'b0 ;
  assign n10298 = n1836 & ~n10297 ;
  assign n10299 = ~n10296 & n10298 ;
  assign n10300 = n10299 ^ n5473 ^ 1'b0 ;
  assign n10301 = n2794 & ~n10300 ;
  assign n10302 = n10293 & n10301 ;
  assign n10309 = ( n3151 & n4190 ) | ( n3151 & n5292 ) | ( n4190 & n5292 ) ;
  assign n10310 = n10309 ^ n7244 ^ 1'b0 ;
  assign n10303 = n647 ^ n291 ^ 1'b0 ;
  assign n10306 = n5199 ^ n1499 ^ n738 ;
  assign n10304 = n3787 ^ n2075 ^ 1'b0 ;
  assign n10305 = ~n4906 & n10304 ;
  assign n10307 = n10306 ^ n10305 ^ n2950 ;
  assign n10308 = n10303 & n10307 ;
  assign n10311 = n10310 ^ n10308 ^ n1136 ;
  assign n10312 = n2568 ^ n1809 ^ n1283 ;
  assign n10313 = n10312 ^ n921 ^ 1'b0 ;
  assign n10314 = n1302 & n10313 ;
  assign n10315 = n10314 ^ n6267 ^ n2953 ;
  assign n10316 = n4668 ^ n4331 ^ n631 ;
  assign n10317 = ( n2810 & n8164 ) | ( n2810 & n10316 ) | ( n8164 & n10316 ) ;
  assign n10324 = ~n431 & n4032 ;
  assign n10325 = n10324 ^ n3071 ^ 1'b0 ;
  assign n10318 = ( ~n1678 & n5305 ) | ( ~n1678 & n8424 ) | ( n5305 & n8424 ) ;
  assign n10319 = n5979 ^ n2993 ^ n1661 ;
  assign n10320 = n600 & ~n10319 ;
  assign n10321 = n5193 & n10320 ;
  assign n10322 = n2220 & n10321 ;
  assign n10323 = n10318 & ~n10322 ;
  assign n10326 = n10325 ^ n10323 ^ 1'b0 ;
  assign n10327 = n10326 ^ n9997 ^ n3842 ;
  assign n10328 = n6621 ^ n2884 ^ n1502 ;
  assign n10329 = ( n10317 & ~n10327 ) | ( n10317 & n10328 ) | ( ~n10327 & n10328 ) ;
  assign n10330 = n10329 ^ n10139 ^ n6206 ;
  assign n10331 = n5391 ^ n2514 ^ n1139 ;
  assign n10332 = ~n8535 & n10331 ;
  assign n10340 = n9177 | n10238 ;
  assign n10341 = n5398 & ~n10340 ;
  assign n10333 = ( n2089 & n2606 ) | ( n2089 & n2923 ) | ( n2606 & n2923 ) ;
  assign n10335 = n3235 ^ n873 ^ 1'b0 ;
  assign n10334 = ( n1118 & n2369 ) | ( n1118 & ~n2631 ) | ( n2369 & ~n2631 ) ;
  assign n10336 = n10335 ^ n10334 ^ n916 ;
  assign n10337 = n10333 & ~n10336 ;
  assign n10338 = n4537 & n10337 ;
  assign n10339 = n10338 ^ n6157 ^ n5246 ;
  assign n10342 = n10341 ^ n10339 ^ n5045 ;
  assign n10345 = n3962 | n8133 ;
  assign n10346 = n10345 ^ n9485 ^ n3740 ;
  assign n10343 = n8474 ^ n7670 ^ n1098 ;
  assign n10344 = n10343 ^ n9020 ^ n8408 ;
  assign n10347 = n10346 ^ n10344 ^ n1351 ;
  assign n10350 = n5628 ^ n622 ^ 1'b0 ;
  assign n10351 = n2788 | n10350 ;
  assign n10348 = ( n1466 & n2120 ) | ( n1466 & ~n6488 ) | ( n2120 & ~n6488 ) ;
  assign n10349 = n10348 ^ n6113 ^ n3693 ;
  assign n10352 = n10351 ^ n10349 ^ 1'b0 ;
  assign n10353 = ~n6887 & n10352 ;
  assign n10355 = n6943 ^ n699 ^ 1'b0 ;
  assign n10356 = ~n6329 & n10355 ;
  assign n10357 = n8406 & n10356 ;
  assign n10358 = n3245 & n10357 ;
  assign n10354 = n890 | n6550 ;
  assign n10359 = n10358 ^ n10354 ^ n7491 ;
  assign n10360 = n861 & n2826 ;
  assign n10361 = n9392 ^ n6743 ^ 1'b0 ;
  assign n10362 = x210 & n10361 ;
  assign n10363 = n10362 ^ n4954 ^ 1'b0 ;
  assign n10364 = n7355 ^ n2683 ^ 1'b0 ;
  assign n10365 = n10364 ^ n1567 ^ 1'b0 ;
  assign n10366 = n3322 & ~n10365 ;
  assign n10367 = ~n5939 & n9072 ;
  assign n10368 = n948 | n10367 ;
  assign n10369 = n2516 ^ n2081 ^ 1'b0 ;
  assign n10370 = n10369 ^ n6839 ^ n6021 ;
  assign n10371 = n8834 ^ n8766 ^ n2654 ;
  assign n10372 = ( ~n1209 & n3715 ) | ( ~n1209 & n10371 ) | ( n3715 & n10371 ) ;
  assign n10373 = n10372 ^ n1529 ^ 1'b0 ;
  assign n10374 = ( ~n5851 & n9758 ) | ( ~n5851 & n10373 ) | ( n9758 & n10373 ) ;
  assign n10375 = ( n8869 & n10370 ) | ( n8869 & ~n10374 ) | ( n10370 & ~n10374 ) ;
  assign n10376 = n1586 | n4551 ;
  assign n10377 = n10376 ^ n1354 ^ 1'b0 ;
  assign n10378 = n9462 ^ n894 ^ 1'b0 ;
  assign n10379 = ( n6964 & ~n10377 ) | ( n6964 & n10378 ) | ( ~n10377 & n10378 ) ;
  assign n10380 = n9863 ^ n1106 ^ 1'b0 ;
  assign n10382 = ~n715 & n7497 ;
  assign n10383 = n1457 & n10382 ;
  assign n10384 = n10383 ^ n8909 ^ n4068 ;
  assign n10381 = n6567 ^ x199 ^ 1'b0 ;
  assign n10385 = n10384 ^ n10381 ^ 1'b0 ;
  assign n10386 = ~n10380 & n10385 ;
  assign n10387 = ( n1990 & n4852 ) | ( n1990 & n6331 ) | ( n4852 & n6331 ) ;
  assign n10388 = n10387 ^ n5992 ^ n5414 ;
  assign n10389 = ( n853 & n2182 ) | ( n853 & ~n2247 ) | ( n2182 & ~n2247 ) ;
  assign n10390 = ( ~n393 & n5766 ) | ( ~n393 & n10389 ) | ( n5766 & n10389 ) ;
  assign n10391 = n1027 | n5246 ;
  assign n10392 = n10391 ^ n6704 ^ 1'b0 ;
  assign n10393 = ( n8267 & ~n10390 ) | ( n8267 & n10392 ) | ( ~n10390 & n10392 ) ;
  assign n10398 = ( ~x47 & n1983 ) | ( ~x47 & n6270 ) | ( n1983 & n6270 ) ;
  assign n10397 = n5322 ^ n1542 ^ n777 ;
  assign n10399 = n10398 ^ n10397 ^ 1'b0 ;
  assign n10394 = n3305 & n5506 ;
  assign n10395 = ( n1038 & ~n1343 ) | ( n1038 & n7216 ) | ( ~n1343 & n7216 ) ;
  assign n10396 = ~n10394 & n10395 ;
  assign n10400 = n10399 ^ n10396 ^ 1'b0 ;
  assign n10401 = n3131 & n4159 ;
  assign n10402 = n10023 | n10401 ;
  assign n10404 = ( ~n599 & n3227 ) | ( ~n599 & n3484 ) | ( n3227 & n3484 ) ;
  assign n10405 = n10404 ^ n8277 ^ n2576 ;
  assign n10406 = n10405 ^ n5852 ^ 1'b0 ;
  assign n10407 = n7601 | n10406 ;
  assign n10408 = n2897 | n10407 ;
  assign n10409 = n9462 | n10408 ;
  assign n10403 = n3363 ^ n3316 ^ n2188 ;
  assign n10410 = n10409 ^ n10403 ^ n1751 ;
  assign n10413 = n1467 ^ n298 ^ 1'b0 ;
  assign n10414 = n3569 & n10413 ;
  assign n10411 = ( n4084 & n4475 ) | ( n4084 & ~n9198 ) | ( n4475 & ~n9198 ) ;
  assign n10412 = n10411 ^ n2282 ^ n340 ;
  assign n10415 = n10414 ^ n10412 ^ 1'b0 ;
  assign n10416 = ( n5517 & ~n10410 ) | ( n5517 & n10415 ) | ( ~n10410 & n10415 ) ;
  assign n10418 = n1893 ^ n1385 ^ n617 ;
  assign n10419 = ( n1769 & ~n2254 ) | ( n1769 & n10418 ) | ( ~n2254 & n10418 ) ;
  assign n10420 = n2719 ^ n1794 ^ n1502 ;
  assign n10421 = n10420 ^ n1416 ^ 1'b0 ;
  assign n10422 = ( n6236 & ~n10419 ) | ( n6236 & n10421 ) | ( ~n10419 & n10421 ) ;
  assign n10417 = ~n1019 & n5400 ;
  assign n10423 = n10422 ^ n10417 ^ 1'b0 ;
  assign n10424 = n3847 ^ n2875 ^ 1'b0 ;
  assign n10425 = n7642 ^ n3088 ^ 1'b0 ;
  assign n10426 = n4197 ^ n755 ^ 1'b0 ;
  assign n10427 = n10426 ^ n2393 ^ 1'b0 ;
  assign n10428 = n6797 & ~n10427 ;
  assign n10431 = ( n484 & ~n2313 ) | ( n484 & n3945 ) | ( ~n2313 & n3945 ) ;
  assign n10432 = n10431 ^ n1119 ^ n366 ;
  assign n10429 = ( n1755 & n4831 ) | ( n1755 & ~n6947 ) | ( n4831 & ~n6947 ) ;
  assign n10430 = n10429 ^ n6552 ^ n861 ;
  assign n10433 = n10432 ^ n10430 ^ n8922 ;
  assign n10434 = n4341 & n6048 ;
  assign n10435 = ( n10148 & n10433 ) | ( n10148 & n10434 ) | ( n10433 & n10434 ) ;
  assign n10436 = n7015 ^ n5237 ^ n2732 ;
  assign n10437 = n8641 ^ n5280 ^ 1'b0 ;
  assign n10438 = x99 & ~n10437 ;
  assign n10451 = n5447 ^ n3125 ^ 1'b0 ;
  assign n10452 = n3697 | n10451 ;
  assign n10441 = n5947 ^ n4822 ^ n2150 ;
  assign n10442 = ( n311 & n3701 ) | ( n311 & ~n10441 ) | ( n3701 & ~n10441 ) ;
  assign n10439 = ~n1323 & n2024 ;
  assign n10440 = n5656 & ~n10439 ;
  assign n10443 = n10442 ^ n10440 ^ 1'b0 ;
  assign n10445 = n3824 ^ n3710 ^ 1'b0 ;
  assign n10446 = n1616 & ~n10445 ;
  assign n10447 = ( n1950 & ~n3500 ) | ( n1950 & n10446 ) | ( ~n3500 & n10446 ) ;
  assign n10444 = n5072 | n5789 ;
  assign n10448 = n10447 ^ n10444 ^ 1'b0 ;
  assign n10449 = ( n2099 & ~n10443 ) | ( n2099 & n10448 ) | ( ~n10443 & n10448 ) ;
  assign n10450 = n7419 & n10449 ;
  assign n10453 = n10452 ^ n10450 ^ 1'b0 ;
  assign n10454 = ( n3155 & ~n5627 ) | ( n3155 & n9931 ) | ( ~n5627 & n9931 ) ;
  assign n10455 = ( n5219 & n5231 ) | ( n5219 & n10454 ) | ( n5231 & n10454 ) ;
  assign n10456 = n6110 | n7597 ;
  assign n10459 = ( n3067 & ~n3435 ) | ( n3067 & n5749 ) | ( ~n3435 & n5749 ) ;
  assign n10460 = n10459 ^ n6946 ^ n5289 ;
  assign n10457 = n1653 & ~n4001 ;
  assign n10458 = ( n3021 & n5566 ) | ( n3021 & ~n10457 ) | ( n5566 & ~n10457 ) ;
  assign n10461 = n10460 ^ n10458 ^ x15 ;
  assign n10462 = ( ~n2839 & n5509 ) | ( ~n2839 & n8889 ) | ( n5509 & n8889 ) ;
  assign n10463 = n10462 ^ n8562 ^ 1'b0 ;
  assign n10464 = n10461 & ~n10463 ;
  assign n10466 = n5358 ^ n2871 ^ n885 ;
  assign n10467 = n10466 ^ n3132 ^ n1592 ;
  assign n10465 = ( n3229 & n4192 ) | ( n3229 & ~n6457 ) | ( n4192 & ~n6457 ) ;
  assign n10468 = n10467 ^ n10465 ^ n9219 ;
  assign n10469 = ~n820 & n5286 ;
  assign n10470 = ~n9447 & n10059 ;
  assign n10471 = n10470 ^ n4348 ^ 1'b0 ;
  assign n10472 = n2617 & ~n10471 ;
  assign n10473 = n10472 ^ n6952 ^ 1'b0 ;
  assign n10474 = ~n1440 & n10473 ;
  assign n10478 = n2281 & ~n4599 ;
  assign n10476 = n6749 ^ n4126 ^ n950 ;
  assign n10475 = n520 | n8273 ;
  assign n10477 = n10476 ^ n10475 ^ 1'b0 ;
  assign n10479 = n10478 ^ n10477 ^ n10174 ;
  assign n10480 = n9982 ^ n4970 ^ 1'b0 ;
  assign n10481 = n5398 | n10480 ;
  assign n10482 = n10481 ^ n4485 ^ 1'b0 ;
  assign n10483 = ~n9294 & n10482 ;
  assign n10484 = n5096 & ~n10023 ;
  assign n10485 = ~n8146 & n10484 ;
  assign n10486 = n773 & n2319 ;
  assign n10487 = n5636 ^ n1042 ^ n268 ;
  assign n10488 = n10487 ^ n8378 ^ n8175 ;
  assign n10489 = ~n3119 & n10488 ;
  assign n10490 = n10486 & n10489 ;
  assign n10494 = n6305 | n6370 ;
  assign n10495 = n6114 | n10494 ;
  assign n10491 = ~n5221 & n6575 ;
  assign n10492 = n10491 ^ n2129 ^ 1'b0 ;
  assign n10493 = ( n1047 & n3286 ) | ( n1047 & ~n10492 ) | ( n3286 & ~n10492 ) ;
  assign n10496 = n10495 ^ n10493 ^ 1'b0 ;
  assign n10497 = n2482 & n10496 ;
  assign n10498 = n10497 ^ n2028 ^ x198 ;
  assign n10499 = ( n8917 & n10490 ) | ( n8917 & ~n10498 ) | ( n10490 & ~n10498 ) ;
  assign n10500 = n7844 ^ n6298 ^ n2955 ;
  assign n10501 = n10500 ^ n6983 ^ n5858 ;
  assign n10502 = n10501 ^ n3126 ^ n1586 ;
  assign n10507 = n6017 ^ n3294 ^ 1'b0 ;
  assign n10503 = n5723 ^ n2848 ^ n2770 ;
  assign n10504 = n10503 ^ n1461 ^ 1'b0 ;
  assign n10505 = n5404 | n10504 ;
  assign n10506 = n10505 ^ n10466 ^ 1'b0 ;
  assign n10508 = n10507 ^ n10506 ^ 1'b0 ;
  assign n10515 = n1241 & ~n4273 ;
  assign n10516 = ~n1164 & n10515 ;
  assign n10510 = n6711 ^ n759 ^ 1'b0 ;
  assign n10511 = ~n8550 & n10510 ;
  assign n10512 = n2184 | n7390 ;
  assign n10513 = n10511 | n10512 ;
  assign n10514 = n10513 ^ n10467 ^ 1'b0 ;
  assign n10509 = ~n3430 & n7098 ;
  assign n10517 = n10516 ^ n10514 ^ n10509 ;
  assign n10518 = n10517 ^ n8569 ^ 1'b0 ;
  assign n10519 = n6389 | n10518 ;
  assign n10520 = ( ~n2366 & n4536 ) | ( ~n2366 & n6578 ) | ( n4536 & n6578 ) ;
  assign n10521 = n9888 ^ n5434 ^ n4661 ;
  assign n10522 = n6806 ^ n3641 ^ 1'b0 ;
  assign n10523 = n3766 & ~n10522 ;
  assign n10524 = n7089 & ~n8635 ;
  assign n10525 = ~n10523 & n10524 ;
  assign n10526 = n5849 ^ n5153 ^ n4309 ;
  assign n10527 = ( n10521 & n10525 ) | ( n10521 & n10526 ) | ( n10525 & n10526 ) ;
  assign n10528 = ~n813 & n9293 ;
  assign n10529 = n4451 & n5260 ;
  assign n10530 = x8 & ~n4003 ;
  assign n10531 = n10530 ^ n4436 ^ n4331 ;
  assign n10532 = n10531 ^ n5681 ^ n3585 ;
  assign n10533 = n5351 ^ n2720 ^ n289 ;
  assign n10534 = ( n2020 & n4357 ) | ( n2020 & n10533 ) | ( n4357 & n10533 ) ;
  assign n10535 = n583 & ~n10534 ;
  assign n10536 = ~n738 & n10535 ;
  assign n10537 = x248 & n700 ;
  assign n10538 = n10537 ^ n2321 ^ 1'b0 ;
  assign n10540 = n6409 ^ n5628 ^ 1'b0 ;
  assign n10539 = n2677 | n5536 ;
  assign n10541 = n10540 ^ n10539 ^ 1'b0 ;
  assign n10542 = ( n3853 & ~n10538 ) | ( n3853 & n10541 ) | ( ~n10538 & n10541 ) ;
  assign n10543 = n778 | n1386 ;
  assign n10544 = x220 & n2988 ;
  assign n10545 = n10544 ^ n1312 ^ 1'b0 ;
  assign n10546 = n10545 ^ n10156 ^ n8806 ;
  assign n10547 = ( ~n2756 & n5498 ) | ( ~n2756 & n9651 ) | ( n5498 & n9651 ) ;
  assign n10548 = ( n1887 & ~n5188 ) | ( n1887 & n10547 ) | ( ~n5188 & n10547 ) ;
  assign n10549 = n6710 ^ n2973 ^ x3 ;
  assign n10550 = x227 | n5248 ;
  assign n10551 = n6373 ^ n2033 ^ 1'b0 ;
  assign n10552 = x36 & ~n10551 ;
  assign n10553 = ( n4598 & n10550 ) | ( n4598 & ~n10552 ) | ( n10550 & ~n10552 ) ;
  assign n10554 = ( n8927 & n10549 ) | ( n8927 & ~n10553 ) | ( n10549 & ~n10553 ) ;
  assign n10555 = n3416 ^ n1482 ^ n1412 ;
  assign n10556 = n6552 ^ n1565 ^ n1070 ;
  assign n10563 = ~n736 & n5454 ;
  assign n10564 = n5300 & n10563 ;
  assign n10565 = ( n755 & n7362 ) | ( n755 & ~n10564 ) | ( n7362 & ~n10564 ) ;
  assign n10562 = ( ~n5185 & n6389 ) | ( ~n5185 & n8195 ) | ( n6389 & n8195 ) ;
  assign n10557 = ( n944 & ~n3379 ) | ( n944 & n7763 ) | ( ~n3379 & n7763 ) ;
  assign n10558 = n7313 ^ n6176 ^ 1'b0 ;
  assign n10559 = n10557 & n10558 ;
  assign n10560 = n10559 ^ n8174 ^ n7173 ;
  assign n10561 = n10560 ^ n10314 ^ n6731 ;
  assign n10566 = n10565 ^ n10562 ^ n10561 ;
  assign n10573 = ( n1897 & ~n2158 ) | ( n1897 & n10072 ) | ( ~n2158 & n10072 ) ;
  assign n10574 = n10573 ^ n3096 ^ n1147 ;
  assign n10572 = ( n476 & ~n716 ) | ( n476 & n6617 ) | ( ~n716 & n6617 ) ;
  assign n10567 = n1293 | n4422 ;
  assign n10568 = n8621 & ~n10567 ;
  assign n10569 = n3126 & n6726 ;
  assign n10570 = ( n7448 & n10568 ) | ( n7448 & n10569 ) | ( n10568 & n10569 ) ;
  assign n10571 = n10570 ^ n5990 ^ n2414 ;
  assign n10575 = n10574 ^ n10572 ^ n10571 ;
  assign n10577 = ~n7802 & n8582 ;
  assign n10576 = n3545 & n5444 ;
  assign n10578 = n10577 ^ n10576 ^ 1'b0 ;
  assign n10579 = n10578 ^ n7253 ^ 1'b0 ;
  assign n10580 = n4704 & n10579 ;
  assign n10581 = n1924 & n4678 ;
  assign n10582 = ( n3065 & n4499 ) | ( n3065 & n9150 ) | ( n4499 & n9150 ) ;
  assign n10583 = ( n1192 & n1983 ) | ( n1192 & ~n6352 ) | ( n1983 & ~n6352 ) ;
  assign n10584 = ( n4496 & ~n9462 ) | ( n4496 & n10583 ) | ( ~n9462 & n10583 ) ;
  assign n10585 = ( n5459 & ~n10582 ) | ( n5459 & n10584 ) | ( ~n10582 & n10584 ) ;
  assign n10586 = n4015 ^ n1808 ^ n1312 ;
  assign n10587 = n6823 ^ n2436 ^ n876 ;
  assign n10588 = n1287 | n3596 ;
  assign n10589 = n10588 ^ n723 ^ 1'b0 ;
  assign n10590 = ( n5085 & n10587 ) | ( n5085 & n10589 ) | ( n10587 & n10589 ) ;
  assign n10591 = ~n8644 & n10590 ;
  assign n10592 = n5440 ^ n5093 ^ 1'b0 ;
  assign n10593 = n6659 ^ n4888 ^ 1'b0 ;
  assign n10594 = n10593 ^ n5598 ^ 1'b0 ;
  assign n10595 = ( ~n6116 & n8270 ) | ( ~n6116 & n10594 ) | ( n8270 & n10594 ) ;
  assign n10596 = n9387 ^ n8099 ^ 1'b0 ;
  assign n10597 = ( n4067 & ~n6739 ) | ( n4067 & n10596 ) | ( ~n6739 & n10596 ) ;
  assign n10598 = n835 | n10597 ;
  assign n10599 = n10598 ^ n4292 ^ n4229 ;
  assign n10600 = ~n3986 & n6745 ;
  assign n10601 = n951 | n3517 ;
  assign n10602 = ( ~n7904 & n9858 ) | ( ~n7904 & n10601 ) | ( n9858 & n10601 ) ;
  assign n10603 = ( n4457 & n10600 ) | ( n4457 & ~n10602 ) | ( n10600 & ~n10602 ) ;
  assign n10604 = ( n1860 & ~n4554 ) | ( n1860 & n6838 ) | ( ~n4554 & n6838 ) ;
  assign n10605 = n282 & n4023 ;
  assign n10606 = ( n452 & ~n2887 ) | ( n452 & n10605 ) | ( ~n2887 & n10605 ) ;
  assign n10607 = ( n8939 & ~n10604 ) | ( n8939 & n10606 ) | ( ~n10604 & n10606 ) ;
  assign n10608 = n2059 ^ n640 ^ 1'b0 ;
  assign n10609 = ~n5307 & n10608 ;
  assign n10610 = n1244 & n2750 ;
  assign n10611 = ~n6270 & n10610 ;
  assign n10612 = ( n710 & n9395 ) | ( n710 & n10611 ) | ( n9395 & n10611 ) ;
  assign n10613 = ( n6590 & n10609 ) | ( n6590 & n10612 ) | ( n10609 & n10612 ) ;
  assign n10616 = ~n400 & n2981 ;
  assign n10617 = ~n6383 & n10616 ;
  assign n10618 = n5089 & n7110 ;
  assign n10619 = ( n1701 & n10617 ) | ( n1701 & n10618 ) | ( n10617 & n10618 ) ;
  assign n10614 = n9122 ^ n2029 ^ 1'b0 ;
  assign n10615 = n5328 | n10614 ;
  assign n10620 = n10619 ^ n10615 ^ n1118 ;
  assign n10635 = n3745 & ~n5190 ;
  assign n10621 = n3966 ^ n1165 ^ 1'b0 ;
  assign n10622 = n3608 | n10621 ;
  assign n10623 = ~n1486 & n2750 ;
  assign n10624 = n10622 & n10623 ;
  assign n10625 = n6346 & ~n10100 ;
  assign n10626 = n1117 & n10625 ;
  assign n10627 = n10626 ^ n2120 ^ 1'b0 ;
  assign n10628 = n10627 ^ n5072 ^ n1134 ;
  assign n10629 = n5050 | n10628 ;
  assign n10630 = n6998 | n10629 ;
  assign n10631 = n10630 ^ n9160 ^ n7540 ;
  assign n10632 = n3198 | n10631 ;
  assign n10633 = n10632 ^ n7700 ^ 1'b0 ;
  assign n10634 = n10624 | n10633 ;
  assign n10636 = n10635 ^ n10634 ^ n8799 ;
  assign n10637 = ~n2428 & n3042 ;
  assign n10638 = n10637 ^ n340 ^ 1'b0 ;
  assign n10639 = n10638 ^ n6796 ^ n837 ;
  assign n10640 = ( ~n566 & n8167 ) | ( ~n566 & n10639 ) | ( n8167 & n10639 ) ;
  assign n10653 = n1679 & n5498 ;
  assign n10654 = n6834 & n10653 ;
  assign n10649 = x181 | n2926 ;
  assign n10650 = n1716 ^ n736 ^ 1'b0 ;
  assign n10651 = ( ~n3628 & n10649 ) | ( ~n3628 & n10650 ) | ( n10649 & n10650 ) ;
  assign n10643 = n8736 ^ n5798 ^ n1962 ;
  assign n10644 = ( n3264 & n3524 ) | ( n3264 & ~n9800 ) | ( n3524 & ~n9800 ) ;
  assign n10645 = ( n4926 & ~n10643 ) | ( n4926 & n10644 ) | ( ~n10643 & n10644 ) ;
  assign n10646 = n5638 ^ n4819 ^ 1'b0 ;
  assign n10647 = n10316 & ~n10646 ;
  assign n10648 = ~n10645 & n10647 ;
  assign n10652 = n10651 ^ n10648 ^ 1'b0 ;
  assign n10641 = n5141 ^ n2353 ^ n424 ;
  assign n10642 = n10641 ^ n10294 ^ n1047 ;
  assign n10655 = n10654 ^ n10652 ^ n10642 ;
  assign n10661 = n3326 & ~n8430 ;
  assign n10659 = n4035 ^ n2635 ^ n344 ;
  assign n10660 = n10659 ^ n2289 ^ n1465 ;
  assign n10656 = ( n5037 & ~n5813 ) | ( n5037 & n6076 ) | ( ~n5813 & n6076 ) ;
  assign n10657 = n2237 | n10656 ;
  assign n10658 = n10657 ^ n9902 ^ n5060 ;
  assign n10662 = n10661 ^ n10660 ^ n10658 ;
  assign n10667 = n10100 ^ n3729 ^ n975 ;
  assign n10665 = n4134 & n6827 ;
  assign n10663 = ( n347 & n1077 ) | ( n347 & n1461 ) | ( n1077 & n1461 ) ;
  assign n10664 = n10663 ^ n8316 ^ n8087 ;
  assign n10666 = n10665 ^ n10664 ^ n7344 ;
  assign n10668 = n10667 ^ n10666 ^ 1'b0 ;
  assign n10669 = n7517 | n10668 ;
  assign n10670 = n460 & ~n2152 ;
  assign n10671 = n1869 & ~n10627 ;
  assign n10672 = n3594 & n10671 ;
  assign n10673 = ( ~n1363 & n10670 ) | ( ~n1363 & n10672 ) | ( n10670 & n10672 ) ;
  assign n10675 = n961 | n4925 ;
  assign n10676 = n1063 & ~n10675 ;
  assign n10674 = ~n639 & n1212 ;
  assign n10677 = n10676 ^ n10674 ^ 1'b0 ;
  assign n10678 = n1412 ^ x110 ^ 1'b0 ;
  assign n10679 = n10134 & n10678 ;
  assign n10680 = ( n5122 & n7553 ) | ( n5122 & n10414 ) | ( n7553 & n10414 ) ;
  assign n10681 = n10680 ^ n318 ^ 1'b0 ;
  assign n10682 = n4852 ^ n2865 ^ x45 ;
  assign n10683 = n10682 ^ n3959 ^ 1'b0 ;
  assign n10684 = ( x13 & n1963 ) | ( x13 & ~n3574 ) | ( n1963 & ~n3574 ) ;
  assign n10688 = n3322 ^ n447 ^ n306 ;
  assign n10689 = n10688 ^ n7729 ^ n912 ;
  assign n10690 = n3753 & n10689 ;
  assign n10685 = ( ~n3381 & n5151 ) | ( ~n3381 & n5976 ) | ( n5151 & n5976 ) ;
  assign n10686 = n6926 ^ n4165 ^ 1'b0 ;
  assign n10687 = n10685 & n10686 ;
  assign n10691 = n10690 ^ n10687 ^ n8814 ;
  assign n10692 = ( n10683 & n10684 ) | ( n10683 & ~n10691 ) | ( n10684 & ~n10691 ) ;
  assign n10693 = n10692 ^ n5864 ^ 1'b0 ;
  assign n10696 = n3031 & n5575 ;
  assign n10697 = n5740 & n10696 ;
  assign n10694 = n2678 ^ n2070 ^ n1492 ;
  assign n10695 = ( n807 & n10672 ) | ( n807 & n10694 ) | ( n10672 & n10694 ) ;
  assign n10698 = n10697 ^ n10695 ^ 1'b0 ;
  assign n10699 = n2964 | n5485 ;
  assign n10700 = n10699 ^ n2057 ^ n1686 ;
  assign n10701 = n5344 ^ n4516 ^ n2792 ;
  assign n10702 = n7601 ^ n4347 ^ n2521 ;
  assign n10703 = ( n7039 & n10701 ) | ( n7039 & ~n10702 ) | ( n10701 & ~n10702 ) ;
  assign n10704 = n4240 ^ n2697 ^ 1'b0 ;
  assign n10705 = ~n10703 & n10704 ;
  assign n10706 = n10700 & n10705 ;
  assign n10707 = n10706 ^ n269 ^ 1'b0 ;
  assign n10708 = ~n10469 & n10707 ;
  assign n10709 = n3789 | n6968 ;
  assign n10710 = n10424 ^ n1869 ^ x37 ;
  assign n10711 = ( ~x113 & n1952 ) | ( ~x113 & n2507 ) | ( n1952 & n2507 ) ;
  assign n10712 = n10711 ^ n786 ^ 1'b0 ;
  assign n10713 = ( n1500 & n2872 ) | ( n1500 & n10712 ) | ( n2872 & n10712 ) ;
  assign n10714 = ( n2331 & ~n3416 ) | ( n2331 & n8754 ) | ( ~n3416 & n8754 ) ;
  assign n10715 = ( n2569 & n6670 ) | ( n2569 & n9254 ) | ( n6670 & n9254 ) ;
  assign n10716 = n4293 ^ n2691 ^ n968 ;
  assign n10717 = n10605 & n10716 ;
  assign n10718 = n10717 ^ n310 ^ 1'b0 ;
  assign n10719 = n10718 ^ n10639 ^ 1'b0 ;
  assign n10720 = ~n2691 & n3350 ;
  assign n10721 = ~n540 & n10720 ;
  assign n10722 = n10721 ^ n6076 ^ n789 ;
  assign n10723 = n10722 ^ n6187 ^ 1'b0 ;
  assign n10724 = n10723 ^ n6749 ^ 1'b0 ;
  assign n10725 = n1097 & ~n10724 ;
  assign n10726 = ( ~n4010 & n7419 ) | ( ~n4010 & n10725 ) | ( n7419 & n10725 ) ;
  assign n10727 = ( n2450 & ~n3510 ) | ( n2450 & n3526 ) | ( ~n3510 & n3526 ) ;
  assign n10728 = ( n3828 & n10726 ) | ( n3828 & n10727 ) | ( n10726 & n10727 ) ;
  assign n10729 = ( ~n395 & n8547 ) | ( ~n395 & n8685 ) | ( n8547 & n8685 ) ;
  assign n10730 = n9258 ^ n408 ^ 1'b0 ;
  assign n10733 = n8001 ^ n3293 ^ n1754 ;
  assign n10731 = n2489 & n10487 ;
  assign n10732 = n2519 & ~n10731 ;
  assign n10734 = n10733 ^ n10732 ^ 1'b0 ;
  assign n10735 = n10734 ^ n3052 ^ n1586 ;
  assign n10736 = ( n1738 & n4510 ) | ( n1738 & ~n9521 ) | ( n4510 & ~n9521 ) ;
  assign n10737 = ( ~n5332 & n5873 ) | ( ~n5332 & n6605 ) | ( n5873 & n6605 ) ;
  assign n10738 = n10737 ^ n1596 ^ n1349 ;
  assign n10739 = n4986 & ~n10738 ;
  assign n10740 = ( n10735 & n10736 ) | ( n10735 & n10739 ) | ( n10736 & n10739 ) ;
  assign n10741 = n3572 ^ n2725 ^ x216 ;
  assign n10742 = n7285 ^ n3860 ^ x115 ;
  assign n10743 = ( n4698 & ~n10741 ) | ( n4698 & n10742 ) | ( ~n10741 & n10742 ) ;
  assign n10744 = n10743 ^ n7368 ^ 1'b0 ;
  assign n10745 = ~n10740 & n10744 ;
  assign n10754 = n3418 | n8494 ;
  assign n10755 = n10754 ^ n295 ^ 1'b0 ;
  assign n10751 = n5367 ^ n5009 ^ n2830 ;
  assign n10752 = n10751 ^ n10444 ^ n3173 ;
  assign n10753 = n10752 ^ n4610 ^ n2643 ;
  assign n10756 = n10755 ^ n10753 ^ n3085 ;
  assign n10748 = n3332 ^ n2488 ^ n1980 ;
  assign n10746 = n9963 ^ n9583 ^ n1516 ;
  assign n10747 = n10746 ^ n2285 ^ n799 ;
  assign n10749 = n10748 ^ n10747 ^ n704 ;
  assign n10750 = n7051 | n10749 ;
  assign n10757 = n10756 ^ n10750 ^ 1'b0 ;
  assign n10758 = n4332 ^ n1209 ^ n812 ;
  assign n10759 = ( n1278 & n6922 ) | ( n1278 & ~n10758 ) | ( n6922 & ~n10758 ) ;
  assign n10760 = n5963 ^ n612 ^ 1'b0 ;
  assign n10761 = n3803 | n10760 ;
  assign n10763 = n3376 ^ n1585 ^ n1497 ;
  assign n10762 = n6260 & ~n6951 ;
  assign n10764 = n10763 ^ n10762 ^ n4348 ;
  assign n10765 = n5352 ^ n2247 ^ 1'b0 ;
  assign n10766 = n10765 ^ n427 ^ x221 ;
  assign n10767 = n10766 ^ n5399 ^ n3028 ;
  assign n10768 = n10764 & ~n10767 ;
  assign n10769 = ~n10764 & n10768 ;
  assign n10770 = n474 | n7673 ;
  assign n10771 = n6338 & ~n10770 ;
  assign n10772 = ( x34 & ~n399 ) | ( x34 & n10771 ) | ( ~n399 & n10771 ) ;
  assign n10773 = n2144 & n3802 ;
  assign n10774 = n10773 ^ n3942 ^ 1'b0 ;
  assign n10775 = n3498 & n10774 ;
  assign n10776 = ~n3915 & n10775 ;
  assign n10777 = n10776 ^ n8792 ^ 1'b0 ;
  assign n10778 = n10777 ^ n5032 ^ x180 ;
  assign n10779 = ( n1177 & n1567 ) | ( n1177 & n9638 ) | ( n1567 & n9638 ) ;
  assign n10780 = ( n6737 & n9810 ) | ( n6737 & n10779 ) | ( n9810 & n10779 ) ;
  assign n10781 = ~n10778 & n10780 ;
  assign n10782 = n2749 ^ n877 ^ 1'b0 ;
  assign n10783 = n9695 | n10782 ;
  assign n10784 = ( n1730 & n5192 ) | ( n1730 & ~n10783 ) | ( n5192 & ~n10783 ) ;
  assign n10785 = ( n8233 & n10659 ) | ( n8233 & n10784 ) | ( n10659 & n10784 ) ;
  assign n10794 = ( ~x84 & n325 ) | ( ~x84 & n5547 ) | ( n325 & n5547 ) ;
  assign n10786 = n1690 ^ n977 ^ 1'b0 ;
  assign n10787 = ( n1901 & ~n7989 ) | ( n1901 & n10786 ) | ( ~n7989 & n10786 ) ;
  assign n10788 = n8242 ^ n5755 ^ 1'b0 ;
  assign n10789 = n3853 & n10788 ;
  assign n10790 = ( n8295 & n10787 ) | ( n8295 & n10789 ) | ( n10787 & n10789 ) ;
  assign n10791 = n4191 ^ n1194 ^ n919 ;
  assign n10792 = n4459 & n10791 ;
  assign n10793 = n10790 & ~n10792 ;
  assign n10795 = n10794 ^ n10793 ^ 1'b0 ;
  assign n10799 = n5162 ^ n2878 ^ n330 ;
  assign n10800 = n4933 & ~n10799 ;
  assign n10796 = n4380 ^ n2791 ^ n1236 ;
  assign n10797 = n6329 ^ n6175 ^ n3350 ;
  assign n10798 = n10796 | n10797 ;
  assign n10801 = n10800 ^ n10798 ^ 1'b0 ;
  assign n10802 = ( n7183 & ~n8584 ) | ( n7183 & n10801 ) | ( ~n8584 & n10801 ) ;
  assign n10803 = n1385 & ~n3654 ;
  assign n10804 = n9335 & n10803 ;
  assign n10805 = n1026 | n10804 ;
  assign n10808 = ( ~n2907 & n3014 ) | ( ~n2907 & n3613 ) | ( n3014 & n3613 ) ;
  assign n10806 = n327 & ~n10765 ;
  assign n10807 = n3244 & n10806 ;
  assign n10809 = n10808 ^ n10807 ^ 1'b0 ;
  assign n10810 = n711 & n9468 ;
  assign n10811 = n10810 ^ n5933 ^ 1'b0 ;
  assign n10812 = n313 ^ x20 ^ 1'b0 ;
  assign n10813 = n10444 ^ n1482 ^ 1'b0 ;
  assign n10814 = ( ~n5580 & n9583 ) | ( ~n5580 & n10813 ) | ( n9583 & n10813 ) ;
  assign n10815 = n10814 ^ n9663 ^ n5922 ;
  assign n10816 = ( ~n9728 & n10812 ) | ( ~n9728 & n10815 ) | ( n10812 & n10815 ) ;
  assign n10817 = ( x243 & n2362 ) | ( x243 & ~n3211 ) | ( n2362 & ~n3211 ) ;
  assign n10818 = ( ~x155 & n5877 ) | ( ~x155 & n10817 ) | ( n5877 & n10817 ) ;
  assign n10819 = n5858 | n10818 ;
  assign n10820 = n2925 & ~n10819 ;
  assign n10821 = n10820 ^ n3838 ^ 1'b0 ;
  assign n10822 = n10821 ^ n5668 ^ n3502 ;
  assign n10823 = ( n1072 & n4730 ) | ( n1072 & ~n9727 ) | ( n4730 & ~n9727 ) ;
  assign n10824 = n10823 ^ n3122 ^ n1521 ;
  assign n10825 = n5310 & ~n10716 ;
  assign n10826 = n10825 ^ n1077 ^ x183 ;
  assign n10827 = n6423 ^ n1784 ^ n1356 ;
  assign n10828 = n5480 | n10827 ;
  assign n10829 = ~n8521 & n10828 ;
  assign n10830 = ~n10826 & n10829 ;
  assign n10831 = n6394 ^ x137 ^ 1'b0 ;
  assign n10832 = n10170 & ~n10831 ;
  assign n10833 = ~n7196 & n7942 ;
  assign n10834 = n10833 ^ n4749 ^ 1'b0 ;
  assign n10835 = ( n1254 & ~n3732 ) | ( n1254 & n5844 ) | ( ~n3732 & n5844 ) ;
  assign n10836 = x101 | n10835 ;
  assign n10837 = n2813 & n10836 ;
  assign n10838 = n10837 ^ n1866 ^ 1'b0 ;
  assign n10839 = n1701 & n10838 ;
  assign n10840 = n10834 & n10839 ;
  assign n10841 = x1 | n3529 ;
  assign n10842 = n10841 ^ n8193 ^ 1'b0 ;
  assign n10843 = ~n10840 & n10842 ;
  assign n10849 = ( ~x198 & n728 ) | ( ~x198 & n1727 ) | ( n728 & n1727 ) ;
  assign n10850 = n9067 & n10849 ;
  assign n10845 = n436 & n3016 ;
  assign n10844 = ( n725 & n3833 ) | ( n725 & ~n5353 ) | ( n3833 & ~n5353 ) ;
  assign n10846 = n10845 ^ n10844 ^ n6730 ;
  assign n10847 = n10418 & n10846 ;
  assign n10848 = n6972 & n10847 ;
  assign n10851 = n10850 ^ n10848 ^ 1'b0 ;
  assign n10852 = n10040 ^ n3672 ^ n3505 ;
  assign n10853 = n10852 ^ n6352 ^ n3538 ;
  assign n10854 = n10853 ^ n3523 ^ 1'b0 ;
  assign n10855 = n4440 | n10854 ;
  assign n10856 = n3010 ^ n2486 ^ n2385 ;
  assign n10857 = n9030 & ~n10856 ;
  assign n10858 = n10857 ^ n8069 ^ 1'b0 ;
  assign n10859 = ( n4991 & n8932 ) | ( n4991 & n10858 ) | ( n8932 & n10858 ) ;
  assign n10860 = ~n5908 & n6383 ;
  assign n10861 = n1905 & n10860 ;
  assign n10862 = ( ~n10855 & n10859 ) | ( ~n10855 & n10861 ) | ( n10859 & n10861 ) ;
  assign n10863 = n4492 ^ n2308 ^ 1'b0 ;
  assign n10864 = ~n1929 & n2202 ;
  assign n10865 = n10864 ^ n944 ^ 1'b0 ;
  assign n10866 = ( n6996 & n10863 ) | ( n6996 & ~n10865 ) | ( n10863 & ~n10865 ) ;
  assign n10867 = n3359 & n3619 ;
  assign n10868 = n10867 ^ n1871 ^ 1'b0 ;
  assign n10869 = n2055 & ~n6613 ;
  assign n10870 = n9096 ^ n995 ^ n861 ;
  assign n10871 = n733 & n6985 ;
  assign n10872 = n7211 & n10871 ;
  assign n10875 = ~n3621 & n4947 ;
  assign n10873 = n5491 ^ n3481 ^ n1424 ;
  assign n10874 = n10873 ^ n6046 ^ n6005 ;
  assign n10876 = n10875 ^ n10874 ^ n5079 ;
  assign n10877 = ( n5002 & ~n6059 ) | ( n5002 & n9251 ) | ( ~n6059 & n9251 ) ;
  assign n10886 = n3601 & ~n9753 ;
  assign n10887 = n8900 ^ n3253 ^ 1'b0 ;
  assign n10888 = ~n10886 & n10887 ;
  assign n10878 = n658 | n2887 ;
  assign n10879 = n10878 ^ n2430 ^ 1'b0 ;
  assign n10880 = ( n434 & n969 ) | ( n434 & n4598 ) | ( n969 & n4598 ) ;
  assign n10881 = n3675 & ~n7897 ;
  assign n10882 = n10775 & ~n10881 ;
  assign n10883 = n10880 & n10882 ;
  assign n10884 = n591 | n10883 ;
  assign n10885 = n10879 | n10884 ;
  assign n10889 = n10888 ^ n10885 ^ n7735 ;
  assign n10890 = ( n817 & n2678 ) | ( n817 & ~n2907 ) | ( n2678 & ~n2907 ) ;
  assign n10891 = ~n1518 & n10890 ;
  assign n10892 = n10891 ^ n1390 ^ 1'b0 ;
  assign n10894 = n6535 ^ n2962 ^ n1958 ;
  assign n10893 = n1264 | n5224 ;
  assign n10895 = n10894 ^ n10893 ^ n7681 ;
  assign n10896 = n7395 ^ n4032 ^ n3173 ;
  assign n10897 = ( n4336 & ~n8529 ) | ( n4336 & n10896 ) | ( ~n8529 & n10896 ) ;
  assign n10898 = ( n6445 & n7144 ) | ( n6445 & ~n10897 ) | ( n7144 & ~n10897 ) ;
  assign n10899 = ( n4626 & n10895 ) | ( n4626 & ~n10898 ) | ( n10895 & ~n10898 ) ;
  assign n10900 = ( n1015 & n10892 ) | ( n1015 & n10899 ) | ( n10892 & n10899 ) ;
  assign n10901 = n360 & n8173 ;
  assign n10902 = ~n3052 & n10901 ;
  assign n10903 = ( n559 & n3439 ) | ( n559 & ~n5000 ) | ( n3439 & ~n5000 ) ;
  assign n10904 = n2268 & n5841 ;
  assign n10905 = n10903 & n10904 ;
  assign n10906 = n10841 ^ n950 ^ x79 ;
  assign n10907 = ( ~n5211 & n6971 ) | ( ~n5211 & n7238 ) | ( n6971 & n7238 ) ;
  assign n10908 = ( n693 & n9264 ) | ( n693 & ~n10907 ) | ( n9264 & ~n10907 ) ;
  assign n10911 = n1129 & n2951 ;
  assign n10912 = n10911 ^ n4230 ^ 1'b0 ;
  assign n10909 = n4970 ^ n3603 ^ 1'b0 ;
  assign n10910 = ~n2560 & n10909 ;
  assign n10913 = n10912 ^ n10910 ^ n4639 ;
  assign n10914 = ( n859 & n2273 ) | ( n859 & n2371 ) | ( n2273 & n2371 ) ;
  assign n10915 = n10914 ^ n9212 ^ n9199 ;
  assign n10916 = n10915 ^ n10093 ^ 1'b0 ;
  assign n10917 = n5054 & n10916 ;
  assign n10918 = n10913 & ~n10917 ;
  assign n10919 = n10918 ^ n8961 ^ n8770 ;
  assign n10920 = n5973 & n10272 ;
  assign n10921 = n6364 ^ n4296 ^ n1020 ;
  assign n10922 = n10921 ^ n3784 ^ n2984 ;
  assign n10923 = ( ~x55 & n4963 ) | ( ~x55 & n7101 ) | ( n4963 & n7101 ) ;
  assign n10924 = ( n5308 & ~n10922 ) | ( n5308 & n10923 ) | ( ~n10922 & n10923 ) ;
  assign n10925 = n9271 ^ n3931 ^ n1842 ;
  assign n10926 = ~n10924 & n10925 ;
  assign n10928 = n6803 ^ n2408 ^ n1202 ;
  assign n10927 = ( n894 & ~n2180 ) | ( n894 & n4049 ) | ( ~n2180 & n4049 ) ;
  assign n10929 = n10928 ^ n10927 ^ n1496 ;
  assign n10930 = n10929 ^ n5205 ^ n589 ;
  assign n10931 = ( n336 & n9584 ) | ( n336 & n10930 ) | ( n9584 & n10930 ) ;
  assign n10932 = n4849 ^ n1316 ^ 1'b0 ;
  assign n10933 = n5118 & n10932 ;
  assign n10934 = ~n1487 & n2260 ;
  assign n10935 = ~n10933 & n10934 ;
  assign n10936 = n10935 ^ n9758 ^ n5265 ;
  assign n10937 = ( ~n8244 & n9919 ) | ( ~n8244 & n10936 ) | ( n9919 & n10936 ) ;
  assign n10959 = n7134 ^ n6062 ^ n4830 ;
  assign n10958 = n3271 ^ n2601 ^ 1'b0 ;
  assign n10960 = n10959 ^ n10958 ^ 1'b0 ;
  assign n10938 = n5759 ^ n3383 ^ 1'b0 ;
  assign n10939 = ~n4673 & n10938 ;
  assign n10940 = n5733 | n10939 ;
  assign n10941 = n6365 ^ n2033 ^ 1'b0 ;
  assign n10942 = n10940 & n10941 ;
  assign n10943 = n3005 ^ n2825 ^ n1924 ;
  assign n10944 = n4093 & ~n5343 ;
  assign n10945 = n10944 ^ n1899 ^ 1'b0 ;
  assign n10946 = n2629 & n10945 ;
  assign n10947 = n4192 & n10946 ;
  assign n10948 = ( ~n3534 & n10943 ) | ( ~n3534 & n10947 ) | ( n10943 & n10947 ) ;
  assign n10949 = n10942 | n10948 ;
  assign n10950 = n2014 | n7566 ;
  assign n10951 = n10950 ^ n3377 ^ 1'b0 ;
  assign n10952 = n5986 ^ n2302 ^ 1'b0 ;
  assign n10953 = ( n1282 & ~n4234 ) | ( n1282 & n10152 ) | ( ~n4234 & n10152 ) ;
  assign n10954 = ( n10951 & n10952 ) | ( n10951 & ~n10953 ) | ( n10952 & ~n10953 ) ;
  assign n10955 = n10954 ^ n5723 ^ n3606 ;
  assign n10956 = n9033 & ~n10955 ;
  assign n10957 = ~n10949 & n10956 ;
  assign n10961 = n10960 ^ n10957 ^ 1'b0 ;
  assign n10962 = n3506 & n4609 ;
  assign n10963 = n10962 ^ n295 ^ 1'b0 ;
  assign n10964 = n10963 ^ n4866 ^ 1'b0 ;
  assign n10965 = n3772 | n10964 ;
  assign n10966 = ( n3668 & n7668 ) | ( n3668 & n10965 ) | ( n7668 & n10965 ) ;
  assign n10967 = n7366 & ~n10966 ;
  assign n10968 = ( ~n6808 & n9725 ) | ( ~n6808 & n10967 ) | ( n9725 & n10967 ) ;
  assign n10969 = ( ~n2441 & n3202 ) | ( ~n2441 & n4147 ) | ( n3202 & n4147 ) ;
  assign n10970 = ( n5249 & n9171 ) | ( n5249 & n10969 ) | ( n9171 & n10969 ) ;
  assign n10971 = ~n2116 & n10970 ;
  assign n10972 = n4012 ^ n2366 ^ n1524 ;
  assign n10973 = n3921 ^ n3508 ^ n2508 ;
  assign n10974 = n6144 & ~n10973 ;
  assign n10975 = x183 & ~n10974 ;
  assign n10976 = ~n3415 & n10975 ;
  assign n10977 = n10972 | n10976 ;
  assign n10978 = n10977 ^ n9012 ^ 1'b0 ;
  assign n10979 = x201 & n4825 ;
  assign n10980 = n4688 ^ n1632 ^ n1612 ;
  assign n10981 = n10980 ^ n9349 ^ n2899 ;
  assign n10982 = ( n4893 & ~n7148 ) | ( n4893 & n10981 ) | ( ~n7148 & n10981 ) ;
  assign n10983 = n5182 ^ n735 ^ 1'b0 ;
  assign n10984 = ~n1826 & n2158 ;
  assign n10985 = n637 & n10984 ;
  assign n10986 = ( n1240 & ~n3737 ) | ( n1240 & n10985 ) | ( ~n3737 & n10985 ) ;
  assign n10987 = ( n3292 & n10983 ) | ( n3292 & ~n10986 ) | ( n10983 & ~n10986 ) ;
  assign n10988 = ( n10979 & n10982 ) | ( n10979 & n10987 ) | ( n10982 & n10987 ) ;
  assign n10989 = ( n1324 & n6394 ) | ( n1324 & n7099 ) | ( n6394 & n7099 ) ;
  assign n10990 = ( ~n1977 & n2995 ) | ( ~n1977 & n3758 ) | ( n2995 & n3758 ) ;
  assign n10991 = n10990 ^ n7261 ^ 1'b0 ;
  assign n10992 = n10991 ^ n7366 ^ 1'b0 ;
  assign n10993 = n7862 & ~n10992 ;
  assign n10994 = n10993 ^ n7979 ^ 1'b0 ;
  assign n10995 = n3452 & ~n10994 ;
  assign n10996 = n6737 ^ n1801 ^ x91 ;
  assign n10997 = ~n10439 & n10996 ;
  assign n10998 = ~n9494 & n10997 ;
  assign n10999 = n4240 ^ n474 ^ 1'b0 ;
  assign n11000 = ~n4571 & n10999 ;
  assign n11001 = ( n3965 & ~n6671 ) | ( n3965 & n11000 ) | ( ~n6671 & n11000 ) ;
  assign n11002 = ( ~n849 & n10998 ) | ( ~n849 & n11001 ) | ( n10998 & n11001 ) ;
  assign n11003 = x68 & ~n7854 ;
  assign n11004 = n11003 ^ n3520 ^ 1'b0 ;
  assign n11005 = ( n3870 & n7292 ) | ( n3870 & ~n11004 ) | ( n7292 & ~n11004 ) ;
  assign n11009 = n7314 ^ n3779 ^ n3670 ;
  assign n11006 = n3552 ^ n2806 ^ 1'b0 ;
  assign n11007 = n11006 ^ n5154 ^ 1'b0 ;
  assign n11008 = ~n8036 & n11007 ;
  assign n11010 = n11009 ^ n11008 ^ n5119 ;
  assign n11011 = n9104 ^ n5129 ^ n4376 ;
  assign n11012 = n5442 | n11011 ;
  assign n11013 = n3538 | n10065 ;
  assign n11014 = n11012 & ~n11013 ;
  assign n11015 = ~n2992 & n3931 ;
  assign n11017 = n2195 ^ n1136 ^ n750 ;
  assign n11020 = n5583 ^ n3738 ^ 1'b0 ;
  assign n11021 = n4410 & n11020 ;
  assign n11018 = n589 | n3554 ;
  assign n11019 = n11018 ^ n1361 ^ 1'b0 ;
  assign n11022 = n11021 ^ n11019 ^ n1848 ;
  assign n11023 = ( ~n3768 & n11017 ) | ( ~n3768 & n11022 ) | ( n11017 & n11022 ) ;
  assign n11016 = ( ~n1435 & n8552 ) | ( ~n1435 & n9878 ) | ( n8552 & n9878 ) ;
  assign n11024 = n11023 ^ n11016 ^ 1'b0 ;
  assign n11025 = ( ~n4623 & n11015 ) | ( ~n4623 & n11024 ) | ( n11015 & n11024 ) ;
  assign n11026 = n10771 ^ n7981 ^ n4229 ;
  assign n11030 = ( ~n903 & n3127 ) | ( ~n903 & n5069 ) | ( n3127 & n5069 ) ;
  assign n11029 = ( n1587 & n4765 ) | ( n1587 & n7214 ) | ( n4765 & n7214 ) ;
  assign n11031 = n11030 ^ n11029 ^ 1'b0 ;
  assign n11027 = n364 | n8810 ;
  assign n11028 = ~n5367 & n11027 ;
  assign n11032 = n11031 ^ n11028 ^ 1'b0 ;
  assign n11033 = x3 & n4014 ;
  assign n11034 = n11033 ^ n1486 ^ 1'b0 ;
  assign n11035 = n11034 ^ n5991 ^ n2631 ;
  assign n11036 = n7971 & ~n11035 ;
  assign n11037 = n4883 ^ n896 ^ 1'b0 ;
  assign n11038 = n11037 ^ n8104 ^ n541 ;
  assign n11039 = n4817 ^ n3636 ^ n1751 ;
  assign n11040 = ( n4310 & n9452 ) | ( n4310 & n11039 ) | ( n9452 & n11039 ) ;
  assign n11041 = n8292 ^ n2011 ^ 1'b0 ;
  assign n11042 = n11040 | n11041 ;
  assign n11044 = ( ~n1957 & n5955 ) | ( ~n1957 & n10335 ) | ( n5955 & n10335 ) ;
  assign n11045 = ( n3724 & n8078 ) | ( n3724 & ~n11044 ) | ( n8078 & ~n11044 ) ;
  assign n11043 = n2740 ^ n2725 ^ 1'b0 ;
  assign n11046 = n11045 ^ n11043 ^ 1'b0 ;
  assign n11052 = n4740 ^ n2024 ^ n1206 ;
  assign n11048 = n2725 | n3441 ;
  assign n11047 = n1278 & ~n3643 ;
  assign n11049 = n11048 ^ n11047 ^ 1'b0 ;
  assign n11050 = n11049 ^ n9212 ^ 1'b0 ;
  assign n11051 = n687 & n11050 ;
  assign n11053 = n11052 ^ n11051 ^ n9405 ;
  assign n11054 = n9552 ^ n3240 ^ 1'b0 ;
  assign n11055 = ~n2989 & n11054 ;
  assign n11056 = ~n11053 & n11055 ;
  assign n11057 = n10054 | n10477 ;
  assign n11058 = n1575 & ~n11057 ;
  assign n11059 = n10910 ^ n7970 ^ n664 ;
  assign n11060 = ( x134 & ~n8916 ) | ( x134 & n11059 ) | ( ~n8916 & n11059 ) ;
  assign n11061 = ( n3643 & n4787 ) | ( n3643 & ~n11060 ) | ( n4787 & ~n11060 ) ;
  assign n11067 = ( n1741 & n2206 ) | ( n1741 & ~n3438 ) | ( n2206 & ~n3438 ) ;
  assign n11065 = ( n1212 & ~n3279 ) | ( n1212 & n3966 ) | ( ~n3279 & n3966 ) ;
  assign n11062 = n4070 ^ n1414 ^ x239 ;
  assign n11063 = n11062 ^ n1722 ^ 1'b0 ;
  assign n11064 = ~n5262 & n11063 ;
  assign n11066 = n11065 ^ n11064 ^ 1'b0 ;
  assign n11068 = n11067 ^ n11066 ^ 1'b0 ;
  assign n11069 = n11068 ^ n10902 ^ n7766 ;
  assign n11078 = ~n508 & n2257 ;
  assign n11070 = n883 & n7151 ;
  assign n11071 = n11070 ^ n3636 ^ 1'b0 ;
  assign n11075 = ( n1058 & n2014 ) | ( n1058 & ~n5293 ) | ( n2014 & ~n5293 ) ;
  assign n11073 = ~n621 & n7611 ;
  assign n11072 = ( x246 & n2645 ) | ( x246 & n8640 ) | ( n2645 & n8640 ) ;
  assign n11074 = n11073 ^ n11072 ^ n2489 ;
  assign n11076 = n11075 ^ n11074 ^ n6653 ;
  assign n11077 = n11071 & n11076 ;
  assign n11079 = n11078 ^ n11077 ^ 1'b0 ;
  assign n11080 = n381 & ~n8014 ;
  assign n11081 = n295 | n11080 ;
  assign n11082 = n951 & n11081 ;
  assign n11085 = n5997 & ~n6049 ;
  assign n11083 = n10212 ^ n8767 ^ n4072 ;
  assign n11084 = n11083 ^ n7202 ^ n6043 ;
  assign n11086 = n11085 ^ n11084 ^ 1'b0 ;
  assign n11087 = ~n4826 & n11086 ;
  assign n11089 = n6704 & n7691 ;
  assign n11088 = n6764 ^ n5743 ^ n4421 ;
  assign n11090 = n11089 ^ n11088 ^ n6775 ;
  assign n11091 = n8019 ^ n7042 ^ x46 ;
  assign n11092 = ( n1871 & ~n5430 ) | ( n1871 & n11091 ) | ( ~n5430 & n11091 ) ;
  assign n11093 = ( n2905 & ~n3646 ) | ( n2905 & n8160 ) | ( ~n3646 & n8160 ) ;
  assign n11094 = n11093 ^ n8690 ^ 1'b0 ;
  assign n11095 = n11092 & n11094 ;
  assign n11096 = n3333 ^ n343 ^ 1'b0 ;
  assign n11097 = n3781 | n11096 ;
  assign n11098 = n11097 ^ n8480 ^ n4638 ;
  assign n11099 = ~n5357 & n8480 ;
  assign n11100 = n11099 ^ n8718 ^ 1'b0 ;
  assign n11101 = ( n7445 & n9109 ) | ( n7445 & n10501 ) | ( n9109 & n10501 ) ;
  assign n11109 = n10091 ^ n4517 ^ 1'b0 ;
  assign n11110 = n552 & ~n11109 ;
  assign n11102 = ( x216 & ~n3040 ) | ( x216 & n4070 ) | ( ~n3040 & n4070 ) ;
  assign n11103 = n987 & n7162 ;
  assign n11104 = ( n1212 & n3860 ) | ( n1212 & ~n10638 ) | ( n3860 & ~n10638 ) ;
  assign n11105 = n11104 ^ n6968 ^ 1'b0 ;
  assign n11106 = n11103 & n11105 ;
  assign n11107 = ( n3397 & n7160 ) | ( n3397 & ~n9019 ) | ( n7160 & ~n9019 ) ;
  assign n11108 = ( n11102 & ~n11106 ) | ( n11102 & n11107 ) | ( ~n11106 & n11107 ) ;
  assign n11111 = n11110 ^ n11108 ^ n3506 ;
  assign n11112 = n2622 & ~n10959 ;
  assign n11113 = n9947 & n11112 ;
  assign n11114 = ( n1265 & n7030 ) | ( n1265 & ~n8169 ) | ( n7030 & ~n8169 ) ;
  assign n11115 = n7060 | n11114 ;
  assign n11116 = n10834 ^ n6216 ^ 1'b0 ;
  assign n11117 = n2348 & n4480 ;
  assign n11118 = n11117 ^ n2614 ^ 1'b0 ;
  assign n11119 = n3885 & ~n7047 ;
  assign n11120 = n11119 ^ n3158 ^ 1'b0 ;
  assign n11121 = n2997 & ~n7968 ;
  assign n11122 = ~n11120 & n11121 ;
  assign n11124 = n10796 ^ x174 ^ 1'b0 ;
  assign n11123 = ~n2053 & n6714 ;
  assign n11125 = n11124 ^ n11123 ^ 1'b0 ;
  assign n11126 = ( ~n344 & n1258 ) | ( ~n344 & n9601 ) | ( n1258 & n9601 ) ;
  assign n11127 = n10487 ^ n2538 ^ 1'b0 ;
  assign n11128 = ( ~n11125 & n11126 ) | ( ~n11125 & n11127 ) | ( n11126 & n11127 ) ;
  assign n11129 = ~n4840 & n11128 ;
  assign n11130 = n11129 ^ n3842 ^ 1'b0 ;
  assign n11131 = x70 & ~x149 ;
  assign n11132 = n7006 | n11131 ;
  assign n11133 = n11132 ^ n6067 ^ 1'b0 ;
  assign n11134 = n11133 ^ n2252 ^ 1'b0 ;
  assign n11135 = ~n11130 & n11134 ;
  assign n11137 = n5823 ^ n5178 ^ n1146 ;
  assign n11138 = n885 | n5932 ;
  assign n11139 = n11138 ^ n5735 ^ 1'b0 ;
  assign n11140 = ( n6994 & ~n7523 ) | ( n6994 & n11139 ) | ( ~n7523 & n11139 ) ;
  assign n11141 = ( n2103 & n8115 ) | ( n2103 & n11140 ) | ( n8115 & n11140 ) ;
  assign n11142 = n11137 | n11141 ;
  assign n11143 = n11142 ^ n1054 ^ 1'b0 ;
  assign n11144 = n11143 ^ n4029 ^ 1'b0 ;
  assign n11136 = ( n7620 & n8304 ) | ( n7620 & n9145 ) | ( n8304 & n9145 ) ;
  assign n11145 = n11144 ^ n11136 ^ 1'b0 ;
  assign n11146 = n4883 | n11145 ;
  assign n11147 = n3931 ^ n3126 ^ n332 ;
  assign n11148 = n11147 ^ n10791 ^ n505 ;
  assign n11149 = n11148 ^ n7283 ^ n1947 ;
  assign n11150 = n3753 & ~n5294 ;
  assign n11151 = n11150 ^ n2889 ^ 1'b0 ;
  assign n11152 = n11151 ^ n2451 ^ n2054 ;
  assign n11153 = n2089 & ~n11152 ;
  assign n11154 = n11153 ^ n8750 ^ 1'b0 ;
  assign n11155 = n11149 | n11154 ;
  assign n11156 = n4665 & ~n10443 ;
  assign n11157 = n7723 & ~n11156 ;
  assign n11158 = n11157 ^ n3920 ^ 1'b0 ;
  assign n11159 = n11155 | n11158 ;
  assign n11160 = ( n336 & n847 ) | ( n336 & ~n5220 ) | ( n847 & ~n5220 ) ;
  assign n11161 = ( ~n5142 & n7294 ) | ( ~n5142 & n11160 ) | ( n7294 & n11160 ) ;
  assign n11164 = n7883 ^ n2452 ^ n1387 ;
  assign n11165 = ( n821 & n6124 ) | ( n821 & n11164 ) | ( n6124 & n11164 ) ;
  assign n11166 = n9253 ^ n2542 ^ 1'b0 ;
  assign n11167 = ( n5870 & ~n11165 ) | ( n5870 & n11166 ) | ( ~n11165 & n11166 ) ;
  assign n11162 = ( ~n4096 & n9576 ) | ( ~n4096 & n10475 ) | ( n9576 & n10475 ) ;
  assign n11163 = ( ~n2525 & n2939 ) | ( ~n2525 & n11162 ) | ( n2939 & n11162 ) ;
  assign n11168 = n11167 ^ n11163 ^ n4550 ;
  assign n11188 = n2960 ^ n2108 ^ n1962 ;
  assign n11187 = n5637 & n6712 ;
  assign n11174 = n4729 ^ n1317 ^ 1'b0 ;
  assign n11175 = n401 & ~n11174 ;
  assign n11183 = n484 ^ x59 ^ 1'b0 ;
  assign n11179 = n5296 & n5790 ;
  assign n11180 = n11179 ^ n6765 ^ 1'b0 ;
  assign n11181 = n8360 & n11180 ;
  assign n11182 = n11181 ^ n4268 ^ 1'b0 ;
  assign n11177 = ( ~n1320 & n1956 ) | ( ~n1320 & n3866 ) | ( n1956 & n3866 ) ;
  assign n11176 = n3158 & n4586 ;
  assign n11178 = n11177 ^ n11176 ^ n4099 ;
  assign n11184 = n11183 ^ n11182 ^ n11178 ;
  assign n11185 = n11184 ^ n10844 ^ 1'b0 ;
  assign n11186 = n11175 & n11185 ;
  assign n11189 = n11188 ^ n11187 ^ n11186 ;
  assign n11169 = n10303 ^ n2152 ^ 1'b0 ;
  assign n11170 = n5620 | n11169 ;
  assign n11171 = x188 | n349 ;
  assign n11172 = n11170 & n11171 ;
  assign n11173 = n4419 | n11172 ;
  assign n11190 = n11189 ^ n11173 ^ 1'b0 ;
  assign n11191 = n6252 ^ n4349 ^ 1'b0 ;
  assign n11192 = ( n3720 & n5948 ) | ( n3720 & ~n6169 ) | ( n5948 & ~n6169 ) ;
  assign n11193 = n11192 ^ n6310 ^ 1'b0 ;
  assign n11194 = n11191 & n11193 ;
  assign n11195 = n1764 | n9969 ;
  assign n11196 = n1402 | n11195 ;
  assign n11197 = n3998 & ~n11196 ;
  assign n11198 = ( n4985 & n6378 ) | ( n4985 & n10371 ) | ( n6378 & n10371 ) ;
  assign n11199 = ( n1845 & n4034 ) | ( n1845 & ~n5207 ) | ( n4034 & ~n5207 ) ;
  assign n11200 = ( n1509 & ~n11198 ) | ( n1509 & n11199 ) | ( ~n11198 & n11199 ) ;
  assign n11201 = n10049 ^ n6917 ^ n5385 ;
  assign n11202 = n5290 & ~n11201 ;
  assign n11203 = n11202 ^ n7110 ^ 1'b0 ;
  assign n11204 = n9272 ^ n7565 ^ n3365 ;
  assign n11206 = n1720 & ~n2531 ;
  assign n11205 = n4466 ^ n3993 ^ n3670 ;
  assign n11207 = n11206 ^ n11205 ^ n10349 ;
  assign n11208 = n6042 ^ n3631 ^ n988 ;
  assign n11209 = n11208 ^ n10940 ^ 1'b0 ;
  assign n11210 = n11209 ^ n9874 ^ n5284 ;
  assign n11211 = ( ~x51 & n5481 ) | ( ~x51 & n11210 ) | ( n5481 & n11210 ) ;
  assign n11212 = n1215 & ~n6794 ;
  assign n11213 = n7465 & n11212 ;
  assign n11214 = n11213 ^ n9957 ^ n3700 ;
  assign n11220 = n2352 ^ n1994 ^ 1'b0 ;
  assign n11221 = n1497 | n11220 ;
  assign n11215 = n571 & n1425 ;
  assign n11216 = n742 & n11215 ;
  assign n11217 = ( n3218 & ~n10154 ) | ( n3218 & n11216 ) | ( ~n10154 & n11216 ) ;
  assign n11218 = ( ~n2589 & n9467 ) | ( ~n2589 & n11217 ) | ( n9467 & n11217 ) ;
  assign n11219 = ~n3530 & n11218 ;
  assign n11222 = n11221 ^ n11219 ^ 1'b0 ;
  assign n11223 = n11214 & ~n11222 ;
  assign n11224 = n4445 ^ x116 ^ 1'b0 ;
  assign n11225 = n3180 & ~n11224 ;
  assign n11226 = n3363 | n5529 ;
  assign n11227 = n11226 ^ n4740 ^ n1012 ;
  assign n11228 = n11227 ^ n11083 ^ 1'b0 ;
  assign n11232 = ~n1194 & n4705 ;
  assign n11233 = n11232 ^ n10791 ^ n3538 ;
  assign n11229 = n3813 & ~n10549 ;
  assign n11230 = n5262 & n11229 ;
  assign n11231 = n11230 ^ n11127 ^ n1217 ;
  assign n11234 = n11233 ^ n11231 ^ n8050 ;
  assign n11235 = n3203 | n8095 ;
  assign n11236 = ( n511 & ~n3730 ) | ( n511 & n5674 ) | ( ~n3730 & n5674 ) ;
  assign n11237 = n8512 & ~n11236 ;
  assign n11238 = ~n7868 & n11237 ;
  assign n11239 = ( n4457 & ~n5399 ) | ( n4457 & n11238 ) | ( ~n5399 & n11238 ) ;
  assign n11240 = n6945 ^ n3678 ^ 1'b0 ;
  assign n11241 = n11240 ^ n6346 ^ n2705 ;
  assign n11242 = n11241 ^ n5887 ^ 1'b0 ;
  assign n11244 = ~n2890 & n3175 ;
  assign n11243 = n4628 & ~n7196 ;
  assign n11245 = n11244 ^ n11243 ^ 1'b0 ;
  assign n11246 = n3977 & n11245 ;
  assign n11247 = n4423 & n11246 ;
  assign n11248 = n11242 | n11247 ;
  assign n11253 = n8692 ^ n4793 ^ n4420 ;
  assign n11249 = ~n697 & n3155 ;
  assign n11250 = n9484 & n11249 ;
  assign n11251 = n11250 ^ n8542 ^ n2926 ;
  assign n11252 = ( n2038 & ~n3858 ) | ( n2038 & n11251 ) | ( ~n3858 & n11251 ) ;
  assign n11254 = n11253 ^ n11252 ^ n5328 ;
  assign n11255 = ( n559 & n2739 ) | ( n559 & n2974 ) | ( n2739 & n2974 ) ;
  assign n11256 = ( ~n747 & n3757 ) | ( ~n747 & n11255 ) | ( n3757 & n11255 ) ;
  assign n11257 = ( n4398 & ~n9101 ) | ( n4398 & n11256 ) | ( ~n9101 & n11256 ) ;
  assign n11258 = n2610 | n3496 ;
  assign n11259 = n11258 ^ n9869 ^ 1'b0 ;
  assign n11260 = ( n9277 & ~n10595 ) | ( n9277 & n11259 ) | ( ~n10595 & n11259 ) ;
  assign n11261 = ( n1240 & n2199 ) | ( n1240 & n3322 ) | ( n2199 & n3322 ) ;
  assign n11262 = ( n4211 & n8939 ) | ( n4211 & n11261 ) | ( n8939 & n11261 ) ;
  assign n11263 = n11262 ^ n2997 ^ n2760 ;
  assign n11264 = n9004 ^ n8839 ^ n7694 ;
  assign n11265 = n11264 ^ n9225 ^ n713 ;
  assign n11266 = n7580 ^ n6766 ^ 1'b0 ;
  assign n11267 = n4886 ^ n3988 ^ n1956 ;
  assign n11268 = n5801 | n11267 ;
  assign n11269 = x134 | n11268 ;
  assign n11270 = n4057 ^ n1560 ^ 1'b0 ;
  assign n11271 = n4420 & ~n11270 ;
  assign n11272 = ~n2256 & n11271 ;
  assign n11273 = ~n11269 & n11272 ;
  assign n11277 = ( n1006 & ~n1638 ) | ( n1006 & n6030 ) | ( ~n1638 & n6030 ) ;
  assign n11278 = ~n2208 & n11277 ;
  assign n11279 = n11278 ^ n1496 ^ 1'b0 ;
  assign n11274 = n2594 ^ x28 ^ 1'b0 ;
  assign n11275 = n4176 & ~n11274 ;
  assign n11276 = ~n4138 & n11275 ;
  assign n11280 = n11279 ^ n11276 ^ 1'b0 ;
  assign n11286 = n2751 & n6905 ;
  assign n11287 = ( n907 & ~n1889 ) | ( n907 & n11286 ) | ( ~n1889 & n11286 ) ;
  assign n11285 = n8732 ^ n7714 ^ n462 ;
  assign n11281 = n3645 ^ n1225 ^ 1'b0 ;
  assign n11282 = ~n901 & n11281 ;
  assign n11283 = n11282 ^ n4075 ^ 1'b0 ;
  assign n11284 = ( n1860 & n4658 ) | ( n1860 & n11283 ) | ( n4658 & n11283 ) ;
  assign n11288 = n11287 ^ n11285 ^ n11284 ;
  assign n11289 = n4653 ^ n3387 ^ 1'b0 ;
  assign n11290 = n1597 | n2810 ;
  assign n11291 = n11290 ^ n389 ^ 1'b0 ;
  assign n11292 = n4928 ^ n1349 ^ n854 ;
  assign n11293 = ( n11289 & ~n11291 ) | ( n11289 & n11292 ) | ( ~n11291 & n11292 ) ;
  assign n11294 = n11293 ^ n9107 ^ 1'b0 ;
  assign n11295 = n360 & n11294 ;
  assign n11296 = n1480 & n7434 ;
  assign n11297 = n3349 & n11296 ;
  assign n11298 = n8877 ^ n8236 ^ n401 ;
  assign n11299 = ( ~n1267 & n2536 ) | ( ~n1267 & n7162 ) | ( n2536 & n7162 ) ;
  assign n11300 = n11299 ^ n3278 ^ n2350 ;
  assign n11301 = n2678 ^ x38 ^ 1'b0 ;
  assign n11302 = n11301 ^ n5328 ^ 1'b0 ;
  assign n11303 = n4636 | n7569 ;
  assign n11304 = n6150 & n11303 ;
  assign n11305 = n11304 ^ n5618 ^ 1'b0 ;
  assign n11306 = ( n1529 & n11302 ) | ( n1529 & n11305 ) | ( n11302 & n11305 ) ;
  assign n11307 = ( n3367 & n11300 ) | ( n3367 & n11306 ) | ( n11300 & n11306 ) ;
  assign n11308 = n9320 | n11307 ;
  assign n11309 = n10429 ^ n1558 ^ n1205 ;
  assign n11320 = ( n1208 & n3408 ) | ( n1208 & ~n5253 ) | ( n3408 & ~n5253 ) ;
  assign n11310 = x191 | n3054 ;
  assign n11311 = n2807 & ~n11310 ;
  assign n11314 = n6666 ^ n4928 ^ n1718 ;
  assign n11315 = ~n1055 & n11314 ;
  assign n11316 = n11315 ^ n845 ^ 1'b0 ;
  assign n11317 = ( x73 & ~n1642 ) | ( x73 & n11316 ) | ( ~n1642 & n11316 ) ;
  assign n11312 = ( n3351 & ~n6831 ) | ( n3351 & n10346 ) | ( ~n6831 & n10346 ) ;
  assign n11313 = ( n676 & n3255 ) | ( n676 & n11312 ) | ( n3255 & n11312 ) ;
  assign n11318 = n11317 ^ n11313 ^ n4288 ;
  assign n11319 = n11311 | n11318 ;
  assign n11321 = n11320 ^ n11319 ^ 1'b0 ;
  assign n11322 = n7603 ^ x202 ^ 1'b0 ;
  assign n11323 = n11322 ^ n8180 ^ n5458 ;
  assign n11324 = n8840 ^ n5774 ^ n1125 ;
  assign n11325 = ( n6081 & ~n11323 ) | ( n6081 & n11324 ) | ( ~n11323 & n11324 ) ;
  assign n11326 = n8804 & ~n11325 ;
  assign n11327 = n11326 ^ n9297 ^ 1'b0 ;
  assign n11328 = n5233 & ~n8551 ;
  assign n11329 = n11328 ^ n9233 ^ n3460 ;
  assign n11330 = ( n1305 & ~n3587 ) | ( n1305 & n4904 ) | ( ~n3587 & n4904 ) ;
  assign n11331 = n11330 ^ n9145 ^ n8519 ;
  assign n11332 = ( ~n5480 & n10688 ) | ( ~n5480 & n11331 ) | ( n10688 & n11331 ) ;
  assign n11333 = n5067 | n9632 ;
  assign n11334 = n11317 ^ x192 ^ x160 ;
  assign n11337 = n1453 & n8926 ;
  assign n11338 = n11337 ^ n2441 ^ 1'b0 ;
  assign n11335 = n10248 ^ n8311 ^ n1401 ;
  assign n11336 = n11335 ^ n5284 ^ n1324 ;
  assign n11339 = n11338 ^ n11336 ^ 1'b0 ;
  assign n11340 = n11334 & n11339 ;
  assign n11342 = n10305 ^ n4668 ^ 1'b0 ;
  assign n11341 = n5512 ^ n2678 ^ 1'b0 ;
  assign n11343 = n11342 ^ n11341 ^ n1123 ;
  assign n11344 = ( n2288 & n10826 ) | ( n2288 & n11343 ) | ( n10826 & n11343 ) ;
  assign n11348 = n9859 ^ n7955 ^ n1219 ;
  assign n11345 = n5994 ^ n4983 ^ 1'b0 ;
  assign n11346 = n8541 & n11345 ;
  assign n11347 = n11346 ^ n10430 ^ 1'b0 ;
  assign n11349 = n11348 ^ n11347 ^ n6345 ;
  assign n11350 = n11349 ^ n3086 ^ 1'b0 ;
  assign n11351 = n8618 | n11350 ;
  assign n11352 = ( n6408 & n7989 ) | ( n6408 & n11191 ) | ( n7989 & n11191 ) ;
  assign n11353 = n2427 | n7133 ;
  assign n11354 = n11353 ^ n1296 ^ 1'b0 ;
  assign n11355 = n11354 ^ n7694 ^ 1'b0 ;
  assign n11356 = ( n7832 & n10879 ) | ( n7832 & ~n11022 ) | ( n10879 & ~n11022 ) ;
  assign n11357 = n4027 & n8338 ;
  assign n11358 = n11357 ^ n856 ^ 1'b0 ;
  assign n11359 = n11356 & ~n11358 ;
  assign n11360 = ( n2777 & n5597 ) | ( n2777 & ~n11359 ) | ( n5597 & ~n11359 ) ;
  assign n11361 = ( n366 & n399 ) | ( n366 & n5421 ) | ( n399 & n5421 ) ;
  assign n11362 = n9226 ^ n797 ^ x49 ;
  assign n11363 = n11362 ^ n4060 ^ n3333 ;
  assign n11364 = n4474 | n11363 ;
  assign n11365 = ( ~n3594 & n7327 ) | ( ~n3594 & n11364 ) | ( n7327 & n11364 ) ;
  assign n11367 = n7328 ^ x141 ^ 1'b0 ;
  assign n11366 = ~n1567 & n5876 ;
  assign n11368 = n11367 ^ n11366 ^ 1'b0 ;
  assign n11369 = n4623 & ~n8338 ;
  assign n11370 = n11369 ^ n1213 ^ 1'b0 ;
  assign n11371 = n11368 & n11370 ;
  assign n11372 = ( n1317 & ~n4945 ) | ( n1317 & n5724 ) | ( ~n4945 & n5724 ) ;
  assign n11373 = ~n3135 & n11017 ;
  assign n11374 = ( n667 & ~n2869 ) | ( n667 & n3569 ) | ( ~n2869 & n3569 ) ;
  assign n11375 = ~n11373 & n11374 ;
  assign n11376 = n11375 ^ n10333 ^ 1'b0 ;
  assign n11377 = n11376 ^ x4 ^ 1'b0 ;
  assign n11378 = n11372 & n11377 ;
  assign n11379 = n11378 ^ n4897 ^ n1915 ;
  assign n11380 = ~n6093 & n11379 ;
  assign n11381 = n11380 ^ n2850 ^ 1'b0 ;
  assign n11383 = n2797 ^ n1848 ^ n1362 ;
  assign n11384 = n11383 ^ n7402 ^ n2163 ;
  assign n11385 = ( n2845 & n3885 ) | ( n2845 & n11384 ) | ( n3885 & n11384 ) ;
  assign n11382 = n6074 ^ n2038 ^ 1'b0 ;
  assign n11386 = n11385 ^ n11382 ^ n4068 ;
  assign n11387 = n1480 & n6400 ;
  assign n11388 = n6221 ^ n6079 ^ n4366 ;
  assign n11389 = ~n304 & n11388 ;
  assign n11390 = ( n5410 & n6659 ) | ( n5410 & ~n11389 ) | ( n6659 & ~n11389 ) ;
  assign n11391 = n4594 & n5190 ;
  assign n11392 = n1871 & n11391 ;
  assign n11393 = ( n6087 & ~n6273 ) | ( n6087 & n11392 ) | ( ~n6273 & n11392 ) ;
  assign n11394 = ~n11390 & n11393 ;
  assign n11395 = n11394 ^ x42 ^ 1'b0 ;
  assign n11397 = n1185 ^ n636 ^ 1'b0 ;
  assign n11396 = n2746 | n6517 ;
  assign n11398 = n11397 ^ n11396 ^ 1'b0 ;
  assign n11400 = n3752 ^ n2021 ^ n716 ;
  assign n11399 = x78 & ~n4641 ;
  assign n11401 = n11400 ^ n11399 ^ 1'b0 ;
  assign n11402 = n4392 ^ n2183 ^ 1'b0 ;
  assign n11403 = ~n11401 & n11402 ;
  assign n11404 = n1233 & ~n3601 ;
  assign n11405 = ( n5596 & n6910 ) | ( n5596 & n11404 ) | ( n6910 & n11404 ) ;
  assign n11406 = ( n1517 & ~n6692 ) | ( n1517 & n8732 ) | ( ~n6692 & n8732 ) ;
  assign n11408 = n9432 ^ n4462 ^ 1'b0 ;
  assign n11407 = n3118 & ~n6282 ;
  assign n11409 = n11408 ^ n11407 ^ 1'b0 ;
  assign n11410 = n11406 & ~n11409 ;
  assign n11423 = ( n474 & n4659 ) | ( n474 & ~n5576 ) | ( n4659 & ~n5576 ) ;
  assign n11420 = n5878 & n9521 ;
  assign n11421 = n11420 ^ n9514 ^ 1'b0 ;
  assign n11416 = n2996 & n9709 ;
  assign n11417 = n11416 ^ n1856 ^ 1'b0 ;
  assign n11418 = n9443 ^ n5187 ^ n1269 ;
  assign n11419 = n11417 | n11418 ;
  assign n11422 = n11421 ^ n11419 ^ 1'b0 ;
  assign n11424 = n11423 ^ n11422 ^ 1'b0 ;
  assign n11411 = n7521 ^ n6223 ^ n1882 ;
  assign n11412 = n2807 ^ n1376 ^ n653 ;
  assign n11413 = n2633 & n11412 ;
  assign n11414 = n11413 ^ n8261 ^ 1'b0 ;
  assign n11415 = ( ~n936 & n11411 ) | ( ~n936 & n11414 ) | ( n11411 & n11414 ) ;
  assign n11425 = n11424 ^ n11415 ^ n11332 ;
  assign n11426 = ( n3245 & ~n7416 ) | ( n3245 & n10589 ) | ( ~n7416 & n10589 ) ;
  assign n11427 = n11426 ^ n8475 ^ 1'b0 ;
  assign n11434 = ( x167 & ~n357 ) | ( x167 & n9601 ) | ( ~n357 & n9601 ) ;
  assign n11428 = n3611 | n3786 ;
  assign n11429 = n11428 ^ n2449 ^ 1'b0 ;
  assign n11430 = n9301 ^ n4241 ^ n3956 ;
  assign n11431 = ~n4332 & n11430 ;
  assign n11432 = n11431 ^ n2987 ^ 1'b0 ;
  assign n11433 = ( n2589 & n11429 ) | ( n2589 & ~n11432 ) | ( n11429 & ~n11432 ) ;
  assign n11435 = n11434 ^ n11433 ^ n6968 ;
  assign n11436 = n366 | n11241 ;
  assign n11437 = n11436 ^ n1948 ^ 1'b0 ;
  assign n11438 = n11437 ^ n2341 ^ 1'b0 ;
  assign n11439 = n4015 | n11438 ;
  assign n11440 = ( n1691 & n3429 ) | ( n1691 & n9441 ) | ( n3429 & n9441 ) ;
  assign n11441 = ~n2957 & n3341 ;
  assign n11442 = ~n3795 & n11441 ;
  assign n11443 = n11442 ^ n7715 ^ n5090 ;
  assign n11444 = ( n8733 & ~n11440 ) | ( n8733 & n11443 ) | ( ~n11440 & n11443 ) ;
  assign n11445 = ( ~x248 & n9881 ) | ( ~x248 & n10683 ) | ( n9881 & n10683 ) ;
  assign n11446 = n2901 & n8842 ;
  assign n11447 = n7234 ^ n3092 ^ n681 ;
  assign n11450 = n9499 ^ n2252 ^ n438 ;
  assign n11448 = n9314 ^ n7566 ^ n1752 ;
  assign n11449 = n1896 | n11448 ;
  assign n11451 = n11450 ^ n11449 ^ 1'b0 ;
  assign n11452 = n11447 & n11451 ;
  assign n11453 = n2022 & n11452 ;
  assign n11460 = n300 | n1766 ;
  assign n11461 = n3919 | n11460 ;
  assign n11462 = n11461 ^ n3245 ^ 1'b0 ;
  assign n11454 = n3204 | n3810 ;
  assign n11455 = n11454 ^ n2208 ^ 1'b0 ;
  assign n11456 = n8062 ^ n5799 ^ n898 ;
  assign n11457 = n5666 & n11456 ;
  assign n11458 = ~n11455 & n11457 ;
  assign n11459 = n3051 & n11458 ;
  assign n11463 = n11462 ^ n11459 ^ n6993 ;
  assign n11464 = n10460 ^ n4721 ^ n339 ;
  assign n11468 = ( n1627 & ~n9144 ) | ( n1627 & n10928 ) | ( ~n9144 & n10928 ) ;
  assign n11469 = n2679 | n11468 ;
  assign n11470 = n11469 ^ n4338 ^ 1'b0 ;
  assign n11471 = n11470 ^ n9056 ^ n8372 ;
  assign n11465 = n4496 & ~n10955 ;
  assign n11466 = n3947 & n11465 ;
  assign n11467 = n801 & n11466 ;
  assign n11472 = n11471 ^ n11467 ^ 1'b0 ;
  assign n11473 = n11472 ^ n10242 ^ n1231 ;
  assign n11477 = n2381 ^ n891 ^ 1'b0 ;
  assign n11476 = n1966 ^ n1499 ^ n1244 ;
  assign n11474 = n1552 & ~n4523 ;
  assign n11475 = ~x196 & n11474 ;
  assign n11478 = n11477 ^ n11476 ^ n11475 ;
  assign n11479 = ( n3416 & n8077 ) | ( n3416 & ~n11478 ) | ( n8077 & ~n11478 ) ;
  assign n11480 = ~n9828 & n11479 ;
  assign n11482 = n4626 & ~n10818 ;
  assign n11483 = n5695 & n11482 ;
  assign n11481 = n6481 ^ n3799 ^ n2356 ;
  assign n11484 = n11483 ^ n11481 ^ n3699 ;
  assign n11485 = n9598 ^ n4334 ^ 1'b0 ;
  assign n11486 = n941 | n5293 ;
  assign n11487 = n2451 & ~n11486 ;
  assign n11488 = n11285 ^ n2064 ^ 1'b0 ;
  assign n11489 = n11487 | n11488 ;
  assign n11493 = ( n2224 & ~n2425 ) | ( n2224 & n3460 ) | ( ~n2425 & n3460 ) ;
  assign n11494 = ( ~n1204 & n2054 ) | ( ~n1204 & n9294 ) | ( n2054 & n9294 ) ;
  assign n11495 = n11494 ^ n870 ^ 1'b0 ;
  assign n11496 = n11493 | n11495 ;
  assign n11491 = n2088 ^ n882 ^ 1'b0 ;
  assign n11490 = n1323 & ~n3608 ;
  assign n11492 = n11491 ^ n11490 ^ 1'b0 ;
  assign n11497 = n11496 ^ n11492 ^ n544 ;
  assign n11498 = n11497 ^ n9405 ^ 1'b0 ;
  assign n11499 = n1661 ^ n684 ^ n537 ;
  assign n11500 = ~n7622 & n11499 ;
  assign n11501 = n11500 ^ n6434 ^ 1'b0 ;
  assign n11502 = n2059 & ~n8612 ;
  assign n11503 = ~n11501 & n11502 ;
  assign n11512 = ~n395 & n10356 ;
  assign n11513 = n2751 & n11512 ;
  assign n11504 = ( n1712 & ~n8349 ) | ( n1712 & n8400 ) | ( ~n8349 & n8400 ) ;
  assign n11505 = n6424 ^ n2535 ^ n481 ;
  assign n11506 = n3820 ^ n3190 ^ 1'b0 ;
  assign n11507 = n11506 ^ n9299 ^ n5922 ;
  assign n11508 = n4736 & ~n11507 ;
  assign n11509 = n11508 ^ n7068 ^ 1'b0 ;
  assign n11510 = n11505 & n11509 ;
  assign n11511 = n11504 & n11510 ;
  assign n11514 = n11513 ^ n11511 ^ 1'b0 ;
  assign n11515 = ~n11503 & n11514 ;
  assign n11517 = n2913 ^ n2378 ^ 1'b0 ;
  assign n11518 = n10478 & ~n11517 ;
  assign n11516 = ( ~n263 & n6708 ) | ( ~n263 & n8659 ) | ( n6708 & n8659 ) ;
  assign n11519 = n11518 ^ n11516 ^ n2875 ;
  assign n11520 = n4641 ^ n3548 ^ n1344 ;
  assign n11521 = n10591 & ~n11520 ;
  assign n11522 = n5492 & n11521 ;
  assign n11525 = n3508 ^ n2809 ^ 1'b0 ;
  assign n11526 = n9533 | n11525 ;
  assign n11524 = ( n3320 & ~n4120 ) | ( n3320 & n4709 ) | ( ~n4120 & n4709 ) ;
  assign n11527 = n11526 ^ n11524 ^ n3800 ;
  assign n11523 = n353 & n6845 ;
  assign n11528 = n11527 ^ n11523 ^ 1'b0 ;
  assign n11529 = n5461 ^ n2778 ^ n914 ;
  assign n11530 = n11529 ^ n6331 ^ n574 ;
  assign n11531 = n11530 ^ n4997 ^ n3249 ;
  assign n11532 = n10795 ^ n10400 ^ n9750 ;
  assign n11533 = n7364 ^ n1107 ^ n367 ;
  assign n11534 = n1077 & ~n11533 ;
  assign n11535 = n6351 & ~n11534 ;
  assign n11536 = n7372 & n11535 ;
  assign n11537 = n2661 & ~n11536 ;
  assign n11538 = n11537 ^ n4502 ^ 1'b0 ;
  assign n11539 = ( n381 & n3639 ) | ( n381 & n5523 ) | ( n3639 & n5523 ) ;
  assign n11540 = n3276 & n8584 ;
  assign n11541 = n9173 & ~n11540 ;
  assign n11542 = n11541 ^ n10189 ^ 1'b0 ;
  assign n11543 = ( n904 & n2801 ) | ( n904 & n3973 ) | ( n2801 & n3973 ) ;
  assign n11544 = n4408 | n11543 ;
  assign n11545 = n4744 | n11544 ;
  assign n11546 = n11545 ^ n11492 ^ n5440 ;
  assign n11547 = n11209 ^ n11004 ^ n10232 ;
  assign n11548 = n9560 & ~n11547 ;
  assign n11549 = ~n7994 & n11548 ;
  assign n11550 = ~n1593 & n11549 ;
  assign n11551 = n535 | n5665 ;
  assign n11552 = n962 & ~n11551 ;
  assign n11558 = n3703 ^ n1261 ^ n1087 ;
  assign n11553 = n983 ^ n489 ^ n343 ;
  assign n11554 = n1983 ^ n356 ^ 1'b0 ;
  assign n11555 = n1548 & ~n11554 ;
  assign n11556 = ~n6169 & n11555 ;
  assign n11557 = n11553 & ~n11556 ;
  assign n11559 = n11558 ^ n11557 ^ 1'b0 ;
  assign n11560 = n6455 & n10364 ;
  assign n11561 = n11560 ^ n9749 ^ n1842 ;
  assign n11563 = ( n802 & n3870 ) | ( n802 & ~n4362 ) | ( n3870 & ~n4362 ) ;
  assign n11562 = n2473 & n5530 ;
  assign n11564 = n11563 ^ n11562 ^ 1'b0 ;
  assign n11565 = n11564 ^ n4537 ^ 1'b0 ;
  assign n11566 = ( n790 & ~n8083 ) | ( n790 & n11565 ) | ( ~n8083 & n11565 ) ;
  assign n11567 = n4537 ^ n1188 ^ 1'b0 ;
  assign n11574 = n3342 ^ n2278 ^ 1'b0 ;
  assign n11575 = n570 | n11574 ;
  assign n11571 = x117 & ~n9212 ;
  assign n11572 = n3327 & n11571 ;
  assign n11568 = ~n5626 & n8062 ;
  assign n11569 = n11568 ^ n702 ^ 1'b0 ;
  assign n11570 = n8862 & ~n11569 ;
  assign n11573 = n11572 ^ n11570 ^ 1'b0 ;
  assign n11576 = n11575 ^ n11573 ^ n6199 ;
  assign n11577 = ( n5188 & n6716 ) | ( n5188 & n7056 ) | ( n6716 & n7056 ) ;
  assign n11578 = ( n11567 & ~n11576 ) | ( n11567 & n11577 ) | ( ~n11576 & n11577 ) ;
  assign n11579 = n1256 & n11578 ;
  assign n11580 = n7494 ^ n934 ^ 1'b0 ;
  assign n11581 = n6076 | n11580 ;
  assign n11582 = n7388 & ~n11581 ;
  assign n11583 = n6668 ^ n4423 ^ 1'b0 ;
  assign n11584 = n9613 | n11583 ;
  assign n11585 = n6697 ^ n6117 ^ 1'b0 ;
  assign n11586 = ( n1532 & n6505 ) | ( n1532 & n11585 ) | ( n6505 & n11585 ) ;
  assign n11587 = ( ~n4033 & n4067 ) | ( ~n4033 & n4510 ) | ( n4067 & n4510 ) ;
  assign n11588 = ( n5802 & n6456 ) | ( n5802 & ~n11587 ) | ( n6456 & ~n11587 ) ;
  assign n11589 = n1897 ^ n997 ^ 1'b0 ;
  assign n11590 = n2301 & ~n11589 ;
  assign n11591 = n10688 ^ n2890 ^ n2843 ;
  assign n11592 = ( ~n3108 & n4472 ) | ( ~n3108 & n11591 ) | ( n4472 & n11591 ) ;
  assign n11593 = n4640 & n11592 ;
  assign n11594 = ~n11590 & n11593 ;
  assign n11598 = x124 & ~n5471 ;
  assign n11599 = n11598 ^ n4531 ^ 1'b0 ;
  assign n11595 = x174 & ~n11049 ;
  assign n11596 = ~n3989 & n11595 ;
  assign n11597 = n11596 ^ n10609 ^ n9746 ;
  assign n11600 = n11599 ^ n11597 ^ n9128 ;
  assign n11601 = ( n3918 & n6507 ) | ( n3918 & n7341 ) | ( n6507 & n7341 ) ;
  assign n11602 = n2875 ^ n735 ^ 1'b0 ;
  assign n11610 = n7298 ^ x251 ^ 1'b0 ;
  assign n11611 = n7821 & ~n11610 ;
  assign n11612 = n11611 ^ x62 ^ 1'b0 ;
  assign n11609 = x21 & ~n635 ;
  assign n11607 = n3132 | n5358 ;
  assign n11603 = n731 ^ x238 ^ x164 ;
  assign n11604 = n5391 & n11603 ;
  assign n11605 = n6698 & n11604 ;
  assign n11606 = n8765 & ~n11605 ;
  assign n11608 = n11607 ^ n11606 ^ 1'b0 ;
  assign n11613 = n11612 ^ n11609 ^ n11608 ;
  assign n11615 = ( n1029 & n2088 ) | ( n1029 & n3872 ) | ( n2088 & n3872 ) ;
  assign n11614 = ( n705 & n3922 ) | ( n705 & n10335 ) | ( n3922 & n10335 ) ;
  assign n11616 = n11615 ^ n11614 ^ n10115 ;
  assign n11617 = ( n2103 & n2948 ) | ( n2103 & n3303 ) | ( n2948 & n3303 ) ;
  assign n11620 = n6616 ^ n1903 ^ n418 ;
  assign n11618 = n8116 ^ n3647 ^ 1'b0 ;
  assign n11619 = n1953 & ~n11618 ;
  assign n11621 = n11620 ^ n11619 ^ n8203 ;
  assign n11622 = ( n4782 & n11617 ) | ( n4782 & ~n11621 ) | ( n11617 & ~n11621 ) ;
  assign n11623 = ~n459 & n6465 ;
  assign n11624 = ~n2226 & n11623 ;
  assign n11628 = n5635 & ~n5912 ;
  assign n11629 = n11628 ^ n3189 ^ 1'b0 ;
  assign n11627 = n2856 & ~n4152 ;
  assign n11630 = n11629 ^ n11627 ^ 1'b0 ;
  assign n11631 = n11630 ^ n5374 ^ n415 ;
  assign n11625 = ( n3429 & n3490 ) | ( n3429 & n11147 ) | ( n3490 & n11147 ) ;
  assign n11626 = ( n8726 & n9614 ) | ( n8726 & ~n11625 ) | ( n9614 & ~n11625 ) ;
  assign n11632 = n11631 ^ n11626 ^ n4372 ;
  assign n11633 = ( n845 & n6755 ) | ( n845 & n9472 ) | ( n6755 & n9472 ) ;
  assign n11634 = n5619 & ~n11633 ;
  assign n11635 = n11634 ^ n3668 ^ x202 ;
  assign n11636 = ( n1264 & n1745 ) | ( n1264 & n5820 ) | ( n1745 & n5820 ) ;
  assign n11637 = n11636 ^ n3724 ^ n2182 ;
  assign n11638 = n2179 & n11637 ;
  assign n11639 = n11638 ^ n1840 ^ 1'b0 ;
  assign n11640 = ( n4634 & ~n9219 ) | ( n4634 & n11639 ) | ( ~n9219 & n11639 ) ;
  assign n11641 = n7035 & n11640 ;
  assign n11642 = n4405 ^ n840 ^ 1'b0 ;
  assign n11643 = n11126 ^ n7570 ^ n987 ;
  assign n11644 = n9085 ^ n3817 ^ 1'b0 ;
  assign n11645 = ~n11643 & n11644 ;
  assign n11646 = n11645 ^ n2252 ^ 1'b0 ;
  assign n11647 = n6359 & ~n11646 ;
  assign n11648 = n11647 ^ n3056 ^ 1'b0 ;
  assign n11649 = n11642 & n11648 ;
  assign n11650 = n1538 & n6785 ;
  assign n11651 = n11650 ^ n933 ^ 1'b0 ;
  assign n11652 = ~n5685 & n11651 ;
  assign n11655 = n3361 ^ n994 ^ 1'b0 ;
  assign n11656 = ~n3925 & n11655 ;
  assign n11657 = ( ~n287 & n2626 ) | ( ~n287 & n11656 ) | ( n2626 & n11656 ) ;
  assign n11658 = ( ~n2786 & n4905 ) | ( ~n2786 & n11657 ) | ( n4905 & n11657 ) ;
  assign n11659 = n705 & n11658 ;
  assign n11660 = ~n2558 & n11659 ;
  assign n11653 = ( x146 & n4482 ) | ( x146 & ~n6331 ) | ( n4482 & ~n6331 ) ;
  assign n11654 = n805 & ~n11653 ;
  assign n11661 = n11660 ^ n11654 ^ 1'b0 ;
  assign n11662 = ~n11652 & n11661 ;
  assign n11663 = n8871 & n10622 ;
  assign n11664 = n4100 ^ n3249 ^ n1309 ;
  assign n11665 = n1418 ^ n785 ^ n326 ;
  assign n11666 = n11665 ^ n3710 ^ 1'b0 ;
  assign n11667 = n11664 & ~n11666 ;
  assign n11668 = ( ~n4351 & n8963 ) | ( ~n4351 & n11667 ) | ( n8963 & n11667 ) ;
  assign n11672 = n1416 & n9385 ;
  assign n11673 = n4257 & n11672 ;
  assign n11674 = ~n3817 & n6474 ;
  assign n11675 = n11673 & n11674 ;
  assign n11671 = ~n3629 & n10643 ;
  assign n11676 = n11675 ^ n11671 ^ 1'b0 ;
  assign n11669 = n1947 & n4744 ;
  assign n11670 = n11669 ^ n6329 ^ n3317 ;
  assign n11677 = n11676 ^ n11670 ^ n7910 ;
  assign n11684 = n2510 & ~n5484 ;
  assign n11685 = n1884 & ~n2516 ;
  assign n11686 = n11684 & n11685 ;
  assign n11681 = n696 ^ x33 ^ 1'b0 ;
  assign n11682 = ~n796 & n11681 ;
  assign n11678 = n1243 ^ n637 ^ n542 ;
  assign n11679 = ( x65 & n939 ) | ( x65 & n11678 ) | ( n939 & n11678 ) ;
  assign n11680 = n11679 ^ n2017 ^ n1120 ;
  assign n11683 = n11682 ^ n11680 ^ n2606 ;
  assign n11687 = n11686 ^ n11683 ^ n5617 ;
  assign n11689 = ( ~n2452 & n3254 ) | ( ~n2452 & n4661 ) | ( n3254 & n4661 ) ;
  assign n11690 = n11689 ^ n6925 ^ n3048 ;
  assign n11688 = n10090 ^ n1730 ^ 1'b0 ;
  assign n11691 = n11690 ^ n11688 ^ n3455 ;
  assign n11692 = n2162 ^ n2122 ^ x109 ;
  assign n11693 = n11692 ^ n3363 ^ 1'b0 ;
  assign n11696 = n321 & ~n4993 ;
  assign n11694 = ( n1070 & n2181 ) | ( n1070 & ~n2213 ) | ( n2181 & ~n2213 ) ;
  assign n11695 = n11694 ^ n8850 ^ n8337 ;
  assign n11697 = n11696 ^ n11695 ^ n9716 ;
  assign n11698 = ( n7881 & n11693 ) | ( n7881 & ~n11697 ) | ( n11693 & ~n11697 ) ;
  assign n11699 = ( n2904 & n5754 ) | ( n2904 & n10723 ) | ( n5754 & n10723 ) ;
  assign n11700 = n9729 & n11699 ;
  assign n11702 = n2427 ^ n2096 ^ n786 ;
  assign n11703 = n11702 ^ n5412 ^ x163 ;
  assign n11701 = n7600 | n8184 ;
  assign n11704 = n11703 ^ n11701 ^ 1'b0 ;
  assign n11705 = n7523 | n11704 ;
  assign n11706 = n4482 | n6271 ;
  assign n11707 = ( n6237 & n9208 ) | ( n6237 & n11706 ) | ( n9208 & n11706 ) ;
  assign n11708 = n2455 & n3035 ;
  assign n11709 = ~n2463 & n11708 ;
  assign n11710 = n1309 & ~n11709 ;
  assign n11711 = ( n478 & n4202 ) | ( n478 & n10481 ) | ( n4202 & n10481 ) ;
  assign n11712 = n11711 ^ n5761 ^ n2770 ;
  assign n11714 = n2216 ^ n1404 ^ 1'b0 ;
  assign n11715 = n557 & n11714 ;
  assign n11713 = n9105 ^ n9050 ^ n1058 ;
  assign n11716 = n11715 ^ n11713 ^ n1078 ;
  assign n11718 = n2774 | n3190 ;
  assign n11719 = ( ~n5209 & n7551 ) | ( ~n5209 & n11718 ) | ( n7551 & n11718 ) ;
  assign n11717 = n4959 | n11389 ;
  assign n11720 = n11719 ^ n11717 ^ 1'b0 ;
  assign n11725 = n1279 ^ n913 ^ n312 ;
  assign n11721 = n3058 & ~n5636 ;
  assign n11722 = n11721 ^ n10441 ^ n3725 ;
  assign n11723 = ~n809 & n11722 ;
  assign n11724 = n11723 ^ n5082 ^ 1'b0 ;
  assign n11726 = n11725 ^ n11724 ^ n8306 ;
  assign n11727 = n6698 ^ n1285 ^ 1'b0 ;
  assign n11728 = ~n3820 & n11727 ;
  assign n11729 = n1137 & n2418 ;
  assign n11730 = n11729 ^ n8534 ^ 1'b0 ;
  assign n11731 = ( n11726 & n11728 ) | ( n11726 & ~n11730 ) | ( n11728 & ~n11730 ) ;
  assign n11732 = n492 & n7783 ;
  assign n11733 = n5213 & n11732 ;
  assign n11734 = n4223 ^ n4080 ^ 1'b0 ;
  assign n11735 = x129 & ~n3752 ;
  assign n11736 = n1119 & n11735 ;
  assign n11737 = n5496 ^ n865 ^ n425 ;
  assign n11738 = ~n4083 & n5566 ;
  assign n11739 = n11737 & n11738 ;
  assign n11740 = n9432 ^ n3072 ^ 1'b0 ;
  assign n11741 = n11739 | n11740 ;
  assign n11742 = n11736 & ~n11741 ;
  assign n11743 = ( n1421 & n2590 ) | ( n1421 & ~n11742 ) | ( n2590 & ~n11742 ) ;
  assign n11744 = ( ~n6850 & n11734 ) | ( ~n6850 & n11743 ) | ( n11734 & n11743 ) ;
  assign n11745 = n4177 ^ n2732 ^ n2192 ;
  assign n11746 = ~n11580 & n11745 ;
  assign n11747 = n11746 ^ n3929 ^ 1'b0 ;
  assign n11757 = n5794 ^ n3706 ^ 1'b0 ;
  assign n11755 = n5602 & n7868 ;
  assign n11756 = n11755 ^ n10504 ^ 1'b0 ;
  assign n11750 = ( n1372 & ~n1717 ) | ( n1372 & n7473 ) | ( ~n1717 & n7473 ) ;
  assign n11751 = n5856 & ~n11750 ;
  assign n11748 = ( n2193 & n6058 ) | ( n2193 & ~n6417 ) | ( n6058 & ~n6417 ) ;
  assign n11749 = n5566 & n11748 ;
  assign n11752 = n11751 ^ n11749 ^ 1'b0 ;
  assign n11753 = n3432 & n4509 ;
  assign n11754 = ~n11752 & n11753 ;
  assign n11758 = n11757 ^ n11756 ^ n11754 ;
  assign n11759 = ( ~n7720 & n11747 ) | ( ~n7720 & n11758 ) | ( n11747 & n11758 ) ;
  assign n11760 = n3424 ^ n2186 ^ n706 ;
  assign n11761 = n4630 & ~n4987 ;
  assign n11762 = ~n1903 & n11761 ;
  assign n11763 = n3866 | n11762 ;
  assign n11764 = n11760 | n11763 ;
  assign n11765 = ( n570 & ~n6678 ) | ( n570 & n7009 ) | ( ~n6678 & n7009 ) ;
  assign n11766 = ( n2708 & n5224 ) | ( n2708 & n11097 ) | ( n5224 & n11097 ) ;
  assign n11767 = n8423 | n11766 ;
  assign n11768 = n11767 ^ x30 ^ 1'b0 ;
  assign n11769 = ( n1622 & n6704 ) | ( n1622 & ~n11768 ) | ( n6704 & ~n11768 ) ;
  assign n11770 = ( n4239 & n6280 ) | ( n4239 & ~n11769 ) | ( n6280 & ~n11769 ) ;
  assign n11771 = ( ~x58 & n6250 ) | ( ~x58 & n11167 ) | ( n6250 & n11167 ) ;
  assign n11773 = ( n2926 & n5261 ) | ( n2926 & n11750 ) | ( n5261 & n11750 ) ;
  assign n11772 = ( n259 & n2463 ) | ( n259 & ~n3691 ) | ( n2463 & ~n3691 ) ;
  assign n11774 = n11773 ^ n11772 ^ x216 ;
  assign n11775 = ( n1643 & ~n3525 ) | ( n1643 & n11774 ) | ( ~n3525 & n11774 ) ;
  assign n11776 = n11775 ^ n7423 ^ 1'b0 ;
  assign n11777 = n8978 ^ n8714 ^ 1'b0 ;
  assign n11778 = n11777 ^ n5067 ^ n4036 ;
  assign n11779 = ( n1016 & n2556 ) | ( n1016 & n3040 ) | ( n2556 & n3040 ) ;
  assign n11781 = n1384 ^ n1198 ^ x23 ;
  assign n11780 = n580 & ~n5832 ;
  assign n11782 = n11781 ^ n11780 ^ n4563 ;
  assign n11783 = ( n11230 & ~n11779 ) | ( n11230 & n11782 ) | ( ~n11779 & n11782 ) ;
  assign n11789 = n11188 ^ n2822 ^ n1464 ;
  assign n11790 = x46 | n11789 ;
  assign n11784 = n3724 & n9800 ;
  assign n11785 = ( n813 & ~n4710 ) | ( n813 & n11784 ) | ( ~n4710 & n11784 ) ;
  assign n11786 = n1368 & n5686 ;
  assign n11787 = n11785 & n11786 ;
  assign n11788 = n2133 | n11787 ;
  assign n11791 = n11790 ^ n11788 ^ 1'b0 ;
  assign n11792 = ( n1071 & n5802 ) | ( n1071 & n11343 ) | ( n5802 & n11343 ) ;
  assign n11793 = n2161 | n11792 ;
  assign n11794 = n8010 ^ n1372 ^ 1'b0 ;
  assign n11795 = ( n1343 & n4940 ) | ( n1343 & n5401 ) | ( n4940 & n5401 ) ;
  assign n11796 = n11794 & n11795 ;
  assign n11797 = n7946 ^ n7556 ^ n4789 ;
  assign n11798 = n4273 ^ n593 ^ 1'b0 ;
  assign n11799 = ( n1267 & n2228 ) | ( n1267 & n11798 ) | ( n2228 & n11798 ) ;
  assign n11800 = ( n2026 & ~n11797 ) | ( n2026 & n11799 ) | ( ~n11797 & n11799 ) ;
  assign n11801 = n11800 ^ n541 ^ 1'b0 ;
  assign n11802 = n7566 ^ n500 ^ 1'b0 ;
  assign n11803 = n11802 ^ n9629 ^ n8247 ;
  assign n11804 = ( ~n327 & n8327 ) | ( ~n327 & n11803 ) | ( n8327 & n11803 ) ;
  assign n11805 = n10115 | n11804 ;
  assign n11806 = n11805 ^ n4257 ^ 1'b0 ;
  assign n11807 = n5934 & n9558 ;
  assign n11808 = ~n7754 & n11807 ;
  assign n11810 = n1940 ^ n571 ^ 1'b0 ;
  assign n11809 = n3267 | n10287 ;
  assign n11811 = n11810 ^ n11809 ^ 1'b0 ;
  assign n11812 = n11811 ^ n1339 ^ 1'b0 ;
  assign n11813 = ~n3860 & n11812 ;
  assign n11814 = n11813 ^ n1879 ^ 1'b0 ;
  assign n11815 = n6645 & n11814 ;
  assign n11816 = n592 & ~n1055 ;
  assign n11817 = n11816 ^ n7653 ^ n5831 ;
  assign n11818 = ~n11768 & n11817 ;
  assign n11819 = ( n2960 & n11343 ) | ( n2960 & n11818 ) | ( n11343 & n11818 ) ;
  assign n11820 = n8537 ^ n8389 ^ n1944 ;
  assign n11821 = n5918 ^ n2997 ^ n2150 ;
  assign n11822 = ( n1629 & n7722 ) | ( n1629 & ~n11821 ) | ( n7722 & ~n11821 ) ;
  assign n11823 = ( n8588 & ~n11820 ) | ( n8588 & n11822 ) | ( ~n11820 & n11822 ) ;
  assign n11824 = ~n727 & n1569 ;
  assign n11825 = n11824 ^ n3603 ^ n3487 ;
  assign n11826 = n6523 ^ n2278 ^ n1066 ;
  assign n11827 = n10016 ^ n9088 ^ x13 ;
  assign n11828 = ( n10741 & n11826 ) | ( n10741 & ~n11827 ) | ( n11826 & ~n11827 ) ;
  assign n11829 = n11825 & n11828 ;
  assign n11830 = n11829 ^ n9075 ^ 1'b0 ;
  assign n11831 = n10879 ^ n6036 ^ 1'b0 ;
  assign n11832 = ( ~n799 & n6770 ) | ( ~n799 & n7428 ) | ( n6770 & n7428 ) ;
  assign n11833 = ( n2345 & n10493 ) | ( n2345 & ~n11832 ) | ( n10493 & ~n11832 ) ;
  assign n11834 = n11833 ^ n11201 ^ 1'b0 ;
  assign n11835 = ~n11831 & n11834 ;
  assign n11836 = n11835 ^ n1794 ^ n1418 ;
  assign n11843 = n2577 | n8308 ;
  assign n11837 = ( ~n1056 & n3868 ) | ( ~n1056 & n4554 ) | ( n3868 & n4554 ) ;
  assign n11838 = n9525 ^ n1735 ^ n1323 ;
  assign n11839 = ( n548 & n6182 ) | ( n548 & ~n11838 ) | ( n6182 & ~n11838 ) ;
  assign n11840 = ( n3725 & ~n11837 ) | ( n3725 & n11839 ) | ( ~n11837 & n11839 ) ;
  assign n11841 = ~n4234 & n11840 ;
  assign n11842 = n11841 ^ n6821 ^ 1'b0 ;
  assign n11844 = n11843 ^ n11842 ^ n3675 ;
  assign n11845 = n508 ^ x120 ^ 1'b0 ;
  assign n11846 = n8674 | n11845 ;
  assign n11847 = n8223 & ~n11846 ;
  assign n11848 = x78 & n9131 ;
  assign n11849 = n2851 ^ n2345 ^ n1402 ;
  assign n11856 = n4325 ^ n3379 ^ n478 ;
  assign n11853 = n3449 ^ n811 ^ 1'b0 ;
  assign n11854 = ~n1436 & n11853 ;
  assign n11855 = n11854 ^ n8548 ^ n3482 ;
  assign n11850 = n1625 | n2255 ;
  assign n11851 = n11850 ^ n1693 ^ 1'b0 ;
  assign n11852 = ( n7910 & n8306 ) | ( n7910 & ~n11851 ) | ( n8306 & ~n11851 ) ;
  assign n11857 = n11856 ^ n11855 ^ n11852 ;
  assign n11858 = ( n1363 & n6301 ) | ( n1363 & ~n6615 ) | ( n6301 & ~n6615 ) ;
  assign n11859 = n11858 ^ n4211 ^ n3076 ;
  assign n11860 = n8561 ^ n6994 ^ n870 ;
  assign n11861 = n1365 & ~n11860 ;
  assign n11862 = n2755 & n11861 ;
  assign n11863 = n11862 ^ n6136 ^ n5269 ;
  assign n11864 = n4507 & n11863 ;
  assign n11865 = n11864 ^ n1019 ^ 1'b0 ;
  assign n11867 = n6546 ^ n1115 ^ 1'b0 ;
  assign n11868 = n7829 & ~n11867 ;
  assign n11866 = ~n2245 & n2254 ;
  assign n11869 = n11868 ^ n11866 ^ 1'b0 ;
  assign n11870 = n8378 ^ n6919 ^ 1'b0 ;
  assign n11871 = n2584 ^ n1373 ^ n312 ;
  assign n11872 = n9232 ^ n5009 ^ 1'b0 ;
  assign n11873 = n11871 & n11872 ;
  assign n11874 = ( n8799 & n11870 ) | ( n8799 & ~n11873 ) | ( n11870 & ~n11873 ) ;
  assign n11875 = n784 & n2263 ;
  assign n11876 = ( n4649 & n8979 ) | ( n4649 & ~n11875 ) | ( n8979 & ~n11875 ) ;
  assign n11877 = n11876 ^ n10642 ^ 1'b0 ;
  assign n11878 = ( x204 & ~n10775 ) | ( x204 & n11577 ) | ( ~n10775 & n11577 ) ;
  assign n11879 = n6586 ^ n2861 ^ x253 ;
  assign n11880 = n1609 & ~n10326 ;
  assign n11881 = n11880 ^ n4621 ^ 1'b0 ;
  assign n11882 = n11879 & n11881 ;
  assign n11895 = n2091 ^ n353 ^ x254 ;
  assign n11896 = n6166 | n11895 ;
  assign n11893 = n10001 ^ n7609 ^ x30 ;
  assign n11891 = ( x44 & n1210 ) | ( x44 & n7539 ) | ( n1210 & n7539 ) ;
  assign n11892 = n11891 ^ n7740 ^ n4338 ;
  assign n11894 = n11893 ^ n11892 ^ n6314 ;
  assign n11888 = n3840 ^ n2283 ^ 1'b0 ;
  assign n11889 = n10875 | n11888 ;
  assign n11883 = ( n3769 & ~n7367 ) | ( n3769 & n8212 ) | ( ~n7367 & n8212 ) ;
  assign n11884 = ( n1879 & n3441 ) | ( n1879 & n7592 ) | ( n3441 & n7592 ) ;
  assign n11885 = n11884 ^ n7262 ^ 1'b0 ;
  assign n11886 = n11883 & ~n11885 ;
  assign n11887 = n2181 & n11886 ;
  assign n11890 = n11889 ^ n11887 ^ 1'b0 ;
  assign n11897 = n11896 ^ n11894 ^ n11890 ;
  assign n11898 = ( n11878 & n11882 ) | ( n11878 & n11897 ) | ( n11882 & n11897 ) ;
  assign n11899 = ( ~n1292 & n3721 ) | ( ~n1292 & n9763 ) | ( n3721 & n9763 ) ;
  assign n11900 = ( n474 & ~n2780 ) | ( n474 & n11899 ) | ( ~n2780 & n11899 ) ;
  assign n11901 = ( n3126 & n3149 ) | ( n3126 & ~n6825 ) | ( n3149 & ~n6825 ) ;
  assign n11902 = n11901 ^ n11586 ^ 1'b0 ;
  assign n11903 = ~n7327 & n11902 ;
  assign n11904 = ( n547 & n1398 ) | ( n547 & ~n4352 ) | ( n1398 & ~n4352 ) ;
  assign n11905 = ( n6923 & n7847 ) | ( n6923 & n9775 ) | ( n7847 & n9775 ) ;
  assign n11906 = ( n3304 & n11904 ) | ( n3304 & n11905 ) | ( n11904 & n11905 ) ;
  assign n11907 = n10335 ^ n1031 ^ 1'b0 ;
  assign n11908 = n11907 ^ n531 ^ 1'b0 ;
  assign n11909 = n4433 ^ n2781 ^ 1'b0 ;
  assign n11910 = n11908 & ~n11909 ;
  assign n11913 = n8733 ^ n3154 ^ 1'b0 ;
  assign n11912 = ~n5620 & n9130 ;
  assign n11914 = n11913 ^ n11912 ^ n6521 ;
  assign n11911 = n509 & n690 ;
  assign n11915 = n11914 ^ n11911 ^ 1'b0 ;
  assign n11916 = n8986 ^ n8971 ^ 1'b0 ;
  assign n11917 = n11916 ^ n8674 ^ 1'b0 ;
  assign n11918 = n11917 ^ n8242 ^ n1529 ;
  assign n11919 = n5950 ^ n2740 ^ n1452 ;
  assign n11920 = ( ~n3989 & n10701 ) | ( ~n3989 & n11919 ) | ( n10701 & n11919 ) ;
  assign n11921 = ~n11918 & n11920 ;
  assign n11922 = ~n11915 & n11921 ;
  assign n11924 = n2904 ^ n365 ^ x10 ;
  assign n11923 = ( x171 & ~n4113 ) | ( x171 & n6505 ) | ( ~n4113 & n6505 ) ;
  assign n11925 = n11924 ^ n11923 ^ 1'b0 ;
  assign n11926 = n6184 & ~n9908 ;
  assign n11927 = ~n5658 & n11926 ;
  assign n11928 = ( n773 & n8738 ) | ( n773 & n11927 ) | ( n8738 & n11927 ) ;
  assign n11929 = ( ~n6437 & n8897 ) | ( ~n6437 & n9601 ) | ( n8897 & n9601 ) ;
  assign n11930 = ( n5133 & n11928 ) | ( n5133 & n11929 ) | ( n11928 & n11929 ) ;
  assign n11931 = ( n3287 & n7355 ) | ( n3287 & n9932 ) | ( n7355 & n9932 ) ;
  assign n11933 = n4647 ^ n2624 ^ 1'b0 ;
  assign n11934 = n10930 & ~n11933 ;
  assign n11935 = n11934 ^ n9613 ^ n1745 ;
  assign n11932 = n1139 & n2218 ;
  assign n11936 = n11935 ^ n11932 ^ 1'b0 ;
  assign n11937 = ( n1123 & n11931 ) | ( n1123 & ~n11936 ) | ( n11931 & ~n11936 ) ;
  assign n11950 = n1179 & n1181 ;
  assign n11951 = ~n4732 & n11950 ;
  assign n11952 = ( ~n9047 & n9952 ) | ( ~n9047 & n11951 ) | ( n9952 & n11951 ) ;
  assign n11939 = n2934 | n5947 ;
  assign n11940 = n11939 ^ n1247 ^ 1'b0 ;
  assign n11941 = ( n2890 & n8569 ) | ( n2890 & ~n11940 ) | ( n8569 & ~n11940 ) ;
  assign n11942 = ( n3467 & n5042 ) | ( n3467 & ~n11941 ) | ( n5042 & ~n11941 ) ;
  assign n11943 = n10736 ^ n8640 ^ n3869 ;
  assign n11944 = n8390 ^ n4586 ^ n4397 ;
  assign n11945 = n11944 ^ n3779 ^ 1'b0 ;
  assign n11946 = n7517 | n11945 ;
  assign n11947 = ( x181 & ~n11943 ) | ( x181 & n11946 ) | ( ~n11943 & n11946 ) ;
  assign n11948 = ( n9666 & n11942 ) | ( n9666 & n11947 ) | ( n11942 & n11947 ) ;
  assign n11938 = n1399 | n11045 ;
  assign n11949 = n11948 ^ n11938 ^ n4653 ;
  assign n11953 = n11952 ^ n11949 ^ 1'b0 ;
  assign n11954 = n995 & n1990 ;
  assign n11955 = n11954 ^ n3791 ^ 1'b0 ;
  assign n11956 = ( n5353 & n6417 ) | ( n5353 & n9946 ) | ( n6417 & n9946 ) ;
  assign n11957 = ~n11955 & n11956 ;
  assign n11958 = n4888 & n9600 ;
  assign n11959 = n8824 ^ n4572 ^ n535 ;
  assign n11960 = ~n5554 & n6193 ;
  assign n11961 = n11959 & n11960 ;
  assign n11962 = ( n3426 & n8166 ) | ( n3426 & ~n11961 ) | ( n8166 & ~n11961 ) ;
  assign n11963 = ~n3016 & n4867 ;
  assign n11964 = n5133 & n11963 ;
  assign n11965 = ( n5343 & n9886 ) | ( n5343 & ~n11964 ) | ( n9886 & ~n11964 ) ;
  assign n11966 = ( ~n3381 & n11962 ) | ( ~n3381 & n11965 ) | ( n11962 & n11965 ) ;
  assign n11967 = n6349 ^ n4072 ^ x15 ;
  assign n11968 = ( n3944 & n11256 ) | ( n3944 & ~n11967 ) | ( n11256 & ~n11967 ) ;
  assign n11969 = n1451 ^ n556 ^ n410 ;
  assign n11970 = ( ~n5060 & n10939 ) | ( ~n5060 & n11969 ) | ( n10939 & n11969 ) ;
  assign n11971 = ( n469 & n3524 ) | ( n469 & n5492 ) | ( n3524 & n5492 ) ;
  assign n11972 = ( n1344 & n7493 ) | ( n1344 & ~n11971 ) | ( n7493 & ~n11971 ) ;
  assign n11973 = ( n7013 & n11970 ) | ( n7013 & ~n11972 ) | ( n11970 & ~n11972 ) ;
  assign n11981 = n9920 ^ n5322 ^ 1'b0 ;
  assign n11982 = ~n2157 & n11981 ;
  assign n11983 = ~n4465 & n11982 ;
  assign n11984 = n11983 ^ n8707 ^ 1'b0 ;
  assign n11985 = n997 | n11984 ;
  assign n11974 = n692 & ~n6012 ;
  assign n11975 = n11974 ^ n4530 ^ n1319 ;
  assign n11976 = n2844 ^ n2140 ^ 1'b0 ;
  assign n11977 = ~x191 & n11976 ;
  assign n11978 = ~n2733 & n11977 ;
  assign n11979 = n6265 | n11978 ;
  assign n11980 = ~n11975 & n11979 ;
  assign n11986 = n11985 ^ n11980 ^ 1'b0 ;
  assign n11988 = n5856 ^ n3227 ^ 1'b0 ;
  assign n11989 = ~n6535 & n11988 ;
  assign n11990 = ( n3384 & n7551 ) | ( n3384 & ~n11989 ) | ( n7551 & ~n11989 ) ;
  assign n11991 = ( n1038 & ~n4215 ) | ( n1038 & n11990 ) | ( ~n4215 & n11990 ) ;
  assign n11992 = ( ~n3925 & n3963 ) | ( ~n3925 & n11991 ) | ( n3963 & n11991 ) ;
  assign n11987 = n4745 | n10179 ;
  assign n11993 = n11992 ^ n11987 ^ n7757 ;
  assign n11994 = n3845 | n6149 ;
  assign n11995 = n1816 | n2173 ;
  assign n11996 = ( n4314 & n6745 ) | ( n4314 & ~n10644 ) | ( n6745 & ~n10644 ) ;
  assign n11997 = n9064 ^ n6112 ^ n2134 ;
  assign n11998 = n3218 | n11997 ;
  assign n12001 = n7920 ^ n7049 ^ n3642 ;
  assign n12002 = ( n3950 & n7313 ) | ( n3950 & ~n7339 ) | ( n7313 & ~n7339 ) ;
  assign n12003 = ( n2161 & n12001 ) | ( n2161 & ~n12002 ) | ( n12001 & ~n12002 ) ;
  assign n11999 = ( n4164 & n4369 ) | ( n4164 & ~n4735 ) | ( n4369 & ~n4735 ) ;
  assign n12000 = n9260 & ~n11999 ;
  assign n12004 = n12003 ^ n12000 ^ n8436 ;
  assign n12005 = n5248 ^ n1024 ^ n904 ;
  assign n12006 = n12004 | n12005 ;
  assign n12012 = n891 | n3051 ;
  assign n12013 = ( n1853 & n4194 ) | ( n1853 & ~n12012 ) | ( n4194 & ~n12012 ) ;
  assign n12014 = n9114 | n12013 ;
  assign n12015 = n3216 & ~n12014 ;
  assign n12016 = n478 | n12015 ;
  assign n12007 = n4780 ^ n1488 ^ n1282 ;
  assign n12008 = ( ~n349 & n3920 ) | ( ~n349 & n12007 ) | ( n3920 & n12007 ) ;
  assign n12009 = n4181 | n8818 ;
  assign n12010 = ( n3550 & ~n12008 ) | ( n3550 & n12009 ) | ( ~n12008 & n12009 ) ;
  assign n12011 = ( n5836 & n10148 ) | ( n5836 & ~n12010 ) | ( n10148 & ~n12010 ) ;
  assign n12017 = n12016 ^ n12011 ^ n4791 ;
  assign n12018 = ( n6954 & n11042 ) | ( n6954 & n12017 ) | ( n11042 & n12017 ) ;
  assign n12019 = n10763 ^ n6012 ^ n2078 ;
  assign n12020 = ( n4673 & ~n6424 ) | ( n4673 & n12019 ) | ( ~n6424 & n12019 ) ;
  assign n12021 = ( n4169 & n10117 ) | ( n4169 & ~n12020 ) | ( n10117 & ~n12020 ) ;
  assign n12022 = n1124 ^ n1088 ^ 1'b0 ;
  assign n12023 = ~n3865 & n12022 ;
  assign n12024 = n7169 ^ n2186 ^ n302 ;
  assign n12025 = n12024 ^ n1758 ^ x137 ;
  assign n12026 = n12025 ^ n4889 ^ 1'b0 ;
  assign n12027 = ( n2660 & ~n10967 ) | ( n2660 & n12026 ) | ( ~n10967 & n12026 ) ;
  assign n12028 = ( ~n2625 & n5251 ) | ( ~n2625 & n7353 ) | ( n5251 & n7353 ) ;
  assign n12029 = n3258 & ~n12028 ;
  assign n12030 = n696 & n11728 ;
  assign n12031 = n12029 & n12030 ;
  assign n12035 = n9164 ^ n7830 ^ n928 ;
  assign n12036 = n8313 ^ n5825 ^ 1'b0 ;
  assign n12037 = n12035 & n12036 ;
  assign n12032 = n11400 ^ n5583 ^ n4445 ;
  assign n12033 = x140 & ~n12032 ;
  assign n12034 = ~n3704 & n12033 ;
  assign n12038 = n12037 ^ n12034 ^ n1186 ;
  assign n12039 = n10500 ^ n4866 ^ n2711 ;
  assign n12040 = ( n474 & n4165 ) | ( n474 & ~n6886 ) | ( n4165 & ~n6886 ) ;
  assign n12041 = ( n4745 & n5466 ) | ( n4745 & ~n12040 ) | ( n5466 & ~n12040 ) ;
  assign n12042 = n12041 ^ n3668 ^ 1'b0 ;
  assign n12043 = n4137 & ~n12042 ;
  assign n12046 = n1184 | n3691 ;
  assign n12047 = n8749 | n12046 ;
  assign n12044 = ( ~n1712 & n1801 ) | ( ~n1712 & n3937 ) | ( n1801 & n3937 ) ;
  assign n12045 = n12044 ^ n4273 ^ n1587 ;
  assign n12048 = n12047 ^ n12045 ^ n8859 ;
  assign n12049 = n1173 & ~n4659 ;
  assign n12050 = n1995 | n2180 ;
  assign n12051 = ~n365 & n12050 ;
  assign n12052 = ~n8135 & n12051 ;
  assign n12053 = n12052 ^ n11639 ^ n9144 ;
  assign n12054 = ( ~x191 & n12049 ) | ( ~x191 & n12053 ) | ( n12049 & n12053 ) ;
  assign n12055 = n12054 ^ n10504 ^ n5969 ;
  assign n12056 = n12055 ^ n11160 ^ n9749 ;
  assign n12057 = ( n3447 & n10224 ) | ( n3447 & n12056 ) | ( n10224 & n12056 ) ;
  assign n12058 = n4983 ^ n3038 ^ n2394 ;
  assign n12069 = ( n1659 & ~n2696 ) | ( n1659 & n3152 ) | ( ~n2696 & n3152 ) ;
  assign n12070 = n12069 ^ n9591 ^ n2106 ;
  assign n12059 = n7043 ^ n5446 ^ n1424 ;
  assign n12060 = ( n1940 & n8054 ) | ( n1940 & ~n12059 ) | ( n8054 & ~n12059 ) ;
  assign n12064 = n6745 | n8726 ;
  assign n12065 = ( n358 & n527 ) | ( n358 & n12064 ) | ( n527 & n12064 ) ;
  assign n12066 = n12065 ^ n4563 ^ n1116 ;
  assign n12061 = ~n1636 & n4438 ;
  assign n12062 = n12061 ^ n2557 ^ 1'b0 ;
  assign n12063 = n1495 | n12062 ;
  assign n12067 = n12066 ^ n12063 ^ 1'b0 ;
  assign n12068 = ~n12060 & n12067 ;
  assign n12071 = n12070 ^ n12068 ^ n7673 ;
  assign n12072 = n5416 | n6626 ;
  assign n12073 = ( ~n6419 & n9991 ) | ( ~n6419 & n12072 ) | ( n9991 & n12072 ) ;
  assign n12074 = ( n3630 & n3832 ) | ( n3630 & n11575 ) | ( n3832 & n11575 ) ;
  assign n12075 = n12074 ^ n8822 ^ 1'b0 ;
  assign n12076 = n6246 & ~n12075 ;
  assign n12077 = n12076 ^ n8651 ^ 1'b0 ;
  assign n12078 = n2836 & ~n12077 ;
  assign n12079 = n12078 ^ n4203 ^ 1'b0 ;
  assign n12080 = n12073 & n12079 ;
  assign n12085 = n10184 ^ n3000 ^ n2687 ;
  assign n12086 = ( n5945 & n7028 ) | ( n5945 & n12085 ) | ( n7028 & n12085 ) ;
  assign n12087 = n7702 | n12086 ;
  assign n12081 = n8326 ^ n5804 ^ 1'b0 ;
  assign n12082 = n2548 & n12081 ;
  assign n12083 = n12082 ^ n6330 ^ 1'b0 ;
  assign n12084 = n1018 & n12083 ;
  assign n12088 = n12087 ^ n12084 ^ n10336 ;
  assign n12089 = n12088 ^ n7417 ^ 1'b0 ;
  assign n12090 = n1567 | n8267 ;
  assign n12091 = n624 ^ n614 ^ 1'b0 ;
  assign n12092 = n2941 & n12091 ;
  assign n12093 = n12092 ^ n1509 ^ 1'b0 ;
  assign n12094 = n9650 ^ n6591 ^ x29 ;
  assign n12095 = ( n4677 & n6903 ) | ( n4677 & ~n12094 ) | ( n6903 & ~n12094 ) ;
  assign n12096 = n8121 ^ n3593 ^ 1'b0 ;
  assign n12097 = n12095 & n12096 ;
  assign n12098 = ( n10808 & n12093 ) | ( n10808 & n12097 ) | ( n12093 & n12097 ) ;
  assign n12099 = ( ~n10921 & n12090 ) | ( ~n10921 & n12098 ) | ( n12090 & n12098 ) ;
  assign n12100 = n495 ^ x141 ^ 1'b0 ;
  assign n12101 = n1067 & ~n12100 ;
  assign n12102 = ( n2055 & n7397 ) | ( n2055 & n12101 ) | ( n7397 & n12101 ) ;
  assign n12103 = ( ~n2932 & n9918 ) | ( ~n2932 & n12102 ) | ( n9918 & n12102 ) ;
  assign n12104 = n12103 ^ n9656 ^ x37 ;
  assign n12106 = n1433 & n2178 ;
  assign n12107 = n12106 ^ n1972 ^ 1'b0 ;
  assign n12105 = n9982 ^ n9956 ^ n6906 ;
  assign n12108 = n12107 ^ n12105 ^ n1777 ;
  assign n12109 = n12108 ^ n6596 ^ n1133 ;
  assign n12110 = n1758 | n12109 ;
  assign n12111 = n10043 ^ n7863 ^ n3956 ;
  assign n12114 = n1233 & n3077 ;
  assign n12112 = ( ~n2197 & n5876 ) | ( ~n2197 & n8173 ) | ( n5876 & n8173 ) ;
  assign n12113 = n987 & n12112 ;
  assign n12115 = n12114 ^ n12113 ^ 1'b0 ;
  assign n12117 = n9552 ^ n6605 ^ 1'b0 ;
  assign n12118 = ( n2411 & n2606 ) | ( n2411 & ~n12117 ) | ( n2606 & ~n12117 ) ;
  assign n12116 = n1995 & n2644 ;
  assign n12119 = n12118 ^ n12116 ^ 1'b0 ;
  assign n12120 = n12119 ^ n3443 ^ 1'b0 ;
  assign n12121 = ( n382 & n2079 ) | ( n382 & n8854 ) | ( n2079 & n8854 ) ;
  assign n12122 = n3349 & ~n12121 ;
  assign n12123 = n11383 | n12122 ;
  assign n12124 = ( n3907 & ~n12120 ) | ( n3907 & n12123 ) | ( ~n12120 & n12123 ) ;
  assign n12126 = n5032 ^ n4538 ^ n2163 ;
  assign n12125 = n11999 ^ n8949 ^ n2381 ;
  assign n12127 = n12126 ^ n12125 ^ 1'b0 ;
  assign n12128 = n8854 & ~n12127 ;
  assign n12129 = n12124 & n12128 ;
  assign n12130 = n9799 & n12129 ;
  assign n12135 = n6056 ^ n5089 ^ n3780 ;
  assign n12136 = n12135 ^ n2608 ^ 1'b0 ;
  assign n12137 = n7032 & ~n12136 ;
  assign n12138 = n1341 & n12137 ;
  assign n12139 = n6589 | n12138 ;
  assign n12133 = n6690 ^ n3998 ^ n2192 ;
  assign n12131 = n10643 ^ n7326 ^ n1726 ;
  assign n12132 = n3211 & n12131 ;
  assign n12134 = n12133 ^ n12132 ^ n994 ;
  assign n12140 = n12139 ^ n12134 ^ 1'b0 ;
  assign n12141 = n11384 ^ n2239 ^ n1346 ;
  assign n12142 = ~n8454 & n12141 ;
  assign n12143 = ( n556 & ~n11401 ) | ( n556 & n12142 ) | ( ~n11401 & n12142 ) ;
  assign n12144 = n12143 ^ n5951 ^ n4164 ;
  assign n12145 = n1017 | n2073 ;
  assign n12146 = n12145 ^ n10082 ^ 1'b0 ;
  assign n12147 = n12146 ^ n4448 ^ n606 ;
  assign n12148 = n4182 & ~n5415 ;
  assign n12149 = n4494 ^ n631 ^ 1'b0 ;
  assign n12150 = n8994 ^ n7883 ^ n1949 ;
  assign n12151 = n5053 ^ n3461 ^ n1457 ;
  assign n12152 = n6269 ^ n5750 ^ n1536 ;
  assign n12153 = n11689 | n12152 ;
  assign n12154 = n12151 & ~n12153 ;
  assign n12155 = n12150 & n12154 ;
  assign n12156 = x68 & ~n7185 ;
  assign n12157 = ( n1856 & n2806 ) | ( n1856 & n2916 ) | ( n2806 & n2916 ) ;
  assign n12158 = ( n4909 & n12156 ) | ( n4909 & n12157 ) | ( n12156 & n12157 ) ;
  assign n12159 = n2275 | n12158 ;
  assign n12160 = n12159 ^ n9986 ^ 1'b0 ;
  assign n12165 = n3676 ^ n2836 ^ 1'b0 ;
  assign n12166 = n7577 & n12165 ;
  assign n12161 = n4492 & ~n9920 ;
  assign n12162 = n12161 ^ n9626 ^ 1'b0 ;
  assign n12163 = ( n4243 & n11824 ) | ( n4243 & ~n12162 ) | ( n11824 & ~n12162 ) ;
  assign n12164 = ~n670 & n12163 ;
  assign n12167 = n12166 ^ n12164 ^ 1'b0 ;
  assign n12168 = ( n3574 & n7452 ) | ( n3574 & n11694 ) | ( n7452 & n11694 ) ;
  assign n12169 = n5270 ^ n3794 ^ 1'b0 ;
  assign n12170 = n12168 & n12169 ;
  assign n12171 = n12170 ^ n4594 ^ n1437 ;
  assign n12172 = ~n8656 & n12171 ;
  assign n12173 = n9946 & n12172 ;
  assign n12174 = ( n12160 & ~n12167 ) | ( n12160 & n12173 ) | ( ~n12167 & n12173 ) ;
  assign n12175 = ( n2001 & n4339 ) | ( n2001 & n8013 ) | ( n4339 & n8013 ) ;
  assign n12176 = n2171 ^ n1225 ^ 1'b0 ;
  assign n12177 = ~n9428 & n12176 ;
  assign n12178 = n2486 & n12177 ;
  assign n12179 = n12178 ^ n8692 ^ 1'b0 ;
  assign n12180 = ( n1482 & n3949 ) | ( n1482 & ~n12073 ) | ( n3949 & ~n12073 ) ;
  assign n12181 = ( n4489 & ~n7211 ) | ( n4489 & n8484 ) | ( ~n7211 & n8484 ) ;
  assign n12182 = n11715 ^ n9781 ^ n6424 ;
  assign n12183 = n12182 ^ n10635 ^ n4879 ;
  assign n12184 = n12086 ^ n10185 ^ 1'b0 ;
  assign n12185 = n1973 | n10140 ;
  assign n12186 = n12184 & ~n12185 ;
  assign n12187 = ( n1131 & n3073 ) | ( n1131 & n10725 ) | ( n3073 & n10725 ) ;
  assign n12188 = n6926 ^ n5406 ^ n2134 ;
  assign n12189 = n12188 ^ n6423 ^ n4812 ;
  assign n12190 = ( n6482 & ~n7192 ) | ( n6482 & n11027 ) | ( ~n7192 & n11027 ) ;
  assign n12191 = ( n2470 & ~n3641 ) | ( n2470 & n4554 ) | ( ~n3641 & n4554 ) ;
  assign n12192 = ( n5350 & ~n12190 ) | ( n5350 & n12191 ) | ( ~n12190 & n12191 ) ;
  assign n12193 = ( n7952 & n12189 ) | ( n7952 & n12192 ) | ( n12189 & n12192 ) ;
  assign n12194 = ( ~n10485 & n12187 ) | ( ~n10485 & n12193 ) | ( n12187 & n12193 ) ;
  assign n12195 = ( ~n3916 & n4283 ) | ( ~n3916 & n11357 ) | ( n4283 & n11357 ) ;
  assign n12196 = n6409 ^ n5033 ^ 1'b0 ;
  assign n12197 = ~n12195 & n12196 ;
  assign n12198 = n12197 ^ n10392 ^ n1132 ;
  assign n12199 = n4730 ^ n2214 ^ n336 ;
  assign n12201 = ~n1082 & n1836 ;
  assign n12202 = n12201 ^ n3002 ^ 1'b0 ;
  assign n12200 = n548 & ~n8593 ;
  assign n12203 = n12202 ^ n12200 ^ n813 ;
  assign n12207 = n5818 & ~n7189 ;
  assign n12204 = n7971 & n9712 ;
  assign n12205 = n12204 ^ n2536 ^ 1'b0 ;
  assign n12206 = ( n5312 & ~n10169 ) | ( n5312 & n12205 ) | ( ~n10169 & n12205 ) ;
  assign n12208 = n12207 ^ n12206 ^ n1369 ;
  assign n12209 = ( ~n4492 & n7641 ) | ( ~n4492 & n7867 ) | ( n7641 & n7867 ) ;
  assign n12210 = n12209 ^ n8223 ^ n2217 ;
  assign n12213 = ( n3059 & n4878 ) | ( n3059 & n6790 ) | ( n4878 & n6790 ) ;
  assign n12211 = n4037 | n5216 ;
  assign n12212 = n12211 ^ n11021 ^ n6677 ;
  assign n12214 = n12213 ^ n12212 ^ n10969 ;
  assign n12215 = n5163 ^ n1444 ^ 1'b0 ;
  assign n12216 = ( n602 & n1583 ) | ( n602 & ~n12119 ) | ( n1583 & ~n12119 ) ;
  assign n12217 = ( ~n6396 & n12215 ) | ( ~n6396 & n12216 ) | ( n12215 & n12216 ) ;
  assign n12218 = n10077 & ~n12217 ;
  assign n12219 = n12218 ^ n5627 ^ 1'b0 ;
  assign n12221 = ( n324 & ~n883 ) | ( n324 & n5897 ) | ( ~n883 & n5897 ) ;
  assign n12220 = ( n728 & n2510 ) | ( n728 & ~n11055 ) | ( n2510 & ~n11055 ) ;
  assign n12222 = n12221 ^ n12220 ^ n11684 ;
  assign n12223 = n12219 & n12222 ;
  assign n12224 = ~n2394 & n12223 ;
  assign n12225 = ~n3593 & n7062 ;
  assign n12226 = n849 & n12225 ;
  assign n12227 = ( n2659 & ~n4047 ) | ( n2659 & n12226 ) | ( ~n4047 & n12226 ) ;
  assign n12228 = ( ~n463 & n2752 ) | ( ~n463 & n4188 ) | ( n2752 & n4188 ) ;
  assign n12229 = n12228 ^ n1278 ^ 1'b0 ;
  assign n12230 = ( n2813 & ~n4453 ) | ( n2813 & n12229 ) | ( ~n4453 & n12229 ) ;
  assign n12231 = ( n600 & n1421 ) | ( n600 & ~n12230 ) | ( n1421 & ~n12230 ) ;
  assign n12232 = ( n10641 & ~n10828 ) | ( n10641 & n12231 ) | ( ~n10828 & n12231 ) ;
  assign n12233 = ( n8718 & ~n12227 ) | ( n8718 & n12232 ) | ( ~n12227 & n12232 ) ;
  assign n12234 = n6667 ^ n3236 ^ n1293 ;
  assign n12235 = n12234 ^ n7443 ^ n3267 ;
  assign n12236 = n1508 ^ n850 ^ 1'b0 ;
  assign n12238 = n2784 ^ n904 ^ 1'b0 ;
  assign n12239 = n8834 | n12238 ;
  assign n12240 = n12239 ^ n11781 ^ n8733 ;
  assign n12237 = n9542 ^ n2108 ^ 1'b0 ;
  assign n12241 = n12240 ^ n12237 ^ n6136 ;
  assign n12242 = ( x86 & ~n486 ) | ( x86 & n1143 ) | ( ~n486 & n1143 ) ;
  assign n12243 = ( n2887 & n5918 ) | ( n2887 & n12242 ) | ( n5918 & n12242 ) ;
  assign n12244 = ( n12236 & ~n12241 ) | ( n12236 & n12243 ) | ( ~n12241 & n12243 ) ;
  assign n12245 = ( ~n4050 & n12235 ) | ( ~n4050 & n12244 ) | ( n12235 & n12244 ) ;
  assign n12246 = n5948 & ~n11682 ;
  assign n12247 = ( n461 & n2099 ) | ( n461 & ~n5293 ) | ( n2099 & ~n5293 ) ;
  assign n12248 = ( ~n1361 & n1385 ) | ( ~n1361 & n12247 ) | ( n1385 & n12247 ) ;
  assign n12249 = ( ~n5579 & n5651 ) | ( ~n5579 & n12248 ) | ( n5651 & n12248 ) ;
  assign n12250 = ( n10430 & ~n12072 ) | ( n10430 & n12249 ) | ( ~n12072 & n12249 ) ;
  assign n12251 = n6239 & ~n12250 ;
  assign n12252 = ~n12246 & n12251 ;
  assign n12253 = n12252 ^ n11274 ^ 1'b0 ;
  assign n12254 = ~n11231 & n12253 ;
  assign n12255 = n4967 & ~n11518 ;
  assign n12260 = n6433 ^ n1944 ^ 1'b0 ;
  assign n12256 = n289 & n3928 ;
  assign n12257 = ~x177 & n12256 ;
  assign n12258 = n12257 ^ n3641 ^ 1'b0 ;
  assign n12259 = n12258 ^ n7092 ^ n1186 ;
  assign n12261 = n12260 ^ n12259 ^ 1'b0 ;
  assign n12262 = ~n1627 & n12261 ;
  assign n12263 = n12262 ^ n7388 ^ n1296 ;
  assign n12264 = ( n350 & n12228 ) | ( n350 & ~n12263 ) | ( n12228 & ~n12263 ) ;
  assign n12265 = n1482 | n1968 ;
  assign n12266 = n5858 & ~n12265 ;
  assign n12267 = n6481 ^ n3180 ^ n828 ;
  assign n12268 = ( ~n3334 & n9264 ) | ( ~n3334 & n12267 ) | ( n9264 & n12267 ) ;
  assign n12269 = n9069 & n10416 ;
  assign n12270 = ~n825 & n12269 ;
  assign n12271 = n12270 ^ n8253 ^ n4834 ;
  assign n12272 = n1817 ^ n1464 ^ 1'b0 ;
  assign n12273 = ( n6018 & n6942 ) | ( n6018 & n12272 ) | ( n6942 & n12272 ) ;
  assign n12282 = ( ~n4263 & n4603 ) | ( ~n4263 & n5386 ) | ( n4603 & n5386 ) ;
  assign n12283 = n7013 & n12282 ;
  assign n12284 = n12283 ^ x209 ^ 1'b0 ;
  assign n12285 = n12284 ^ n10623 ^ n9785 ;
  assign n12279 = n2365 ^ n790 ^ 1'b0 ;
  assign n12280 = ~n2311 & n12279 ;
  assign n12281 = ( n1920 & n8555 ) | ( n1920 & ~n12280 ) | ( n8555 & ~n12280 ) ;
  assign n12286 = n12285 ^ n12281 ^ n1743 ;
  assign n12287 = n11376 | n12286 ;
  assign n12274 = n6716 ^ n3632 ^ 1'b0 ;
  assign n12275 = n12274 ^ n10319 ^ n8833 ;
  assign n12276 = n12275 ^ n3270 ^ n3067 ;
  assign n12277 = ( x140 & ~n9312 ) | ( x140 & n12276 ) | ( ~n9312 & n12276 ) ;
  assign n12278 = ~n11026 & n12277 ;
  assign n12288 = n12287 ^ n12278 ^ 1'b0 ;
  assign n12289 = n6232 ^ x140 ^ 1'b0 ;
  assign n12290 = n5155 & n12289 ;
  assign n12291 = n12290 ^ n9955 ^ 1'b0 ;
  assign n12292 = n10701 ^ n4300 ^ x38 ;
  assign n12293 = ( x191 & n4729 ) | ( x191 & n12249 ) | ( n4729 & n12249 ) ;
  assign n12294 = ( n1804 & ~n3157 ) | ( n1804 & n8825 ) | ( ~n3157 & n8825 ) ;
  assign n12295 = n10282 ^ n3571 ^ 1'b0 ;
  assign n12296 = n5352 | n12295 ;
  assign n12297 = ~n12294 & n12296 ;
  assign n12298 = n12293 & n12297 ;
  assign n12299 = ~n795 & n856 ;
  assign n12300 = ( ~n2031 & n6342 ) | ( ~n2031 & n9007 ) | ( n6342 & n9007 ) ;
  assign n12301 = ( n1788 & n12299 ) | ( n1788 & ~n12300 ) | ( n12299 & ~n12300 ) ;
  assign n12302 = ( n8889 & n9677 ) | ( n8889 & ~n12301 ) | ( n9677 & ~n12301 ) ;
  assign n12303 = n10154 ^ n3979 ^ x64 ;
  assign n12304 = ( n3209 & n4787 ) | ( n3209 & ~n12303 ) | ( n4787 & ~n12303 ) ;
  assign n12305 = n12302 & n12304 ;
  assign n12307 = n5640 ^ n4302 ^ n1308 ;
  assign n12308 = ( n3870 & n10318 ) | ( n3870 & n12307 ) | ( n10318 & n12307 ) ;
  assign n12306 = n4201 & ~n6840 ;
  assign n12309 = n12308 ^ n12306 ^ n9464 ;
  assign n12310 = n8259 ^ n4196 ^ n3777 ;
  assign n12311 = n7982 ^ n3136 ^ 1'b0 ;
  assign n12312 = n12310 | n12311 ;
  assign n12313 = n12312 ^ n10886 ^ 1'b0 ;
  assign n12314 = n12309 & ~n12313 ;
  assign n12315 = n4265 | n12314 ;
  assign n12316 = n9835 ^ n6951 ^ n2763 ;
  assign n12317 = n12316 ^ n997 ^ 1'b0 ;
  assign n12318 = n9602 | n12317 ;
  assign n12319 = n5130 ^ n4838 ^ n3591 ;
  assign n12320 = n6028 & ~n7105 ;
  assign n12321 = ( n10779 & ~n12319 ) | ( n10779 & n12320 ) | ( ~n12319 & n12320 ) ;
  assign n12322 = ( ~n5079 & n12318 ) | ( ~n5079 & n12321 ) | ( n12318 & n12321 ) ;
  assign n12323 = n8573 ^ n2383 ^ n310 ;
  assign n12324 = n2997 & n12323 ;
  assign n12325 = n11101 ^ n4349 ^ n3859 ;
  assign n12326 = n3307 & n5560 ;
  assign n12327 = n3987 ^ n3847 ^ 1'b0 ;
  assign n12328 = ~n1643 & n12327 ;
  assign n12329 = n2592 & n12328 ;
  assign n12330 = n5941 ^ n1955 ^ n1460 ;
  assign n12331 = ( n2415 & n12242 ) | ( n2415 & ~n12330 ) | ( n12242 & ~n12330 ) ;
  assign n12332 = n10953 ^ n7667 ^ n2449 ;
  assign n12333 = n7199 & ~n11703 ;
  assign n12334 = ~n6376 & n12333 ;
  assign n12336 = ~n2738 & n3798 ;
  assign n12335 = n6161 ^ n3566 ^ 1'b0 ;
  assign n12337 = n12336 ^ n12335 ^ 1'b0 ;
  assign n12340 = x115 | n341 ;
  assign n12338 = n537 ^ x45 ^ 1'b0 ;
  assign n12339 = ~n2958 & n12338 ;
  assign n12341 = n12340 ^ n12339 ^ n992 ;
  assign n12342 = n12341 ^ n349 ^ 1'b0 ;
  assign n12343 = ~n12337 & n12342 ;
  assign n12344 = ( ~n777 & n9533 ) | ( ~n777 & n12343 ) | ( n9533 & n12343 ) ;
  assign n12349 = n2740 | n6517 ;
  assign n12350 = n12349 ^ n622 ^ 1'b0 ;
  assign n12345 = ~n2339 & n2913 ;
  assign n12346 = n6560 ^ n4651 ^ n522 ;
  assign n12347 = n12345 & n12346 ;
  assign n12348 = ~n7062 & n12347 ;
  assign n12351 = n12350 ^ n12348 ^ n2884 ;
  assign n12352 = n12344 & n12351 ;
  assign n12353 = n12352 ^ n4011 ^ 1'b0 ;
  assign n12354 = n2778 ^ n333 ^ 1'b0 ;
  assign n12355 = n5745 | n12354 ;
  assign n12356 = n2176 ^ n360 ^ 1'b0 ;
  assign n12357 = n4635 & n12356 ;
  assign n12358 = ~n3905 & n12357 ;
  assign n12359 = n2352 ^ n1344 ^ 1'b0 ;
  assign n12360 = n425 & n12359 ;
  assign n12361 = n10309 ^ n3921 ^ 1'b0 ;
  assign n12362 = ( n2400 & ~n12360 ) | ( n2400 & n12361 ) | ( ~n12360 & n12361 ) ;
  assign n12368 = ( n2034 & ~n2853 ) | ( n2034 & n5951 ) | ( ~n2853 & n5951 ) ;
  assign n12364 = n1397 & n11400 ;
  assign n12365 = n12364 ^ n4152 ^ 1'b0 ;
  assign n12363 = ( n5316 & ~n5912 ) | ( n5316 & n7861 ) | ( ~n5912 & n7861 ) ;
  assign n12366 = n12365 ^ n12363 ^ n5002 ;
  assign n12367 = ( n2842 & n4559 ) | ( n2842 & n12366 ) | ( n4559 & n12366 ) ;
  assign n12369 = n12368 ^ n12367 ^ 1'b0 ;
  assign n12370 = ~n12362 & n12369 ;
  assign n12371 = ( n5484 & ~n12358 ) | ( n5484 & n12370 ) | ( ~n12358 & n12370 ) ;
  assign n12372 = ~n12355 & n12371 ;
  assign n12373 = ( n12334 & ~n12353 ) | ( n12334 & n12372 ) | ( ~n12353 & n12372 ) ;
  assign n12374 = ( n1278 & n2888 ) | ( n1278 & ~n4190 ) | ( n2888 & ~n4190 ) ;
  assign n12375 = n12374 ^ x70 ^ 1'b0 ;
  assign n12376 = n8933 ^ n7596 ^ n874 ;
  assign n12377 = ( n4355 & n12375 ) | ( n4355 & n12376 ) | ( n12375 & n12376 ) ;
  assign n12385 = n562 | n5964 ;
  assign n12386 = n9350 ^ n6430 ^ n5230 ;
  assign n12387 = ( n1309 & n12385 ) | ( n1309 & n12386 ) | ( n12385 & n12386 ) ;
  assign n12384 = n2952 & n2962 ;
  assign n12388 = n12387 ^ n12384 ^ 1'b0 ;
  assign n12378 = x232 & n1195 ;
  assign n12379 = n12378 ^ n4651 ^ 1'b0 ;
  assign n12380 = n10921 ^ n5233 ^ 1'b0 ;
  assign n12381 = n12379 | n12380 ;
  assign n12382 = ( n687 & ~n11835 ) | ( n687 & n12381 ) | ( ~n11835 & n12381 ) ;
  assign n12383 = n11045 | n12382 ;
  assign n12389 = n12388 ^ n12383 ^ 1'b0 ;
  assign n12396 = ( ~n1636 & n1814 ) | ( ~n1636 & n1875 ) | ( n1814 & n1875 ) ;
  assign n12397 = n3157 ^ n903 ^ 1'b0 ;
  assign n12398 = n12396 & n12397 ;
  assign n12399 = n12398 ^ n4044 ^ 1'b0 ;
  assign n12400 = ~n3967 & n12399 ;
  assign n12401 = ( n1309 & n2750 ) | ( n1309 & ~n12400 ) | ( n2750 & ~n12400 ) ;
  assign n12392 = n5818 ^ n3008 ^ n2960 ;
  assign n12393 = n12392 ^ n270 ^ 1'b0 ;
  assign n12394 = ~n3449 & n12393 ;
  assign n12395 = n6920 | n12394 ;
  assign n12402 = n12401 ^ n12395 ^ 1'b0 ;
  assign n12403 = ( n1023 & n8023 ) | ( n1023 & ~n12402 ) | ( n8023 & ~n12402 ) ;
  assign n12390 = n9586 ^ n7171 ^ 1'b0 ;
  assign n12391 = n12390 ^ n3617 ^ x212 ;
  assign n12404 = n12403 ^ n12391 ^ n1713 ;
  assign n12405 = n10121 ^ n4431 ^ n1095 ;
  assign n12406 = n12405 ^ n4810 ^ n1226 ;
  assign n12407 = n7330 & n12406 ;
  assign n12408 = n6971 ^ n5800 ^ 1'b0 ;
  assign n12409 = ~n2651 & n12408 ;
  assign n12410 = n10582 ^ n1657 ^ 1'b0 ;
  assign n12411 = n12409 & ~n12410 ;
  assign n12412 = n6111 ^ n1821 ^ 1'b0 ;
  assign n12413 = ( ~n5738 & n7732 ) | ( ~n5738 & n12412 ) | ( n7732 & n12412 ) ;
  assign n12414 = ( n1981 & n8522 ) | ( n1981 & n12413 ) | ( n8522 & n12413 ) ;
  assign n12415 = ( n8096 & n10476 ) | ( n8096 & ~n12103 ) | ( n10476 & ~n12103 ) ;
  assign n12416 = n12415 ^ n3213 ^ n2016 ;
  assign n12417 = x13 & ~n9895 ;
  assign n12418 = ~n2607 & n12417 ;
  assign n12419 = ( x68 & n664 ) | ( x68 & n8630 ) | ( n664 & n8630 ) ;
  assign n12420 = ( n1188 & ~n3129 ) | ( n1188 & n12419 ) | ( ~n3129 & n12419 ) ;
  assign n12421 = n10924 ^ n9310 ^ n6684 ;
  assign n12422 = ( ~n2550 & n12420 ) | ( ~n2550 & n12421 ) | ( n12420 & n12421 ) ;
  assign n12423 = ( n5761 & n7158 ) | ( n5761 & ~n11049 ) | ( n7158 & ~n11049 ) ;
  assign n12424 = n12423 ^ n2737 ^ n1357 ;
  assign n12425 = ( n1560 & n6732 ) | ( n1560 & ~n12424 ) | ( n6732 & ~n12424 ) ;
  assign n12427 = ( ~n756 & n2066 ) | ( ~n756 & n2756 ) | ( n2066 & n2756 ) ;
  assign n12426 = n2993 & ~n3548 ;
  assign n12428 = n12427 ^ n12426 ^ 1'b0 ;
  assign n12429 = n6851 ^ n3721 ^ 1'b0 ;
  assign n12430 = n10697 ^ n3461 ^ n1137 ;
  assign n12431 = n760 & n4738 ;
  assign n12432 = n12430 & n12431 ;
  assign n12433 = n12307 ^ n11942 ^ n5480 ;
  assign n12434 = ( n12429 & ~n12432 ) | ( n12429 & n12433 ) | ( ~n12432 & n12433 ) ;
  assign n12436 = ~n385 & n4608 ;
  assign n12435 = x247 & n7766 ;
  assign n12437 = n12436 ^ n12435 ^ 1'b0 ;
  assign n12438 = n12234 ^ n298 ^ x32 ;
  assign n12439 = n10650 ^ n5040 ^ 1'b0 ;
  assign n12440 = ( n12437 & ~n12438 ) | ( n12437 & n12439 ) | ( ~n12438 & n12439 ) ;
  assign n12441 = n1479 & ~n1626 ;
  assign n12442 = n12441 ^ n604 ^ 1'b0 ;
  assign n12443 = ( ~n3933 & n5534 ) | ( ~n3933 & n10883 ) | ( n5534 & n10883 ) ;
  assign n12444 = ( n2447 & n12442 ) | ( n2447 & n12443 ) | ( n12442 & n12443 ) ;
  assign n12445 = n12444 ^ n1838 ^ n1230 ;
  assign n12446 = ( n2648 & n8970 ) | ( n2648 & ~n11969 ) | ( n8970 & ~n11969 ) ;
  assign n12447 = ( n2080 & n6697 ) | ( n2080 & ~n12446 ) | ( n6697 & ~n12446 ) ;
  assign n12448 = n9039 ^ n5177 ^ n3681 ;
  assign n12449 = n3654 ^ n942 ^ 1'b0 ;
  assign n12450 = n2696 & n12449 ;
  assign n12451 = n12450 ^ n945 ^ x15 ;
  assign n12452 = n12451 ^ n8387 ^ 1'b0 ;
  assign n12453 = ( n3870 & n12448 ) | ( n3870 & ~n12452 ) | ( n12448 & ~n12452 ) ;
  assign n12454 = ( n2045 & ~n6997 ) | ( n2045 & n11526 ) | ( ~n6997 & n11526 ) ;
  assign n12455 = n4057 ^ n628 ^ n300 ;
  assign n12456 = ( n5742 & n7454 ) | ( n5742 & ~n12455 ) | ( n7454 & ~n12455 ) ;
  assign n12457 = n5514 & n12456 ;
  assign n12458 = n12454 & n12457 ;
  assign n12459 = ~n8100 & n11545 ;
  assign n12460 = n1631 & n12459 ;
  assign n12461 = n5983 & n12460 ;
  assign n12462 = n3397 ^ n2019 ^ n508 ;
  assign n12463 = n5291 ^ n3485 ^ n1692 ;
  assign n12464 = ( n8241 & n12462 ) | ( n8241 & ~n12463 ) | ( n12462 & ~n12463 ) ;
  assign n12465 = n9118 ^ n5614 ^ n5131 ;
  assign n12466 = ( n1139 & ~n12464 ) | ( n1139 & n12465 ) | ( ~n12464 & n12465 ) ;
  assign n12467 = n8880 ^ n6110 ^ n3931 ;
  assign n12468 = n575 ^ n382 ^ 1'b0 ;
  assign n12469 = n12468 ^ n3219 ^ n2428 ;
  assign n12470 = ( n2557 & ~n12467 ) | ( n2557 & n12469 ) | ( ~n12467 & n12469 ) ;
  assign n12471 = n10627 ^ n620 ^ 1'b0 ;
  assign n12472 = n336 & ~n2561 ;
  assign n12473 = ~n2499 & n12472 ;
  assign n12474 = n5915 & ~n12473 ;
  assign n12475 = n12474 ^ n3989 ^ 1'b0 ;
  assign n12476 = n12475 ^ n2194 ^ n796 ;
  assign n12477 = n12476 ^ n8923 ^ n978 ;
  assign n12478 = x144 & n6602 ;
  assign n12479 = n12307 & n12478 ;
  assign n12482 = n4894 ^ n2667 ^ 1'b0 ;
  assign n12483 = n687 & ~n12482 ;
  assign n12484 = ~n8155 & n12483 ;
  assign n12480 = n425 & n5614 ;
  assign n12481 = ~n2101 & n12480 ;
  assign n12485 = n12484 ^ n12481 ^ n2181 ;
  assign n12486 = ( ~n6769 & n12479 ) | ( ~n6769 & n12485 ) | ( n12479 & n12485 ) ;
  assign n12488 = n8522 ^ n4225 ^ n1902 ;
  assign n12487 = ~n5066 & n9669 ;
  assign n12489 = n12488 ^ n12487 ^ 1'b0 ;
  assign n12490 = n12489 ^ n11826 ^ n6762 ;
  assign n12491 = ~n1626 & n3351 ;
  assign n12492 = ( n5719 & n7243 ) | ( n5719 & ~n7939 ) | ( n7243 & ~n7939 ) ;
  assign n12493 = ( x103 & ~n1637 ) | ( x103 & n12492 ) | ( ~n1637 & n12492 ) ;
  assign n12494 = n12493 ^ n8606 ^ 1'b0 ;
  assign n12495 = ~n6338 & n12494 ;
  assign n12499 = n7642 ^ n4644 ^ 1'b0 ;
  assign n12496 = n5132 & n10398 ;
  assign n12497 = ~n282 & n12496 ;
  assign n12498 = ( ~n1899 & n6970 ) | ( ~n1899 & n12497 ) | ( n6970 & n12497 ) ;
  assign n12500 = n12499 ^ n12498 ^ n5322 ;
  assign n12501 = n7594 ^ n2367 ^ 1'b0 ;
  assign n12502 = ~n5335 & n12501 ;
  assign n12503 = ( ~n4003 & n12453 ) | ( ~n4003 & n12502 ) | ( n12453 & n12502 ) ;
  assign n12504 = n12267 ^ n5639 ^ 1'b0 ;
  assign n12505 = n5354 & ~n12504 ;
  assign n12506 = n3936 ^ n2703 ^ 1'b0 ;
  assign n12507 = n2417 | n12506 ;
  assign n12508 = ( n4396 & ~n9062 ) | ( n4396 & n12507 ) | ( ~n9062 & n12507 ) ;
  assign n12512 = n11854 ^ n3460 ^ n3138 ;
  assign n12509 = ( n530 & n3441 ) | ( n530 & n9907 ) | ( n3441 & n9907 ) ;
  assign n12510 = n12050 ^ n9001 ^ n7037 ;
  assign n12511 = n12509 & ~n12510 ;
  assign n12513 = n12512 ^ n12511 ^ 1'b0 ;
  assign n12515 = x30 & ~n5769 ;
  assign n12516 = n12515 ^ n6389 ^ 1'b0 ;
  assign n12517 = n4009 ^ n2305 ^ 1'b0 ;
  assign n12518 = n5407 | n12517 ;
  assign n12519 = ( n8923 & n12516 ) | ( n8923 & ~n12518 ) | ( n12516 & ~n12518 ) ;
  assign n12514 = ~n3481 & n4339 ;
  assign n12520 = n12519 ^ n12514 ^ 1'b0 ;
  assign n12524 = ( n429 & ~n1804 ) | ( n429 & n2278 ) | ( ~n1804 & n2278 ) ;
  assign n12525 = ~n4521 & n12524 ;
  assign n12526 = n12525 ^ n4485 ^ 1'b0 ;
  assign n12521 = ( ~n1797 & n2699 ) | ( ~n1797 & n11183 ) | ( n2699 & n11183 ) ;
  assign n12522 = n9883 ^ n4579 ^ 1'b0 ;
  assign n12523 = n12521 | n12522 ;
  assign n12527 = n12526 ^ n12523 ^ 1'b0 ;
  assign n12528 = n10414 | n12527 ;
  assign n12529 = n12528 ^ n9927 ^ n5111 ;
  assign n12530 = n10270 ^ n4570 ^ 1'b0 ;
  assign n12531 = n9930 | n10691 ;
  assign n12532 = n1383 & ~n2933 ;
  assign n12533 = n11773 & n12532 ;
  assign n12534 = n12533 ^ n10955 ^ n2951 ;
  assign n12535 = n12534 ^ n3318 ^ 1'b0 ;
  assign n12536 = n12535 ^ n6771 ^ n4424 ;
  assign n12538 = n6356 & ~n11884 ;
  assign n12539 = n6323 & n12538 ;
  assign n12537 = n3490 & n7322 ;
  assign n12540 = n12539 ^ n12537 ^ 1'b0 ;
  assign n12541 = ( n858 & ~n2875 ) | ( n858 & n5055 ) | ( ~n2875 & n5055 ) ;
  assign n12542 = n12541 ^ n8302 ^ n3747 ;
  assign n12545 = n10059 ^ n7493 ^ n2462 ;
  assign n12543 = n12360 ^ n7523 ^ n2097 ;
  assign n12544 = ( n5303 & ~n10185 ) | ( n5303 & n12543 ) | ( ~n10185 & n12543 ) ;
  assign n12546 = n12545 ^ n12544 ^ n3658 ;
  assign n12547 = n1334 ^ x139 ^ 1'b0 ;
  assign n12548 = n12547 ^ n10140 ^ 1'b0 ;
  assign n12552 = n702 & ~n2907 ;
  assign n12553 = ~x77 & n12552 ;
  assign n12550 = n4640 ^ n4166 ^ n4156 ;
  assign n12551 = ~n4911 & n12550 ;
  assign n12554 = n12553 ^ n12551 ^ n1995 ;
  assign n12549 = n7582 & ~n10109 ;
  assign n12555 = n12554 ^ n12549 ^ 1'b0 ;
  assign n12561 = n3919 ^ n3260 ^ n877 ;
  assign n12560 = ( n4744 & n8188 ) | ( n4744 & ~n10762 ) | ( n8188 & ~n10762 ) ;
  assign n12557 = n4502 ^ n1999 ^ n1883 ;
  assign n12558 = n12557 ^ n6887 ^ n1759 ;
  assign n12556 = ~n376 & n4744 ;
  assign n12559 = n12558 ^ n12556 ^ 1'b0 ;
  assign n12562 = n12561 ^ n12560 ^ n12559 ;
  assign n12565 = n3899 ^ n1229 ^ 1'b0 ;
  assign n12566 = n6535 | n12565 ;
  assign n12563 = ( ~x101 & n1672 ) | ( ~x101 & n1997 ) | ( n1672 & n1997 ) ;
  assign n12564 = n12563 ^ n5219 ^ n4559 ;
  assign n12567 = n12566 ^ n12564 ^ n920 ;
  assign n12568 = n12567 ^ n871 ^ 1'b0 ;
  assign n12569 = n12562 & n12568 ;
  assign n12570 = n4982 ^ n2381 ^ n2230 ;
  assign n12571 = n12570 ^ n6579 ^ n4897 ;
  assign n12572 = n7023 ^ n4548 ^ 1'b0 ;
  assign n12573 = ( n5452 & ~n12571 ) | ( n5452 & n12572 ) | ( ~n12571 & n12572 ) ;
  assign n12579 = n2625 ^ n2329 ^ 1'b0 ;
  assign n12574 = ( n340 & n1177 ) | ( n340 & ~n5697 ) | ( n1177 & ~n5697 ) ;
  assign n12575 = ( n1009 & n2939 ) | ( n1009 & ~n12574 ) | ( n2939 & ~n12574 ) ;
  assign n12576 = ( n2060 & n2079 ) | ( n2060 & n9349 ) | ( n2079 & n9349 ) ;
  assign n12577 = ( n691 & ~n6863 ) | ( n691 & n12576 ) | ( ~n6863 & n12576 ) ;
  assign n12578 = ( n12427 & n12575 ) | ( n12427 & n12577 ) | ( n12575 & n12577 ) ;
  assign n12580 = n12579 ^ n12578 ^ n650 ;
  assign n12583 = n7417 ^ n2918 ^ 1'b0 ;
  assign n12584 = n8755 | n12583 ;
  assign n12582 = n2806 & n3044 ;
  assign n12581 = ( ~n4191 & n7429 ) | ( ~n4191 & n12206 ) | ( n7429 & n12206 ) ;
  assign n12585 = n12584 ^ n12582 ^ n12581 ;
  assign n12586 = n6627 ^ n5981 ^ n5152 ;
  assign n12587 = n5144 & ~n12586 ;
  assign n12588 = n12587 ^ n7907 ^ 1'b0 ;
  assign n12589 = n9812 & ~n12588 ;
  assign n12590 = ~n6027 & n12589 ;
  assign n12591 = n1261 & ~n7104 ;
  assign n12599 = n7858 ^ n2412 ^ 1'b0 ;
  assign n12600 = n3942 & n12599 ;
  assign n12593 = ( n1639 & ~n2887 ) | ( n1639 & n3525 ) | ( ~n2887 & n3525 ) ;
  assign n12594 = n8252 ^ n6906 ^ 1'b0 ;
  assign n12595 = n1037 | n12594 ;
  assign n12596 = ( ~n1778 & n12593 ) | ( ~n1778 & n12595 ) | ( n12593 & n12595 ) ;
  assign n12592 = n5323 ^ n4388 ^ n3262 ;
  assign n12597 = n12596 ^ n12592 ^ 1'b0 ;
  assign n12598 = n2695 & ~n12597 ;
  assign n12601 = n12600 ^ n12598 ^ 1'b0 ;
  assign n12602 = n7171 ^ n5635 ^ n4965 ;
  assign n12603 = n5480 ^ n621 ^ 1'b0 ;
  assign n12604 = n4010 & ~n12603 ;
  assign n12605 = ~n12602 & n12604 ;
  assign n12606 = n4787 & n6340 ;
  assign n12607 = n6915 ^ n5425 ^ n4109 ;
  assign n12608 = ( n12387 & n12606 ) | ( n12387 & n12607 ) | ( n12606 & n12607 ) ;
  assign n12609 = ( n4769 & n7057 ) | ( n4769 & n11727 ) | ( n7057 & n11727 ) ;
  assign n12610 = n12609 ^ n10935 ^ n1020 ;
  assign n12611 = ( n983 & n2029 ) | ( n983 & ~n8436 ) | ( n2029 & ~n8436 ) ;
  assign n12612 = ( n540 & ~n3125 ) | ( n540 & n5428 ) | ( ~n3125 & n5428 ) ;
  assign n12613 = n12612 ^ n11789 ^ 1'b0 ;
  assign n12614 = n1206 & ~n12613 ;
  assign n12615 = n12614 ^ n9100 ^ 1'b0 ;
  assign n12616 = n12611 & ~n12615 ;
  assign n12617 = n4323 ^ n3792 ^ n2786 ;
  assign n12618 = n12617 ^ n12301 ^ n3791 ;
  assign n12619 = ( n1914 & ~n12072 ) | ( n1914 & n12618 ) | ( ~n12072 & n12618 ) ;
  assign n12630 = n9279 ^ n7369 ^ n3325 ;
  assign n12620 = ( n2397 & n9344 ) | ( n2397 & ~n11037 ) | ( n9344 & ~n11037 ) ;
  assign n12623 = n620 | n2835 ;
  assign n12624 = n12623 ^ x46 ^ 1'b0 ;
  assign n12621 = x211 & n1031 ;
  assign n12622 = n12621 ^ n5679 ^ 1'b0 ;
  assign n12625 = n12624 ^ n12622 ^ 1'b0 ;
  assign n12626 = n12625 ^ n8983 ^ 1'b0 ;
  assign n12627 = ( n7121 & ~n12620 ) | ( n7121 & n12626 ) | ( ~n12620 & n12626 ) ;
  assign n12628 = ( n4852 & n5764 ) | ( n4852 & ~n12627 ) | ( n5764 & ~n12627 ) ;
  assign n12629 = ~n1014 & n12628 ;
  assign n12631 = n12630 ^ n12629 ^ n10775 ;
  assign n12637 = ~n1833 & n5543 ;
  assign n12632 = n1896 & ~n2353 ;
  assign n12633 = n12073 ^ n463 ^ 1'b0 ;
  assign n12634 = n6253 & n12633 ;
  assign n12635 = n12634 ^ n9067 ^ 1'b0 ;
  assign n12636 = n12632 | n12635 ;
  assign n12638 = n12637 ^ n12636 ^ 1'b0 ;
  assign n12639 = n5571 & n10844 ;
  assign n12640 = n8628 ^ n2684 ^ 1'b0 ;
  assign n12641 = n1595 | n12640 ;
  assign n12642 = n4295 | n12641 ;
  assign n12643 = n8041 & n12642 ;
  assign n12644 = n12643 ^ n3990 ^ 1'b0 ;
  assign n12645 = ~n4365 & n12644 ;
  assign n12646 = n12645 ^ n3167 ^ 1'b0 ;
  assign n12647 = n12646 ^ n1122 ^ 1'b0 ;
  assign n12648 = n10148 & ~n12647 ;
  assign n12649 = n12229 ^ n11760 ^ n11279 ;
  assign n12650 = n12649 ^ n8842 ^ 1'b0 ;
  assign n12651 = n9771 & ~n12650 ;
  assign n12652 = n11747 ^ n5564 ^ n603 ;
  assign n12653 = n8659 & ~n12652 ;
  assign n12654 = n12653 ^ n12592 ^ 1'b0 ;
  assign n12660 = n1974 ^ n1564 ^ n1559 ;
  assign n12661 = n4877 | n12660 ;
  assign n12662 = ~n4120 & n12661 ;
  assign n12663 = n7485 & n12662 ;
  assign n12655 = x184 & n2813 ;
  assign n12656 = ~n1372 & n12655 ;
  assign n12657 = n2743 | n3505 ;
  assign n12658 = n12657 ^ n3000 ^ 1'b0 ;
  assign n12659 = ( n6456 & n12656 ) | ( n6456 & ~n12658 ) | ( n12656 & ~n12658 ) ;
  assign n12664 = n12663 ^ n12659 ^ n673 ;
  assign n12666 = n433 | n5429 ;
  assign n12665 = ~n8593 & n11125 ;
  assign n12667 = n12666 ^ n12665 ^ n2948 ;
  assign n12668 = ( n1283 & n4891 ) | ( n1283 & ~n7917 ) | ( n4891 & ~n7917 ) ;
  assign n12669 = n6535 ^ n6092 ^ n4893 ;
  assign n12670 = n9189 & ~n12669 ;
  assign n12671 = n12670 ^ n12216 ^ n9165 ;
  assign n12672 = n4051 & n5698 ;
  assign n12673 = n11619 ^ n3094 ^ 1'b0 ;
  assign n12674 = ~n1697 & n12673 ;
  assign n12675 = n12438 ^ n10738 ^ 1'b0 ;
  assign n12678 = n5738 ^ n2674 ^ 1'b0 ;
  assign n12679 = n3720 | n7982 ;
  assign n12680 = n12678 | n12679 ;
  assign n12676 = n691 & ~n9536 ;
  assign n12677 = n12676 ^ n4169 ^ 1'b0 ;
  assign n12681 = n12680 ^ n12677 ^ n5412 ;
  assign n12682 = n12675 & ~n12681 ;
  assign n12683 = ( n2686 & n4150 ) | ( n2686 & n5163 ) | ( n4150 & n5163 ) ;
  assign n12684 = ~n7553 & n12683 ;
  assign n12685 = n4934 & n12684 ;
  assign n12686 = n3922 | n7401 ;
  assign n12687 = ( n3031 & ~n12685 ) | ( n3031 & n12686 ) | ( ~n12685 & n12686 ) ;
  assign n12688 = ( n2527 & n3310 ) | ( n2527 & ~n8872 ) | ( n3310 & ~n8872 ) ;
  assign n12689 = n7860 ^ n5199 ^ 1'b0 ;
  assign n12690 = ( n9027 & ~n10226 ) | ( n9027 & n11085 ) | ( ~n10226 & n11085 ) ;
  assign n12691 = ( n12688 & ~n12689 ) | ( n12688 & n12690 ) | ( ~n12689 & n12690 ) ;
  assign n12692 = ( ~n9341 & n12687 ) | ( ~n9341 & n12691 ) | ( n12687 & n12691 ) ;
  assign n12693 = n12692 ^ n1305 ^ 1'b0 ;
  assign n12694 = n6695 | n12693 ;
  assign n12695 = ( ~n2223 & n6351 ) | ( ~n2223 & n6433 ) | ( n6351 & n6433 ) ;
  assign n12696 = ( n452 & n10601 ) | ( n452 & ~n11696 ) | ( n10601 & ~n11696 ) ;
  assign n12697 = n10389 ^ n870 ^ n583 ;
  assign n12698 = n1362 ^ n1262 ^ 1'b0 ;
  assign n12699 = n12697 & n12698 ;
  assign n12700 = n6494 & n12699 ;
  assign n12701 = n486 & n12700 ;
  assign n12702 = ( n1095 & n12696 ) | ( n1095 & n12701 ) | ( n12696 & n12701 ) ;
  assign n12703 = n9910 ^ n1850 ^ 1'b0 ;
  assign n12704 = ( ~n5058 & n5953 ) | ( ~n5058 & n12703 ) | ( n5953 & n12703 ) ;
  assign n12705 = n4307 & n12704 ;
  assign n12706 = ( ~n5294 & n12702 ) | ( ~n5294 & n12705 ) | ( n12702 & n12705 ) ;
  assign n12710 = n6130 & ~n6498 ;
  assign n12711 = n12710 ^ n6205 ^ 1'b0 ;
  assign n12707 = n6990 ^ n4570 ^ n442 ;
  assign n12708 = n7721 ^ n3708 ^ 1'b0 ;
  assign n12709 = ( n6954 & ~n12707 ) | ( n6954 & n12708 ) | ( ~n12707 & n12708 ) ;
  assign n12712 = n12711 ^ n12709 ^ n4749 ;
  assign n12713 = n5506 ^ n2837 ^ 1'b0 ;
  assign n12714 = n12712 | n12713 ;
  assign n12715 = ( ~n4205 & n8582 ) | ( ~n4205 & n12360 ) | ( n8582 & n12360 ) ;
  assign n12719 = n6193 & n11715 ;
  assign n12720 = ( n468 & ~n854 ) | ( n468 & n12719 ) | ( ~n854 & n12719 ) ;
  assign n12717 = n5488 ^ n4772 ^ n1900 ;
  assign n12716 = n7184 ^ n5034 ^ n4400 ;
  assign n12718 = n12717 ^ n12716 ^ 1'b0 ;
  assign n12721 = n12720 ^ n12718 ^ n9524 ;
  assign n12722 = ( ~n2318 & n5169 ) | ( ~n2318 & n6232 ) | ( n5169 & n6232 ) ;
  assign n12723 = n12722 ^ n1264 ^ 1'b0 ;
  assign n12724 = n7732 | n12723 ;
  assign n12725 = n10156 ^ n5777 ^ n2825 ;
  assign n12726 = n4866 ^ n1331 ^ 1'b0 ;
  assign n12727 = n4074 ^ n2450 ^ n1191 ;
  assign n12728 = n1706 | n6544 ;
  assign n12729 = n12727 & ~n12728 ;
  assign n12730 = ~n12726 & n12729 ;
  assign n12731 = ( n12724 & n12725 ) | ( n12724 & ~n12730 ) | ( n12725 & ~n12730 ) ;
  assign n12732 = n2871 & ~n5022 ;
  assign n12733 = n12732 ^ n1541 ^ 1'b0 ;
  assign n12734 = n12733 ^ n3494 ^ 1'b0 ;
  assign n12735 = n12731 & n12734 ;
  assign n12736 = ( n2319 & n5213 ) | ( n2319 & ~n10912 ) | ( n5213 & ~n10912 ) ;
  assign n12737 = ( n3956 & ~n8588 ) | ( n3956 & n12736 ) | ( ~n8588 & n12736 ) ;
  assign n12739 = n2347 & ~n2371 ;
  assign n12740 = n1717 & ~n12739 ;
  assign n12741 = n4588 & n12740 ;
  assign n12738 = ( ~n2341 & n7856 ) | ( ~n2341 & n9907 ) | ( n7856 & n9907 ) ;
  assign n12742 = n12741 ^ n12738 ^ n5471 ;
  assign n12743 = n12742 ^ n8085 ^ x24 ;
  assign n12744 = n12743 ^ n7437 ^ 1'b0 ;
  assign n12754 = n1107 & ~n7183 ;
  assign n12755 = ~n3181 & n12754 ;
  assign n12753 = n12575 ^ n11802 ^ n5315 ;
  assign n12756 = n12755 ^ n12753 ^ n8688 ;
  assign n12757 = n12756 ^ n4634 ^ n2370 ;
  assign n12748 = n6398 & ~n10383 ;
  assign n12749 = n12748 ^ n6362 ^ 1'b0 ;
  assign n12746 = n7703 ^ n5754 ^ n1899 ;
  assign n12747 = n8844 & ~n12746 ;
  assign n12750 = n12749 ^ n12747 ^ 1'b0 ;
  assign n12745 = n4128 ^ n476 ^ 1'b0 ;
  assign n12751 = n12750 ^ n12745 ^ 1'b0 ;
  assign n12752 = n10574 & n12751 ;
  assign n12758 = n12757 ^ n12752 ^ 1'b0 ;
  assign n12759 = n4070 | n12758 ;
  assign n12760 = n6347 & ~n10638 ;
  assign n12761 = ( n11712 & n12759 ) | ( n11712 & ~n12760 ) | ( n12759 & ~n12760 ) ;
  assign n12764 = n9056 ^ n3082 ^ 1'b0 ;
  assign n12762 = ( n1159 & n4106 ) | ( n1159 & ~n4502 ) | ( n4106 & ~n4502 ) ;
  assign n12763 = ( n3505 & ~n11284 ) | ( n3505 & n12762 ) | ( ~n11284 & n12762 ) ;
  assign n12765 = n12764 ^ n12763 ^ 1'b0 ;
  assign n12766 = ~n8059 & n12765 ;
  assign n12767 = n9535 ^ n7939 ^ 1'b0 ;
  assign n12768 = n5616 & n12767 ;
  assign n12769 = ~n12122 & n12768 ;
  assign n12770 = n12769 ^ n3643 ^ 1'b0 ;
  assign n12771 = n12738 & n12770 ;
  assign n12772 = ~n4671 & n5640 ;
  assign n12773 = n355 & n12772 ;
  assign n12774 = n12773 ^ n7006 ^ 1'b0 ;
  assign n12775 = ( n7826 & n9525 ) | ( n7826 & n12774 ) | ( n9525 & n12774 ) ;
  assign n12776 = ~n3966 & n7185 ;
  assign n12777 = n8931 & ~n12776 ;
  assign n12778 = n288 | n12777 ;
  assign n12779 = ( n5084 & n7644 ) | ( n5084 & ~n8092 ) | ( n7644 & ~n8092 ) ;
  assign n12780 = n3908 ^ n3851 ^ n1076 ;
  assign n12781 = ( ~n9313 & n12598 ) | ( ~n9313 & n12780 ) | ( n12598 & n12780 ) ;
  assign n12782 = n5209 ^ n707 ^ 1'b0 ;
  assign n12783 = ( ~n409 & n12781 ) | ( ~n409 & n12782 ) | ( n12781 & n12782 ) ;
  assign n12784 = n10317 ^ n6558 ^ n1595 ;
  assign n12785 = ( n1131 & n8210 ) | ( n1131 & ~n12784 ) | ( n8210 & ~n12784 ) ;
  assign n12786 = ( n3860 & n3956 ) | ( n3860 & ~n10983 ) | ( n3956 & ~n10983 ) ;
  assign n12787 = n12786 ^ n5555 ^ n5284 ;
  assign n12788 = n4616 & ~n12310 ;
  assign n12789 = n12788 ^ n2422 ^ 1'b0 ;
  assign n12790 = n12789 ^ n1142 ^ 1'b0 ;
  assign n12791 = n5204 & n12790 ;
  assign n12792 = ~n5302 & n12791 ;
  assign n12793 = ( n11476 & n12787 ) | ( n11476 & n12792 ) | ( n12787 & n12792 ) ;
  assign n12794 = n12793 ^ n12586 ^ 1'b0 ;
  assign n12795 = n3065 & n9349 ;
  assign n12796 = ( n2964 & n8371 ) | ( n2964 & n12795 ) | ( n8371 & n12795 ) ;
  assign n12797 = n7569 & ~n12796 ;
  assign n12798 = n12797 ^ n7072 ^ 1'b0 ;
  assign n12805 = ~n2273 & n4130 ;
  assign n12806 = n9294 & n12805 ;
  assign n12807 = n5046 & n8827 ;
  assign n12808 = ( ~n4564 & n12806 ) | ( ~n4564 & n12807 ) | ( n12806 & n12807 ) ;
  assign n12799 = ~n574 & n5847 ;
  assign n12800 = n4089 & n12799 ;
  assign n12801 = n5017 ^ n4037 ^ n653 ;
  assign n12802 = n537 & n12272 ;
  assign n12803 = ( n12800 & ~n12801 ) | ( n12800 & n12802 ) | ( ~n12801 & n12802 ) ;
  assign n12804 = n12803 ^ n282 ^ 1'b0 ;
  assign n12809 = n12808 ^ n12804 ^ n3340 ;
  assign n12811 = n987 & ~n6245 ;
  assign n12812 = n12811 ^ n1883 ^ 1'b0 ;
  assign n12810 = ~n4322 & n11499 ;
  assign n12813 = n12812 ^ n12810 ^ 1'b0 ;
  assign n12816 = ( ~n2257 & n5599 ) | ( ~n2257 & n7949 ) | ( n5599 & n7949 ) ;
  assign n12815 = n10211 ^ n7574 ^ n5491 ;
  assign n12814 = n8443 ^ n5990 ^ n4352 ;
  assign n12817 = n12816 ^ n12815 ^ n12814 ;
  assign n12820 = ( n2864 & n3074 ) | ( n2864 & ~n6555 ) | ( n3074 & ~n6555 ) ;
  assign n12818 = n6272 ^ n4305 ^ n1274 ;
  assign n12819 = n2326 & n12818 ;
  assign n12821 = n12820 ^ n12819 ^ n336 ;
  assign n12822 = ( n5010 & n12460 ) | ( n5010 & n12707 ) | ( n12460 & n12707 ) ;
  assign n12823 = n9248 ^ n1385 ^ 1'b0 ;
  assign n12824 = n4570 & ~n5755 ;
  assign n12825 = n12823 & n12824 ;
  assign n12826 = ( ~n11298 & n11361 ) | ( ~n11298 & n12825 ) | ( n11361 & n12825 ) ;
  assign n12827 = n5118 & n11093 ;
  assign n12828 = ~n6422 & n12827 ;
  assign n12829 = ~n3557 & n6473 ;
  assign n12830 = n12829 ^ n1371 ^ 1'b0 ;
  assign n12831 = ( n7866 & ~n8523 ) | ( n7866 & n12830 ) | ( ~n8523 & n12830 ) ;
  assign n12832 = n12831 ^ n5218 ^ n3987 ;
  assign n12833 = n10672 ^ n4933 ^ 1'b0 ;
  assign n12834 = n12833 ^ n5815 ^ 1'b0 ;
  assign n12835 = n5030 & ~n11304 ;
  assign n12836 = n12835 ^ n5251 ^ 1'b0 ;
  assign n12837 = n12836 ^ n4137 ^ n3061 ;
  assign n12838 = n9962 ^ n7402 ^ n6437 ;
  assign n12839 = ~n7575 & n12838 ;
  assign n12840 = n10255 ^ n2186 ^ 1'b0 ;
  assign n12856 = n7774 ^ n6067 ^ 1'b0 ;
  assign n12857 = n4536 & n12856 ;
  assign n12848 = ( n860 & n1873 ) | ( n860 & n4510 ) | ( n1873 & n4510 ) ;
  assign n12849 = n12848 ^ n10437 ^ n9387 ;
  assign n12850 = n5465 ^ n5233 ^ n3368 ;
  assign n12851 = n12849 | n12850 ;
  assign n12852 = n6307 ^ n5638 ^ x54 ;
  assign n12853 = n12852 ^ n10189 ^ n6622 ;
  assign n12854 = n12851 & ~n12853 ;
  assign n12855 = n12854 ^ n5138 ^ 1'b0 ;
  assign n12844 = n7645 ^ n3170 ^ 1'b0 ;
  assign n12845 = n12844 ^ n5897 ^ n4812 ;
  assign n12846 = n12845 ^ n8194 ^ n5293 ;
  assign n12842 = n10951 ^ n6490 ^ n3786 ;
  assign n12843 = n12842 ^ n491 ^ x108 ;
  assign n12841 = ( n2475 & ~n2630 ) | ( n2475 & n3658 ) | ( ~n2630 & n3658 ) ;
  assign n12847 = n12846 ^ n12843 ^ n12841 ;
  assign n12858 = n12857 ^ n12855 ^ n12847 ;
  assign n12859 = ( n1152 & n12840 ) | ( n1152 & n12858 ) | ( n12840 & n12858 ) ;
  assign n12860 = n11534 ^ n8324 ^ n2372 ;
  assign n12863 = n10074 ^ n5367 ^ n395 ;
  assign n12862 = n2302 & n4035 ;
  assign n12864 = n12863 ^ n12862 ^ 1'b0 ;
  assign n12861 = n6277 & ~n7279 ;
  assign n12865 = n12864 ^ n12861 ^ 1'b0 ;
  assign n12866 = ~n12860 & n12865 ;
  assign n12867 = n12193 ^ n7065 ^ 1'b0 ;
  assign n12868 = n12867 ^ n8612 ^ n370 ;
  assign n12869 = n4226 & ~n6841 ;
  assign n12870 = n3307 & n12869 ;
  assign n12871 = n9886 & n12870 ;
  assign n12876 = n666 & ~n11311 ;
  assign n12877 = n3220 | n12876 ;
  assign n12878 = n3209 | n12877 ;
  assign n12879 = n421 & n12878 ;
  assign n12880 = n12879 ^ n6139 ^ 1'b0 ;
  assign n12881 = n10540 ^ n5736 ^ 1'b0 ;
  assign n12882 = ~n6937 & n12881 ;
  assign n12883 = n12246 ^ n4046 ^ n2341 ;
  assign n12884 = ( n12880 & ~n12882 ) | ( n12880 & n12883 ) | ( ~n12882 & n12883 ) ;
  assign n12872 = n1552 & ~n6640 ;
  assign n12873 = n3907 & n12872 ;
  assign n12874 = n12873 ^ n6849 ^ 1'b0 ;
  assign n12875 = ( ~n2699 & n2793 ) | ( ~n2699 & n12874 ) | ( n2793 & n12874 ) ;
  assign n12885 = n12884 ^ n12875 ^ 1'b0 ;
  assign n12890 = n2369 ^ n1386 ^ n899 ;
  assign n12888 = n7815 ^ n1143 ^ 1'b0 ;
  assign n12889 = n1319 & n12888 ;
  assign n12886 = n6270 | n8002 ;
  assign n12887 = ( n8146 & ~n8752 ) | ( n8146 & n12886 ) | ( ~n8752 & n12886 ) ;
  assign n12891 = n12890 ^ n12889 ^ n12887 ;
  assign n12892 = n9857 | n10896 ;
  assign n12893 = n2740 & ~n12892 ;
  assign n12894 = n12893 ^ n12234 ^ 1'b0 ;
  assign n12895 = n12894 ^ n11485 ^ n6029 ;
  assign n12896 = n2854 & ~n6456 ;
  assign n12897 = ~n4032 & n12896 ;
  assign n12899 = n869 ^ n452 ^ x201 ;
  assign n12900 = n633 & ~n1597 ;
  assign n12901 = ~n2517 & n12900 ;
  assign n12902 = ( n4631 & n12899 ) | ( n4631 & ~n12901 ) | ( n12899 & ~n12901 ) ;
  assign n12898 = ( n1852 & n3171 ) | ( n1852 & ~n5476 ) | ( n3171 & ~n5476 ) ;
  assign n12903 = n12902 ^ n12898 ^ 1'b0 ;
  assign n12906 = n10797 ^ n7884 ^ n7163 ;
  assign n12907 = ( n6768 & n7185 ) | ( n6768 & n12906 ) | ( n7185 & n12906 ) ;
  assign n12904 = n7728 ^ n2096 ^ 1'b0 ;
  assign n12905 = n438 | n12904 ;
  assign n12908 = n12907 ^ n12905 ^ 1'b0 ;
  assign n12909 = x10 & ~n12908 ;
  assign n12910 = n8027 | n12909 ;
  assign n12911 = ( ~n9877 & n12903 ) | ( ~n9877 & n12910 ) | ( n12903 & n12910 ) ;
  assign n12912 = n9256 ^ n6789 ^ 1'b0 ;
  assign n12913 = n4003 & n5146 ;
  assign n12914 = n12913 ^ n1358 ^ 1'b0 ;
  assign n12915 = n12914 ^ n10267 ^ 1'b0 ;
  assign n12916 = n12239 ^ x241 ^ 1'b0 ;
  assign n12920 = n2566 ^ n1377 ^ n1117 ;
  assign n12917 = n8139 ^ n2943 ^ 1'b0 ;
  assign n12918 = n12917 ^ n5923 ^ 1'b0 ;
  assign n12919 = n6465 | n12918 ;
  assign n12921 = n12920 ^ n12919 ^ n5258 ;
  assign n12925 = n433 & ~n1868 ;
  assign n12926 = n12925 ^ n1653 ^ 1'b0 ;
  assign n12923 = n8844 & ~n11599 ;
  assign n12924 = n1532 & n12923 ;
  assign n12927 = n12926 ^ n12924 ^ n3814 ;
  assign n12922 = n3575 ^ n2058 ^ n556 ;
  assign n12928 = n12927 ^ n12922 ^ 1'b0 ;
  assign n12929 = n12928 ^ n5671 ^ n1982 ;
  assign n12930 = n12929 ^ n7149 ^ n1090 ;
  assign n12931 = ( n4844 & ~n7400 ) | ( n4844 & n12146 ) | ( ~n7400 & n12146 ) ;
  assign n12932 = n5311 & n8328 ;
  assign n12933 = ( n11892 & n12931 ) | ( n11892 & ~n12932 ) | ( n12931 & ~n12932 ) ;
  assign n12934 = ~n2994 & n12328 ;
  assign n12935 = ~n1104 & n12934 ;
  assign n12936 = ( n2020 & n9251 ) | ( n2020 & ~n10399 ) | ( n9251 & ~n10399 ) ;
  assign n12937 = n12936 ^ n12512 ^ n5797 ;
  assign n12939 = n1496 | n7813 ;
  assign n12940 = n12939 ^ n5309 ^ n562 ;
  assign n12938 = n12649 ^ n1198 ^ n913 ;
  assign n12941 = n12940 ^ n12938 ^ 1'b0 ;
  assign n12942 = n578 & ~n6545 ;
  assign n12943 = ~n6908 & n12942 ;
  assign n12956 = ~n988 & n3271 ;
  assign n12958 = ~n740 & n6132 ;
  assign n12959 = n12958 ^ n2999 ^ 1'b0 ;
  assign n12957 = n8156 ^ n6557 ^ 1'b0 ;
  assign n12960 = n12959 ^ n12957 ^ 1'b0 ;
  assign n12961 = ~n8882 & n12960 ;
  assign n12962 = n12956 & n12961 ;
  assign n12963 = ~n4306 & n12962 ;
  assign n12946 = n5307 ^ n4158 ^ n1866 ;
  assign n12949 = ( n733 & n1586 ) | ( n733 & ~n1634 ) | ( n1586 & ~n1634 ) ;
  assign n12947 = n3096 & n6073 ;
  assign n12948 = n12947 ^ n4069 ^ n2719 ;
  assign n12950 = n12949 ^ n12948 ^ n4849 ;
  assign n12951 = n12950 ^ n8138 ^ 1'b0 ;
  assign n12952 = ( n2132 & n10139 ) | ( n2132 & n12951 ) | ( n10139 & n12951 ) ;
  assign n12953 = n2362 & n7504 ;
  assign n12954 = ( n3888 & n12952 ) | ( n3888 & n12953 ) | ( n12952 & n12953 ) ;
  assign n12955 = ( ~n12187 & n12946 ) | ( ~n12187 & n12954 ) | ( n12946 & n12954 ) ;
  assign n12944 = n5593 ^ n3617 ^ n1124 ;
  assign n12945 = ( n6461 & n6886 ) | ( n6461 & n12944 ) | ( n6886 & n12944 ) ;
  assign n12964 = n12963 ^ n12955 ^ n12945 ;
  assign n12966 = n11631 ^ n8539 ^ n501 ;
  assign n12965 = n11433 ^ n2488 ^ 1'b0 ;
  assign n12967 = n12966 ^ n12965 ^ n12461 ;
  assign n12969 = n7353 ^ n6607 ^ 1'b0 ;
  assign n12970 = n12969 ^ n4935 ^ n3707 ;
  assign n12971 = n3452 & ~n12970 ;
  assign n12972 = n12971 ^ n6810 ^ 1'b0 ;
  assign n12968 = n11940 ^ n6164 ^ x6 ;
  assign n12973 = n12972 ^ n12968 ^ n12424 ;
  assign n12974 = n6109 ^ n1868 ^ 1'b0 ;
  assign n12975 = n12948 | n12974 ;
  assign n12979 = ( ~n664 & n2719 ) | ( ~n664 & n8014 ) | ( n2719 & n8014 ) ;
  assign n12976 = n6888 ^ n431 ^ 1'b0 ;
  assign n12977 = ~n10229 & n12976 ;
  assign n12978 = ~n5955 & n12977 ;
  assign n12980 = n12979 ^ n12978 ^ 1'b0 ;
  assign n12981 = ~n12975 & n12980 ;
  assign n12982 = n12981 ^ n9348 ^ 1'b0 ;
  assign n12983 = n6018 & ~n6268 ;
  assign n12984 = n3679 ^ n3152 ^ n912 ;
  assign n12985 = n12984 ^ n4067 ^ 1'b0 ;
  assign n12987 = ~n1848 & n8360 ;
  assign n12986 = n11356 ^ n3399 ^ n1823 ;
  assign n12988 = n12987 ^ n12986 ^ n786 ;
  assign n12989 = ( n490 & ~n12985 ) | ( n490 & n12988 ) | ( ~n12985 & n12988 ) ;
  assign n12990 = n1454 & n11024 ;
  assign n12991 = n9361 & n12990 ;
  assign n12992 = n5418 ^ n2522 ^ n708 ;
  assign n12996 = n8264 ^ n3192 ^ 1'b0 ;
  assign n12997 = ~n6558 & n12996 ;
  assign n12994 = n6394 ^ n2803 ^ 1'b0 ;
  assign n12995 = n969 & n12994 ;
  assign n12993 = n12105 ^ n11320 ^ 1'b0 ;
  assign n12998 = n12997 ^ n12995 ^ n12993 ;
  assign n12999 = ( n6592 & ~n12992 ) | ( n6592 & n12998 ) | ( ~n12992 & n12998 ) ;
  assign n13000 = n4933 ^ n4623 ^ n2995 ;
  assign n13001 = n5457 ^ n5020 ^ 1'b0 ;
  assign n13002 = n9815 ^ n7218 ^ 1'b0 ;
  assign n13003 = ( n13000 & n13001 ) | ( n13000 & ~n13002 ) | ( n13001 & ~n13002 ) ;
  assign n13004 = n7001 ^ n4006 ^ 1'b0 ;
  assign n13005 = ~n13003 & n13004 ;
  assign n13006 = n3679 | n9502 ;
  assign n13007 = ( n575 & n2058 ) | ( n575 & ~n5525 ) | ( n2058 & ~n5525 ) ;
  assign n13008 = n13007 ^ n11999 ^ x156 ;
  assign n13009 = n12236 ^ n6817 ^ x34 ;
  assign n13010 = ~n11742 & n13009 ;
  assign n13011 = n13008 & n13010 ;
  assign n13012 = n2004 | n9698 ;
  assign n13013 = n9701 & n13012 ;
  assign n13014 = n8839 & n9911 ;
  assign n13015 = ~n10431 & n13014 ;
  assign n13016 = n1055 | n2334 ;
  assign n13017 = n13016 ^ n12320 ^ n1391 ;
  assign n13018 = ( n2515 & n13015 ) | ( n2515 & ~n13017 ) | ( n13015 & ~n13017 ) ;
  assign n13020 = ( n865 & n4190 ) | ( n865 & ~n6149 ) | ( n4190 & ~n6149 ) ;
  assign n13021 = x226 & n13020 ;
  assign n13022 = n13021 ^ n3512 ^ 1'b0 ;
  assign n13019 = n6383 ^ n5280 ^ n2849 ;
  assign n13023 = n13022 ^ n13019 ^ n3331 ;
  assign n13024 = n13023 ^ n5256 ^ n1573 ;
  assign n13025 = ( ~n4161 & n7281 ) | ( ~n4161 & n11942 ) | ( n7281 & n11942 ) ;
  assign n13026 = ( ~n3722 & n4601 ) | ( ~n3722 & n5259 ) | ( n4601 & n5259 ) ;
  assign n13027 = ( n3598 & n5892 ) | ( n3598 & n13026 ) | ( n5892 & n13026 ) ;
  assign n13028 = n13027 ^ n3900 ^ n1652 ;
  assign n13029 = ~n3291 & n6136 ;
  assign n13030 = n13029 ^ n6453 ^ 1'b0 ;
  assign n13031 = n12146 ^ n6488 ^ n903 ;
  assign n13032 = n13031 ^ n5538 ^ n2941 ;
  assign n13033 = ( ~n13028 & n13030 ) | ( ~n13028 & n13032 ) | ( n13030 & n13032 ) ;
  assign n13034 = ( n331 & ~n7827 ) | ( n331 & n13033 ) | ( ~n7827 & n13033 ) ;
  assign n13035 = n10815 ^ n7685 ^ n2960 ;
  assign n13036 = ~n1695 & n4179 ;
  assign n13037 = n13036 ^ n3950 ^ 1'b0 ;
  assign n13038 = n2402 ^ n1219 ^ n716 ;
  assign n13039 = n7568 & n13038 ;
  assign n13040 = n13037 & n13039 ;
  assign n13046 = n7053 | n8866 ;
  assign n13047 = n1769 | n13046 ;
  assign n13041 = ~n1625 & n6855 ;
  assign n13042 = ~x42 & n13041 ;
  assign n13043 = n13042 ^ n6654 ^ x234 ;
  assign n13044 = n13043 ^ n7416 ^ 1'b0 ;
  assign n13045 = ~n1882 & n13044 ;
  assign n13048 = n13047 ^ n13045 ^ x100 ;
  assign n13049 = n10561 ^ n6997 ^ 1'b0 ;
  assign n13050 = ( ~n2103 & n5583 ) | ( ~n2103 & n8206 ) | ( n5583 & n8206 ) ;
  assign n13051 = ( n501 & n8613 ) | ( n501 & n13050 ) | ( n8613 & n13050 ) ;
  assign n13056 = x134 & n4601 ;
  assign n13057 = n11244 & n13056 ;
  assign n13052 = n8519 ^ n1897 ^ 1'b0 ;
  assign n13053 = n13052 ^ n3381 ^ 1'b0 ;
  assign n13054 = ~n11411 & n12350 ;
  assign n13055 = ~n13053 & n13054 ;
  assign n13058 = n13057 ^ n13055 ^ n9660 ;
  assign n13059 = ( n6887 & n13042 ) | ( n6887 & n13058 ) | ( n13042 & n13058 ) ;
  assign n13060 = ( n1366 & ~n5119 ) | ( n1366 & n6167 ) | ( ~n5119 & n6167 ) ;
  assign n13061 = n13060 ^ n5654 ^ 1'b0 ;
  assign n13062 = ~n7563 & n13061 ;
  assign n13063 = n8962 ^ n6283 ^ 1'b0 ;
  assign n13064 = ( n10721 & n13062 ) | ( n10721 & ~n13063 ) | ( n13062 & ~n13063 ) ;
  assign n13065 = n8813 ^ n6577 ^ n2070 ;
  assign n13066 = n1946 | n13065 ;
  assign n13067 = ( n8242 & n9650 ) | ( n8242 & n13066 ) | ( n9650 & n13066 ) ;
  assign n13068 = n13067 ^ n1173 ^ 1'b0 ;
  assign n13073 = n9039 & ~n9273 ;
  assign n13074 = n13073 ^ n2927 ^ 1'b0 ;
  assign n13072 = n11886 ^ n11533 ^ n6666 ;
  assign n13069 = ( x92 & ~n1463 ) | ( x92 & n1915 ) | ( ~n1463 & n1915 ) ;
  assign n13070 = n13069 ^ x207 ^ 1'b0 ;
  assign n13071 = ( n2465 & n5957 ) | ( n2465 & n13070 ) | ( n5957 & n13070 ) ;
  assign n13075 = n13074 ^ n13072 ^ n13071 ;
  assign n13079 = ( ~n527 & n10021 ) | ( ~n527 & n11780 ) | ( n10021 & n11780 ) ;
  assign n13080 = n13079 ^ n4457 ^ 1'b0 ;
  assign n13076 = ( n3180 & ~n4017 ) | ( n3180 & n9230 ) | ( ~n4017 & n9230 ) ;
  assign n13077 = ( n523 & n10022 ) | ( n523 & n13076 ) | ( n10022 & n13076 ) ;
  assign n13078 = n13077 ^ n11840 ^ n8900 ;
  assign n13081 = n13080 ^ n13078 ^ 1'b0 ;
  assign n13082 = n1093 & ~n7671 ;
  assign n13083 = ( n7461 & n9019 ) | ( n7461 & n13082 ) | ( n9019 & n13082 ) ;
  assign n13084 = n9579 ^ n2085 ^ n1052 ;
  assign n13085 = ( n7568 & ~n10947 ) | ( n7568 & n13084 ) | ( ~n10947 & n13084 ) ;
  assign n13086 = n2080 ^ n384 ^ 1'b0 ;
  assign n13087 = n12438 | n13086 ;
  assign n13088 = n2823 & ~n13087 ;
  assign n13089 = n504 & ~n4109 ;
  assign n13090 = n1431 & n13089 ;
  assign n13091 = ( n2552 & n3251 ) | ( n2552 & ~n4880 ) | ( n3251 & ~n4880 ) ;
  assign n13092 = n4762 & ~n13091 ;
  assign n13093 = n7022 ^ n284 ^ 1'b0 ;
  assign n13094 = ~n2888 & n13093 ;
  assign n13095 = ~n13092 & n13094 ;
  assign n13096 = n13090 & n13095 ;
  assign n13097 = n3391 & ~n13096 ;
  assign n13098 = n317 & n6869 ;
  assign n13099 = ( n1278 & n11599 ) | ( n1278 & n13098 ) | ( n11599 & n13098 ) ;
  assign n13100 = ( n1599 & ~n3508 ) | ( n1599 & n8694 ) | ( ~n3508 & n8694 ) ;
  assign n13101 = ( n6351 & n9083 ) | ( n6351 & n13100 ) | ( n9083 & n13100 ) ;
  assign n13102 = ~n3327 & n11591 ;
  assign n13103 = ~x21 & n13102 ;
  assign n13104 = x41 & ~n8367 ;
  assign n13105 = ~n13103 & n13104 ;
  assign n13106 = ~n11378 & n13105 ;
  assign n13107 = ( n5078 & n11427 ) | ( n5078 & n13106 ) | ( n11427 & n13106 ) ;
  assign n13108 = n2717 & ~n12975 ;
  assign n13109 = n2797 & n13108 ;
  assign n13110 = n13109 ^ n562 ^ 1'b0 ;
  assign n13111 = ( ~n1771 & n8232 ) | ( ~n1771 & n13110 ) | ( n8232 & n13110 ) ;
  assign n13112 = n11004 & n13111 ;
  assign n13113 = n13112 ^ n2437 ^ 1'b0 ;
  assign n13114 = ( ~n2162 & n3082 ) | ( ~n2162 & n12280 ) | ( n3082 & n12280 ) ;
  assign n13115 = n5955 | n13114 ;
  assign n13116 = n13115 ^ n10808 ^ 1'b0 ;
  assign n13117 = ( n4541 & n6752 ) | ( n4541 & n13116 ) | ( n6752 & n13116 ) ;
  assign n13118 = n13117 ^ n9962 ^ n7569 ;
  assign n13119 = n6602 | n11969 ;
  assign n13120 = ( ~n1085 & n4161 ) | ( ~n1085 & n10807 ) | ( n4161 & n10807 ) ;
  assign n13121 = n5164 ^ n4026 ^ x135 ;
  assign n13122 = ( n8235 & n12898 ) | ( n8235 & n13121 ) | ( n12898 & n13121 ) ;
  assign n13123 = n9490 ^ n5347 ^ n4815 ;
  assign n13124 = n13123 ^ n10467 ^ n962 ;
  assign n13125 = ( n6759 & n9589 ) | ( n6759 & n11959 ) | ( n9589 & n11959 ) ;
  assign n13126 = n9931 | n13125 ;
  assign n13127 = n13126 ^ n2462 ^ 1'b0 ;
  assign n13128 = n13127 ^ n5282 ^ n1581 ;
  assign n13129 = n8369 ^ n1131 ^ 1'b0 ;
  assign n13135 = n11639 ^ n5351 ^ n3722 ;
  assign n13136 = n13135 ^ n2422 ^ x131 ;
  assign n13130 = ( n5000 & n7457 ) | ( n5000 & ~n8455 ) | ( n7457 & ~n8455 ) ;
  assign n13131 = ( ~n4147 & n6670 ) | ( ~n4147 & n13130 ) | ( n6670 & n13130 ) ;
  assign n13132 = x48 & n13131 ;
  assign n13133 = n6184 & ~n11317 ;
  assign n13134 = ~n13132 & n13133 ;
  assign n13137 = n13136 ^ n13134 ^ 1'b0 ;
  assign n13138 = n1653 ^ n1246 ^ 1'b0 ;
  assign n13139 = ( ~n3381 & n9794 ) | ( ~n3381 & n13138 ) | ( n9794 & n13138 ) ;
  assign n13140 = n6669 ^ n5802 ^ x193 ;
  assign n13141 = ( n6825 & n13139 ) | ( n6825 & ~n13140 ) | ( n13139 & ~n13140 ) ;
  assign n13142 = n5149 & n11323 ;
  assign n13143 = n13142 ^ n4029 ^ 1'b0 ;
  assign n13151 = n2018 | n7389 ;
  assign n13152 = n4574 & ~n13151 ;
  assign n13145 = ( ~n563 & n2525 ) | ( ~n563 & n9106 ) | ( n2525 & n9106 ) ;
  assign n13146 = n3629 | n7382 ;
  assign n13147 = n7808 & ~n9023 ;
  assign n13148 = n13146 & n13147 ;
  assign n13149 = ( n8088 & n13145 ) | ( n8088 & n13148 ) | ( n13145 & n13148 ) ;
  assign n13144 = n12310 ^ n8265 ^ n4781 ;
  assign n13150 = n13149 ^ n13144 ^ n6103 ;
  assign n13153 = n13152 ^ n13150 ^ 1'b0 ;
  assign n13154 = n11045 ^ n3786 ^ n1095 ;
  assign n13155 = ( n6646 & n8936 ) | ( n6646 & n13154 ) | ( n8936 & n13154 ) ;
  assign n13156 = n2055 & n3728 ;
  assign n13157 = n5202 & n13156 ;
  assign n13158 = n12786 ^ n2538 ^ 1'b0 ;
  assign n13159 = n4256 | n13158 ;
  assign n13160 = ~n2332 & n8971 ;
  assign n13161 = ~n1539 & n13160 ;
  assign n13162 = ( n1064 & n4322 ) | ( n1064 & n13161 ) | ( n4322 & n13161 ) ;
  assign n13163 = ( n1653 & ~n7509 ) | ( n1653 & n13162 ) | ( ~n7509 & n13162 ) ;
  assign n13164 = n11266 & ~n13163 ;
  assign n13165 = n13159 & n13164 ;
  assign n13166 = n1345 ^ n1305 ^ 1'b0 ;
  assign n13167 = ( ~n1312 & n9569 ) | ( ~n1312 & n13166 ) | ( n9569 & n13166 ) ;
  assign n13168 = n12111 ^ n2422 ^ 1'b0 ;
  assign n13169 = n7891 | n13168 ;
  assign n13172 = n3550 ^ n2664 ^ n1079 ;
  assign n13171 = ( n2893 & n3767 ) | ( n2893 & n6803 ) | ( n3767 & n6803 ) ;
  assign n13173 = n13172 ^ n13171 ^ n9639 ;
  assign n13170 = n2189 ^ n1576 ^ x243 ;
  assign n13174 = n13173 ^ n13170 ^ n6130 ;
  assign n13177 = ~n2610 & n8370 ;
  assign n13178 = ~n2118 & n13177 ;
  assign n13179 = ( n5478 & ~n7713 ) | ( n5478 & n13178 ) | ( ~n7713 & n13178 ) ;
  assign n13175 = ~n4376 & n10418 ;
  assign n13176 = n13175 ^ n2066 ^ 1'b0 ;
  assign n13180 = n13179 ^ n13176 ^ n11029 ;
  assign n13181 = n10303 ^ n1130 ^ 1'b0 ;
  assign n13182 = n3488 | n13181 ;
  assign n13183 = n11774 | n13182 ;
  assign n13184 = ( n2193 & ~n8944 ) | ( n2193 & n13183 ) | ( ~n8944 & n13183 ) ;
  assign n13185 = ( n8000 & n13180 ) | ( n8000 & ~n13184 ) | ( n13180 & ~n13184 ) ;
  assign n13186 = n9811 ^ n1248 ^ n620 ;
  assign n13187 = n13186 ^ n10152 ^ n9901 ;
  assign n13188 = ( n3411 & ~n12757 ) | ( n3411 & n13187 ) | ( ~n12757 & n13187 ) ;
  assign n13189 = n6944 ^ n5864 ^ 1'b0 ;
  assign n13195 = n10152 ^ x43 ^ 1'b0 ;
  assign n13192 = n8372 ^ n1513 ^ 1'b0 ;
  assign n13193 = n7176 & ~n13192 ;
  assign n13190 = n6781 ^ n6632 ^ 1'b0 ;
  assign n13191 = ( n2996 & n9223 ) | ( n2996 & ~n13190 ) | ( n9223 & ~n13190 ) ;
  assign n13194 = n13193 ^ n13191 ^ n12132 ;
  assign n13196 = n13195 ^ n13194 ^ n1855 ;
  assign n13197 = ( ~n4438 & n9012 ) | ( ~n4438 & n13196 ) | ( n9012 & n13196 ) ;
  assign n13198 = n13189 & ~n13197 ;
  assign n13199 = ( n2705 & n6387 ) | ( n2705 & ~n8519 ) | ( n6387 & ~n8519 ) ;
  assign n13203 = ( n3184 & n3486 ) | ( n3184 & ~n12191 ) | ( n3486 & ~n12191 ) ;
  assign n13200 = ( n1077 & n2788 ) | ( n1077 & ~n10835 ) | ( n2788 & ~n10835 ) ;
  assign n13201 = n13200 ^ n5950 ^ 1'b0 ;
  assign n13202 = ~n8577 & n13201 ;
  assign n13204 = n13203 ^ n13202 ^ 1'b0 ;
  assign n13213 = ( n2882 & n6887 ) | ( n2882 & ~n8239 ) | ( n6887 & ~n8239 ) ;
  assign n13209 = n2589 & n5174 ;
  assign n13210 = ( n4330 & n10703 ) | ( n4330 & n13209 ) | ( n10703 & n13209 ) ;
  assign n13211 = n8383 ^ n6583 ^ 1'b0 ;
  assign n13212 = n13210 | n13211 ;
  assign n13205 = n4627 ^ n1801 ^ 1'b0 ;
  assign n13206 = ( n3443 & ~n9449 ) | ( n3443 & n11274 ) | ( ~n9449 & n11274 ) ;
  assign n13207 = n13206 ^ n9917 ^ n4902 ;
  assign n13208 = ( ~n318 & n13205 ) | ( ~n318 & n13207 ) | ( n13205 & n13207 ) ;
  assign n13214 = n13213 ^ n13212 ^ n13208 ;
  assign n13215 = n7758 & n12427 ;
  assign n13216 = ~n2382 & n6361 ;
  assign n13217 = n13216 ^ n3482 ^ 1'b0 ;
  assign n13218 = n12739 | n13217 ;
  assign n13219 = n3092 | n13218 ;
  assign n13220 = n9131 ^ n5267 ^ n4216 ;
  assign n13221 = n13220 ^ n8406 ^ n8348 ;
  assign n13222 = ( x173 & n13219 ) | ( x173 & ~n13221 ) | ( n13219 & ~n13221 ) ;
  assign n13223 = ~n473 & n5562 ;
  assign n13224 = ( ~n902 & n4925 ) | ( ~n902 & n13223 ) | ( n4925 & n13223 ) ;
  assign n13225 = n13224 ^ n6644 ^ 1'b0 ;
  assign n13226 = ( n2824 & n10200 ) | ( n2824 & n13225 ) | ( n10200 & n13225 ) ;
  assign n13227 = n10954 ^ n1310 ^ 1'b0 ;
  assign n13228 = n8561 & n13227 ;
  assign n13229 = ( n1132 & ~n2010 ) | ( n1132 & n13228 ) | ( ~n2010 & n13228 ) ;
  assign n13230 = n12156 ^ n4136 ^ 1'b0 ;
  assign n13231 = n11073 & ~n13230 ;
  assign n13232 = n13231 ^ n12484 ^ n995 ;
  assign n13233 = ( n6468 & ~n11929 ) | ( n6468 & n13232 ) | ( ~n11929 & n13232 ) ;
  assign n13234 = n353 | n3280 ;
  assign n13235 = n5184 | n13234 ;
  assign n13236 = n13235 ^ n9669 ^ 1'b0 ;
  assign n13237 = n8130 & ~n10453 ;
  assign n13238 = n8267 ^ n6983 ^ n805 ;
  assign n13249 = ( n3051 & n9040 ) | ( n3051 & n10394 ) | ( n9040 & n10394 ) ;
  assign n13250 = ( n4323 & n8383 ) | ( n4323 & ~n13249 ) | ( n8383 & ~n13249 ) ;
  assign n13241 = n13231 ^ n1605 ^ 1'b0 ;
  assign n13242 = ~n3204 & n13241 ;
  assign n13240 = ~n5576 & n10150 ;
  assign n13243 = n13242 ^ n13240 ^ 1'b0 ;
  assign n13239 = n2666 & ~n5637 ;
  assign n13244 = n13243 ^ n13239 ^ 1'b0 ;
  assign n13245 = n6193 & ~n7814 ;
  assign n13246 = n11533 & n13245 ;
  assign n13247 = n13246 ^ n7523 ^ 1'b0 ;
  assign n13248 = ( n11214 & ~n13244 ) | ( n11214 & n13247 ) | ( ~n13244 & n13247 ) ;
  assign n13251 = n13250 ^ n13248 ^ n1901 ;
  assign n13252 = n13238 & n13251 ;
  assign n13253 = ~n615 & n13252 ;
  assign n13258 = ( n757 & n1452 ) | ( n757 & n3747 ) | ( n1452 & n3747 ) ;
  assign n13254 = n1189 ^ n423 ^ 1'b0 ;
  assign n13255 = n2010 & n13254 ;
  assign n13256 = ~n1122 & n13255 ;
  assign n13257 = n2865 & n13256 ;
  assign n13259 = n13258 ^ n13257 ^ 1'b0 ;
  assign n13260 = n4067 | n13259 ;
  assign n13261 = ~n983 & n4921 ;
  assign n13262 = ( n8089 & ~n10041 ) | ( n8089 & n12807 ) | ( ~n10041 & n12807 ) ;
  assign n13284 = n4470 ^ n3806 ^ 1'b0 ;
  assign n13283 = ~n3054 & n12002 ;
  assign n13285 = n13284 ^ n13283 ^ 1'b0 ;
  assign n13286 = n13285 ^ n13208 ^ 1'b0 ;
  assign n13279 = ( ~n1475 & n4115 ) | ( ~n1475 & n8096 ) | ( n4115 & n8096 ) ;
  assign n13269 = n460 & ~n2515 ;
  assign n13270 = n13269 ^ n5147 ^ 1'b0 ;
  assign n13271 = n4000 & n5201 ;
  assign n13272 = n13270 & n13271 ;
  assign n13273 = n13272 ^ n4203 ^ n3385 ;
  assign n13274 = ( n7544 & n8034 ) | ( n7544 & ~n13273 ) | ( n8034 & ~n13273 ) ;
  assign n13275 = ( ~n5411 & n12230 ) | ( ~n5411 & n13274 ) | ( n12230 & n13274 ) ;
  assign n13276 = n13275 ^ n1325 ^ 1'b0 ;
  assign n13277 = n866 & n13276 ;
  assign n13278 = n12551 & n13277 ;
  assign n13280 = n13279 ^ n13278 ^ 1'b0 ;
  assign n13281 = n13280 ^ n10034 ^ 1'b0 ;
  assign n13282 = n6118 & n13281 ;
  assign n13263 = n6653 ^ n4576 ^ n1481 ;
  assign n13264 = n4282 ^ n1764 ^ 1'b0 ;
  assign n13265 = ( n7635 & n13263 ) | ( n7635 & ~n13264 ) | ( n13263 & ~n13264 ) ;
  assign n13266 = ( n1218 & n4064 ) | ( n1218 & ~n13020 ) | ( n4064 & ~n13020 ) ;
  assign n13267 = n6405 & ~n13266 ;
  assign n13268 = ( n12221 & n13265 ) | ( n12221 & n13267 ) | ( n13265 & n13267 ) ;
  assign n13287 = n13286 ^ n13282 ^ n13268 ;
  assign n13288 = n8525 ^ n5581 ^ n907 ;
  assign n13289 = ( n6136 & n8882 ) | ( n6136 & ~n9379 ) | ( n8882 & ~n9379 ) ;
  assign n13298 = n5777 ^ n4760 ^ 1'b0 ;
  assign n13290 = ~n802 & n2621 ;
  assign n13291 = n13290 ^ n1983 ^ 1'b0 ;
  assign n13292 = ( n1534 & n1736 ) | ( n1534 & ~n4060 ) | ( n1736 & ~n4060 ) ;
  assign n13293 = ~n1695 & n13292 ;
  assign n13294 = n10619 & n13293 ;
  assign n13295 = n4994 ^ n4902 ^ 1'b0 ;
  assign n13296 = ~n13294 & n13295 ;
  assign n13297 = ~n13291 & n13296 ;
  assign n13299 = n13298 ^ n13297 ^ 1'b0 ;
  assign n13300 = n10792 | n13299 ;
  assign n13301 = n13300 ^ n6918 ^ 1'b0 ;
  assign n13304 = n2021 & n2618 ;
  assign n13302 = n5231 ^ n3754 ^ 1'b0 ;
  assign n13303 = ( n2980 & ~n3659 ) | ( n2980 & n13302 ) | ( ~n3659 & n13302 ) ;
  assign n13305 = n13304 ^ n13303 ^ n3583 ;
  assign n13310 = n10446 ^ n3530 ^ n1453 ;
  assign n13308 = ( n2860 & n6373 ) | ( n2860 & n10101 ) | ( n6373 & n10101 ) ;
  assign n13306 = n6937 | n9283 ;
  assign n13307 = ( n1537 & n3999 ) | ( n1537 & ~n13306 ) | ( n3999 & ~n13306 ) ;
  assign n13309 = n13308 ^ n13307 ^ n7075 ;
  assign n13311 = n13310 ^ n13309 ^ n10230 ;
  assign n13312 = n13310 ^ n9830 ^ n8860 ;
  assign n13313 = n507 & ~n5880 ;
  assign n13314 = ~n9357 & n13313 ;
  assign n13315 = n5905 ^ n3633 ^ n895 ;
  assign n13316 = ~n13314 & n13315 ;
  assign n13317 = n9154 & n13316 ;
  assign n13319 = n4685 ^ x242 ^ 1'b0 ;
  assign n13320 = n12073 | n13319 ;
  assign n13321 = n13320 ^ n1050 ^ 1'b0 ;
  assign n13318 = n7056 & ~n8169 ;
  assign n13322 = n13321 ^ n13318 ^ n7980 ;
  assign n13323 = ( ~n5147 & n12447 ) | ( ~n5147 & n13322 ) | ( n12447 & n13322 ) ;
  assign n13324 = n665 & ~n2442 ;
  assign n13325 = n5175 & n13324 ;
  assign n13326 = ( n4451 & n10684 ) | ( n4451 & n13325 ) | ( n10684 & n13325 ) ;
  assign n13327 = n7783 ^ n5380 ^ 1'b0 ;
  assign n13328 = ( n458 & n1794 ) | ( n458 & ~n11832 ) | ( n1794 & ~n11832 ) ;
  assign n13329 = n9614 & ~n12363 ;
  assign n13330 = n1740 & n13329 ;
  assign n13342 = ~n295 & n10670 ;
  assign n13343 = ( ~n9479 & n12764 ) | ( ~n9479 & n13342 ) | ( n12764 & n13342 ) ;
  assign n13337 = n3859 & n5937 ;
  assign n13338 = n13337 ^ n2958 ^ 1'b0 ;
  assign n13335 = n3795 ^ n3532 ^ 1'b0 ;
  assign n13334 = ( x254 & n1141 ) | ( x254 & ~n3482 ) | ( n1141 & ~n3482 ) ;
  assign n13336 = n13335 ^ n13334 ^ 1'b0 ;
  assign n13339 = n13338 ^ n13336 ^ 1'b0 ;
  assign n13340 = n13339 ^ n11734 ^ n9174 ;
  assign n13341 = n13340 ^ n12940 ^ 1'b0 ;
  assign n13331 = n3765 ^ n3004 ^ n795 ;
  assign n13332 = n13331 ^ n1518 ^ x106 ;
  assign n13333 = ( n3983 & n8586 ) | ( n3983 & n13332 ) | ( n8586 & n13332 ) ;
  assign n13344 = n13343 ^ n13341 ^ n13333 ;
  assign n13346 = n4841 ^ n422 ^ 1'b0 ;
  assign n13347 = ~n5151 & n13346 ;
  assign n13348 = n10240 ^ n1387 ^ n431 ;
  assign n13349 = ( n12190 & ~n13347 ) | ( n12190 & n13348 ) | ( ~n13347 & n13348 ) ;
  assign n13345 = n9451 ^ n6054 ^ 1'b0 ;
  assign n13350 = n13349 ^ n13345 ^ n3345 ;
  assign n13351 = ( n3547 & ~n3550 ) | ( n3547 & n12150 ) | ( ~n3550 & n12150 ) ;
  assign n13352 = ( ~n3635 & n8549 ) | ( ~n3635 & n13351 ) | ( n8549 & n13351 ) ;
  assign n13353 = ~n3777 & n8893 ;
  assign n13354 = n13353 ^ n576 ^ 1'b0 ;
  assign n13355 = n3088 ^ n375 ^ 1'b0 ;
  assign n13356 = n13355 ^ n5196 ^ n5130 ;
  assign n13357 = ( ~n6005 & n9344 ) | ( ~n6005 & n10292 ) | ( n9344 & n10292 ) ;
  assign n13358 = ( n13354 & n13356 ) | ( n13354 & ~n13357 ) | ( n13356 & ~n13357 ) ;
  assign n13359 = n13358 ^ n3967 ^ 1'b0 ;
  assign n13360 = n13359 ^ n4239 ^ 1'b0 ;
  assign n13361 = n5505 ^ n3514 ^ n2775 ;
  assign n13362 = n13361 ^ n5834 ^ n4674 ;
  assign n13363 = ~n8687 & n13362 ;
  assign n13364 = n5628 | n13363 ;
  assign n13365 = ( n4878 & ~n5256 ) | ( n4878 & n13364 ) | ( ~n5256 & n13364 ) ;
  assign n13366 = n4630 ^ n708 ^ 1'b0 ;
  assign n13367 = ( n555 & n1957 ) | ( n555 & ~n13366 ) | ( n1957 & ~n13366 ) ;
  assign n13369 = ~n5141 & n5829 ;
  assign n13370 = n10879 ^ n3192 ^ 1'b0 ;
  assign n13371 = n13370 ^ n10082 ^ n2765 ;
  assign n13372 = ~n633 & n13371 ;
  assign n13373 = n13372 ^ n2315 ^ 1'b0 ;
  assign n13374 = n13373 ^ n4475 ^ n2667 ;
  assign n13375 = ( ~n5241 & n13369 ) | ( ~n5241 & n13374 ) | ( n13369 & n13374 ) ;
  assign n13368 = ( n2226 & n8450 ) | ( n2226 & n9406 ) | ( n8450 & n9406 ) ;
  assign n13376 = n13375 ^ n13368 ^ 1'b0 ;
  assign n13377 = n13367 | n13376 ;
  assign n13379 = ~n1060 & n1784 ;
  assign n13380 = n6937 & n13379 ;
  assign n13381 = ( n7095 & ~n9017 ) | ( n7095 & n13380 ) | ( ~n9017 & n13380 ) ;
  assign n13378 = n7922 | n9452 ;
  assign n13382 = n13381 ^ n13378 ^ 1'b0 ;
  assign n13383 = ~n5628 & n13382 ;
  assign n13384 = ( n2555 & n2856 ) | ( n2555 & ~n5147 ) | ( n2856 & ~n5147 ) ;
  assign n13385 = ( x102 & ~n706 ) | ( x102 & n2362 ) | ( ~n706 & n2362 ) ;
  assign n13386 = n13385 ^ n9995 ^ n6592 ;
  assign n13387 = ( ~n13138 & n13384 ) | ( ~n13138 & n13386 ) | ( n13384 & n13386 ) ;
  assign n13388 = n7457 ^ n2803 ^ 1'b0 ;
  assign n13389 = ~n13387 & n13388 ;
  assign n13390 = n7342 | n9123 ;
  assign n13397 = n4976 ^ n2967 ^ 1'b0 ;
  assign n13395 = n1623 & n3549 ;
  assign n13393 = ~x70 & n883 ;
  assign n13391 = n7379 & n12634 ;
  assign n13392 = n13391 ^ n1131 ^ 1'b0 ;
  assign n13394 = n13393 ^ n13392 ^ n8845 ;
  assign n13396 = n13395 ^ n13394 ^ n10915 ;
  assign n13398 = n13397 ^ n13396 ^ n6891 ;
  assign n13399 = n13398 ^ n10783 ^ n10245 ;
  assign n13400 = n13399 ^ n12476 ^ 1'b0 ;
  assign n13401 = ~n13390 & n13400 ;
  assign n13402 = n10459 & n11860 ;
  assign n13411 = n2816 ^ n573 ^ 1'b0 ;
  assign n13412 = x43 & n13411 ;
  assign n13413 = n13412 ^ n4570 ^ n3722 ;
  assign n13414 = ( ~n1906 & n6143 ) | ( ~n1906 & n13413 ) | ( n6143 & n13413 ) ;
  assign n13410 = ( ~n1185 & n3908 ) | ( ~n1185 & n8902 ) | ( n3908 & n8902 ) ;
  assign n13415 = n13414 ^ n13410 ^ 1'b0 ;
  assign n13416 = n4066 & n13415 ;
  assign n13417 = n13416 ^ n13065 ^ n11011 ;
  assign n13418 = n13417 ^ n8324 ^ n5908 ;
  assign n13403 = n883 ^ n367 ^ 1'b0 ;
  assign n13404 = ~n1154 & n12462 ;
  assign n13405 = n13404 ^ n3452 ^ 1'b0 ;
  assign n13406 = n13405 ^ n1486 ^ n1124 ;
  assign n13407 = ( n4613 & ~n13403 ) | ( n4613 & n13406 ) | ( ~n13403 & n13406 ) ;
  assign n13408 = ( n4798 & n5339 ) | ( n4798 & ~n13407 ) | ( n5339 & ~n13407 ) ;
  assign n13409 = n11078 | n13408 ;
  assign n13419 = n13418 ^ n13409 ^ 1'b0 ;
  assign n13420 = n13419 ^ n9714 ^ n3014 ;
  assign n13421 = x191 & ~n1768 ;
  assign n13422 = n13421 ^ n10201 ^ n7563 ;
  assign n13423 = n13422 ^ n5585 ^ n502 ;
  assign n13424 = n666 ^ x121 ^ 1'b0 ;
  assign n13425 = n1578 & ~n13424 ;
  assign n13426 = n4850 ^ n2981 ^ 1'b0 ;
  assign n13427 = ( ~x217 & n13425 ) | ( ~x217 & n13426 ) | ( n13425 & n13426 ) ;
  assign n13428 = n5222 & ~n13427 ;
  assign n13429 = n13428 ^ n4168 ^ 1'b0 ;
  assign n13430 = n5832 & ~n13375 ;
  assign n13431 = ~n13429 & n13430 ;
  assign n13432 = n8750 ^ n764 ^ n704 ;
  assign n13433 = ~n2222 & n4749 ;
  assign n13434 = n13433 ^ n11642 ^ 1'b0 ;
  assign n13435 = n2594 | n8169 ;
  assign n13436 = ( n7228 & n13434 ) | ( n7228 & ~n13435 ) | ( n13434 & ~n13435 ) ;
  assign n13437 = x17 & ~n1272 ;
  assign n13438 = n13436 & n13437 ;
  assign n13439 = n4446 & ~n13438 ;
  assign n13440 = n13439 ^ n7590 ^ 1'b0 ;
  assign n13442 = n1683 ^ n1241 ^ x149 ;
  assign n13441 = ( n1564 & n1884 ) | ( n1564 & n2463 ) | ( n1884 & n2463 ) ;
  assign n13443 = n13442 ^ n13441 ^ n8554 ;
  assign n13444 = n13443 ^ n6960 ^ n1175 ;
  assign n13445 = n10627 & n13255 ;
  assign n13446 = n10490 ^ n8947 ^ 1'b0 ;
  assign n13447 = ~n6158 & n11331 ;
  assign n13448 = n4574 & n13447 ;
  assign n13449 = n13448 ^ n9392 ^ 1'b0 ;
  assign n13450 = ( n2926 & ~n5463 ) | ( n2926 & n12692 ) | ( ~n5463 & n12692 ) ;
  assign n13451 = ~n3923 & n13450 ;
  assign n13452 = n13449 & n13451 ;
  assign n13453 = ~n11475 & n11824 ;
  assign n13454 = n1933 & n13453 ;
  assign n13455 = n2517 ^ n2051 ^ x173 ;
  assign n13456 = n13455 ^ n12059 ^ 1'b0 ;
  assign n13457 = n3614 & n9295 ;
  assign n13458 = n1097 & ~n3974 ;
  assign n13459 = n13458 ^ n10306 ^ n4116 ;
  assign n13460 = ( n959 & n1591 ) | ( n959 & ~n7088 ) | ( n1591 & ~n7088 ) ;
  assign n13461 = ( n1665 & n5703 ) | ( n1665 & n13460 ) | ( n5703 & n13460 ) ;
  assign n13462 = ~n13459 & n13461 ;
  assign n13464 = ( ~n552 & n2334 ) | ( ~n552 & n6535 ) | ( n2334 & n6535 ) ;
  assign n13463 = n266 | n4050 ;
  assign n13465 = n13464 ^ n13463 ^ 1'b0 ;
  assign n13477 = ~n936 & n12419 ;
  assign n13474 = ( n501 & n1537 ) | ( n501 & n5745 ) | ( n1537 & n5745 ) ;
  assign n13475 = n2973 | n13474 ;
  assign n13476 = n10022 | n13475 ;
  assign n13466 = n11468 ^ n5312 ^ 1'b0 ;
  assign n13467 = n7858 | n13466 ;
  assign n13468 = n683 | n13467 ;
  assign n13469 = ( ~n1714 & n5986 ) | ( ~n1714 & n13468 ) | ( n5986 & n13468 ) ;
  assign n13470 = ( ~n1750 & n3773 ) | ( ~n1750 & n13469 ) | ( n3773 & n13469 ) ;
  assign n13471 = ( n604 & n7128 ) | ( n604 & n11591 ) | ( n7128 & n11591 ) ;
  assign n13472 = n13470 & ~n13471 ;
  assign n13473 = n5381 & n13472 ;
  assign n13478 = n13477 ^ n13476 ^ n13473 ;
  assign n13479 = ( n11496 & ~n13465 ) | ( n11496 & n13478 ) | ( ~n13465 & n13478 ) ;
  assign n13480 = n8014 ^ n4848 ^ n3684 ;
  assign n13481 = n13480 ^ n9524 ^ n4417 ;
  assign n13482 = ( n1836 & n2876 ) | ( n1836 & ~n8871 ) | ( n2876 & ~n8871 ) ;
  assign n13483 = n13482 ^ n4720 ^ n3138 ;
  assign n13484 = n13481 | n13483 ;
  assign n13485 = n13484 ^ n9140 ^ n3933 ;
  assign n13487 = n10074 ^ n4613 ^ n585 ;
  assign n13488 = n516 | n7493 ;
  assign n13489 = ( n10279 & n13487 ) | ( n10279 & n13488 ) | ( n13487 & n13488 ) ;
  assign n13490 = n13489 ^ n12966 ^ n4606 ;
  assign n13486 = ( x236 & n2904 ) | ( x236 & ~n4553 ) | ( n2904 & ~n4553 ) ;
  assign n13491 = n13490 ^ n13486 ^ n1909 ;
  assign n13493 = ( n2508 & ~n3976 ) | ( n2508 & n4945 ) | ( ~n3976 & n4945 ) ;
  assign n13494 = n13493 ^ n4903 ^ n4870 ;
  assign n13492 = ~n1188 & n5517 ;
  assign n13495 = n13494 ^ n13492 ^ 1'b0 ;
  assign n13503 = n6644 ^ x246 ^ 1'b0 ;
  assign n13504 = ( n360 & n1796 ) | ( n360 & n13503 ) | ( n1796 & n13503 ) ;
  assign n13505 = ( n1463 & n2581 ) | ( n1463 & ~n10701 ) | ( n2581 & ~n10701 ) ;
  assign n13506 = ( ~n267 & n13504 ) | ( ~n267 & n13505 ) | ( n13504 & n13505 ) ;
  assign n13501 = n11139 ^ n8230 ^ 1'b0 ;
  assign n13496 = n8119 ^ n4729 ^ n1500 ;
  assign n13497 = ( x232 & n1509 ) | ( x232 & n7306 ) | ( n1509 & n7306 ) ;
  assign n13498 = n13497 ^ n6851 ^ 1'b0 ;
  assign n13499 = ~n13496 & n13498 ;
  assign n13500 = n13499 ^ n3415 ^ 1'b0 ;
  assign n13502 = n13501 ^ n13500 ^ 1'b0 ;
  assign n13507 = n13506 ^ n13502 ^ n3849 ;
  assign n13508 = n9132 ^ n5195 ^ n1605 ;
  assign n13509 = n13508 ^ n7022 ^ 1'b0 ;
  assign n13513 = n2984 | n8071 ;
  assign n13510 = n10969 ^ n6955 ^ n538 ;
  assign n13511 = ( n376 & n6716 ) | ( n376 & n13510 ) | ( n6716 & n13510 ) ;
  assign n13512 = n13511 ^ n2250 ^ n581 ;
  assign n13514 = n13513 ^ n13512 ^ n6540 ;
  assign n13515 = n13514 ^ n13361 ^ n3267 ;
  assign n13516 = ( n4225 & ~n6050 ) | ( n4225 & n6182 ) | ( ~n6050 & n6182 ) ;
  assign n13517 = n13516 ^ n13118 ^ x157 ;
  assign n13518 = n12320 ^ n9014 ^ n895 ;
  assign n13519 = n13518 ^ n7832 ^ n4448 ;
  assign n13520 = n9062 ^ n3938 ^ n787 ;
  assign n13521 = n1518 | n7694 ;
  assign n13522 = ( n3663 & ~n8750 ) | ( n3663 & n11689 ) | ( ~n8750 & n11689 ) ;
  assign n13523 = n13522 ^ n2995 ^ 1'b0 ;
  assign n13524 = ( ~n289 & n9193 ) | ( ~n289 & n13523 ) | ( n9193 & n13523 ) ;
  assign n13525 = n13524 ^ n9181 ^ 1'b0 ;
  assign n13526 = ~n13521 & n13525 ;
  assign n13527 = n3931 & ~n12322 ;
  assign n13528 = n7878 & n13527 ;
  assign n13529 = n2394 & ~n4257 ;
  assign n13530 = ~n3459 & n13529 ;
  assign n13531 = n13530 ^ n1972 ^ n541 ;
  assign n13532 = n13531 ^ n13116 ^ n12683 ;
  assign n13533 = n8833 ^ n7155 ^ 1'b0 ;
  assign n13534 = ( ~n3236 & n13532 ) | ( ~n3236 & n13533 ) | ( n13532 & n13533 ) ;
  assign n13535 = n9313 ^ n8815 ^ n7469 ;
  assign n13540 = ( n1583 & ~n5607 ) | ( n1583 & n10488 ) | ( ~n5607 & n10488 ) ;
  assign n13536 = ( n559 & n2310 ) | ( n559 & n5074 ) | ( n2310 & n5074 ) ;
  assign n13537 = ~n7124 & n13536 ;
  assign n13538 = n869 & n13537 ;
  assign n13539 = n4774 & n13538 ;
  assign n13541 = n13540 ^ n13539 ^ n9746 ;
  assign n13542 = ~n3607 & n5639 ;
  assign n13543 = n13542 ^ n3525 ^ 1'b0 ;
  assign n13544 = n13543 ^ n9861 ^ n8111 ;
  assign n13545 = n3951 ^ n3437 ^ n1734 ;
  assign n13546 = n13545 ^ n13279 ^ 1'b0 ;
  assign n13547 = ~n5492 & n7883 ;
  assign n13548 = n13547 ^ n12901 ^ n7607 ;
  assign n13549 = ( n2240 & n13546 ) | ( n2240 & ~n13548 ) | ( n13546 & ~n13548 ) ;
  assign n13550 = ( n2241 & ~n3928 ) | ( n2241 & n6230 ) | ( ~n3928 & n6230 ) ;
  assign n13553 = n7286 | n7633 ;
  assign n13554 = n4772 & ~n13553 ;
  assign n13551 = n12543 ^ n3901 ^ n1659 ;
  assign n13552 = n7822 & n13551 ;
  assign n13555 = n13554 ^ n13552 ^ 1'b0 ;
  assign n13556 = ( n7611 & n13550 ) | ( n7611 & ~n13555 ) | ( n13550 & ~n13555 ) ;
  assign n13557 = ( n4591 & ~n7605 ) | ( n4591 & n13556 ) | ( ~n7605 & n13556 ) ;
  assign n13558 = ( ~n1090 & n3058 ) | ( ~n1090 & n13001 ) | ( n3058 & n13001 ) ;
  assign n13559 = n12935 | n13558 ;
  assign n13560 = n3266 | n13559 ;
  assign n13561 = n10981 ^ n4548 ^ n1207 ;
  assign n13562 = n2894 & ~n11311 ;
  assign n13563 = ( ~n791 & n12576 ) | ( ~n791 & n12617 ) | ( n12576 & n12617 ) ;
  assign n13564 = ( n610 & ~n1940 ) | ( n610 & n7883 ) | ( ~n1940 & n7883 ) ;
  assign n13565 = n13564 ^ n3044 ^ n524 ;
  assign n13566 = n3005 & ~n13565 ;
  assign n13567 = ( n6437 & ~n13563 ) | ( n6437 & n13566 ) | ( ~n13563 & n13566 ) ;
  assign n13568 = ( n6505 & n13562 ) | ( n6505 & n13567 ) | ( n13562 & n13567 ) ;
  assign n13569 = n1620 | n8125 ;
  assign n13570 = n13568 & ~n13569 ;
  assign n13571 = n907 ^ n446 ^ 1'b0 ;
  assign n13582 = n4984 & n9160 ;
  assign n13577 = ~n1769 & n4678 ;
  assign n13578 = n2717 | n5192 ;
  assign n13579 = ~n2145 & n13578 ;
  assign n13580 = n6049 & n13579 ;
  assign n13581 = ( ~n11506 & n13577 ) | ( ~n11506 & n13580 ) | ( n13577 & n13580 ) ;
  assign n13572 = ~n430 & n2882 ;
  assign n13573 = n13270 & n13572 ;
  assign n13574 = n8782 | n13573 ;
  assign n13575 = n13574 ^ x44 ^ 1'b0 ;
  assign n13576 = n13575 ^ n2127 ^ n848 ;
  assign n13583 = n13582 ^ n13581 ^ n13576 ;
  assign n13588 = n3044 & ~n7152 ;
  assign n13589 = n13588 ^ n3647 ^ 1'b0 ;
  assign n13586 = n4305 ^ n3736 ^ n624 ;
  assign n13584 = ( n628 & ~n6507 ) | ( n628 & n13547 ) | ( ~n6507 & n13547 ) ;
  assign n13585 = n13584 ^ n10853 ^ 1'b0 ;
  assign n13587 = n13586 ^ n13585 ^ n7163 ;
  assign n13590 = n13589 ^ n13587 ^ 1'b0 ;
  assign n13591 = ~n13583 & n13590 ;
  assign n13597 = n6434 ^ n3025 ^ n942 ;
  assign n13593 = x109 & ~n7400 ;
  assign n13594 = n13593 ^ n6079 ^ 1'b0 ;
  assign n13595 = n11320 & ~n13338 ;
  assign n13596 = ( n3767 & n13594 ) | ( n3767 & ~n13595 ) | ( n13594 & ~n13595 ) ;
  assign n13592 = n6970 & ~n12029 ;
  assign n13598 = n13597 ^ n13596 ^ n13592 ;
  assign n13599 = ( n2055 & n6804 ) | ( n2055 & n11880 ) | ( n6804 & n11880 ) ;
  assign n13602 = n941 | n12045 ;
  assign n13603 = n5952 & ~n13602 ;
  assign n13600 = ( ~n586 & n3962 ) | ( ~n586 & n4593 ) | ( n3962 & n4593 ) ;
  assign n13601 = n11136 | n13600 ;
  assign n13604 = n13603 ^ n13601 ^ 1'b0 ;
  assign n13605 = ( ~n6648 & n7368 ) | ( ~n6648 & n10631 ) | ( n7368 & n10631 ) ;
  assign n13606 = n12668 & n13605 ;
  assign n13607 = n13606 ^ n1719 ^ 1'b0 ;
  assign n13608 = n5450 ^ n3245 ^ n899 ;
  assign n13609 = n13608 ^ n10215 ^ n8164 ;
  assign n13610 = n13609 ^ n8784 ^ n7531 ;
  assign n13611 = n4666 & n5040 ;
  assign n13612 = ( n1238 & n13610 ) | ( n1238 & ~n13611 ) | ( n13610 & ~n13611 ) ;
  assign n13613 = n13371 ^ n8692 ^ n1865 ;
  assign n13614 = ( x62 & n1725 ) | ( x62 & ~n4118 ) | ( n1725 & ~n4118 ) ;
  assign n13615 = ~n4423 & n13614 ;
  assign n13616 = n3149 ^ n1061 ^ 1'b0 ;
  assign n13617 = n13615 & ~n13616 ;
  assign n13618 = ( ~n1916 & n4794 ) | ( ~n1916 & n7442 ) | ( n4794 & n7442 ) ;
  assign n13619 = ( ~n434 & n2809 ) | ( ~n434 & n13618 ) | ( n2809 & n13618 ) ;
  assign n13620 = ( ~n13613 & n13617 ) | ( ~n13613 & n13619 ) | ( n13617 & n13619 ) ;
  assign n13621 = x30 & n3102 ;
  assign n13622 = ~x134 & n13621 ;
  assign n13623 = n13261 & n13622 ;
  assign n13624 = ~n1362 & n11803 ;
  assign n13625 = n13624 ^ n2417 ^ 1'b0 ;
  assign n13626 = n13625 ^ n10405 ^ n994 ;
  assign n13627 = n11713 ^ n6854 ^ 1'b0 ;
  assign n13628 = ( ~n2430 & n9712 ) | ( ~n2430 & n13627 ) | ( n9712 & n13627 ) ;
  assign n13629 = ( n11633 & n13626 ) | ( n11633 & ~n13628 ) | ( n13626 & ~n13628 ) ;
  assign n13630 = ~n1665 & n2432 ;
  assign n13631 = ~n461 & n13630 ;
  assign n13632 = n2073 & ~n13631 ;
  assign n13633 = n13632 ^ n1928 ^ 1'b0 ;
  assign n13634 = ( n4460 & n4722 ) | ( n4460 & ~n5373 ) | ( n4722 & ~n5373 ) ;
  assign n13635 = n736 | n13634 ;
  assign n13636 = ~n3276 & n7815 ;
  assign n13637 = n13635 | n13636 ;
  assign n13638 = n10219 & ~n13637 ;
  assign n13639 = n4381 ^ n3518 ^ x9 ;
  assign n13640 = ( ~x173 & n7302 ) | ( ~x173 & n13639 ) | ( n7302 & n13639 ) ;
  assign n13641 = n13640 ^ n11748 ^ n2004 ;
  assign n13642 = ( n495 & n8649 ) | ( n495 & n8694 ) | ( n8649 & n8694 ) ;
  assign n13643 = ( n3518 & n13641 ) | ( n3518 & ~n13642 ) | ( n13641 & ~n13642 ) ;
  assign n13645 = n8549 ^ n4271 ^ n1567 ;
  assign n13644 = n3180 & n7578 ;
  assign n13646 = n13645 ^ n13644 ^ 1'b0 ;
  assign n13647 = ( n5478 & n11843 ) | ( n5478 & n13646 ) | ( n11843 & n13646 ) ;
  assign n13648 = ~n11197 & n13647 ;
  assign n13649 = n13648 ^ n8982 ^ 1'b0 ;
  assign n13650 = n4827 | n5348 ;
  assign n13651 = n13650 ^ n1849 ^ 1'b0 ;
  assign n13652 = n10011 & ~n13651 ;
  assign n13653 = ( n7803 & n12928 ) | ( n7803 & n13652 ) | ( n12928 & n13652 ) ;
  assign n13654 = n6074 ^ n5833 ^ 1'b0 ;
  assign n13655 = n2011 & ~n13654 ;
  assign n13656 = n6158 & n13655 ;
  assign n13657 = ~n3572 & n5938 ;
  assign n13658 = n13657 ^ n2801 ^ 1'b0 ;
  assign n13659 = ( n2295 & ~n4680 ) | ( n2295 & n13658 ) | ( ~n4680 & n13658 ) ;
  assign n13660 = n2905 | n5600 ;
  assign n13661 = n13660 ^ n13412 ^ n5804 ;
  assign n13662 = ~n8822 & n13661 ;
  assign n13663 = ( ~n1517 & n7895 ) | ( ~n1517 & n9113 ) | ( n7895 & n9113 ) ;
  assign n13664 = ( n627 & ~n3154 ) | ( n627 & n7467 ) | ( ~n3154 & n7467 ) ;
  assign n13665 = n13664 ^ n8825 ^ n353 ;
  assign n13667 = n3024 ^ n794 ^ 1'b0 ;
  assign n13666 = n9249 ^ n3132 ^ n2459 ;
  assign n13668 = n13667 ^ n13666 ^ n10356 ;
  assign n13669 = n13665 | n13668 ;
  assign n13670 = n582 ^ x134 ^ 1'b0 ;
  assign n13671 = ~n4976 & n13670 ;
  assign n13672 = n13671 ^ n5901 ^ n3086 ;
  assign n13673 = x143 & ~n3591 ;
  assign n13674 = n462 & n13673 ;
  assign n13675 = ( n4874 & n5367 ) | ( n4874 & ~n13674 ) | ( n5367 & ~n13674 ) ;
  assign n13676 = ( n10690 & n13672 ) | ( n10690 & ~n13675 ) | ( n13672 & ~n13675 ) ;
  assign n13677 = n6757 ^ n1789 ^ n280 ;
  assign n13678 = ( n3203 & n5635 ) | ( n3203 & ~n13677 ) | ( n5635 & ~n13677 ) ;
  assign n13679 = n13678 ^ n9716 ^ n4533 ;
  assign n13680 = ( n5671 & ~n13676 ) | ( n5671 & n13679 ) | ( ~n13676 & n13679 ) ;
  assign n13681 = x250 | n641 ;
  assign n13682 = ( n5084 & ~n10048 ) | ( n5084 & n13681 ) | ( ~n10048 & n13681 ) ;
  assign n13683 = n13682 ^ n5516 ^ n2241 ;
  assign n13684 = n13683 ^ n10976 ^ n8777 ;
  assign n13685 = ( n3360 & n8733 ) | ( n3360 & ~n13684 ) | ( n8733 & ~n13684 ) ;
  assign n13686 = ( ~n1329 & n7416 ) | ( ~n1329 & n8285 ) | ( n7416 & n8285 ) ;
  assign n13687 = ( n2020 & n8970 ) | ( n2020 & n13686 ) | ( n8970 & n13686 ) ;
  assign n13688 = ( n348 & n2643 ) | ( n348 & n4630 ) | ( n2643 & n4630 ) ;
  assign n13689 = n809 & n13688 ;
  assign n13692 = ( n1264 & n3151 ) | ( n1264 & ~n3588 ) | ( n3151 & ~n3588 ) ;
  assign n13690 = ~n2008 & n4110 ;
  assign n13691 = n13460 & n13690 ;
  assign n13693 = n13692 ^ n13691 ^ n5671 ;
  assign n13694 = ( n11748 & n13689 ) | ( n11748 & ~n13693 ) | ( n13689 & ~n13693 ) ;
  assign n13695 = n13687 & n13694 ;
  assign n13696 = n13695 ^ n2315 ^ 1'b0 ;
  assign n13697 = n12681 & n13696 ;
  assign n13698 = n12833 & n13697 ;
  assign n13699 = n5945 ^ n5387 ^ 1'b0 ;
  assign n13700 = ( n3209 & n9251 ) | ( n3209 & n11076 ) | ( n9251 & n11076 ) ;
  assign n13701 = ( n2199 & n13699 ) | ( n2199 & ~n13700 ) | ( n13699 & ~n13700 ) ;
  assign n13702 = ( ~n7234 & n8015 ) | ( ~n7234 & n13701 ) | ( n8015 & n13701 ) ;
  assign n13703 = ( n931 & n2262 ) | ( n931 & ~n3998 ) | ( n2262 & ~n3998 ) ;
  assign n13704 = n3993 & n8986 ;
  assign n13705 = ~n13703 & n13704 ;
  assign n13706 = n13705 ^ n9644 ^ n7113 ;
  assign n13707 = n13706 ^ n8948 ^ n1273 ;
  assign n13708 = n13707 ^ n9040 ^ 1'b0 ;
  assign n13712 = n12008 ^ n6465 ^ n1387 ;
  assign n13709 = n6836 | n13000 ;
  assign n13710 = ( n5023 & n5132 ) | ( n5023 & n10072 ) | ( n5132 & n10072 ) ;
  assign n13711 = ( n9729 & n13709 ) | ( n9729 & ~n13710 ) | ( n13709 & ~n13710 ) ;
  assign n13713 = n13712 ^ n13711 ^ n971 ;
  assign n13714 = ( n9684 & n11156 ) | ( n9684 & ~n13713 ) | ( n11156 & ~n13713 ) ;
  assign n13715 = n3500 ^ n2306 ^ 1'b0 ;
  assign n13716 = n9352 & n13715 ;
  assign n13717 = n13716 ^ n1629 ^ 1'b0 ;
  assign n13722 = n11983 ^ n825 ^ 1'b0 ;
  assign n13723 = n5316 | n13722 ;
  assign n13724 = ( ~n8967 & n12403 ) | ( ~n8967 & n13723 ) | ( n12403 & n13723 ) ;
  assign n13725 = n2123 | n13724 ;
  assign n13726 = ~n5157 & n13725 ;
  assign n13718 = n13073 ^ n10335 ^ n7144 ;
  assign n13719 = n5349 ^ n2174 ^ n1990 ;
  assign n13720 = ( ~n1889 & n10380 ) | ( ~n1889 & n13719 ) | ( n10380 & n13719 ) ;
  assign n13721 = n13718 | n13720 ;
  assign n13727 = n13726 ^ n13721 ^ 1'b0 ;
  assign n13728 = n13727 ^ n12340 ^ n5210 ;
  assign n13729 = n5962 | n6188 ;
  assign n13736 = ( n7883 & n9744 ) | ( n7883 & ~n10194 ) | ( n9744 & ~n10194 ) ;
  assign n13737 = n13736 ^ n4777 ^ n2158 ;
  assign n13730 = ( n2244 & ~n2603 ) | ( n2244 & n2740 ) | ( ~n2603 & n2740 ) ;
  assign n13731 = ( n3802 & n4074 ) | ( n3802 & ~n10892 ) | ( n4074 & ~n10892 ) ;
  assign n13732 = ( n3019 & n8273 ) | ( n3019 & ~n13731 ) | ( n8273 & ~n13731 ) ;
  assign n13733 = ( n1830 & n3073 ) | ( n1830 & ~n13732 ) | ( n3073 & ~n13732 ) ;
  assign n13734 = n13733 ^ x83 ^ 1'b0 ;
  assign n13735 = n13730 | n13734 ;
  assign n13738 = n13737 ^ n13735 ^ 1'b0 ;
  assign n13740 = n1530 & n8682 ;
  assign n13741 = n6847 ^ n2273 ^ 1'b0 ;
  assign n13742 = n13740 | n13741 ;
  assign n13739 = ( n2326 & n2620 ) | ( n2326 & n4633 ) | ( n2620 & n4633 ) ;
  assign n13743 = n13742 ^ n13739 ^ n13608 ;
  assign n13746 = ( n1436 & n6992 ) | ( n1436 & n8560 ) | ( n6992 & n8560 ) ;
  assign n13747 = n13746 ^ n5911 ^ 1'b0 ;
  assign n13744 = ~n5034 & n7618 ;
  assign n13745 = ~n1217 & n13744 ;
  assign n13748 = n13747 ^ n13745 ^ 1'b0 ;
  assign n13749 = n2345 ^ n1437 ^ n1309 ;
  assign n13750 = ( n5587 & ~n11715 ) | ( n5587 & n13749 ) | ( ~n11715 & n13749 ) ;
  assign n13751 = n2418 ^ n1246 ^ 1'b0 ;
  assign n13752 = n4771 | n13751 ;
  assign n13753 = n12524 | n13752 ;
  assign n13754 = n7505 ^ n7297 ^ 1'b0 ;
  assign n13755 = n4392 ^ n1416 ^ 1'b0 ;
  assign n13757 = x133 & ~n768 ;
  assign n13756 = n12236 ^ n6924 ^ n1697 ;
  assign n13758 = n13757 ^ n13756 ^ n10676 ;
  assign n13759 = n8406 ^ n7911 ^ 1'b0 ;
  assign n13760 = ( n12593 & n13758 ) | ( n12593 & n13759 ) | ( n13758 & n13759 ) ;
  assign n13761 = n10601 ^ n6110 ^ n1578 ;
  assign n13762 = n13761 ^ n3489 ^ n1312 ;
  assign n13763 = n7424 & n13762 ;
  assign n13764 = n4436 ^ n2904 ^ 1'b0 ;
  assign n13765 = n5421 & ~n13764 ;
  assign n13766 = n10348 ^ n9829 ^ 1'b0 ;
  assign n13767 = n13765 & n13766 ;
  assign n13768 = ~n13763 & n13767 ;
  assign n13769 = n13768 ^ n5775 ^ 1'b0 ;
  assign n13770 = ~n9335 & n13769 ;
  assign n13771 = ( n2163 & n2545 ) | ( n2163 & ~n8158 ) | ( n2545 & ~n8158 ) ;
  assign n13772 = n12470 ^ n10609 ^ 1'b0 ;
  assign n13773 = ( n2228 & n3195 ) | ( n2228 & n5973 ) | ( n3195 & n5973 ) ;
  assign n13774 = n13773 ^ n5384 ^ 1'b0 ;
  assign n13775 = n634 & ~n13774 ;
  assign n13776 = n2694 & ~n13609 ;
  assign n13777 = ( n2857 & ~n3525 ) | ( n2857 & n8360 ) | ( ~n3525 & n8360 ) ;
  assign n13778 = ( ~n7665 & n13776 ) | ( ~n7665 & n13777 ) | ( n13776 & n13777 ) ;
  assign n13789 = ( n7347 & ~n7603 ) | ( n7347 & n13073 ) | ( ~n7603 & n13073 ) ;
  assign n13784 = n13578 ^ n2378 ^ n1209 ;
  assign n13785 = n13784 ^ n5069 ^ 1'b0 ;
  assign n13786 = n11768 & n13785 ;
  assign n13787 = ( ~n1224 & n12596 ) | ( ~n1224 & n13786 ) | ( n12596 & n13786 ) ;
  assign n13779 = ( ~x106 & x161 ) | ( ~x106 & n800 ) | ( x161 & n800 ) ;
  assign n13780 = n1481 & ~n13779 ;
  assign n13781 = n8682 | n13780 ;
  assign n13782 = n13781 ^ n615 ^ 1'b0 ;
  assign n13783 = ~n6579 & n13782 ;
  assign n13788 = n13787 ^ n13783 ^ 1'b0 ;
  assign n13790 = n13789 ^ n13788 ^ 1'b0 ;
  assign n13791 = n4101 ^ n1636 ^ 1'b0 ;
  assign n13792 = n8046 & n13791 ;
  assign n13793 = ( x22 & ~n487 ) | ( x22 & n3067 ) | ( ~n487 & n3067 ) ;
  assign n13794 = n13793 ^ n6104 ^ n2455 ;
  assign n13795 = n13794 ^ n3927 ^ n547 ;
  assign n13796 = ( n3575 & ~n13792 ) | ( n3575 & n13795 ) | ( ~n13792 & n13795 ) ;
  assign n13797 = n13796 ^ n2750 ^ 1'b0 ;
  assign n13798 = n6017 ^ n5611 ^ n2715 ;
  assign n13799 = ~n1957 & n10459 ;
  assign n13800 = ( n8917 & ~n13798 ) | ( n8917 & n13799 ) | ( ~n13798 & n13799 ) ;
  assign n13801 = ( n1813 & n11974 ) | ( n1813 & n13800 ) | ( n11974 & n13800 ) ;
  assign n13802 = n13801 ^ n10322 ^ 1'b0 ;
  assign n13803 = x67 & ~n4866 ;
  assign n13804 = n9283 & n13803 ;
  assign n13805 = n13804 ^ n12211 ^ 1'b0 ;
  assign n13806 = n13805 ^ n6667 ^ 1'b0 ;
  assign n13807 = n11053 & ~n13806 ;
  assign n13808 = n10391 ^ n5957 ^ n5451 ;
  assign n13809 = n13808 ^ n11228 ^ n3485 ;
  assign n13810 = n2027 | n4523 ;
  assign n13811 = n2357 | n13810 ;
  assign n13812 = ~n2559 & n9007 ;
  assign n13813 = ~n4230 & n13812 ;
  assign n13814 = ( n3597 & ~n4564 ) | ( n3597 & n13813 ) | ( ~n4564 & n13813 ) ;
  assign n13815 = n13811 | n13814 ;
  assign n13816 = ( n2884 & n11186 ) | ( n2884 & ~n13815 ) | ( n11186 & ~n13815 ) ;
  assign n13818 = ( n3663 & n7077 ) | ( n3663 & ~n13131 ) | ( n7077 & ~n13131 ) ;
  assign n13817 = ( n5037 & n7822 ) | ( n5037 & n13341 ) | ( n7822 & n13341 ) ;
  assign n13819 = n13818 ^ n13817 ^ 1'b0 ;
  assign n13820 = n5828 ^ n3288 ^ n829 ;
  assign n13821 = n1860 & n4263 ;
  assign n13822 = n3287 & ~n4118 ;
  assign n13823 = n13822 ^ n4826 ^ 1'b0 ;
  assign n13824 = n13823 ^ n4937 ^ n1416 ;
  assign n13825 = n13824 ^ n713 ^ 1'b0 ;
  assign n13826 = ~n2305 & n13825 ;
  assign n13827 = n13826 ^ n5187 ^ n1451 ;
  assign n13828 = ( x92 & ~n13821 ) | ( x92 & n13827 ) | ( ~n13821 & n13827 ) ;
  assign n13829 = n13828 ^ n11501 ^ 1'b0 ;
  assign n13830 = ~n2009 & n13829 ;
  assign n13831 = n7793 ^ n4366 ^ 1'b0 ;
  assign n13832 = ( n4567 & n8194 ) | ( n4567 & ~n13831 ) | ( n8194 & ~n13831 ) ;
  assign n13833 = n13832 ^ n5991 ^ 1'b0 ;
  assign n13834 = ~n9402 & n13833 ;
  assign n13835 = ( n1376 & n7479 ) | ( n1376 & ~n13834 ) | ( n7479 & ~n13834 ) ;
  assign n13836 = ( n989 & n992 ) | ( n989 & ~n7388 ) | ( n992 & ~n7388 ) ;
  assign n13837 = n10488 ^ n5287 ^ 1'b0 ;
  assign n13838 = n7041 & ~n13837 ;
  assign n13839 = n13838 ^ n11816 ^ n708 ;
  assign n13840 = ( n1475 & n3012 ) | ( n1475 & n7263 ) | ( n3012 & n7263 ) ;
  assign n13841 = ( n13836 & n13839 ) | ( n13836 & n13840 ) | ( n13839 & n13840 ) ;
  assign n13843 = x117 & ~n3744 ;
  assign n13844 = n13843 ^ n2390 ^ 1'b0 ;
  assign n13842 = x80 & n11051 ;
  assign n13845 = n13844 ^ n13842 ^ 1'b0 ;
  assign n13846 = n348 | n13845 ;
  assign n13847 = ( x211 & n6261 ) | ( x211 & n7783 ) | ( n6261 & n7783 ) ;
  assign n13848 = n4653 | n13847 ;
  assign n13851 = n7965 ^ n566 ^ 1'b0 ;
  assign n13852 = ~n2828 & n13851 ;
  assign n13849 = ( ~n2521 & n9769 ) | ( ~n2521 & n10380 ) | ( n9769 & n10380 ) ;
  assign n13850 = n13849 ^ n12158 ^ n905 ;
  assign n13853 = n13852 ^ n13850 ^ n5010 ;
  assign n13855 = n9717 | n11348 ;
  assign n13856 = n4165 | n13855 ;
  assign n13854 = n3873 ^ n3811 ^ 1'b0 ;
  assign n13857 = n13856 ^ n13854 ^ n3041 ;
  assign n13864 = n8679 ^ n3487 ^ n2411 ;
  assign n13861 = n383 & n1195 ;
  assign n13862 = n3841 & n13861 ;
  assign n13863 = ( n668 & ~n10471 ) | ( n668 & n13862 ) | ( ~n10471 & n13862 ) ;
  assign n13865 = n13864 ^ n13863 ^ n1764 ;
  assign n13858 = n4691 ^ n1329 ^ 1'b0 ;
  assign n13859 = n2043 ^ n831 ^ n778 ;
  assign n13860 = ~n13858 & n13859 ;
  assign n13866 = n13865 ^ n13860 ^ 1'b0 ;
  assign n13867 = n4135 | n7824 ;
  assign n13868 = n13867 ^ n3690 ^ 1'b0 ;
  assign n13869 = n4758 ^ n2985 ^ x138 ;
  assign n13870 = n9422 ^ n7490 ^ x19 ;
  assign n13871 = n13870 ^ n12371 ^ 1'b0 ;
  assign n13872 = ~n13869 & n13871 ;
  assign n13878 = ( n7327 & n13139 ) | ( n7327 & n13405 ) | ( n13139 & n13405 ) ;
  assign n13879 = n13878 ^ n2321 ^ 1'b0 ;
  assign n13873 = n8521 ^ n6161 ^ 1'b0 ;
  assign n13874 = n5841 & ~n13873 ;
  assign n13875 = n8718 ^ n5947 ^ n2445 ;
  assign n13876 = ( n3524 & n13504 ) | ( n3524 & ~n13875 ) | ( n13504 & ~n13875 ) ;
  assign n13877 = n13874 & n13876 ;
  assign n13880 = n13879 ^ n13877 ^ 1'b0 ;
  assign n13881 = ( n4320 & n10923 ) | ( n4320 & ~n13880 ) | ( n10923 & ~n13880 ) ;
  assign n13882 = ~n1893 & n3536 ;
  assign n13883 = n13882 ^ n3723 ^ 1'b0 ;
  assign n13884 = n6469 ^ n4249 ^ x74 ;
  assign n13885 = n13883 & ~n13884 ;
  assign n13886 = n13885 ^ n280 ^ 1'b0 ;
  assign n13887 = ( n7217 & n7856 ) | ( n7217 & ~n8075 ) | ( n7856 & ~n8075 ) ;
  assign n13889 = ( n861 & n1102 ) | ( n861 & n1730 ) | ( n1102 & n1730 ) ;
  assign n13888 = ( ~x102 & x103 ) | ( ~x102 & n1258 ) | ( x103 & n1258 ) ;
  assign n13890 = n13889 ^ n13888 ^ n7068 ;
  assign n13891 = n13890 ^ n6622 ^ n5531 ;
  assign n13894 = n7681 ^ n3686 ^ n973 ;
  assign n13895 = n13894 ^ n12975 ^ n6509 ;
  assign n13892 = n6582 ^ n5844 ^ 1'b0 ;
  assign n13893 = ~n4401 & n13892 ;
  assign n13896 = n13895 ^ n13893 ^ 1'b0 ;
  assign n13897 = n13896 ^ n11316 ^ 1'b0 ;
  assign n13898 = n10649 & n11893 ;
  assign n13899 = n13223 ^ n9639 ^ n4017 ;
  assign n13900 = n13899 ^ n8145 ^ 1'b0 ;
  assign n13901 = n13419 ^ n7981 ^ n5021 ;
  assign n13902 = n11956 ^ n835 ^ 1'b0 ;
  assign n13903 = ~n13471 & n13902 ;
  assign n13904 = n4192 ^ n2528 ^ x16 ;
  assign n13905 = ( n1883 & n4427 ) | ( n1883 & ~n13904 ) | ( n4427 & ~n13904 ) ;
  assign n13906 = ( n5236 & n5466 ) | ( n5236 & n9171 ) | ( n5466 & n9171 ) ;
  assign n13907 = n13906 ^ n10133 ^ 1'b0 ;
  assign n13908 = ( n752 & n2372 ) | ( n752 & n4623 ) | ( n2372 & n4623 ) ;
  assign n13909 = n13908 ^ n2310 ^ 1'b0 ;
  assign n13910 = n7339 ^ n5766 ^ n4512 ;
  assign n13911 = n7949 & ~n13910 ;
  assign n13912 = n6701 & n13911 ;
  assign n13913 = n8096 ^ x133 ^ 1'b0 ;
  assign n13914 = n5023 & n13913 ;
  assign n13915 = ( ~n13909 & n13912 ) | ( ~n13909 & n13914 ) | ( n13912 & n13914 ) ;
  assign n13921 = n2862 ^ n2263 ^ n748 ;
  assign n13922 = n795 & n1645 ;
  assign n13923 = x129 & n13922 ;
  assign n13924 = n846 & ~n13923 ;
  assign n13925 = n13921 & ~n13924 ;
  assign n13926 = ( n4657 & n6739 ) | ( n4657 & n13925 ) | ( n6739 & n13925 ) ;
  assign n13916 = n7588 ^ n4792 ^ 1'b0 ;
  assign n13917 = n9485 ^ n9186 ^ n1902 ;
  assign n13918 = ( n6806 & n13916 ) | ( n6806 & ~n13917 ) | ( n13916 & ~n13917 ) ;
  assign n13919 = n2090 & ~n13918 ;
  assign n13920 = ~n11944 & n13919 ;
  assign n13927 = n13926 ^ n13920 ^ 1'b0 ;
  assign n13929 = x178 & ~n785 ;
  assign n13930 = ( x47 & n9273 ) | ( x47 & n9903 ) | ( n9273 & n9903 ) ;
  assign n13932 = ( n793 & ~n2635 ) | ( n793 & n6979 ) | ( ~n2635 & n6979 ) ;
  assign n13933 = n13932 ^ n6789 ^ n3250 ;
  assign n13931 = n2997 & n8172 ;
  assign n13934 = n13933 ^ n13931 ^ n7580 ;
  assign n13935 = n13934 ^ n9040 ^ n2480 ;
  assign n13936 = ( n13929 & ~n13930 ) | ( n13929 & n13935 ) | ( ~n13930 & n13935 ) ;
  assign n13928 = ~n2018 & n5504 ;
  assign n13937 = n13936 ^ n13928 ^ n1380 ;
  assign n13941 = n9952 ^ n304 ^ 1'b0 ;
  assign n13938 = n2869 & n5532 ;
  assign n13939 = n7835 & ~n13938 ;
  assign n13940 = ~n7740 & n13939 ;
  assign n13942 = n13941 ^ n13940 ^ x109 ;
  assign n13943 = n11803 & ~n13942 ;
  assign n13944 = n6451 & ~n7301 ;
  assign n13945 = n5461 ^ n1753 ^ x201 ;
  assign n13946 = n13944 | n13945 ;
  assign n13947 = ~n693 & n1017 ;
  assign n13948 = n1463 | n3340 ;
  assign n13949 = ( n3518 & n13844 ) | ( n3518 & ~n13948 ) | ( n13844 & ~n13948 ) ;
  assign n13950 = ( n811 & n1592 ) | ( n811 & ~n13949 ) | ( n1592 & ~n13949 ) ;
  assign n13951 = n13950 ^ n5870 ^ n4908 ;
  assign n13952 = n13951 ^ n9712 ^ 1'b0 ;
  assign n13956 = x19 & n10702 ;
  assign n13957 = n7328 & n13956 ;
  assign n13953 = n2144 & ~n2252 ;
  assign n13954 = n13953 ^ n568 ^ 1'b0 ;
  assign n13955 = n10676 | n13954 ;
  assign n13958 = n13957 ^ n13955 ^ n7928 ;
  assign n13959 = n13958 ^ n9687 ^ n8974 ;
  assign n13960 = n1793 ^ n1539 ^ n1164 ;
  assign n13961 = n7635 ^ n2305 ^ 1'b0 ;
  assign n13962 = n5904 ^ n4608 ^ x200 ;
  assign n13963 = n13962 ^ n7229 ^ 1'b0 ;
  assign n13964 = n13961 & ~n13963 ;
  assign n13965 = ( n7521 & n13960 ) | ( n7521 & n13964 ) | ( n13960 & n13964 ) ;
  assign n13966 = n10345 ^ n2522 ^ 1'b0 ;
  assign n13967 = ~n4890 & n13966 ;
  assign n13968 = n7075 & n9535 ;
  assign n13969 = n13968 ^ n2695 ^ 1'b0 ;
  assign n13970 = n13969 ^ n13079 ^ 1'b0 ;
  assign n13971 = ( ~n5638 & n13967 ) | ( ~n5638 & n13970 ) | ( n13967 & n13970 ) ;
  assign n13972 = ( ~n1419 & n2319 ) | ( ~n1419 & n13971 ) | ( n2319 & n13971 ) ;
  assign n13973 = ( ~n4005 & n12077 ) | ( ~n4005 & n12812 ) | ( n12077 & n12812 ) ;
  assign n13980 = x20 & x106 ;
  assign n13981 = ~n1629 & n13980 ;
  assign n13982 = n13981 ^ n9315 ^ n4570 ;
  assign n13974 = n13573 ^ n385 ^ 1'b0 ;
  assign n13975 = ~n2069 & n2232 ;
  assign n13976 = n13975 ^ n6621 ^ 1'b0 ;
  assign n13977 = ( n639 & n9078 ) | ( n639 & ~n13976 ) | ( n9078 & ~n13976 ) ;
  assign n13978 = ( n12726 & ~n13974 ) | ( n12726 & n13977 ) | ( ~n13974 & n13977 ) ;
  assign n13979 = n10762 & ~n13978 ;
  assign n13983 = n13982 ^ n13979 ^ 1'b0 ;
  assign n13984 = n12168 ^ n6024 ^ 1'b0 ;
  assign n13985 = n9733 & ~n13984 ;
  assign n13986 = n13985 ^ n3747 ^ 1'b0 ;
  assign n13987 = n10476 ^ n3865 ^ 1'b0 ;
  assign n13988 = n8458 | n13987 ;
  assign n13989 = n11773 ^ n427 ^ x19 ;
  assign n13990 = ( ~n10464 & n13988 ) | ( ~n10464 & n13989 ) | ( n13988 & n13989 ) ;
  assign n13991 = n8991 ^ n5008 ^ n2417 ;
  assign n13992 = ( n1553 & n4836 ) | ( n1553 & n13991 ) | ( n4836 & n13991 ) ;
  assign n13993 = n13992 ^ n12842 ^ n2619 ;
  assign n13994 = n6280 ^ n1805 ^ n1211 ;
  assign n13995 = n7667 & ~n13994 ;
  assign n13996 = n13995 ^ n1080 ^ 1'b0 ;
  assign n13997 = n13996 ^ n360 ^ x49 ;
  assign n13998 = n3862 & ~n4600 ;
  assign n13999 = ~n1913 & n13998 ;
  assign n14000 = ( n1397 & n7021 ) | ( n1397 & ~n13999 ) | ( n7021 & ~n13999 ) ;
  assign n14001 = n10663 ^ n10342 ^ n3688 ;
  assign n14002 = ( n4456 & n8041 ) | ( n4456 & ~n14001 ) | ( n8041 & ~n14001 ) ;
  assign n14003 = ( n6430 & n12462 ) | ( n6430 & n14002 ) | ( n12462 & n14002 ) ;
  assign n14004 = n6652 ^ n6344 ^ 1'b0 ;
  assign n14009 = x192 & ~n1214 ;
  assign n14010 = n14009 ^ n5302 ^ 1'b0 ;
  assign n14011 = n14010 ^ n11397 ^ n2427 ;
  assign n14005 = n919 | n3280 ;
  assign n14006 = n14005 ^ n676 ^ 1'b0 ;
  assign n14007 = ( ~n6064 & n13410 ) | ( ~n6064 & n14006 ) | ( n13410 & n14006 ) ;
  assign n14008 = n1577 & n14007 ;
  assign n14012 = n14011 ^ n14008 ^ n9607 ;
  assign n14013 = ( n9802 & ~n11711 ) | ( n9802 & n14012 ) | ( ~n11711 & n14012 ) ;
  assign n14017 = n4789 ^ n4051 ^ n3227 ;
  assign n14014 = n8680 ^ n7733 ^ n5450 ;
  assign n14015 = n2502 | n14014 ;
  assign n14016 = n2933 & ~n14015 ;
  assign n14018 = n14017 ^ n14016 ^ 1'b0 ;
  assign n14019 = n2404 & n4973 ;
  assign n14020 = n1635 & n14019 ;
  assign n14021 = ( ~n1527 & n8197 ) | ( ~n1527 & n14020 ) | ( n8197 & n14020 ) ;
  assign n14022 = n14021 ^ n9476 ^ 1'b0 ;
  assign n14023 = n7107 & n10893 ;
  assign n14024 = n14023 ^ n4260 ^ n511 ;
  assign n14025 = n7272 ^ n3999 ^ 1'b0 ;
  assign n14026 = n14024 | n14025 ;
  assign n14027 = n8487 & ~n14026 ;
  assign n14028 = n3813 & n14027 ;
  assign n14039 = n3536 & n7905 ;
  assign n14040 = n14039 ^ n814 ^ 1'b0 ;
  assign n14036 = n4208 ^ n3515 ^ 1'b0 ;
  assign n14037 = x156 & ~n14036 ;
  assign n14038 = n14037 ^ n4211 ^ 1'b0 ;
  assign n14033 = ( n2278 & n3668 ) | ( n2278 & n4423 ) | ( n3668 & n4423 ) ;
  assign n14029 = ( n779 & ~n3965 ) | ( n779 & n9064 ) | ( ~n3965 & n9064 ) ;
  assign n14030 = n14029 ^ n9122 ^ n4547 ;
  assign n14031 = ( n873 & ~n9344 ) | ( n873 & n14030 ) | ( ~n9344 & n14030 ) ;
  assign n14032 = n6772 | n14031 ;
  assign n14034 = n14033 ^ n14032 ^ 1'b0 ;
  assign n14035 = n14034 ^ n8108 ^ n1020 ;
  assign n14041 = n14040 ^ n14038 ^ n14035 ;
  assign n14042 = n12906 ^ n4147 ^ n2064 ;
  assign n14043 = n14042 ^ n10469 ^ 1'b0 ;
  assign n14044 = n607 & ~n1599 ;
  assign n14048 = ( n6305 & n6687 ) | ( n6305 & n8926 ) | ( n6687 & n8926 ) ;
  assign n14045 = n7277 ^ n2777 ^ 1'b0 ;
  assign n14046 = ( n3151 & ~n3384 ) | ( n3151 & n5171 ) | ( ~n3384 & n5171 ) ;
  assign n14047 = ( n4466 & ~n14045 ) | ( n4466 & n14046 ) | ( ~n14045 & n14046 ) ;
  assign n14049 = n14048 ^ n14047 ^ n10734 ;
  assign n14050 = ( n11906 & n14044 ) | ( n11906 & ~n14049 ) | ( n14044 & ~n14049 ) ;
  assign n14051 = ( n1709 & n4651 ) | ( n1709 & ~n14050 ) | ( n4651 & ~n14050 ) ;
  assign n14052 = n14051 ^ n3353 ^ 1'b0 ;
  assign n14054 = n7580 ^ n2659 ^ n863 ;
  assign n14053 = ( n3416 & n9601 ) | ( n3416 & ~n9921 ) | ( n9601 & ~n9921 ) ;
  assign n14055 = n14054 ^ n14053 ^ n3274 ;
  assign n14056 = n13556 ^ n5440 ^ n4651 ;
  assign n14057 = n8412 ^ n6126 ^ n1480 ;
  assign n14064 = n9371 ^ n1526 ^ 1'b0 ;
  assign n14058 = n7044 ^ n963 ^ n757 ;
  assign n14059 = n11989 & n14058 ;
  assign n14060 = n14059 ^ n1111 ^ 1'b0 ;
  assign n14061 = n7570 | n11931 ;
  assign n14062 = n14060 | n14061 ;
  assign n14063 = ~n7732 & n14062 ;
  assign n14065 = n14064 ^ n14063 ^ n11971 ;
  assign n14066 = ~n13908 & n14065 ;
  assign n14067 = ~n5447 & n14066 ;
  assign n14068 = ( n3624 & ~n14057 ) | ( n3624 & n14067 ) | ( ~n14057 & n14067 ) ;
  assign n14069 = ( n5095 & n5906 ) | ( n5095 & n6669 ) | ( n5906 & n6669 ) ;
  assign n14070 = n1774 & n5344 ;
  assign n14071 = n1349 & n14070 ;
  assign n14072 = n1101 & n12768 ;
  assign n14073 = n14072 ^ n8414 ^ 1'b0 ;
  assign n14074 = ( n8767 & ~n14071 ) | ( n8767 & n14073 ) | ( ~n14071 & n14073 ) ;
  assign n14075 = n14074 ^ n9383 ^ 1'b0 ;
  assign n14076 = n14069 & ~n14075 ;
  assign n14077 = n2773 & n11279 ;
  assign n14078 = n12248 ^ n5086 ^ x111 ;
  assign n14079 = ( n612 & ~n2011 ) | ( n612 & n14078 ) | ( ~n2011 & n14078 ) ;
  assign n14080 = n7222 & n11198 ;
  assign n14081 = n5391 ^ x0 ^ 1'b0 ;
  assign n14082 = n14080 & n14081 ;
  assign n14083 = n14079 & n14082 ;
  assign n14084 = ( n1027 & n6397 ) | ( n1027 & ~n6442 ) | ( n6397 & ~n6442 ) ;
  assign n14085 = n14084 ^ n12802 ^ n6529 ;
  assign n14086 = n4078 & n12483 ;
  assign n14087 = n2224 & n14086 ;
  assign n14088 = n13875 & ~n14087 ;
  assign n14089 = n14088 ^ n3071 ^ 1'b0 ;
  assign n14090 = ( x93 & n2476 ) | ( x93 & ~n13441 ) | ( n2476 & ~n13441 ) ;
  assign n14091 = ( ~n14085 & n14089 ) | ( ~n14085 & n14090 ) | ( n14089 & n14090 ) ;
  assign n14093 = n621 | n1935 ;
  assign n14094 = n3668 | n14093 ;
  assign n14095 = ( n4060 & n6363 ) | ( n4060 & n14094 ) | ( n6363 & n14094 ) ;
  assign n14096 = n14095 ^ n7766 ^ n6435 ;
  assign n14092 = ~n3949 & n5975 ;
  assign n14097 = n14096 ^ n14092 ^ 1'b0 ;
  assign n14098 = n8431 ^ n3710 ^ n2622 ;
  assign n14099 = n14098 ^ n11657 ^ n7696 ;
  assign n14100 = ( n9749 & n14097 ) | ( n9749 & ~n14099 ) | ( n14097 & ~n14099 ) ;
  assign n14101 = n5886 ^ n317 ^ 1'b0 ;
  assign n14102 = ~n8503 & n11153 ;
  assign n14103 = n14102 ^ x217 ^ 1'b0 ;
  assign n14106 = ( n3225 & n8136 ) | ( n3225 & n13503 ) | ( n8136 & n13503 ) ;
  assign n14104 = n2868 & n6222 ;
  assign n14105 = n3711 & n14104 ;
  assign n14107 = n14106 ^ n14105 ^ n10068 ;
  assign n14111 = ~n3844 & n6136 ;
  assign n14112 = n14111 ^ x35 ^ 1'b0 ;
  assign n14109 = n11558 ^ n4040 ^ n981 ;
  assign n14110 = n2442 | n14109 ;
  assign n14108 = n280 & n5115 ;
  assign n14113 = n14112 ^ n14110 ^ n14108 ;
  assign n14114 = n7758 ^ n2640 ^ n2573 ;
  assign n14115 = n14114 ^ n7732 ^ 1'b0 ;
  assign n14116 = n1139 & n14115 ;
  assign n14117 = n14116 ^ n7842 ^ 1'b0 ;
  assign n14118 = n10628 | n14117 ;
  assign n14119 = n4789 ^ n3152 ^ 1'b0 ;
  assign n14120 = n2070 & n14119 ;
  assign n14121 = n6431 | n7300 ;
  assign n14122 = n14121 ^ n4134 ^ 1'b0 ;
  assign n14123 = ( n8187 & ~n14120 ) | ( n8187 & n14122 ) | ( ~n14120 & n14122 ) ;
  assign n14124 = ~n14118 & n14123 ;
  assign n14125 = n14124 ^ n12567 ^ 1'b0 ;
  assign n14126 = ( ~n1003 & n5965 ) | ( ~n1003 & n7574 ) | ( n5965 & n7574 ) ;
  assign n14127 = ( n7189 & ~n12901 ) | ( n7189 & n14126 ) | ( ~n12901 & n14126 ) ;
  assign n14128 = n8338 | n14127 ;
  assign n14138 = n787 & n6914 ;
  assign n14139 = n14138 ^ n2931 ^ 1'b0 ;
  assign n14140 = ~x66 & n14139 ;
  assign n14141 = n12409 | n14140 ;
  assign n14142 = n1580 & ~n2728 ;
  assign n14143 = ~n692 & n14142 ;
  assign n14144 = ( n2673 & ~n4721 ) | ( n2673 & n14143 ) | ( ~n4721 & n14143 ) ;
  assign n14145 = n14144 ^ n14071 ^ n12310 ;
  assign n14146 = ( n8882 & n14141 ) | ( n8882 & n14145 ) | ( n14141 & n14145 ) ;
  assign n14136 = ( ~n4362 & n4880 ) | ( ~n4362 & n10834 ) | ( n4880 & n10834 ) ;
  assign n14137 = n14136 ^ n7038 ^ n6716 ;
  assign n14129 = n7292 ^ n5621 ^ n3005 ;
  assign n14130 = n1076 | n7907 ;
  assign n14131 = n14130 ^ n4950 ^ 1'b0 ;
  assign n14132 = n8743 ^ n7972 ^ n7002 ;
  assign n14133 = n14131 & n14132 ;
  assign n14134 = ( n13921 & ~n14129 ) | ( n13921 & n14133 ) | ( ~n14129 & n14133 ) ;
  assign n14135 = n14134 ^ n5619 ^ 1'b0 ;
  assign n14147 = n14146 ^ n14137 ^ n14135 ;
  assign n14148 = n7957 ^ n5220 ^ 1'b0 ;
  assign n14150 = ( n2309 & n5211 ) | ( n2309 & n5294 ) | ( n5211 & n5294 ) ;
  assign n14151 = ~n1112 & n10641 ;
  assign n14152 = ( n1212 & ~n14150 ) | ( n1212 & n14151 ) | ( ~n14150 & n14151 ) ;
  assign n14149 = ( n2413 & n3002 ) | ( n2413 & n5743 ) | ( n3002 & n5743 ) ;
  assign n14153 = n14152 ^ n14149 ^ n7690 ;
  assign n14154 = n4555 ^ n1134 ^ 1'b0 ;
  assign n14155 = n6988 & n14154 ;
  assign n14156 = n834 & n8201 ;
  assign n14157 = n3438 & n14156 ;
  assign n14158 = ( n8492 & ~n8612 ) | ( n8492 & n14157 ) | ( ~n8612 & n14157 ) ;
  assign n14159 = ( n1502 & ~n2657 ) | ( n1502 & n14158 ) | ( ~n2657 & n14158 ) ;
  assign n14160 = n5141 ^ n3504 ^ 1'b0 ;
  assign n14161 = n14160 ^ n12206 ^ n8892 ;
  assign n14162 = ( n14155 & ~n14159 ) | ( n14155 & n14161 ) | ( ~n14159 & n14161 ) ;
  assign n14163 = n14153 & ~n14162 ;
  assign n14182 = ( n5529 & ~n7599 ) | ( n5529 & n7863 ) | ( ~n7599 & n7863 ) ;
  assign n14174 = ( ~n5420 & n6926 ) | ( ~n5420 & n7051 ) | ( n6926 & n7051 ) ;
  assign n14175 = n10694 | n14174 ;
  assign n14176 = n14175 ^ n10101 ^ 1'b0 ;
  assign n14177 = n414 & n14176 ;
  assign n14178 = n14177 ^ n7136 ^ 1'b0 ;
  assign n14179 = n6859 & ~n14178 ;
  assign n14180 = n14179 ^ n11931 ^ n3623 ;
  assign n14181 = n14180 ^ n8263 ^ n3871 ;
  assign n14172 = ( ~n1529 & n1728 ) | ( ~n1529 & n3845 ) | ( n1728 & n3845 ) ;
  assign n14164 = n4987 | n5348 ;
  assign n14165 = n8912 | n14164 ;
  assign n14166 = n7542 ^ n2544 ^ n556 ;
  assign n14167 = n14166 ^ n8961 ^ n6329 ;
  assign n14168 = n4236 ^ n1701 ^ 1'b0 ;
  assign n14169 = n14167 | n14168 ;
  assign n14170 = ( n11487 & n11664 ) | ( n11487 & n14169 ) | ( n11664 & n14169 ) ;
  assign n14171 = n14165 & ~n14170 ;
  assign n14173 = n14172 ^ n14171 ^ 1'b0 ;
  assign n14183 = n14182 ^ n14181 ^ n14173 ;
  assign n14184 = n12360 ^ n3639 ^ n708 ;
  assign n14185 = n3120 & n5776 ;
  assign n14186 = n14185 ^ n5448 ^ 1'b0 ;
  assign n14187 = ( n2675 & n7306 ) | ( n2675 & n14186 ) | ( n7306 & n14186 ) ;
  assign n14188 = n9120 | n14187 ;
  assign n14189 = n11800 | n14188 ;
  assign n14190 = ( n5642 & n14184 ) | ( n5642 & ~n14189 ) | ( n14184 & ~n14189 ) ;
  assign n14191 = x151 & ~n9822 ;
  assign n14192 = n14191 ^ n5506 ^ 1'b0 ;
  assign n14193 = ( ~x10 & n13949 ) | ( ~x10 & n14192 ) | ( n13949 & n14192 ) ;
  assign n14197 = n7850 ^ n1331 ^ n1003 ;
  assign n14196 = n8488 ^ n5249 ^ n1880 ;
  assign n14194 = ( n3041 & ~n5309 ) | ( n3041 & n5824 ) | ( ~n5309 & n5824 ) ;
  assign n14195 = n14194 ^ n8174 ^ n482 ;
  assign n14198 = n14197 ^ n14196 ^ n14195 ;
  assign n14199 = ( n715 & ~n801 ) | ( n715 & n12468 ) | ( ~n801 & n12468 ) ;
  assign n14200 = n854 & ~n6355 ;
  assign n14201 = n382 & n14200 ;
  assign n14202 = n2576 | n12279 ;
  assign n14203 = ( n5328 & ~n14201 ) | ( n5328 & n14202 ) | ( ~n14201 & n14202 ) ;
  assign n14204 = n5344 ^ n2989 ^ 1'b0 ;
  assign n14205 = n9072 ^ n6063 ^ n4750 ;
  assign n14206 = ( n12626 & ~n14204 ) | ( n12626 & n14205 ) | ( ~n14204 & n14205 ) ;
  assign n14207 = ( n14199 & n14203 ) | ( n14199 & ~n14206 ) | ( n14203 & ~n14206 ) ;
  assign n14209 = n8178 ^ n6480 ^ n973 ;
  assign n14208 = n13104 ^ n6090 ^ 1'b0 ;
  assign n14210 = n14209 ^ n14208 ^ 1'b0 ;
  assign n14211 = n11726 ^ n2436 ^ x19 ;
  assign n14212 = ( n885 & n1416 ) | ( n885 & ~n5468 ) | ( n1416 & ~n5468 ) ;
  assign n14213 = n14212 ^ n9193 ^ 1'b0 ;
  assign n14214 = n5240 ^ n4517 ^ 1'b0 ;
  assign n14215 = n7073 | n14214 ;
  assign n14216 = n1307 | n3754 ;
  assign n14217 = n14216 ^ n4910 ^ 1'b0 ;
  assign n14218 = ~n14215 & n14217 ;
  assign n14219 = n14218 ^ n9871 ^ 1'b0 ;
  assign n14221 = ( ~n7813 & n10897 ) | ( ~n7813 & n13405 ) | ( n10897 & n13405 ) ;
  assign n14222 = n14221 ^ n7884 ^ 1'b0 ;
  assign n14223 = n7971 ^ n6238 ^ 1'b0 ;
  assign n14224 = n1072 & n4842 ;
  assign n14225 = ~n12707 & n14224 ;
  assign n14226 = ( n8854 & n14223 ) | ( n8854 & n14225 ) | ( n14223 & n14225 ) ;
  assign n14227 = n14222 & n14226 ;
  assign n14220 = n10670 | n13659 ;
  assign n14228 = n14227 ^ n14220 ^ 1'b0 ;
  assign n14229 = n10085 ^ n7952 ^ n373 ;
  assign n14230 = ( n4924 & n5932 ) | ( n4924 & ~n11480 ) | ( n5932 & ~n11480 ) ;
  assign n14231 = ~n1960 & n14230 ;
  assign n14232 = n9557 ^ n4022 ^ n2632 ;
  assign n14233 = ( n5737 & ~n12437 ) | ( n5737 & n14232 ) | ( ~n12437 & n14232 ) ;
  assign n14234 = n13730 ^ n772 ^ 1'b0 ;
  assign n14235 = ~n14233 & n14234 ;
  assign n14237 = ~n4192 & n9366 ;
  assign n14236 = n11089 ^ n6564 ^ 1'b0 ;
  assign n14238 = n14237 ^ n14236 ^ 1'b0 ;
  assign n14239 = n14235 & n14238 ;
  assign n14240 = ( ~n4248 & n4757 ) | ( ~n4248 & n6872 ) | ( n4757 & n6872 ) ;
  assign n14241 = n6105 & ~n14240 ;
  assign n14246 = n8740 ^ n5932 ^ n1412 ;
  assign n14242 = ( ~n4434 & n5919 ) | ( ~n4434 & n6334 ) | ( n5919 & n6334 ) ;
  assign n14243 = n1745 & ~n14242 ;
  assign n14244 = n14243 ^ n5530 ^ n4198 ;
  assign n14245 = n271 & ~n14244 ;
  assign n14247 = n14246 ^ n14245 ^ 1'b0 ;
  assign n14248 = n12578 ^ n5487 ^ n2124 ;
  assign n14249 = n5443 | n7813 ;
  assign n14250 = n2676 | n14249 ;
  assign n14251 = n482 & n14250 ;
  assign n14252 = n3699 | n3877 ;
  assign n14253 = ( ~n4764 & n14251 ) | ( ~n4764 & n14252 ) | ( n14251 & n14252 ) ;
  assign n14257 = ( n836 & n5465 ) | ( n836 & n5829 ) | ( n5465 & n5829 ) ;
  assign n14258 = ( n2021 & n3181 ) | ( n2021 & n14257 ) | ( n3181 & n14257 ) ;
  assign n14254 = n4937 & n7141 ;
  assign n14255 = n14254 ^ n6707 ^ 1'b0 ;
  assign n14256 = n14255 ^ n12015 ^ n5811 ;
  assign n14259 = n14258 ^ n14256 ^ n12060 ;
  assign n14260 = ( n3873 & n7378 ) | ( n3873 & ~n8058 ) | ( n7378 & ~n8058 ) ;
  assign n14261 = n14260 ^ n5138 ^ 1'b0 ;
  assign n14262 = n3311 | n14261 ;
  assign n14263 = n2547 | n5246 ;
  assign n14264 = n14263 ^ n13583 ^ 1'b0 ;
  assign n14265 = n14262 | n14264 ;
  assign n14270 = n8389 ^ n3927 ^ n916 ;
  assign n14267 = ( x228 & n378 ) | ( x228 & ~n711 ) | ( n378 & ~n711 ) ;
  assign n14266 = ( n3781 & ~n7768 ) | ( n3781 & n9917 ) | ( ~n7768 & n9917 ) ;
  assign n14268 = n14267 ^ n14266 ^ n10952 ;
  assign n14269 = n12784 | n14268 ;
  assign n14271 = n14270 ^ n14269 ^ 1'b0 ;
  assign n14272 = ( n5656 & n10695 ) | ( n5656 & n14271 ) | ( n10695 & n14271 ) ;
  assign n14273 = ~n1124 & n10813 ;
  assign n14274 = ~n3965 & n14273 ;
  assign n14275 = n2414 & n3151 ;
  assign n14276 = x112 & ~n4521 ;
  assign n14277 = n14275 & n14276 ;
  assign n14278 = n2652 & ~n3383 ;
  assign n14279 = ( n3865 & n7981 ) | ( n3865 & n14278 ) | ( n7981 & n14278 ) ;
  assign n14280 = x146 & ~n3247 ;
  assign n14284 = ( n4300 & n6097 ) | ( n4300 & n6141 ) | ( n6097 & n6141 ) ;
  assign n14281 = n5964 ^ n1718 ^ 1'b0 ;
  assign n14282 = n9847 | n14281 ;
  assign n14283 = n14282 ^ n12944 ^ n911 ;
  assign n14285 = n14284 ^ n14283 ^ n12062 ;
  assign n14286 = n14285 ^ n10112 ^ n2021 ;
  assign n14287 = n14280 & n14286 ;
  assign n14288 = n14287 ^ x235 ^ 1'b0 ;
  assign n14289 = ( n324 & n14279 ) | ( n324 & ~n14288 ) | ( n14279 & ~n14288 ) ;
  assign n14290 = n2590 & ~n8477 ;
  assign n14291 = n14290 ^ n8197 ^ n7339 ;
  assign n14292 = ~n11520 & n12036 ;
  assign n14293 = ( n3125 & n6076 ) | ( n3125 & n14292 ) | ( n6076 & n14292 ) ;
  assign n14294 = n7925 ^ n3500 ^ n1377 ;
  assign n14295 = x230 & n534 ;
  assign n14296 = n14295 ^ n5054 ^ 1'b0 ;
  assign n14297 = ( ~n6301 & n7515 ) | ( ~n6301 & n14296 ) | ( n7515 & n14296 ) ;
  assign n14298 = n14297 ^ n13479 ^ 1'b0 ;
  assign n14299 = n6657 ^ n4539 ^ n1548 ;
  assign n14314 = ( n617 & ~n7901 ) | ( n617 & n11182 ) | ( ~n7901 & n11182 ) ;
  assign n14310 = n3296 ^ n2168 ^ n1025 ;
  assign n14311 = ( n725 & ~n7042 ) | ( n725 & n14310 ) | ( ~n7042 & n14310 ) ;
  assign n14312 = n10862 & ~n14311 ;
  assign n14313 = n9092 & n14312 ;
  assign n14300 = n5354 ^ n790 ^ 1'b0 ;
  assign n14301 = n3695 & n5974 ;
  assign n14302 = n14301 ^ n4102 ^ 1'b0 ;
  assign n14303 = ( n3371 & n3488 ) | ( n3371 & n14302 ) | ( n3488 & n14302 ) ;
  assign n14304 = ( n6311 & n14197 ) | ( n6311 & n14303 ) | ( n14197 & n14303 ) ;
  assign n14305 = ( ~n5362 & n14300 ) | ( ~n5362 & n14304 ) | ( n14300 & n14304 ) ;
  assign n14306 = n3973 ^ x226 ^ 1'b0 ;
  assign n14307 = n14306 ^ n6862 ^ 1'b0 ;
  assign n14308 = n9733 & ~n14307 ;
  assign n14309 = n14305 & n14308 ;
  assign n14315 = n14314 ^ n14313 ^ n14309 ;
  assign n14316 = n2880 & ~n8170 ;
  assign n14317 = n4883 | n14316 ;
  assign n14318 = n14317 ^ n13448 ^ 1'b0 ;
  assign n14319 = n10737 & n14318 ;
  assign n14320 = ~n2989 & n6207 ;
  assign n14321 = n14320 ^ n8388 ^ 1'b0 ;
  assign n14322 = ( n5003 & n8105 ) | ( n5003 & n14321 ) | ( n8105 & n14321 ) ;
  assign n14323 = n12409 ^ n1367 ^ 1'b0 ;
  assign n14324 = ~n2753 & n14323 ;
  assign n14325 = ( n261 & n10447 ) | ( n261 & ~n14324 ) | ( n10447 & ~n14324 ) ;
  assign n14326 = n14325 ^ n295 ^ 1'b0 ;
  assign n14327 = n10953 & n14326 ;
  assign n14328 = n12357 ^ n5916 ^ 1'b0 ;
  assign n14329 = n11897 ^ n4432 ^ 1'b0 ;
  assign n14330 = ( x114 & n14328 ) | ( x114 & ~n14329 ) | ( n14328 & ~n14329 ) ;
  assign n14331 = n6816 & ~n12006 ;
  assign n14332 = n14331 ^ n9857 ^ 1'b0 ;
  assign n14333 = n10359 & ~n12461 ;
  assign n14334 = ( n353 & ~n5210 ) | ( n353 & n5654 ) | ( ~n5210 & n5654 ) ;
  assign n14335 = n1882 | n14334 ;
  assign n14337 = n1184 ^ n1111 ^ 1'b0 ;
  assign n14338 = ~n1276 & n14337 ;
  assign n14339 = n14338 ^ n866 ^ 1'b0 ;
  assign n14340 = ( n4109 & n8010 ) | ( n4109 & ~n14339 ) | ( n8010 & ~n14339 ) ;
  assign n14336 = ( n2627 & ~n4445 ) | ( n2627 & n9232 ) | ( ~n4445 & n9232 ) ;
  assign n14341 = n14340 ^ n14336 ^ n3004 ;
  assign n14342 = ( n6680 & n14335 ) | ( n6680 & ~n14341 ) | ( n14335 & ~n14341 ) ;
  assign n14343 = ( x182 & n1197 ) | ( x182 & ~n4589 ) | ( n1197 & ~n4589 ) ;
  assign n14344 = n5022 ^ n3365 ^ n2273 ;
  assign n14345 = n14344 ^ n429 ^ 1'b0 ;
  assign n14346 = n14345 ^ n4402 ^ 1'b0 ;
  assign n14347 = n14343 & ~n14346 ;
  assign n14349 = ( n1906 & n4933 ) | ( n1906 & n7781 ) | ( n4933 & n7781 ) ;
  assign n14348 = n12142 ^ n4796 ^ n2145 ;
  assign n14350 = n14349 ^ n14348 ^ 1'b0 ;
  assign n14351 = ( ~n7676 & n14170 ) | ( ~n7676 & n14350 ) | ( n14170 & n14350 ) ;
  assign n14352 = n2774 ^ n502 ^ 1'b0 ;
  assign n14353 = n3195 | n14352 ;
  assign n14354 = n8675 | n14353 ;
  assign n14355 = n11609 ^ n5859 ^ n4258 ;
  assign n14356 = ( n8775 & ~n13438 ) | ( n8775 & n14355 ) | ( ~n13438 & n14355 ) ;
  assign n14357 = ( n1173 & ~n1916 ) | ( n1173 & n2430 ) | ( ~n1916 & n2430 ) ;
  assign n14358 = n14357 ^ n9600 ^ n4464 ;
  assign n14359 = ( x195 & ~n5582 ) | ( x195 & n13090 ) | ( ~n5582 & n13090 ) ;
  assign n14360 = n14359 ^ n7050 ^ 1'b0 ;
  assign n14361 = n12192 | n14360 ;
  assign n14362 = n8208 & ~n14361 ;
  assign n14363 = ~n11702 & n14362 ;
  assign n14364 = n9077 ^ n8477 ^ n917 ;
  assign n14365 = ~n8470 & n14364 ;
  assign n14367 = ( n1659 & n6205 ) | ( n1659 & n13674 ) | ( n6205 & n13674 ) ;
  assign n14366 = ( n585 & n6509 ) | ( n585 & ~n9810 ) | ( n6509 & ~n9810 ) ;
  assign n14368 = n14367 ^ n14366 ^ n4935 ;
  assign n14369 = n1625 | n11040 ;
  assign n14370 = n13090 | n14369 ;
  assign n14372 = n12392 ^ n10352 ^ n1061 ;
  assign n14371 = n3743 | n13018 ;
  assign n14373 = n14372 ^ n14371 ^ 1'b0 ;
  assign n14374 = n2583 & ~n10319 ;
  assign n14375 = n14374 ^ n12114 ^ n8726 ;
  assign n14379 = n2750 ^ n1569 ^ n1106 ;
  assign n14380 = n14379 ^ x92 ^ 1'b0 ;
  assign n14381 = n12702 | n14380 ;
  assign n14376 = n2185 & n2243 ;
  assign n14377 = ( n280 & ~n8150 ) | ( n280 & n14376 ) | ( ~n8150 & n14376 ) ;
  assign n14378 = n7077 & n14377 ;
  assign n14382 = n14381 ^ n14378 ^ 1'b0 ;
  assign n14383 = n5245 ^ n2619 ^ n571 ;
  assign n14384 = n14383 ^ n10599 ^ n7720 ;
  assign n14385 = ( n14375 & n14382 ) | ( n14375 & ~n14384 ) | ( n14382 & ~n14384 ) ;
  assign n14386 = n10529 ^ x248 ^ 1'b0 ;
  assign n14387 = n10513 ^ n8923 ^ 1'b0 ;
  assign n14388 = n1719 | n14387 ;
  assign n14389 = n1553 | n14388 ;
  assign n14390 = n14334 ^ n11092 ^ n1622 ;
  assign n14391 = n14390 ^ n6985 ^ n1028 ;
  assign n14392 = n14391 ^ n9690 ^ 1'b0 ;
  assign n14393 = n14389 | n14392 ;
  assign n14394 = ( x153 & n7024 ) | ( x153 & n9888 ) | ( n7024 & n9888 ) ;
  assign n14395 = n13834 ^ n9799 ^ n2266 ;
  assign n14396 = ( ~n9235 & n11629 ) | ( ~n9235 & n14395 ) | ( n11629 & n14395 ) ;
  assign n14400 = n9251 | n12366 ;
  assign n14401 = n14400 ^ n12029 ^ 1'b0 ;
  assign n14402 = n14401 ^ n892 ^ 1'b0 ;
  assign n14397 = n4685 ^ n2255 ^ n1034 ;
  assign n14398 = n1487 & ~n14397 ;
  assign n14399 = n14398 ^ n10444 ^ n825 ;
  assign n14403 = n14402 ^ n14399 ^ n2006 ;
  assign n14406 = ( n2214 & n2851 ) | ( n2214 & n10431 ) | ( n2851 & n10431 ) ;
  assign n14404 = n2696 & ~n8261 ;
  assign n14405 = n14404 ^ n13191 ^ 1'b0 ;
  assign n14407 = n14406 ^ n14405 ^ n6712 ;
  assign n14408 = n1927 ^ n522 ^ 1'b0 ;
  assign n14409 = n5596 & n14344 ;
  assign n14410 = n14409 ^ n1395 ^ 1'b0 ;
  assign n14411 = ( n3458 & n14408 ) | ( n3458 & n14410 ) | ( n14408 & n14410 ) ;
  assign n14412 = n14411 ^ n12111 ^ n11794 ;
  assign n14413 = n6340 ^ n2135 ^ n1407 ;
  assign n14414 = n14413 ^ n2615 ^ 1'b0 ;
  assign n14415 = ( n8844 & ~n10476 ) | ( n8844 & n14414 ) | ( ~n10476 & n14414 ) ;
  assign n14416 = ~n598 & n2664 ;
  assign n14417 = n7351 & n14416 ;
  assign n14418 = ~n7149 & n8881 ;
  assign n14423 = n14281 ^ n11448 ^ 1'b0 ;
  assign n14424 = ~n9023 & n14423 ;
  assign n14419 = ( ~n1873 & n3139 ) | ( ~n1873 & n8047 ) | ( n3139 & n8047 ) ;
  assign n14420 = n14419 ^ n6463 ^ n5827 ;
  assign n14421 = ( n2546 & ~n7355 ) | ( n2546 & n14420 ) | ( ~n7355 & n14420 ) ;
  assign n14422 = ~n10129 & n14421 ;
  assign n14425 = n14424 ^ n14422 ^ 1'b0 ;
  assign n14426 = ~n4965 & n9964 ;
  assign n14427 = n14426 ^ n12476 ^ x39 ;
  assign n14430 = n13608 & n13875 ;
  assign n14428 = n8630 ^ n5339 ^ 1'b0 ;
  assign n14429 = n13784 & n14428 ;
  assign n14431 = n14430 ^ n14429 ^ 1'b0 ;
  assign n14432 = n4608 ^ n3254 ^ x214 ;
  assign n14433 = ( n4520 & n12212 ) | ( n4520 & ~n14432 ) | ( n12212 & ~n14432 ) ;
  assign n14437 = n5613 ^ n3249 ^ x197 ;
  assign n14435 = n10398 ^ n6711 ^ n6184 ;
  assign n14436 = ( ~n1503 & n5935 ) | ( ~n1503 & n14435 ) | ( n5935 & n14435 ) ;
  assign n14434 = ( n4921 & n12386 ) | ( n4921 & n12675 ) | ( n12386 & n12675 ) ;
  assign n14438 = n14437 ^ n14436 ^ n14434 ;
  assign n14439 = n14438 ^ n14209 ^ 1'b0 ;
  assign n14440 = n1808 ^ n469 ^ 1'b0 ;
  assign n14441 = n14440 ^ n7654 ^ 1'b0 ;
  assign n14442 = ~n603 & n14441 ;
  assign n14443 = n6205 ^ n6119 ^ 1'b0 ;
  assign n14444 = ( n2203 & n4001 ) | ( n2203 & n6627 ) | ( n4001 & n6627 ) ;
  assign n14445 = n14444 ^ n1675 ^ n667 ;
  assign n14446 = n14445 ^ n1820 ^ x238 ;
  assign n14447 = n2197 & ~n6079 ;
  assign n14448 = n14447 ^ n13405 ^ n1292 ;
  assign n14449 = n14448 ^ n8235 ^ 1'b0 ;
  assign n14450 = ( n14443 & n14446 ) | ( n14443 & n14449 ) | ( n14446 & n14449 ) ;
  assign n14451 = n1818 & n8541 ;
  assign n14452 = ~n3265 & n14451 ;
  assign n14454 = ~n2457 & n4086 ;
  assign n14455 = n14454 ^ n3508 ^ 1'b0 ;
  assign n14453 = n14302 ^ n1444 ^ x92 ;
  assign n14456 = n14455 ^ n14453 ^ 1'b0 ;
  assign n14457 = n9077 & ~n14456 ;
  assign n14458 = n9679 ^ n7489 ^ n5339 ;
  assign n14459 = ( n8310 & n11893 ) | ( n8310 & ~n14458 ) | ( n11893 & ~n14458 ) ;
  assign n14460 = ~n1548 & n14459 ;
  assign n14461 = n6271 | n14460 ;
  assign n14462 = n9225 & ~n14461 ;
  assign n14463 = ( ~n8344 & n13582 ) | ( ~n8344 & n14462 ) | ( n13582 & n14462 ) ;
  assign n14464 = n7934 ^ n5830 ^ 1'b0 ;
  assign n14465 = ( x59 & n3986 ) | ( x59 & ~n8310 ) | ( n3986 & ~n8310 ) ;
  assign n14466 = n13410 ^ n5565 ^ 1'b0 ;
  assign n14467 = n5432 | n14466 ;
  assign n14468 = n7466 & n9316 ;
  assign n14469 = n14374 ^ n1117 ^ 1'b0 ;
  assign n14470 = n12867 | n14469 ;
  assign n14471 = ( n5111 & n8236 ) | ( n5111 & n14470 ) | ( n8236 & n14470 ) ;
  assign n14472 = ~n539 & n7585 ;
  assign n14473 = ~n2784 & n14472 ;
  assign n14474 = n14473 ^ n6827 ^ n390 ;
  assign n14475 = n7804 & ~n14474 ;
  assign n14476 = n14475 ^ n11277 ^ n7607 ;
  assign n14477 = ( n14468 & ~n14471 ) | ( n14468 & n14476 ) | ( ~n14471 & n14476 ) ;
  assign n14478 = ( n3002 & n14467 ) | ( n3002 & ~n14477 ) | ( n14467 & ~n14477 ) ;
  assign n14482 = n8618 ^ n5884 ^ n425 ;
  assign n14483 = n14482 ^ n5166 ^ 1'b0 ;
  assign n14484 = n2070 & n14483 ;
  assign n14485 = ( n486 & ~n7804 ) | ( n486 & n8226 ) | ( ~n7804 & n8226 ) ;
  assign n14486 = n14485 ^ n10216 ^ 1'b0 ;
  assign n14487 = n14484 & ~n14486 ;
  assign n14479 = ( n3207 & n12780 ) | ( n3207 & ~n14343 ) | ( n12780 & ~n14343 ) ;
  assign n14480 = n14479 ^ n9735 ^ n3538 ;
  assign n14481 = n1656 | n14480 ;
  assign n14488 = n14487 ^ n14481 ^ 1'b0 ;
  assign n14489 = n1319 & ~n4331 ;
  assign n14490 = n14489 ^ n2743 ^ 1'b0 ;
  assign n14491 = n14490 ^ n11962 ^ n3555 ;
  assign n14492 = n14491 ^ n4693 ^ 1'b0 ;
  assign n14493 = ~n6318 & n14492 ;
  assign n14494 = ~n12764 & n14493 ;
  assign n14495 = ( x68 & n3255 ) | ( x68 & n7180 ) | ( n3255 & n7180 ) ;
  assign n14496 = ( n2755 & n13545 ) | ( n2755 & ~n14495 ) | ( n13545 & ~n14495 ) ;
  assign n14497 = ( n1653 & n1661 ) | ( n1653 & n4281 ) | ( n1661 & n4281 ) ;
  assign n14498 = n14497 ^ n6985 ^ n3926 ;
  assign n14499 = ( n2612 & n7357 ) | ( n2612 & n14498 ) | ( n7357 & n14498 ) ;
  assign n14500 = ~n8307 & n9479 ;
  assign n14501 = n14500 ^ n13061 ^ x163 ;
  assign n14502 = n3676 ^ n1991 ^ 1'b0 ;
  assign n14503 = n14502 ^ n10430 ^ n5723 ;
  assign n14504 = n661 | n4388 ;
  assign n14505 = n14504 ^ n7531 ^ n547 ;
  assign n14506 = n14505 ^ n14268 ^ 1'b0 ;
  assign n14507 = ( x8 & ~n4851 ) | ( x8 & n9232 ) | ( ~n4851 & n9232 ) ;
  assign n14508 = n2542 ^ n1553 ^ n1395 ;
  assign n14509 = n3017 & n14508 ;
  assign n14510 = n14509 ^ n6328 ^ n836 ;
  assign n14511 = ( ~n13884 & n14507 ) | ( ~n13884 & n14510 ) | ( n14507 & n14510 ) ;
  assign n14512 = n5220 ^ n1033 ^ n529 ;
  assign n14513 = ~n5994 & n6285 ;
  assign n14514 = ( n10367 & ~n14512 ) | ( n10367 & n14513 ) | ( ~n14512 & n14513 ) ;
  assign n14523 = n8991 ^ n5171 ^ n1251 ;
  assign n14521 = n9281 ^ n5831 ^ 1'b0 ;
  assign n14515 = ( n666 & n959 ) | ( n666 & n1821 ) | ( n959 & n1821 ) ;
  assign n14516 = n5624 ^ n3299 ^ n649 ;
  assign n14517 = n9991 | n14516 ;
  assign n14518 = n14515 | n14517 ;
  assign n14519 = ~n1935 & n10371 ;
  assign n14520 = n14518 & n14519 ;
  assign n14522 = n14521 ^ n14520 ^ 1'b0 ;
  assign n14524 = n14523 ^ n14522 ^ n1572 ;
  assign n14525 = n11679 ^ n2667 ^ x68 ;
  assign n14526 = ~n470 & n10216 ;
  assign n14527 = n14526 ^ n10996 ^ 1'b0 ;
  assign n14528 = ( ~n6974 & n14525 ) | ( ~n6974 & n14527 ) | ( n14525 & n14527 ) ;
  assign n14529 = n12173 | n14528 ;
  assign n14530 = n14529 ^ n347 ^ 1'b0 ;
  assign n14535 = n7853 & n7982 ;
  assign n14536 = ~n5546 & n9746 ;
  assign n14537 = n14535 & n14536 ;
  assign n14532 = ( n2564 & n4156 ) | ( n2564 & n13642 ) | ( n4156 & n13642 ) ;
  assign n14531 = n9275 | n9787 ;
  assign n14533 = n14532 ^ n14531 ^ 1'b0 ;
  assign n14534 = n11266 & ~n14533 ;
  assign n14538 = n14537 ^ n14534 ^ 1'b0 ;
  assign n14540 = n9174 ^ n7176 ^ n3107 ;
  assign n14539 = ( n628 & ~n3623 ) | ( n628 & n10564 ) | ( ~n3623 & n10564 ) ;
  assign n14541 = n14540 ^ n14539 ^ n5035 ;
  assign n14542 = ( n5324 & n7082 ) | ( n5324 & n10310 ) | ( n7082 & n10310 ) ;
  assign n14545 = n4631 ^ n1420 ^ x63 ;
  assign n14544 = n4728 ^ n2704 ^ 1'b0 ;
  assign n14543 = ( n2516 & n4469 ) | ( n2516 & n6733 ) | ( n4469 & n6733 ) ;
  assign n14546 = n14545 ^ n14544 ^ n14543 ;
  assign n14547 = n14546 ^ n8750 ^ 1'b0 ;
  assign n14551 = ~n3478 & n13874 ;
  assign n14552 = ~n808 & n14551 ;
  assign n14548 = x23 & ~n2099 ;
  assign n14549 = ~n1862 & n14548 ;
  assign n14550 = n14549 ^ n10688 ^ 1'b0 ;
  assign n14553 = n14552 ^ n14550 ^ n5175 ;
  assign n14554 = n794 | n1394 ;
  assign n14555 = n1629 | n14554 ;
  assign n14556 = n10568 & n14555 ;
  assign n14557 = n5931 & n11031 ;
  assign n14558 = n14556 & n14557 ;
  assign n14559 = ( n4260 & n11207 ) | ( n4260 & ~n14558 ) | ( n11207 & ~n14558 ) ;
  assign n14561 = n11556 | n12558 ;
  assign n14560 = ~n1500 & n11071 ;
  assign n14562 = n14561 ^ n14560 ^ n1210 ;
  assign n14563 = n10106 ^ n4348 ^ n4289 ;
  assign n14564 = ( n1133 & ~n13351 ) | ( n1133 & n14563 ) | ( ~n13351 & n14563 ) ;
  assign n14565 = n14564 ^ n5058 ^ n2527 ;
  assign n14566 = n6527 & ~n10734 ;
  assign n14567 = ~n13395 & n14566 ;
  assign n14568 = n14567 ^ n14428 ^ n7252 ;
  assign n14571 = ( ~n2864 & n8588 ) | ( ~n2864 & n13007 ) | ( n8588 & n13007 ) ;
  assign n14572 = ( ~n10490 & n12436 ) | ( ~n10490 & n14571 ) | ( n12436 & n14571 ) ;
  assign n14573 = n14572 ^ n10461 ^ n3647 ;
  assign n14569 = n5212 & ~n8686 ;
  assign n14570 = n13808 & n14569 ;
  assign n14574 = n14573 ^ n14570 ^ 1'b0 ;
  assign n14581 = n11150 ^ n4973 ^ 1'b0 ;
  assign n14578 = n2227 & ~n3636 ;
  assign n14579 = n3552 & n14578 ;
  assign n14580 = n14579 ^ n12001 ^ 1'b0 ;
  assign n14575 = ( n574 & ~n1534 ) | ( n574 & n2877 ) | ( ~n1534 & n2877 ) ;
  assign n14576 = ( x164 & n10112 ) | ( x164 & n14575 ) | ( n10112 & n14575 ) ;
  assign n14577 = n14576 ^ n9382 ^ n1589 ;
  assign n14582 = n14581 ^ n14580 ^ n14577 ;
  assign n14589 = ( n1915 & n3031 ) | ( n1915 & ~n4479 ) | ( n3031 & ~n4479 ) ;
  assign n14587 = n7962 & n12502 ;
  assign n14588 = n14587 ^ n971 ^ 1'b0 ;
  assign n14583 = n13186 ^ n4449 ^ n2883 ;
  assign n14584 = n14583 ^ n5524 ^ n3659 ;
  assign n14585 = n3083 | n14584 ;
  assign n14586 = n6285 | n14585 ;
  assign n14590 = n14589 ^ n14588 ^ n14586 ;
  assign n14591 = n5921 | n14590 ;
  assign n14592 = n8590 & ~n12903 ;
  assign n14593 = ( n3337 & n8455 ) | ( n3337 & ~n8854 ) | ( n8455 & ~n8854 ) ;
  assign n14594 = n14593 ^ n14512 ^ n595 ;
  assign n14595 = ~n8434 & n11811 ;
  assign n14596 = ( n3002 & n14594 ) | ( n3002 & ~n14595 ) | ( n14594 & ~n14595 ) ;
  assign n14597 = ( n12276 & n14592 ) | ( n12276 & n14596 ) | ( n14592 & n14596 ) ;
  assign n14598 = n11144 ^ n6906 ^ 1'b0 ;
  assign n14606 = n10861 & n11269 ;
  assign n14600 = n6828 ^ n2763 ^ x65 ;
  assign n14601 = n14600 ^ n10644 ^ n10139 ;
  assign n14599 = n5942 | n6680 ;
  assign n14602 = n14601 ^ n14599 ^ n12800 ;
  assign n14603 = ( ~n3029 & n4109 ) | ( ~n3029 & n4536 ) | ( n4109 & n4536 ) ;
  assign n14604 = n14602 & n14603 ;
  assign n14605 = ( ~n7341 & n11719 ) | ( ~n7341 & n14604 ) | ( n11719 & n14604 ) ;
  assign n14607 = n14606 ^ n14605 ^ n2452 ;
  assign n14608 = ( n2508 & n3556 ) | ( n2508 & ~n3826 ) | ( n3556 & ~n3826 ) ;
  assign n14609 = n14608 ^ n14571 ^ n2106 ;
  assign n14612 = n5992 ^ x5 ^ 1'b0 ;
  assign n14613 = n14201 | n14612 ;
  assign n14610 = n12997 ^ n12102 ^ n9621 ;
  assign n14611 = n14610 ^ n13131 ^ n4147 ;
  assign n14614 = n14613 ^ n14611 ^ x223 ;
  assign n14615 = ~n419 & n1776 ;
  assign n14616 = n2329 & n14615 ;
  assign n14617 = ( ~n10167 & n13892 ) | ( ~n10167 & n14616 ) | ( n13892 & n14616 ) ;
  assign n14618 = ( n2014 & n4213 ) | ( n2014 & ~n11943 ) | ( n4213 & ~n11943 ) ;
  assign n14619 = n14618 ^ n8825 ^ x84 ;
  assign n14620 = n4191 ^ n1706 ^ 1'b0 ;
  assign n14621 = n14620 ^ n3836 ^ 1'b0 ;
  assign n14622 = n14621 ^ n4323 ^ 1'b0 ;
  assign n14623 = n14619 | n14622 ;
  assign n14624 = n6433 ^ n4467 ^ 1'b0 ;
  assign n14625 = n3572 | n14624 ;
  assign n14626 = n14625 ^ n5973 ^ 1'b0 ;
  assign n14627 = ( n11859 & ~n14623 ) | ( n11859 & n14626 ) | ( ~n14623 & n14626 ) ;
  assign n14628 = ( n348 & n2303 ) | ( n348 & ~n6222 ) | ( n2303 & ~n6222 ) ;
  assign n14629 = n14628 ^ n5450 ^ n410 ;
  assign n14630 = ( n1455 & ~n6069 ) | ( n1455 & n14629 ) | ( ~n6069 & n14629 ) ;
  assign n14631 = n11322 ^ n6730 ^ 1'b0 ;
  assign n14632 = ( n3802 & n3844 ) | ( n3802 & ~n14631 ) | ( n3844 & ~n14631 ) ;
  assign n14633 = ~n13849 & n14632 ;
  assign n14634 = n5521 ^ n3387 ^ n766 ;
  assign n14635 = n5112 | n14634 ;
  assign n14636 = ( n14630 & n14633 ) | ( n14630 & n14635 ) | ( n14633 & n14635 ) ;
  assign n14637 = n9777 | n9901 ;
  assign n14638 = n12085 & ~n14637 ;
  assign n14639 = ( x130 & ~n4099 ) | ( x130 & n4666 ) | ( ~n4099 & n4666 ) ;
  assign n14640 = n8186 & n14639 ;
  assign n14641 = ( n3813 & ~n5098 ) | ( n3813 & n9141 ) | ( ~n5098 & n9141 ) ;
  assign n14642 = n14641 ^ n8061 ^ 1'b0 ;
  assign n14643 = n11147 ^ n5147 ^ n279 ;
  assign n14644 = ( ~n3781 & n10783 ) | ( ~n3781 & n14643 ) | ( n10783 & n14643 ) ;
  assign n14645 = n14526 ^ n9763 ^ 1'b0 ;
  assign n14646 = ( n4902 & ~n14644 ) | ( n4902 & n14645 ) | ( ~n14644 & n14645 ) ;
  assign n14647 = n1714 & ~n3538 ;
  assign n14649 = n9151 ^ n5171 ^ x111 ;
  assign n14648 = ( ~n6560 & n12670 ) | ( ~n6560 & n14320 ) | ( n12670 & n14320 ) ;
  assign n14650 = n14649 ^ n14648 ^ 1'b0 ;
  assign n14651 = ~n1391 & n14650 ;
  assign n14652 = n1732 & n10609 ;
  assign n14653 = n7735 ^ n4873 ^ n3342 ;
  assign n14654 = ( n2801 & ~n9473 ) | ( n2801 & n14653 ) | ( ~n9473 & n14653 ) ;
  assign n14655 = n2062 & ~n3520 ;
  assign n14656 = n10486 & n14655 ;
  assign n14657 = n6019 ^ n3715 ^ 1'b0 ;
  assign n14658 = n6619 ^ n3269 ^ 1'b0 ;
  assign n14659 = n14657 | n14658 ;
  assign n14660 = ( n3338 & n4710 ) | ( n3338 & ~n7378 ) | ( n4710 & ~n7378 ) ;
  assign n14661 = ~n602 & n14660 ;
  assign n14662 = ( ~n3207 & n4130 ) | ( ~n3207 & n14661 ) | ( n4130 & n14661 ) ;
  assign n14663 = ( n11641 & n12350 ) | ( n11641 & n14662 ) | ( n12350 & n14662 ) ;
  assign n14664 = n9797 | n13538 ;
  assign n14665 = n14664 ^ n8020 ^ 1'b0 ;
  assign n14666 = n676 | n10699 ;
  assign n14667 = n14666 ^ n5110 ^ 1'b0 ;
  assign n14668 = ~n5710 & n14667 ;
  assign n14669 = n2064 & n14668 ;
  assign n14670 = n11282 | n14669 ;
  assign n14671 = ( n14213 & ~n14665 ) | ( n14213 & n14670 ) | ( ~n14665 & n14670 ) ;
  assign n14672 = n12456 ^ n9794 ^ 1'b0 ;
  assign n14673 = n9830 & n12534 ;
  assign n14674 = n2882 & n3158 ;
  assign n14675 = n14674 ^ n7342 ^ n2035 ;
  assign n14676 = n3750 & n14675 ;
  assign n14677 = n14673 & n14676 ;
  assign n14681 = n1433 ^ n1146 ^ n430 ;
  assign n14682 = ( n3894 & n10235 ) | ( n3894 & n14681 ) | ( n10235 & n14681 ) ;
  assign n14683 = n3653 ^ x217 ^ 1'b0 ;
  assign n14684 = ~n4703 & n14683 ;
  assign n14685 = n14682 & n14684 ;
  assign n14679 = ( n2185 & n4776 ) | ( n2185 & n8078 ) | ( n4776 & n8078 ) ;
  assign n14678 = ( n4357 & n7353 ) | ( n4357 & ~n14047 ) | ( n7353 & ~n14047 ) ;
  assign n14680 = n14679 ^ n14678 ^ n1477 ;
  assign n14686 = n14685 ^ n14680 ^ 1'b0 ;
  assign n14687 = n4477 ^ n2519 ^ n874 ;
  assign n14688 = n7856 | n14687 ;
  assign n14689 = n4934 & n14688 ;
  assign n14690 = n8250 & ~n10947 ;
  assign n14691 = n14690 ^ n10650 ^ 1'b0 ;
  assign n14692 = ~n8621 & n14691 ;
  assign n14693 = n14692 ^ n9260 ^ 1'b0 ;
  assign n14694 = n2998 | n12816 ;
  assign n14695 = n3338 & n9224 ;
  assign n14696 = ~n5820 & n14695 ;
  assign n14697 = ( n1503 & ~n12439 ) | ( n1503 & n14696 ) | ( ~n12439 & n14696 ) ;
  assign n14698 = n13942 & ~n14697 ;
  assign n14704 = ~n4279 & n4923 ;
  assign n14705 = n3713 & n14704 ;
  assign n14699 = n4245 & ~n9864 ;
  assign n14700 = n14699 ^ n1487 ^ x46 ;
  assign n14701 = n1970 | n2222 ;
  assign n14702 = n14701 ^ n12242 ^ 1'b0 ;
  assign n14703 = ( n12013 & ~n14700 ) | ( n12013 & n14702 ) | ( ~n14700 & n14702 ) ;
  assign n14706 = n14705 ^ n14703 ^ n10781 ;
  assign n14707 = n5435 ^ n3017 ^ 1'b0 ;
  assign n14708 = n278 | n7686 ;
  assign n14711 = n6770 ^ x80 ^ 1'b0 ;
  assign n14710 = n7043 & n10951 ;
  assign n14712 = n14711 ^ n14710 ^ 1'b0 ;
  assign n14709 = n3280 | n5166 ;
  assign n14713 = n14712 ^ n14709 ^ 1'b0 ;
  assign n14714 = n14713 ^ n5384 ^ 1'b0 ;
  assign n14715 = n14708 & ~n14714 ;
  assign n14716 = n14715 ^ n11955 ^ 1'b0 ;
  assign n14717 = n14707 & ~n14716 ;
  assign n14718 = ( n8013 & n9042 ) | ( n8013 & ~n14717 ) | ( n9042 & ~n14717 ) ;
  assign n14720 = ( n1084 & ~n1842 ) | ( n1084 & n8220 ) | ( ~n1842 & n8220 ) ;
  assign n14721 = ( n4026 & n4282 ) | ( n4026 & n14720 ) | ( n4282 & n14720 ) ;
  assign n14722 = n14721 ^ n8599 ^ n3524 ;
  assign n14723 = ( ~n4235 & n10163 ) | ( ~n4235 & n14722 ) | ( n10163 & n14722 ) ;
  assign n14719 = ~n5293 & n11298 ;
  assign n14724 = n14723 ^ n14719 ^ n7182 ;
  assign n14725 = n4371 ^ n2502 ^ n2461 ;
  assign n14726 = n1611 & ~n3617 ;
  assign n14727 = n14726 ^ n8513 ^ 1'b0 ;
  assign n14728 = n8001 ^ n6638 ^ 1'b0 ;
  assign n14729 = n14727 | n14728 ;
  assign n14730 = n4752 & n4965 ;
  assign n14731 = n14730 ^ n5218 ^ 1'b0 ;
  assign n14732 = n14731 ^ n9479 ^ 1'b0 ;
  assign n14733 = n14729 | n14732 ;
  assign n14734 = ( n9771 & ~n14725 ) | ( n9771 & n14733 ) | ( ~n14725 & n14733 ) ;
  assign n14735 = n13564 ^ n5347 ^ 1'b0 ;
  assign n14736 = n289 & ~n14735 ;
  assign n14737 = ~n5903 & n11034 ;
  assign n14738 = n14737 ^ n9859 ^ 1'b0 ;
  assign n14739 = n396 & n14738 ;
  assign n14740 = n14739 ^ n13694 ^ 1'b0 ;
  assign n14741 = n14736 & ~n14740 ;
  assign n14742 = n3213 ^ n2186 ^ n561 ;
  assign n14743 = n14742 ^ n3851 ^ 1'b0 ;
  assign n14744 = ~n5740 & n14743 ;
  assign n14745 = n7290 ^ n5637 ^ x43 ;
  assign n14746 = ( n1746 & n12041 ) | ( n1746 & ~n14745 ) | ( n12041 & ~n14745 ) ;
  assign n14747 = n14744 & ~n14746 ;
  assign n14748 = n4036 & n14747 ;
  assign n14749 = n8119 & ~n11322 ;
  assign n14750 = ( n882 & n3858 ) | ( n882 & n14749 ) | ( n3858 & n14749 ) ;
  assign n14751 = n5928 & ~n14750 ;
  assign n14752 = n14751 ^ n11242 ^ 1'b0 ;
  assign n14753 = ( n1529 & ~n9264 ) | ( n1529 & n14752 ) | ( ~n9264 & n14752 ) ;
  assign n14754 = n632 | n7515 ;
  assign n14755 = n2014 & ~n14754 ;
  assign n14756 = n9170 & ~n14755 ;
  assign n14757 = n6490 & n14756 ;
  assign n14758 = ( n1385 & n14753 ) | ( n1385 & n14757 ) | ( n14753 & n14757 ) ;
  assign n14759 = n1224 & ~n1564 ;
  assign n14760 = n14759 ^ n5185 ^ n4524 ;
  assign n14761 = n2804 | n14760 ;
  assign n14762 = ( n465 & ~n2509 ) | ( n465 & n10570 ) | ( ~n2509 & n10570 ) ;
  assign n14763 = ( ~n8699 & n14761 ) | ( ~n8699 & n14762 ) | ( n14761 & n14762 ) ;
  assign n14764 = n14763 ^ n10283 ^ 1'b0 ;
  assign n14765 = n4263 | n7457 ;
  assign n14766 = ( n1730 & n2427 ) | ( n1730 & n7100 ) | ( n2427 & n7100 ) ;
  assign n14767 = n9745 ^ n8123 ^ n5308 ;
  assign n14768 = n14767 ^ n1149 ^ 1'b0 ;
  assign n14769 = n14766 | n14768 ;
  assign n14770 = n561 | n14769 ;
  assign n14771 = n11611 | n14770 ;
  assign n14772 = n13773 ^ n7844 ^ n5393 ;
  assign n14773 = n14772 ^ n3980 ^ n1928 ;
  assign n14774 = n14773 ^ n14288 ^ n4460 ;
  assign n14777 = n5609 | n14084 ;
  assign n14775 = n13982 ^ n2533 ^ x57 ;
  assign n14776 = n14775 ^ n4866 ^ 1'b0 ;
  assign n14778 = n14777 ^ n14776 ^ n1813 ;
  assign n14779 = n1784 & ~n3852 ;
  assign n14780 = n14779 ^ n14572 ^ n3987 ;
  assign n14781 = n1437 | n2192 ;
  assign n14782 = n14781 ^ n9443 ^ 1'b0 ;
  assign n14783 = n6453 ^ n1093 ^ n841 ;
  assign n14784 = ( n5206 & ~n14782 ) | ( n5206 & n14783 ) | ( ~n14782 & n14783 ) ;
  assign n14785 = ( n2156 & n2233 ) | ( n2156 & ~n14784 ) | ( n2233 & ~n14784 ) ;
  assign n14788 = ( n2657 & n3268 ) | ( n2657 & n12876 ) | ( n3268 & n12876 ) ;
  assign n14789 = n10791 & n14788 ;
  assign n14786 = x164 & n4891 ;
  assign n14787 = n9061 & n14786 ;
  assign n14790 = n14789 ^ n14787 ^ n8780 ;
  assign n14791 = ( n8023 & n14785 ) | ( n8023 & ~n14790 ) | ( n14785 & ~n14790 ) ;
  assign n14792 = n3838 ^ n2506 ^ n1873 ;
  assign n14793 = n14792 ^ n14302 ^ n10418 ;
  assign n14794 = n14793 ^ n9385 ^ 1'b0 ;
  assign n14795 = n14794 ^ n14165 ^ n7581 ;
  assign n14796 = n7389 ^ n5689 ^ 1'b0 ;
  assign n14797 = n14795 & n14796 ;
  assign n14798 = ~n3851 & n8799 ;
  assign n14799 = n7202 & n14798 ;
  assign n14800 = n13345 | n14799 ;
  assign n14801 = ( n2947 & n7907 ) | ( n2947 & ~n8048 ) | ( n7907 & ~n8048 ) ;
  assign n14802 = n12346 & ~n13106 ;
  assign n14803 = n5762 | n8663 ;
  assign n14804 = n2008 & ~n14803 ;
  assign n14805 = ( n1707 & n9643 ) | ( n1707 & n12678 ) | ( n9643 & n12678 ) ;
  assign n14806 = n5176 & n14805 ;
  assign n14807 = n1890 | n11496 ;
  assign n14808 = n14807 ^ n5915 ^ 1'b0 ;
  assign n14809 = n10582 ^ n1762 ^ x112 ;
  assign n14810 = n5088 & n14809 ;
  assign n14811 = ~n14808 & n14810 ;
  assign n14812 = n12310 ^ n7949 ^ n3547 ;
  assign n14814 = ~n5731 & n9863 ;
  assign n14815 = n14814 ^ n6732 ^ 1'b0 ;
  assign n14813 = n8410 ^ n881 ^ 1'b0 ;
  assign n14816 = n14815 ^ n14813 ^ 1'b0 ;
  assign n14817 = ~n841 & n7251 ;
  assign n14818 = n14817 ^ n8462 ^ 1'b0 ;
  assign n14819 = n13895 ^ n1961 ^ 1'b0 ;
  assign n14824 = n12085 ^ n3316 ^ 1'b0 ;
  assign n14825 = n2883 & n14824 ;
  assign n14820 = n9621 ^ n3547 ^ 1'b0 ;
  assign n14821 = n5809 | n14820 ;
  assign n14822 = n14150 ^ n6535 ^ 1'b0 ;
  assign n14823 = ( n11383 & ~n14821 ) | ( n11383 & n14822 ) | ( ~n14821 & n14822 ) ;
  assign n14826 = n14825 ^ n14823 ^ n7705 ;
  assign n14827 = n13614 ^ n7290 ^ n4330 ;
  assign n14830 = ( n4348 & ~n4591 ) | ( n4348 & n6790 ) | ( ~n4591 & n6790 ) ;
  assign n14828 = n2044 & ~n5446 ;
  assign n14829 = n14828 ^ n3232 ^ 1'b0 ;
  assign n14831 = n14830 ^ n14829 ^ 1'b0 ;
  assign n14832 = n14827 & ~n14831 ;
  assign n14833 = n13110 ^ n11693 ^ 1'b0 ;
  assign n14835 = ( n3007 & n3936 ) | ( n3007 & ~n5257 ) | ( n3936 & ~n5257 ) ;
  assign n14836 = n14835 ^ n3826 ^ 1'b0 ;
  assign n14834 = n6648 ^ n951 ^ 1'b0 ;
  assign n14837 = n14836 ^ n14834 ^ n7769 ;
  assign n14838 = ( n492 & n3128 ) | ( n492 & ~n14837 ) | ( n3128 & ~n14837 ) ;
  assign n14839 = n13079 & ~n14838 ;
  assign n14840 = n14839 ^ n8744 ^ 1'b0 ;
  assign n14846 = n12483 ^ n5727 ^ 1'b0 ;
  assign n14847 = n8203 ^ n6760 ^ 1'b0 ;
  assign n14848 = n4283 | n14847 ;
  assign n14849 = n14846 & ~n14848 ;
  assign n14841 = n11188 ^ n1883 ^ 1'b0 ;
  assign n14842 = n3566 & ~n14841 ;
  assign n14843 = ( ~n6021 & n7045 ) | ( ~n6021 & n8844 ) | ( n7045 & n8844 ) ;
  assign n14844 = n14843 ^ n7988 ^ n5107 ;
  assign n14845 = n14842 & n14844 ;
  assign n14850 = n14849 ^ n14845 ^ 1'b0 ;
  assign n14851 = ( n3942 & n11673 ) | ( n3942 & n14002 ) | ( n11673 & n14002 ) ;
  assign n14852 = ~n1844 & n14851 ;
  assign n14853 = ( n11534 & n13395 ) | ( n11534 & n14852 ) | ( n13395 & n14852 ) ;
  assign n14854 = ( ~n4025 & n8506 ) | ( ~n4025 & n8866 ) | ( n8506 & n8866 ) ;
  assign n14855 = n5668 ^ n4346 ^ n459 ;
  assign n14856 = n6937 ^ n3449 ^ n683 ;
  assign n14857 = n14856 ^ n12420 ^ n2774 ;
  assign n14858 = n1717 & n9301 ;
  assign n14859 = n14857 & n14858 ;
  assign n14860 = ( ~n8674 & n11088 ) | ( ~n8674 & n14859 ) | ( n11088 & n14859 ) ;
  assign n14864 = ~n2729 & n3904 ;
  assign n14865 = n14864 ^ n6794 ^ 1'b0 ;
  assign n14866 = n14865 ^ n12844 ^ n10547 ;
  assign n14861 = n11429 ^ n4072 ^ n813 ;
  assign n14862 = n4005 ^ n894 ^ 1'b0 ;
  assign n14863 = ( n6565 & ~n14861 ) | ( n6565 & n14862 ) | ( ~n14861 & n14862 ) ;
  assign n14867 = n14866 ^ n14863 ^ n3352 ;
  assign n14868 = n9639 ^ n1612 ^ 1'b0 ;
  assign n14869 = n11856 ^ n7785 ^ n6122 ;
  assign n14870 = ( ~n3226 & n4449 ) | ( ~n3226 & n4634 ) | ( n4449 & n4634 ) ;
  assign n14871 = n14870 ^ n6933 ^ n1970 ;
  assign n14872 = n14871 ^ n6763 ^ n1422 ;
  assign n14873 = n8037 ^ n5609 ^ 1'b0 ;
  assign n14874 = n3795 & ~n14873 ;
  assign n14875 = ( n9007 & n14872 ) | ( n9007 & ~n14874 ) | ( n14872 & ~n14874 ) ;
  assign n14876 = n13075 ^ n9958 ^ n5435 ;
  assign n14877 = n11657 ^ n9101 ^ n1805 ;
  assign n14878 = n9411 ^ n5621 ^ 1'b0 ;
  assign n14879 = n14878 ^ n11063 ^ n8859 ;
  assign n14880 = ~n14877 & n14879 ;
  assign n14881 = ( n344 & n463 ) | ( n344 & n13132 ) | ( n463 & n13132 ) ;
  assign n14882 = n14881 ^ n535 ^ 1'b0 ;
  assign n14883 = n6955 ^ n2960 ^ n2075 ;
  assign n14884 = n14883 ^ n14635 ^ n836 ;
  assign n14885 = n4411 ^ n3239 ^ n1646 ;
  assign n14887 = n2726 ^ n2523 ^ n892 ;
  assign n14886 = n6541 | n12249 ;
  assign n14888 = n14887 ^ n14886 ^ 1'b0 ;
  assign n14889 = n11300 ^ n7581 ^ n6806 ;
  assign n14890 = n14889 ^ n9835 ^ n1867 ;
  assign n14891 = ( ~n10708 & n14888 ) | ( ~n10708 & n14890 ) | ( n14888 & n14890 ) ;
  assign n14892 = ( n2558 & n3009 ) | ( n2558 & n5755 ) | ( n3009 & n5755 ) ;
  assign n14893 = n984 & n2659 ;
  assign n14894 = n14893 ^ n2272 ^ 1'b0 ;
  assign n14895 = n14892 & n14894 ;
  assign n14896 = ( n931 & ~n4548 ) | ( n931 & n4777 ) | ( ~n4548 & n4777 ) ;
  assign n14897 = n14896 ^ n6095 ^ n676 ;
  assign n14898 = ( n2164 & ~n3429 ) | ( n2164 & n14897 ) | ( ~n3429 & n14897 ) ;
  assign n14900 = n11760 ^ n6990 ^ n666 ;
  assign n14899 = ( ~n352 & n1600 ) | ( ~n352 & n14098 ) | ( n1600 & n14098 ) ;
  assign n14901 = n14900 ^ n14899 ^ n674 ;
  assign n14902 = n14898 & ~n14901 ;
  assign n14903 = n14902 ^ n366 ^ 1'b0 ;
  assign n14904 = n14903 ^ n13942 ^ n4510 ;
  assign n14905 = ( n10442 & n10620 ) | ( n10442 & ~n14904 ) | ( n10620 & ~n14904 ) ;
  assign n14906 = n3255 ^ n697 ^ 1'b0 ;
  assign n14907 = n14906 ^ n3452 ^ 1'b0 ;
  assign n14908 = n14907 ^ n13441 ^ n4087 ;
  assign n14909 = n14908 ^ n12836 ^ n1542 ;
  assign n14910 = ( n492 & ~n9683 ) | ( n492 & n14909 ) | ( ~n9683 & n14909 ) ;
  assign n14911 = ( ~n565 & n11232 ) | ( ~n565 & n14455 ) | ( n11232 & n14455 ) ;
  assign n14912 = ( ~n9765 & n13443 ) | ( ~n9765 & n14911 ) | ( n13443 & n14911 ) ;
  assign n14913 = n7569 & ~n14912 ;
  assign n14914 = n14913 ^ n9932 ^ 1'b0 ;
  assign n14915 = n3427 ^ n1706 ^ n1466 ;
  assign n14916 = ~n5010 & n8075 ;
  assign n14917 = ~n7219 & n14916 ;
  assign n14918 = n14917 ^ n356 ^ 1'b0 ;
  assign n14919 = n14915 | n14918 ;
  assign n14920 = n2527 | n10303 ;
  assign n14921 = n600 | n14920 ;
  assign n14922 = n9128 & ~n10189 ;
  assign n14923 = n13236 ^ n6951 ^ 1'b0 ;
  assign n14924 = n5583 | n14923 ;
  assign n14928 = n484 | n7428 ;
  assign n14929 = n9135 & ~n14928 ;
  assign n14927 = n11384 ^ n8393 ^ 1'b0 ;
  assign n14925 = n627 ^ x118 ^ 1'b0 ;
  assign n14926 = n3732 & ~n14925 ;
  assign n14930 = n14929 ^ n14927 ^ n14926 ;
  assign n14931 = n14930 ^ n3902 ^ n2884 ;
  assign n14932 = ( ~n4715 & n6386 ) | ( ~n4715 & n14931 ) | ( n6386 & n14931 ) ;
  assign n14933 = ( n1343 & ~n13693 ) | ( n1343 & n14932 ) | ( ~n13693 & n14932 ) ;
  assign n14934 = n6849 ^ n5597 ^ n4328 ;
  assign n14935 = n14934 ^ n10030 ^ 1'b0 ;
  assign n14936 = n9439 & n14935 ;
  assign n14937 = n1172 & n14936 ;
  assign n14938 = n14937 ^ n2871 ^ 1'b0 ;
  assign n14939 = ( n8885 & ~n14933 ) | ( n8885 & n14938 ) | ( ~n14933 & n14938 ) ;
  assign n14940 = n1708 ^ x244 ^ 1'b0 ;
  assign n14945 = n6193 ^ n3819 ^ 1'b0 ;
  assign n14946 = ( n4118 & ~n8130 ) | ( n4118 & n14945 ) | ( ~n8130 & n14945 ) ;
  assign n14941 = ( n2859 & n3270 ) | ( n2859 & n5935 ) | ( n3270 & n5935 ) ;
  assign n14942 = n10407 ^ n1664 ^ 1'b0 ;
  assign n14943 = ~n14941 & n14942 ;
  assign n14944 = ( n3794 & n3931 ) | ( n3794 & ~n14943 ) | ( n3931 & ~n14943 ) ;
  assign n14947 = n14946 ^ n14944 ^ n12147 ;
  assign n14948 = n12696 ^ n6470 ^ 1'b0 ;
  assign n14950 = n8462 ^ n916 ^ 1'b0 ;
  assign n14949 = ~n495 & n8240 ;
  assign n14951 = n14950 ^ n14949 ^ 1'b0 ;
  assign n14952 = ( n3460 & n6963 ) | ( n3460 & ~n11780 ) | ( n6963 & ~n11780 ) ;
  assign n14953 = n12379 ^ n5916 ^ 1'b0 ;
  assign n14954 = n14952 & ~n14953 ;
  assign n14959 = n2525 & ~n4279 ;
  assign n14960 = n14959 ^ n6392 ^ 1'b0 ;
  assign n14958 = ~n1808 & n6651 ;
  assign n14956 = n2635 ^ n2558 ^ n1169 ;
  assign n14955 = ( n1028 & ~n3298 ) | ( n1028 & n12442 ) | ( ~n3298 & n12442 ) ;
  assign n14957 = n14956 ^ n14955 ^ n7617 ;
  assign n14961 = n14960 ^ n14958 ^ n14957 ;
  assign n14962 = n14242 ^ n7769 ^ n727 ;
  assign n14963 = ( n1484 & n5922 ) | ( n1484 & ~n11751 ) | ( n5922 & ~n11751 ) ;
  assign n14964 = ( n574 & ~n801 ) | ( n574 & n3899 ) | ( ~n801 & n3899 ) ;
  assign n14965 = ~n13007 & n14964 ;
  assign n14966 = ~n9371 & n14965 ;
  assign n14967 = n7054 ^ n4415 ^ n1233 ;
  assign n14968 = ( n12578 & n14966 ) | ( n12578 & ~n14967 ) | ( n14966 & ~n14967 ) ;
  assign n14969 = ( n12211 & ~n12257 ) | ( n12211 & n14968 ) | ( ~n12257 & n14968 ) ;
  assign n14970 = x227 | n8031 ;
  assign n14971 = n14970 ^ n8302 ^ 1'b0 ;
  assign n14972 = n315 & n4496 ;
  assign n14973 = n10164 & n14972 ;
  assign n14974 = n13262 | n14973 ;
  assign n14975 = n14974 ^ n5113 ^ 1'b0 ;
  assign n14976 = ( ~n2983 & n10212 ) | ( ~n2983 & n11976 ) | ( n10212 & n11976 ) ;
  assign n14977 = n582 & n14976 ;
  assign n14978 = n14977 ^ n4772 ^ 1'b0 ;
  assign n14979 = ( n2728 & n5464 ) | ( n2728 & ~n7558 ) | ( n5464 & ~n7558 ) ;
  assign n14980 = n11974 ^ n4990 ^ 1'b0 ;
  assign n14981 = n2075 & n14980 ;
  assign n14982 = n9598 & n14981 ;
  assign n14983 = n14979 & n14982 ;
  assign n14984 = ~n5762 & n8406 ;
  assign n14985 = n4942 & n14984 ;
  assign n14992 = n14508 ^ n3696 ^ n754 ;
  assign n14991 = n3717 & ~n4256 ;
  assign n14986 = ( n2106 & ~n5188 ) | ( n2106 & n7920 ) | ( ~n5188 & n7920 ) ;
  assign n14987 = n12578 ^ n3656 ^ 1'b0 ;
  assign n14988 = n14986 & n14987 ;
  assign n14989 = n1091 & ~n6442 ;
  assign n14990 = ~n14988 & n14989 ;
  assign n14993 = n14992 ^ n14991 ^ n14990 ;
  assign n14994 = ( n10506 & n12442 ) | ( n10506 & ~n14993 ) | ( n12442 & ~n14993 ) ;
  assign n14995 = ( n3147 & n10389 ) | ( n3147 & n12697 ) | ( n10389 & n12697 ) ;
  assign n14996 = n1896 & n14995 ;
  assign n14997 = n14996 ^ n14477 ^ 1'b0 ;
  assign n14998 = n6692 ^ n4306 ^ x201 ;
  assign n14999 = n14998 ^ n10497 ^ n2022 ;
  assign n15000 = n14999 ^ n4957 ^ x187 ;
  assign n15001 = n11291 ^ n4445 ^ 1'b0 ;
  assign n15002 = n8282 ^ n3966 ^ 1'b0 ;
  assign n15003 = ( n1356 & ~n5963 ) | ( n1356 & n15002 ) | ( ~n5963 & n15002 ) ;
  assign n15004 = ( n4245 & n5726 ) | ( n4245 & ~n15003 ) | ( n5726 & ~n15003 ) ;
  assign n15005 = ~n14090 & n15004 ;
  assign n15008 = n4337 | n5372 ;
  assign n15009 = n15008 ^ n5765 ^ 1'b0 ;
  assign n15010 = n15009 ^ n5594 ^ n1096 ;
  assign n15006 = n10016 ^ n461 ^ 1'b0 ;
  assign n15007 = n13823 & ~n15006 ;
  assign n15011 = n15010 ^ n15007 ^ n6167 ;
  assign n15012 = ~n4543 & n6644 ;
  assign n15013 = n5912 & n15012 ;
  assign n15014 = ~n2271 & n7047 ;
  assign n15015 = n15013 & n15014 ;
  assign n15016 = n15015 ^ n10665 ^ n5380 ;
  assign n15017 = n8803 ^ n8000 ^ 1'b0 ;
  assign n15018 = ( ~n779 & n15016 ) | ( ~n779 & n15017 ) | ( n15016 & n15017 ) ;
  assign n15019 = n9311 ^ n4944 ^ 1'b0 ;
  assign n15020 = n615 & ~n15019 ;
  assign n15021 = n15020 ^ n7572 ^ 1'b0 ;
  assign n15022 = n11475 | n15021 ;
  assign n15023 = n8946 & n14060 ;
  assign n15024 = x26 | n610 ;
  assign n15025 = ( n5727 & ~n13584 ) | ( n5727 & n15024 ) | ( ~n13584 & n15024 ) ;
  assign n15026 = n14215 ^ n7162 ^ 1'b0 ;
  assign n15027 = n15025 | n15026 ;
  assign n15028 = n15023 | n15027 ;
  assign n15029 = n3621 & n15028 ;
  assign n15030 = n6872 ^ n3808 ^ n1764 ;
  assign n15031 = n12842 ^ n1977 ^ 1'b0 ;
  assign n15032 = n15030 | n15031 ;
  assign n15033 = n4219 ^ n3376 ^ 1'b0 ;
  assign n15034 = n7890 | n15033 ;
  assign n15035 = ( n4239 & n10903 ) | ( n4239 & n15034 ) | ( n10903 & n15034 ) ;
  assign n15036 = ( n6008 & n10477 ) | ( n6008 & n15035 ) | ( n10477 & n15035 ) ;
  assign n15037 = n3524 ^ n2055 ^ n901 ;
  assign n15038 = ( n5065 & n13935 ) | ( n5065 & n15037 ) | ( n13935 & n15037 ) ;
  assign n15039 = ( ~n15032 & n15036 ) | ( ~n15032 & n15038 ) | ( n15036 & n15038 ) ;
  assign n15040 = ~n12969 & n15039 ;
  assign n15041 = n14244 ^ n6639 ^ n5703 ;
  assign n15042 = ( n1382 & n4436 ) | ( n1382 & n6985 ) | ( n4436 & n6985 ) ;
  assign n15043 = n15042 ^ n7965 ^ n6184 ;
  assign n15044 = ~n11532 & n15043 ;
  assign n15045 = n15044 ^ n6764 ^ 1'b0 ;
  assign n15046 = ~n15041 & n15045 ;
  assign n15047 = n14078 ^ n11640 ^ n3649 ;
  assign n15048 = ~n2289 & n5857 ;
  assign n15049 = n15048 ^ n988 ^ 1'b0 ;
  assign n15050 = n287 | n15049 ;
  assign n15051 = ( n3965 & ~n11209 ) | ( n3965 & n15050 ) | ( ~n11209 & n15050 ) ;
  assign n15052 = n7760 & n15051 ;
  assign n15053 = x50 & ~n465 ;
  assign n15054 = ~n2315 & n15053 ;
  assign n15056 = n6598 ^ n3259 ^ x57 ;
  assign n15055 = n728 & ~n3356 ;
  assign n15057 = n15056 ^ n15055 ^ 1'b0 ;
  assign n15058 = ~n15054 & n15057 ;
  assign n15059 = ( n6828 & n8133 ) | ( n6828 & ~n12656 ) | ( n8133 & ~n12656 ) ;
  assign n15060 = n15059 ^ n4272 ^ n3684 ;
  assign n15061 = ( n2213 & ~n4383 ) | ( n2213 & n7818 ) | ( ~n4383 & n7818 ) ;
  assign n15062 = ( n4326 & n5981 ) | ( n4326 & ~n15061 ) | ( n5981 & ~n15061 ) ;
  assign n15063 = ( n598 & n987 ) | ( n598 & n15062 ) | ( n987 & n15062 ) ;
  assign n15064 = n15063 ^ n12254 ^ 1'b0 ;
  assign n15065 = n14280 ^ n8126 ^ x181 ;
  assign n15066 = n15065 ^ n4910 ^ n4748 ;
  assign n15067 = n11810 ^ n6796 ^ 1'b0 ;
  assign n15068 = ~n2826 & n15067 ;
  assign n15069 = n15068 ^ n3791 ^ 1'b0 ;
  assign n15070 = n1970 ^ n396 ^ 1'b0 ;
  assign n15071 = n6901 | n15070 ;
  assign n15072 = n14297 & ~n15071 ;
  assign n15073 = n15069 | n15072 ;
  assign n15074 = n6162 ^ n5162 ^ n2012 ;
  assign n15075 = n3881 & ~n15074 ;
  assign n15076 = ( n10791 & n13813 ) | ( n10791 & ~n15075 ) | ( n13813 & ~n15075 ) ;
  assign n15077 = n12243 ^ n7339 ^ 1'b0 ;
  assign n15078 = ~n6286 & n15077 ;
  assign n15079 = n15078 ^ n5673 ^ n4787 ;
  assign n15080 = n13043 ^ n8048 ^ n5883 ;
  assign n15081 = ~n7774 & n15080 ;
  assign n15082 = n1623 & ~n11210 ;
  assign n15083 = n15082 ^ n3181 ^ 1'b0 ;
  assign n15084 = n3155 & n11083 ;
  assign n15085 = n14519 & ~n15084 ;
  assign n15086 = ( n561 & n1740 ) | ( n561 & n4894 ) | ( n1740 & n4894 ) ;
  assign n15087 = n15086 ^ n11485 ^ n2818 ;
  assign n15088 = ( n2146 & ~n6755 ) | ( n2146 & n8856 ) | ( ~n6755 & n8856 ) ;
  assign n15089 = ( n1181 & n1945 ) | ( n1181 & ~n6987 ) | ( n1945 & ~n6987 ) ;
  assign n15090 = n15089 ^ n4074 ^ n858 ;
  assign n15091 = ( n2329 & ~n12858 ) | ( n2329 & n15090 ) | ( ~n12858 & n15090 ) ;
  assign n15092 = n9669 ^ n6337 ^ n4776 ;
  assign n15093 = ( n4400 & n6191 ) | ( n4400 & ~n15092 ) | ( n6191 & ~n15092 ) ;
  assign n15094 = n15093 ^ n11516 ^ n9769 ;
  assign n15095 = n1759 & ~n10082 ;
  assign n15096 = n15095 ^ n854 ^ 1'b0 ;
  assign n15097 = n15096 ^ n6018 ^ 1'b0 ;
  assign n15098 = n4226 & n15097 ;
  assign n15099 = n7213 & n15098 ;
  assign n15100 = n15099 ^ n11012 ^ 1'b0 ;
  assign n15101 = n3446 & n10404 ;
  assign n15102 = n15101 ^ n3219 ^ 1'b0 ;
  assign n15103 = n14267 ^ n7273 ^ 1'b0 ;
  assign n15104 = n1068 & n15103 ;
  assign n15105 = n9222 & n15104 ;
  assign n15106 = n15102 & n15105 ;
  assign n15109 = ( n4794 & n8820 ) | ( n4794 & n11048 ) | ( n8820 & n11048 ) ;
  assign n15110 = n15109 ^ n12947 ^ n3377 ;
  assign n15111 = n5524 & ~n15110 ;
  assign n15112 = n10287 & n15111 ;
  assign n15119 = n13412 ^ n2729 ^ n986 ;
  assign n15120 = ( n9890 & ~n10840 ) | ( n9890 & n15119 ) | ( ~n10840 & n15119 ) ;
  assign n15113 = x99 | n684 ;
  assign n15114 = ( x175 & n2244 ) | ( x175 & n15113 ) | ( n2244 & n15113 ) ;
  assign n15115 = n15114 ^ n6618 ^ n470 ;
  assign n15116 = n15115 ^ n3943 ^ n3936 ;
  assign n15117 = n15116 ^ n6507 ^ 1'b0 ;
  assign n15118 = n8024 | n15117 ;
  assign n15121 = n15120 ^ n15118 ^ n1258 ;
  assign n15122 = ~n15112 & n15121 ;
  assign n15123 = n796 & n15122 ;
  assign n15124 = n963 & n8047 ;
  assign n15125 = n15123 | n15124 ;
  assign n15107 = ~n415 & n1365 ;
  assign n15108 = n8375 & n15107 ;
  assign n15126 = n15125 ^ n15108 ^ 1'b0 ;
  assign n15127 = n14358 | n15126 ;
  assign n15129 = ( ~n5385 & n7402 ) | ( ~n5385 & n11045 ) | ( n7402 & n11045 ) ;
  assign n15128 = ( n1693 & n5503 ) | ( n1693 & n7562 ) | ( n5503 & n7562 ) ;
  assign n15130 = n15129 ^ n15128 ^ 1'b0 ;
  assign n15136 = n10241 ^ n4215 ^ 1'b0 ;
  assign n15131 = n7268 ^ n2729 ^ 1'b0 ;
  assign n15132 = ~n8428 & n15131 ;
  assign n15133 = n15132 ^ n6087 ^ n2981 ;
  assign n15134 = ( n6617 & n13589 ) | ( n6617 & n15133 ) | ( n13589 & n15133 ) ;
  assign n15135 = ~n1390 & n15134 ;
  assign n15137 = n15136 ^ n15135 ^ 1'b0 ;
  assign n15138 = n14560 ^ n13244 ^ 1'b0 ;
  assign n15139 = n9255 ^ n2685 ^ 1'b0 ;
  assign n15141 = n6131 ^ n5658 ^ n3732 ;
  assign n15140 = ( ~n749 & n6585 ) | ( ~n749 & n12182 ) | ( n6585 & n12182 ) ;
  assign n15142 = n15141 ^ n15140 ^ n14277 ;
  assign n15146 = n13405 ^ n7025 ^ n2764 ;
  assign n15145 = n12050 ^ n3270 ^ n597 ;
  assign n15147 = n15146 ^ n15145 ^ n2903 ;
  assign n15144 = n6828 ^ n4804 ^ n348 ;
  assign n15143 = ( ~n1372 & n1406 ) | ( ~n1372 & n9969 ) | ( n1406 & n9969 ) ;
  assign n15148 = n15147 ^ n15144 ^ n15143 ;
  assign n15149 = ( n5261 & n12151 ) | ( n5261 & n14460 ) | ( n12151 & n14460 ) ;
  assign n15150 = n9216 | n15149 ;
  assign n15151 = n15150 ^ n7373 ^ 1'b0 ;
  assign n15152 = n15148 | n15151 ;
  assign n15153 = ( n950 & n3209 ) | ( n950 & n11843 ) | ( n3209 & n11843 ) ;
  assign n15154 = ( n667 & n4642 ) | ( n667 & n15153 ) | ( n4642 & n15153 ) ;
  assign n15155 = n5174 ^ n1761 ^ n488 ;
  assign n15156 = n2141 & n7432 ;
  assign n15157 = n4583 & n15156 ;
  assign n15158 = n15157 ^ n13493 ^ n4300 ;
  assign n15159 = ( n882 & ~n967 ) | ( n882 & n15158 ) | ( ~n967 & n15158 ) ;
  assign n15160 = ( n12080 & n15155 ) | ( n12080 & n15159 ) | ( n15155 & n15159 ) ;
  assign n15161 = n2774 ^ n1096 ^ x201 ;
  assign n15162 = n15161 ^ n9118 ^ n2960 ;
  assign n15163 = n15162 ^ n7515 ^ n427 ;
  assign n15165 = n12479 ^ n4529 ^ 1'b0 ;
  assign n15166 = n1125 | n15165 ;
  assign n15164 = n4005 ^ n3536 ^ n3312 ;
  assign n15167 = n15166 ^ n15164 ^ 1'b0 ;
  assign n15168 = n15167 ^ n14722 ^ n10492 ;
  assign n15169 = n6605 ^ n5830 ^ n4279 ;
  assign n15170 = n15169 ^ n9328 ^ n4735 ;
  assign n15171 = n11778 ^ n7137 ^ 1'b0 ;
  assign n15172 = n15171 ^ n13801 ^ n7340 ;
  assign n15173 = n10985 ^ n6037 ^ n3711 ;
  assign n15174 = n11802 ^ n4327 ^ 1'b0 ;
  assign n15175 = ( n639 & n5918 ) | ( n639 & ~n15174 ) | ( n5918 & ~n15174 ) ;
  assign n15176 = ( n507 & n15173 ) | ( n507 & ~n15175 ) | ( n15173 & ~n15175 ) ;
  assign n15177 = n10684 ^ n4664 ^ n2471 ;
  assign n15178 = ( n4881 & n5861 ) | ( n4881 & n15177 ) | ( n5861 & n15177 ) ;
  assign n15179 = n15178 ^ n8571 ^ n5082 ;
  assign n15180 = ( ~n4526 & n4560 ) | ( ~n4526 & n8754 ) | ( n4560 & n8754 ) ;
  assign n15181 = n10162 ^ n5629 ^ n5238 ;
  assign n15182 = n15181 ^ n14543 ^ 1'b0 ;
  assign n15183 = ( n10783 & ~n12815 ) | ( n10783 & n15182 ) | ( ~n12815 & n15182 ) ;
  assign n15184 = n6640 ^ x71 ^ 1'b0 ;
  assign n15185 = n8062 ^ n4180 ^ 1'b0 ;
  assign n15186 = ~n1106 & n15185 ;
  assign n15187 = n15186 ^ n7337 ^ n1212 ;
  assign n15188 = ( n9864 & n10348 ) | ( n9864 & n15187 ) | ( n10348 & n15187 ) ;
  assign n15191 = n470 ^ x0 ^ 1'b0 ;
  assign n15192 = ( n4798 & n9022 ) | ( n4798 & n15191 ) | ( n9022 & n15191 ) ;
  assign n15193 = ( n7218 & ~n13258 ) | ( n7218 & n15192 ) | ( ~n13258 & n15192 ) ;
  assign n15189 = ~n715 & n3014 ;
  assign n15190 = n10030 & ~n15189 ;
  assign n15194 = n15193 ^ n15190 ^ 1'b0 ;
  assign n15195 = n5685 ^ n453 ^ x21 ;
  assign n15196 = ( ~n4889 & n11934 ) | ( ~n4889 & n15195 ) | ( n11934 & n15195 ) ;
  assign n15197 = ( n8570 & n11155 ) | ( n8570 & n15196 ) | ( n11155 & n15196 ) ;
  assign n15198 = n1788 & ~n3130 ;
  assign n15199 = n15198 ^ n5146 ^ 1'b0 ;
  assign n15200 = n3173 & n8752 ;
  assign n15201 = n15199 & n15200 ;
  assign n15202 = n542 & n1673 ;
  assign n15203 = ~n12213 & n15202 ;
  assign n15204 = n3483 | n15203 ;
  assign n15205 = n15204 ^ n7263 ^ 1'b0 ;
  assign n15206 = n9625 ^ n2521 ^ 1'b0 ;
  assign n15207 = n5778 & ~n7500 ;
  assign n15208 = n15207 ^ n3989 ^ n334 ;
  assign n15209 = n2491 ^ n800 ^ 1'b0 ;
  assign n15210 = n15208 | n15209 ;
  assign n15212 = ~n1109 & n2638 ;
  assign n15213 = ( n6917 & n7977 ) | ( n6917 & n15212 ) | ( n7977 & n15212 ) ;
  assign n15211 = n8419 & n10019 ;
  assign n15214 = n15213 ^ n15211 ^ 1'b0 ;
  assign n15215 = n15214 ^ n8446 ^ n1641 ;
  assign n15216 = n508 & ~n3244 ;
  assign n15217 = ~n8480 & n15216 ;
  assign n15218 = n15217 ^ n7425 ^ n7420 ;
  assign n15219 = n15218 ^ n4626 ^ 1'b0 ;
  assign n15220 = n11101 & n15219 ;
  assign n15221 = ( n9671 & ~n14232 ) | ( n9671 & n14896 ) | ( ~n14232 & n14896 ) ;
  assign n15222 = n659 & n779 ;
  assign n15223 = n15222 ^ n6898 ^ 1'b0 ;
  assign n15224 = n15221 & ~n15223 ;
  assign n15225 = ( ~n5994 & n9105 ) | ( ~n5994 & n15224 ) | ( n9105 & n15224 ) ;
  assign n15226 = n2068 ^ n1561 ^ 1'b0 ;
  assign n15227 = ~n3620 & n15226 ;
  assign n15228 = ( n4029 & n11802 ) | ( n4029 & n15227 ) | ( n11802 & n15227 ) ;
  assign n15229 = n6632 ^ n1953 ^ n959 ;
  assign n15230 = n15228 & n15229 ;
  assign n15231 = n15225 & n15230 ;
  assign n15232 = ( ~n9571 & n10625 ) | ( ~n9571 & n15231 ) | ( n10625 & n15231 ) ;
  assign n15233 = ( ~n12257 & n15167 ) | ( ~n12257 & n15232 ) | ( n15167 & n15232 ) ;
  assign n15234 = n15233 ^ n12708 ^ n282 ;
  assign n15235 = n13394 ^ n11342 ^ 1'b0 ;
  assign n15236 = n5617 ^ n4501 ^ n4023 ;
  assign n15237 = n8019 | n13243 ;
  assign n15238 = n15236 | n15237 ;
  assign n15239 = n15238 ^ n2203 ^ 1'b0 ;
  assign n15240 = n2345 & n15239 ;
  assign n15241 = n5562 ^ n1787 ^ x21 ;
  assign n15242 = n15240 & n15241 ;
  assign n15243 = ( n7776 & ~n12728 ) | ( n7776 & n13459 ) | ( ~n12728 & n13459 ) ;
  assign n15244 = ~n7448 & n14376 ;
  assign n15245 = n15244 ^ n2306 ^ 1'b0 ;
  assign n15246 = ( n3980 & ~n14898 ) | ( n3980 & n15245 ) | ( ~n14898 & n15245 ) ;
  assign n15247 = n12950 ^ n9105 ^ n7066 ;
  assign n15248 = n13371 ^ x77 ^ 1'b0 ;
  assign n15249 = ( n7563 & n15247 ) | ( n7563 & ~n15248 ) | ( n15247 & ~n15248 ) ;
  assign n15250 = n4388 & n15249 ;
  assign n15251 = n12168 ^ n7313 ^ n4722 ;
  assign n15252 = n15251 ^ n5588 ^ 1'b0 ;
  assign n15253 = n15252 ^ n14863 ^ 1'b0 ;
  assign n15254 = n2428 & n13265 ;
  assign n15255 = n1791 & n6939 ;
  assign n15256 = ( n14321 & n15254 ) | ( n14321 & n15255 ) | ( n15254 & n15255 ) ;
  assign n15257 = ( n1877 & n13342 ) | ( n1877 & n15256 ) | ( n13342 & n15256 ) ;
  assign n15258 = n14711 ^ n7682 ^ 1'b0 ;
  assign n15259 = ~n2051 & n15258 ;
  assign n15261 = ( x146 & n2084 ) | ( x146 & ~n9778 ) | ( n2084 & ~n9778 ) ;
  assign n15262 = n348 & n14270 ;
  assign n15263 = ~n5165 & n15262 ;
  assign n15264 = n15263 ^ n13777 ^ n3950 ;
  assign n15268 = n2762 & n9288 ;
  assign n15265 = ( n1957 & n5732 ) | ( n1957 & ~n6362 ) | ( n5732 & ~n6362 ) ;
  assign n15266 = n15265 ^ n8002 ^ n1394 ;
  assign n15267 = n7500 & n15266 ;
  assign n15269 = n15268 ^ n15267 ^ 1'b0 ;
  assign n15270 = n15269 ^ n1230 ^ 1'b0 ;
  assign n15271 = ( n15261 & n15264 ) | ( n15261 & n15270 ) | ( n15264 & n15270 ) ;
  assign n15260 = n13688 & n14135 ;
  assign n15272 = n15271 ^ n15260 ^ 1'b0 ;
  assign n15273 = n13631 ^ n476 ^ 1'b0 ;
  assign n15274 = ( n286 & ~n8016 ) | ( n286 & n11373 ) | ( ~n8016 & n11373 ) ;
  assign n15275 = n11871 ^ n3731 ^ n2341 ;
  assign n15276 = ( n4721 & n15274 ) | ( n4721 & ~n15275 ) | ( n15274 & ~n15275 ) ;
  assign n15277 = n15273 & ~n15276 ;
  assign n15282 = n2489 | n2612 ;
  assign n15283 = n15282 ^ n4581 ^ 1'b0 ;
  assign n15284 = n15283 ^ n8710 ^ 1'b0 ;
  assign n15278 = n885 & ~n1136 ;
  assign n15279 = n491 & ~n15278 ;
  assign n15280 = n8145 & n15279 ;
  assign n15281 = ( n7222 & ~n10497 ) | ( n7222 & n15280 ) | ( ~n10497 & n15280 ) ;
  assign n15285 = n15284 ^ n15281 ^ n2070 ;
  assign n15286 = n6515 ^ n3691 ^ 1'b0 ;
  assign n15287 = n6453 | n15286 ;
  assign n15288 = n5798 & ~n15287 ;
  assign n15289 = ( n3845 & ~n11182 ) | ( n3845 & n15288 ) | ( ~n11182 & n15288 ) ;
  assign n15290 = ~n2626 & n15252 ;
  assign n15300 = n8068 ^ n1769 ^ x246 ;
  assign n15299 = n3943 ^ n2575 ^ 1'b0 ;
  assign n15298 = n14589 ^ n13380 ^ n5737 ;
  assign n15301 = n15300 ^ n15299 ^ n15298 ;
  assign n15302 = n15301 ^ n4419 ^ n1711 ;
  assign n15291 = n5612 ^ n1457 ^ n819 ;
  assign n15292 = ~n3217 & n15291 ;
  assign n15293 = n3514 & n15292 ;
  assign n15294 = n15293 ^ n2001 ^ 1'b0 ;
  assign n15295 = n10031 ^ n5181 ^ 1'b0 ;
  assign n15296 = n8774 | n15295 ;
  assign n15297 = ( ~n5501 & n15294 ) | ( ~n5501 & n15296 ) | ( n15294 & n15296 ) ;
  assign n15303 = n15302 ^ n15297 ^ n6500 ;
  assign n15304 = n1514 & n15303 ;
  assign n15305 = ~n15290 & n15304 ;
  assign n15306 = n13776 ^ n8684 ^ 1'b0 ;
  assign n15307 = n6491 | n9251 ;
  assign n15308 = n1307 | n15307 ;
  assign n15310 = n14473 ^ n12634 ^ n4824 ;
  assign n15311 = n5449 ^ n1327 ^ n917 ;
  assign n15312 = ~n15310 & n15311 ;
  assign n15313 = ~n2104 & n15312 ;
  assign n15309 = n7464 ^ n3757 ^ n2785 ;
  assign n15314 = n15313 ^ n15309 ^ n8160 ;
  assign n15315 = n2870 & ~n4256 ;
  assign n15316 = ( n5450 & ~n6281 ) | ( n5450 & n15315 ) | ( ~n6281 & n15315 ) ;
  assign n15317 = ( ~n748 & n7164 ) | ( ~n748 & n9593 ) | ( n7164 & n9593 ) ;
  assign n15318 = ( n2619 & ~n5526 ) | ( n2619 & n5607 ) | ( ~n5526 & n5607 ) ;
  assign n15319 = ~n1725 & n15318 ;
  assign n15320 = n15319 ^ n3393 ^ 1'b0 ;
  assign n15321 = n846 | n15320 ;
  assign n15322 = n15321 ^ n6424 ^ n3973 ;
  assign n15323 = ~n15317 & n15322 ;
  assign n15324 = n15323 ^ n5262 ^ 1'b0 ;
  assign n15325 = n2630 ^ x88 ^ 1'b0 ;
  assign n15326 = n15324 & n15325 ;
  assign n15327 = n15326 ^ n6668 ^ n4279 ;
  assign n15328 = n15316 & n15327 ;
  assign n15329 = n7498 ^ n7147 ^ n5286 ;
  assign n15330 = n15329 ^ n4972 ^ n2779 ;
  assign n15331 = ( n6414 & ~n8067 ) | ( n6414 & n9993 ) | ( ~n8067 & n9993 ) ;
  assign n15332 = n7103 ^ n5500 ^ n4100 ;
  assign n15333 = ( n7850 & ~n13818 ) | ( n7850 & n15332 ) | ( ~n13818 & n15332 ) ;
  assign n15334 = n15318 ^ n2825 ^ 1'b0 ;
  assign n15335 = ( n10007 & n15333 ) | ( n10007 & n15334 ) | ( n15333 & n15334 ) ;
  assign n15336 = n15335 ^ n15193 ^ 1'b0 ;
  assign n15337 = n5216 | n15336 ;
  assign n15338 = n15337 ^ n13399 ^ n2797 ;
  assign n15339 = ( ~n8976 & n15331 ) | ( ~n8976 & n15338 ) | ( n15331 & n15338 ) ;
  assign n15340 = n1797 & n6454 ;
  assign n15341 = n3806 & n15340 ;
  assign n15344 = n9626 ^ n4479 ^ 1'b0 ;
  assign n15345 = n9334 & ~n15344 ;
  assign n15342 = n2422 | n6363 ;
  assign n15343 = n11762 & ~n15342 ;
  assign n15346 = n15345 ^ n15343 ^ 1'b0 ;
  assign n15347 = n11567 ^ n10007 ^ 1'b0 ;
  assign n15348 = n4294 & n5948 ;
  assign n15349 = n10759 | n15348 ;
  assign n15350 = n15347 | n15349 ;
  assign n15351 = n8581 & n10086 ;
  assign n15352 = n13929 ^ n11183 ^ n1871 ;
  assign n15353 = n15352 ^ n2997 ^ 1'b0 ;
  assign n15354 = n15351 | n15353 ;
  assign n15355 = n9656 & ~n15354 ;
  assign n15356 = n15355 ^ n6544 ^ 1'b0 ;
  assign n15357 = ~n1440 & n2948 ;
  assign n15358 = ~n4248 & n15357 ;
  assign n15359 = n8641 ^ n2866 ^ 1'b0 ;
  assign n15360 = x51 & n717 ;
  assign n15361 = ~n15359 & n15360 ;
  assign n15362 = ( n2538 & n15358 ) | ( n2538 & ~n15361 ) | ( n15358 & ~n15361 ) ;
  assign n15363 = n15362 ^ n11856 ^ n8479 ;
  assign n15364 = n6985 | n10296 ;
  assign n15365 = n15364 ^ n5554 ^ n2556 ;
  assign n15366 = ~n11392 & n15365 ;
  assign n15367 = n15363 & n15366 ;
  assign n15368 = ( n529 & n2599 ) | ( n529 & n7779 ) | ( n2599 & n7779 ) ;
  assign n15369 = n13109 ^ n4579 ^ 1'b0 ;
  assign n15370 = n396 & ~n15369 ;
  assign n15371 = ( ~n8705 & n15368 ) | ( ~n8705 & n15370 ) | ( n15368 & n15370 ) ;
  assign n15372 = ~n4628 & n15371 ;
  assign n15373 = n15372 ^ n12268 ^ n10587 ;
  assign n15381 = n13681 ^ n13483 ^ n1363 ;
  assign n15377 = ( ~n3356 & n7651 ) | ( ~n3356 & n15352 ) | ( n7651 & n15352 ) ;
  assign n15378 = ( ~n829 & n6137 ) | ( ~n829 & n15377 ) | ( n6137 & n15377 ) ;
  assign n15379 = n15378 ^ n7653 ^ n4397 ;
  assign n15374 = n4042 | n10152 ;
  assign n15375 = n15374 ^ n5291 ^ 1'b0 ;
  assign n15376 = n10561 & n15375 ;
  assign n15380 = n15379 ^ n15376 ^ n1283 ;
  assign n15382 = n15381 ^ n15380 ^ n10740 ;
  assign n15383 = n4474 ^ n1044 ^ 1'b0 ;
  assign n15384 = n10321 ^ n4232 ^ 1'b0 ;
  assign n15385 = n15384 ^ n582 ^ 1'b0 ;
  assign n15386 = ~n15383 & n15385 ;
  assign n15387 = ~n668 & n2430 ;
  assign n15388 = n15387 ^ n5145 ^ n2128 ;
  assign n15389 = n14232 & ~n15388 ;
  assign n15390 = ( n2389 & n2676 ) | ( n2389 & ~n15389 ) | ( n2676 & ~n15389 ) ;
  assign n15391 = n15390 ^ n13715 ^ n12451 ;
  assign n15392 = n11216 ^ n5592 ^ n749 ;
  assign n15393 = n15392 ^ n4701 ^ n3429 ;
  assign n15394 = n6505 ^ n2867 ^ 1'b0 ;
  assign n15395 = n404 & ~n15394 ;
  assign n15396 = ( n6965 & ~n7903 ) | ( n6965 & n15395 ) | ( ~n7903 & n15395 ) ;
  assign n15397 = ( n6009 & n15393 ) | ( n6009 & n15396 ) | ( n15393 & n15396 ) ;
  assign n15398 = ( n1739 & n7613 ) | ( n1739 & ~n15397 ) | ( n7613 & ~n15397 ) ;
  assign n15399 = n3369 | n9902 ;
  assign n15400 = n15398 | n15399 ;
  assign n15401 = ( ~n5766 & n10913 ) | ( ~n5766 & n14761 ) | ( n10913 & n14761 ) ;
  assign n15402 = n11696 ^ n1762 ^ n1717 ;
  assign n15403 = n15402 ^ n3614 ^ 1'b0 ;
  assign n15404 = n4722 ^ n4260 ^ 1'b0 ;
  assign n15405 = n2659 & ~n15404 ;
  assign n15406 = n15405 ^ n12899 ^ 1'b0 ;
  assign n15407 = n15406 ^ n3481 ^ x141 ;
  assign n15408 = n15407 ^ n9586 ^ n4583 ;
  assign n15409 = n5896 & ~n15408 ;
  assign n15410 = n11147 ^ n1245 ^ 1'b0 ;
  assign n15411 = n15115 & ~n15410 ;
  assign n15412 = ( n1230 & ~n4553 ) | ( n1230 & n9774 ) | ( ~n4553 & n9774 ) ;
  assign n15413 = ~n3448 & n8978 ;
  assign n15414 = ~n4746 & n15413 ;
  assign n15415 = ( ~n261 & n15412 ) | ( ~n261 & n15414 ) | ( n15412 & n15414 ) ;
  assign n15416 = ( ~n8710 & n15411 ) | ( ~n8710 & n15415 ) | ( n15411 & n15415 ) ;
  assign n15417 = ( n2930 & n9778 ) | ( n2930 & n15416 ) | ( n9778 & n15416 ) ;
  assign n15420 = n9744 ^ n3083 ^ 1'b0 ;
  assign n15421 = n2971 | n15420 ;
  assign n15422 = ( n2739 & ~n4533 ) | ( n2739 & n15421 ) | ( ~n4533 & n15421 ) ;
  assign n15418 = n14779 ^ n5411 ^ 1'b0 ;
  assign n15419 = n10186 | n15418 ;
  assign n15423 = n15422 ^ n15419 ^ n8319 ;
  assign n15424 = n7063 ^ n6865 ^ 1'b0 ;
  assign n15425 = n306 & ~n1016 ;
  assign n15426 = n15424 & n15425 ;
  assign n15427 = n15426 ^ n14109 ^ 1'b0 ;
  assign n15430 = n6051 ^ n5815 ^ n5088 ;
  assign n15428 = n10199 ^ n6186 ^ 1'b0 ;
  assign n15429 = n10101 & ~n15428 ;
  assign n15431 = n15430 ^ n15429 ^ n1527 ;
  assign n15432 = n15431 ^ n7415 ^ n4519 ;
  assign n15433 = n1144 | n4853 ;
  assign n15434 = n4908 & ~n15433 ;
  assign n15435 = ( n4808 & n5662 ) | ( n4808 & n15434 ) | ( n5662 & n15434 ) ;
  assign n15436 = n3044 ^ n1594 ^ x144 ;
  assign n15437 = n15436 ^ n3948 ^ n1842 ;
  assign n15438 = ( n7589 & ~n11768 ) | ( n7589 & n15437 ) | ( ~n11768 & n15437 ) ;
  assign n15439 = n5858 | n15438 ;
  assign n15440 = ( n12527 & ~n15435 ) | ( n12527 & n15439 ) | ( ~n15435 & n15439 ) ;
  assign n15441 = n10694 ^ n2784 ^ 1'b0 ;
  assign n15442 = ( ~n3614 & n5134 ) | ( ~n3614 & n15441 ) | ( n5134 & n15441 ) ;
  assign n15443 = n15442 ^ n5724 ^ n1323 ;
  assign n15444 = ( n507 & ~n4611 ) | ( n507 & n10115 ) | ( ~n4611 & n10115 ) ;
  assign n15445 = n15444 ^ n2847 ^ 1'b0 ;
  assign n15446 = ~n5675 & n15445 ;
  assign n15447 = n15446 ^ n8085 ^ 1'b0 ;
  assign n15448 = n10890 ^ n2471 ^ 1'b0 ;
  assign n15449 = n10885 ^ n2481 ^ n1827 ;
  assign n15450 = n15449 ^ n15067 ^ 1'b0 ;
  assign n15451 = ( n6694 & n15448 ) | ( n6694 & ~n15450 ) | ( n15448 & ~n15450 ) ;
  assign n15452 = n754 & ~n9586 ;
  assign n15453 = n15452 ^ n15016 ^ n1668 ;
  assign n15454 = ( n2866 & n6309 ) | ( n2866 & ~n6732 ) | ( n6309 & ~n6732 ) ;
  assign n15460 = n647 & ~n1754 ;
  assign n15461 = n2882 & n15460 ;
  assign n15462 = n15461 ^ n6269 ^ 1'b0 ;
  assign n15455 = n5638 & ~n12281 ;
  assign n15456 = ( x25 & ~n1018 ) | ( x25 & n3268 ) | ( ~n1018 & n3268 ) ;
  assign n15457 = n15456 ^ n10346 ^ n1868 ;
  assign n15458 = ( n598 & n5812 ) | ( n598 & ~n15457 ) | ( n5812 & ~n15457 ) ;
  assign n15459 = ~n15455 & n15458 ;
  assign n15463 = n15462 ^ n15459 ^ n7326 ;
  assign n15464 = n5675 & n14406 ;
  assign n15465 = ~n2256 & n13516 ;
  assign n15466 = n15464 & n15465 ;
  assign n15467 = n15466 ^ n14963 ^ 1'b0 ;
  assign n15468 = n13922 & n15467 ;
  assign n15469 = n7965 ^ n2445 ^ n871 ;
  assign n15470 = n15469 ^ n4994 ^ n3963 ;
  assign n15471 = ( ~n2227 & n3198 ) | ( ~n2227 & n11779 ) | ( n3198 & n11779 ) ;
  assign n15472 = n1451 ^ n713 ^ 1'b0 ;
  assign n15473 = n2712 & ~n15472 ;
  assign n15474 = n15473 ^ n4784 ^ 1'b0 ;
  assign n15475 = n9439 & ~n15474 ;
  assign n15476 = ( ~n6511 & n15471 ) | ( ~n6511 & n15475 ) | ( n15471 & n15475 ) ;
  assign n15477 = ( n1127 & ~n15470 ) | ( n1127 & n15476 ) | ( ~n15470 & n15476 ) ;
  assign n15478 = ( n2126 & ~n2885 ) | ( n2126 & n14713 ) | ( ~n2885 & n14713 ) ;
  assign n15479 = n2226 & n15478 ;
  assign n15480 = n13921 ^ n6855 ^ n5213 ;
  assign n15481 = ~n9729 & n10963 ;
  assign n15482 = n15481 ^ n14857 ^ n2733 ;
  assign n15483 = n5725 ^ n678 ^ 1'b0 ;
  assign n15484 = n15483 ^ n13084 ^ n3115 ;
  assign n15485 = ( n9538 & ~n9596 ) | ( n9538 & n12015 ) | ( ~n9596 & n12015 ) ;
  assign n15486 = n15485 ^ n5407 ^ n3244 ;
  assign n15487 = ( n2450 & n9769 ) | ( n2450 & n15486 ) | ( n9769 & n15486 ) ;
  assign n15488 = n5351 & n7947 ;
  assign n15489 = n5917 & n15488 ;
  assign n15490 = ( n9216 & n12790 ) | ( n9216 & ~n15489 ) | ( n12790 & ~n15489 ) ;
  assign n15491 = n326 & n1866 ;
  assign n15492 = ( n1312 & n10041 ) | ( n1312 & n15491 ) | ( n10041 & n15491 ) ;
  assign n15495 = ~n9131 & n15321 ;
  assign n15496 = n8184 & n15495 ;
  assign n15493 = n11426 ^ n1439 ^ 1'b0 ;
  assign n15494 = n15493 ^ n12249 ^ n3555 ;
  assign n15497 = n15496 ^ n15494 ^ n1271 ;
  assign n15498 = ( n1688 & n1743 ) | ( n1688 & n5576 ) | ( n1743 & n5576 ) ;
  assign n15499 = ( n5132 & n7888 ) | ( n5132 & n15498 ) | ( n7888 & n15498 ) ;
  assign n15500 = ~n2605 & n15499 ;
  assign n15501 = n15397 & n15500 ;
  assign n15502 = n2905 ^ n2430 ^ 1'b0 ;
  assign n15503 = n15502 ^ n4414 ^ 1'b0 ;
  assign n15504 = n14296 ^ n7520 ^ 1'b0 ;
  assign n15505 = n12035 | n15504 ;
  assign n15506 = n15505 ^ n14515 ^ 1'b0 ;
  assign n15507 = n15506 ^ n13699 ^ 1'b0 ;
  assign n15508 = n15507 ^ n387 ^ 1'b0 ;
  assign n15509 = n7985 | n15508 ;
  assign n15510 = ( ~n5976 & n15503 ) | ( ~n5976 & n15509 ) | ( n15503 & n15509 ) ;
  assign n15511 = ( n8898 & n10654 ) | ( n8898 & ~n15510 ) | ( n10654 & ~n15510 ) ;
  assign n15512 = ( n10840 & ~n13766 ) | ( n10840 & n14366 ) | ( ~n13766 & n14366 ) ;
  assign n15518 = n1753 & n4080 ;
  assign n15516 = n4697 ^ n2187 ^ 1'b0 ;
  assign n15514 = ~n3369 & n6728 ;
  assign n15515 = n15514 ^ n632 ^ 1'b0 ;
  assign n15517 = n15516 ^ n15515 ^ n1260 ;
  assign n15513 = ~n323 & n1826 ;
  assign n15519 = n15518 ^ n15517 ^ n15513 ;
  assign n15520 = n15519 ^ n5622 ^ n775 ;
  assign n15521 = n6355 | n7525 ;
  assign n15522 = n3483 ^ n2502 ^ n2042 ;
  assign n15523 = n5447 ^ n2746 ^ 1'b0 ;
  assign n15524 = n8348 | n15523 ;
  assign n15525 = ( n8634 & n15522 ) | ( n8634 & ~n15524 ) | ( n15522 & ~n15524 ) ;
  assign n15526 = n14029 ^ n11300 ^ n3206 ;
  assign n15527 = n7711 ^ n6825 ^ 1'b0 ;
  assign n15528 = ~n15526 & n15527 ;
  assign n15536 = ~n1714 & n14725 ;
  assign n15537 = n15536 ^ n5158 ^ 1'b0 ;
  assign n15535 = ( x140 & n4837 ) | ( x140 & n12072 ) | ( n4837 & n12072 ) ;
  assign n15532 = ~n2737 & n15161 ;
  assign n15533 = n15532 ^ n2950 ^ 1'b0 ;
  assign n15531 = n555 & n7297 ;
  assign n15529 = n8285 ^ n4807 ^ 1'b0 ;
  assign n15530 = n8971 & ~n15529 ;
  assign n15534 = n15533 ^ n15531 ^ n15530 ;
  assign n15538 = n15537 ^ n15535 ^ n15534 ;
  assign n15539 = ( ~n6031 & n6400 ) | ( ~n6031 & n10026 ) | ( n6400 & n10026 ) ;
  assign n15540 = n5461 & n9549 ;
  assign n15541 = n8016 ^ n3319 ^ 1'b0 ;
  assign n15542 = n15541 ^ n10232 ^ n8616 ;
  assign n15543 = n15540 & n15542 ;
  assign n15544 = ( ~n4248 & n6428 ) | ( ~n4248 & n10813 ) | ( n6428 & n10813 ) ;
  assign n15545 = ( n5572 & n15543 ) | ( n5572 & n15544 ) | ( n15543 & n15544 ) ;
  assign n15546 = n482 & n12840 ;
  assign n15547 = n13284 | n13651 ;
  assign n15548 = ( n14078 & n15546 ) | ( n14078 & n15547 ) | ( n15546 & n15547 ) ;
  assign n15549 = n3858 | n5251 ;
  assign n15550 = n381 | n15549 ;
  assign n15551 = ~n1950 & n15550 ;
  assign n15552 = n15551 ^ n4594 ^ 1'b0 ;
  assign n15553 = n15552 ^ n13210 ^ n498 ;
  assign n15554 = ( n4698 & n15548 ) | ( n4698 & n15553 ) | ( n15548 & n15553 ) ;
  assign n15555 = n8906 ^ n8501 ^ n7749 ;
  assign n15557 = n3116 & n3952 ;
  assign n15558 = n15557 ^ n4758 ^ 1'b0 ;
  assign n15559 = n15558 ^ n2868 ^ 1'b0 ;
  assign n15560 = ~n3016 & n15559 ;
  assign n15561 = n15560 ^ n13070 ^ n12008 ;
  assign n15556 = n15384 ^ n7949 ^ n1398 ;
  assign n15562 = n15561 ^ n15556 ^ n13737 ;
  assign n15563 = ( ~n14619 & n15555 ) | ( ~n14619 & n15562 ) | ( n15555 & n15562 ) ;
  assign n15564 = n1785 & n1820 ;
  assign n15565 = ~n11611 & n15564 ;
  assign n15567 = n10982 ^ n4062 ^ n3485 ;
  assign n15566 = ( n3526 & n6077 ) | ( n3526 & n9494 ) | ( n6077 & n9494 ) ;
  assign n15568 = n15567 ^ n15566 ^ n13932 ;
  assign n15569 = n15568 ^ n14581 ^ 1'b0 ;
  assign n15570 = ~n12983 & n15569 ;
  assign n15571 = n12745 ^ n11726 ^ n10424 ;
  assign n15572 = n15571 ^ n6122 ^ 1'b0 ;
  assign n15573 = n9739 ^ n9045 ^ n3416 ;
  assign n15574 = n3744 ^ n2728 ^ x240 ;
  assign n15575 = ( n3010 & n13109 ) | ( n3010 & ~n15574 ) | ( n13109 & ~n15574 ) ;
  assign n15576 = n15575 ^ n6119 ^ 1'b0 ;
  assign n15577 = ~n15573 & n15576 ;
  assign n15578 = n15577 ^ n12614 ^ 1'b0 ;
  assign n15579 = n6520 & n15578 ;
  assign n15580 = ~n431 & n13615 ;
  assign n15581 = n15580 ^ n9940 ^ 1'b0 ;
  assign n15582 = ( n1542 & n2393 ) | ( n1542 & n3920 ) | ( n2393 & n3920 ) ;
  assign n15583 = ~n1022 & n9538 ;
  assign n15584 = n7010 | n15583 ;
  assign n15585 = n2912 & ~n15584 ;
  assign n15586 = n15582 | n15585 ;
  assign n15587 = n15581 & ~n15586 ;
  assign n15589 = n10856 ^ n2964 ^ 1'b0 ;
  assign n15588 = n13586 ^ n8222 ^ n6403 ;
  assign n15590 = n15589 ^ n15588 ^ n323 ;
  assign n15591 = n2173 & n13170 ;
  assign n15593 = n4102 ^ n3078 ^ n1120 ;
  assign n15592 = ( n360 & n4113 ) | ( n360 & n4951 ) | ( n4113 & n4951 ) ;
  assign n15594 = n15593 ^ n15592 ^ n2717 ;
  assign n15595 = n15594 ^ n3540 ^ n348 ;
  assign n15596 = n5515 & n7574 ;
  assign n15597 = n9128 | n15596 ;
  assign n15598 = ( ~n15591 & n15595 ) | ( ~n15591 & n15597 ) | ( n15595 & n15597 ) ;
  assign n15599 = ( n3240 & n3960 ) | ( n3240 & ~n11682 ) | ( n3960 & ~n11682 ) ;
  assign n15600 = ( n6195 & n9686 ) | ( n6195 & n15599 ) | ( n9686 & n15599 ) ;
  assign n15601 = ( n6026 & ~n11137 ) | ( n6026 & n15600 ) | ( ~n11137 & n15600 ) ;
  assign n15602 = ( n10741 & n14094 ) | ( n10741 & n15601 ) | ( n14094 & n15601 ) ;
  assign n15603 = ( n2135 & n15524 ) | ( n2135 & ~n15602 ) | ( n15524 & ~n15602 ) ;
  assign n15604 = ( ~x151 & n9061 ) | ( ~x151 & n13012 ) | ( n9061 & n13012 ) ;
  assign n15605 = n6915 & ~n9515 ;
  assign n15606 = n15604 & n15605 ;
  assign n15607 = n4201 ^ x102 ^ 1'b0 ;
  assign n15608 = n14029 & n15607 ;
  assign n15609 = n15608 ^ n12003 ^ 1'b0 ;
  assign n15611 = ( ~n848 & n8391 ) | ( ~n848 & n13950 ) | ( n8391 & n13950 ) ;
  assign n15610 = n13291 ^ n7608 ^ 1'b0 ;
  assign n15612 = n15611 ^ n15610 ^ 1'b0 ;
  assign n15613 = n3107 & n15612 ;
  assign n15614 = n2960 & n7458 ;
  assign n15615 = n15614 ^ n11990 ^ 1'b0 ;
  assign n15616 = ( ~n8410 & n9603 ) | ( ~n8410 & n13065 ) | ( n9603 & n13065 ) ;
  assign n15617 = ( n7140 & n15470 ) | ( n7140 & n15616 ) | ( n15470 & n15616 ) ;
  assign n15618 = n15617 ^ n3512 ^ 1'b0 ;
  assign n15619 = n15615 & ~n15618 ;
  assign n15620 = n15619 ^ n10758 ^ n6677 ;
  assign n15625 = n5651 ^ n5251 ^ n525 ;
  assign n15626 = n15625 ^ n15436 ^ n5795 ;
  assign n15621 = n13458 ^ n10881 ^ n4574 ;
  assign n15622 = n15621 ^ n3495 ^ n1639 ;
  assign n15623 = ~n1493 & n15622 ;
  assign n15624 = n15623 ^ n12117 ^ 1'b0 ;
  assign n15627 = n15626 ^ n15624 ^ n7447 ;
  assign n15628 = ( n2663 & n3031 ) | ( n2663 & n6348 ) | ( n3031 & n6348 ) ;
  assign n15629 = n3624 & n5316 ;
  assign n15630 = ( n9118 & n15208 ) | ( n9118 & ~n15629 ) | ( n15208 & ~n15629 ) ;
  assign n15631 = ( n14396 & n15628 ) | ( n14396 & n15630 ) | ( n15628 & n15630 ) ;
  assign n15635 = ( x119 & ~x213 ) | ( x119 & n467 ) | ( ~x213 & n467 ) ;
  assign n15632 = n8232 ^ n2558 ^ n529 ;
  assign n15633 = n11338 ^ n9881 ^ n7609 ;
  assign n15634 = ( n1244 & n15632 ) | ( n1244 & ~n15633 ) | ( n15632 & ~n15633 ) ;
  assign n15636 = n15635 ^ n15634 ^ n11892 ;
  assign n15637 = n5737 ^ n5703 ^ 1'b0 ;
  assign n15638 = n15637 ^ n11151 ^ n3983 ;
  assign n15639 = ( n8908 & n15636 ) | ( n8908 & n15638 ) | ( n15636 & n15638 ) ;
  assign n15641 = n7500 ^ n2381 ^ 1'b0 ;
  assign n15640 = n468 & ~n5964 ;
  assign n15642 = n15641 ^ n15640 ^ n7330 ;
  assign n15643 = n15642 ^ n7801 ^ 1'b0 ;
  assign n15644 = ~n12093 & n15643 ;
  assign n15645 = n15644 ^ n15478 ^ 1'b0 ;
  assign n15646 = ~n3892 & n8722 ;
  assign n15647 = n15646 ^ n10095 ^ 1'b0 ;
  assign n15648 = n14930 | n15647 ;
  assign n15649 = x69 | n15648 ;
  assign n15650 = ( n1175 & n5832 ) | ( n1175 & n10763 ) | ( n5832 & n10763 ) ;
  assign n15651 = n14927 ^ n7462 ^ n2016 ;
  assign n15652 = ( n4600 & ~n6762 ) | ( n4600 & n15651 ) | ( ~n6762 & n15651 ) ;
  assign n15653 = ( n1677 & n15650 ) | ( n1677 & ~n15652 ) | ( n15650 & ~n15652 ) ;
  assign n15655 = x10 & ~n12812 ;
  assign n15656 = n15655 ^ n2123 ^ 1'b0 ;
  assign n15657 = n15656 ^ n5776 ^ x194 ;
  assign n15654 = n3128 ^ n1998 ^ 1'b0 ;
  assign n15658 = n15657 ^ n15654 ^ n6765 ;
  assign n15659 = n1437 ^ n1179 ^ n680 ;
  assign n15660 = ( n2080 & ~n3369 ) | ( n2080 & n10432 ) | ( ~n3369 & n10432 ) ;
  assign n15661 = ( n2539 & n9343 ) | ( n2539 & ~n15660 ) | ( n9343 & ~n15660 ) ;
  assign n15662 = n15659 | n15661 ;
  assign n15663 = n15658 | n15662 ;
  assign n15664 = n11590 ^ n2648 ^ 1'b0 ;
  assign n15665 = n15664 ^ n4010 ^ n3494 ;
  assign n15666 = ~n7195 & n8677 ;
  assign n15667 = n494 & n15666 ;
  assign n15668 = n15667 ^ n9854 ^ 1'b0 ;
  assign n15669 = n13627 & ~n15668 ;
  assign n15670 = n6653 ^ n5961 ^ 1'b0 ;
  assign n15671 = n15669 & n15670 ;
  assign n15672 = ( n4805 & ~n7025 ) | ( n4805 & n10369 ) | ( ~n7025 & n10369 ) ;
  assign n15673 = n15672 ^ n13737 ^ n3005 ;
  assign n15674 = n5533 & ~n13063 ;
  assign n15675 = n15674 ^ n10711 ^ n10650 ;
  assign n15676 = n9895 ^ n7950 ^ 1'b0 ;
  assign n15677 = n1014 & n3244 ;
  assign n15678 = ( n783 & ~n1783 ) | ( n783 & n4998 ) | ( ~n1783 & n4998 ) ;
  assign n15679 = n15678 ^ n3937 ^ n2958 ;
  assign n15680 = n13784 ^ n13247 ^ 1'b0 ;
  assign n15681 = ~n3106 & n15680 ;
  assign n15682 = n13205 ^ n2362 ^ 1'b0 ;
  assign n15683 = n8336 | n15682 ;
  assign n15684 = n15683 ^ n8905 ^ n8751 ;
  assign n15685 = ~n14227 & n15684 ;
  assign n15686 = ~n15681 & n15685 ;
  assign n15687 = n6933 ^ n6644 ^ n4738 ;
  assign n15688 = n15687 ^ n15456 ^ n10976 ;
  assign n15689 = n8754 & ~n15688 ;
  assign n15690 = n10303 ^ n9100 ^ n5312 ;
  assign n15691 = n9565 ^ n9142 ^ n7667 ;
  assign n15692 = ( ~n15689 & n15690 ) | ( ~n15689 & n15691 ) | ( n15690 & n15691 ) ;
  assign n15693 = ~x39 & n5462 ;
  assign n15694 = n4249 | n15693 ;
  assign n15695 = n5782 | n6824 ;
  assign n15696 = n13689 & ~n15695 ;
  assign n15697 = ( n5503 & ~n6991 ) | ( n5503 & n15696 ) | ( ~n6991 & n15696 ) ;
  assign n15698 = ( n7109 & n15694 ) | ( n7109 & ~n15697 ) | ( n15694 & ~n15697 ) ;
  assign n15699 = ( x192 & n9662 ) | ( x192 & n10826 ) | ( n9662 & n10826 ) ;
  assign n15700 = ~n13367 & n15699 ;
  assign n15701 = ~n14784 & n15700 ;
  assign n15702 = n12337 ^ n4965 ^ 1'b0 ;
  assign n15703 = n15701 | n15702 ;
  assign n15704 = n15703 ^ n2523 ^ 1'b0 ;
  assign n15705 = n4285 & n15704 ;
  assign n15706 = n6976 ^ n2085 ^ 1'b0 ;
  assign n15707 = ~n9171 & n15706 ;
  assign n15711 = n8002 ^ n4451 ^ 1'b0 ;
  assign n15710 = n12588 & ~n13482 ;
  assign n15712 = n15711 ^ n15710 ^ 1'b0 ;
  assign n15708 = n12577 ^ n4884 ^ 1'b0 ;
  assign n15709 = n11567 & n15708 ;
  assign n15713 = n15712 ^ n15709 ^ 1'b0 ;
  assign n15714 = n5203 & n15713 ;
  assign n15715 = n2680 & ~n4652 ;
  assign n15716 = n15715 ^ n14725 ^ n9396 ;
  assign n15717 = ( n2695 & ~n12070 ) | ( n2695 & n15716 ) | ( ~n12070 & n15716 ) ;
  assign n15718 = n2560 & n15717 ;
  assign n15721 = n8964 ^ n7132 ^ n6348 ;
  assign n15719 = ( n3213 & n3736 ) | ( n3213 & n6017 ) | ( n3736 & n6017 ) ;
  assign n15720 = n4657 | n15719 ;
  assign n15722 = n15721 ^ n15720 ^ n4697 ;
  assign n15723 = n12961 ^ n908 ^ 1'b0 ;
  assign n15733 = n5820 ^ n355 ^ 1'b0 ;
  assign n15734 = n508 & ~n15733 ;
  assign n15735 = n3916 & n15734 ;
  assign n15736 = ~n2052 & n15735 ;
  assign n15737 = n15736 ^ n15368 ^ n6035 ;
  assign n15731 = ( n1771 & n3532 ) | ( n1771 & n10947 ) | ( n3532 & n10947 ) ;
  assign n15732 = n15731 ^ n13521 ^ 1'b0 ;
  assign n15726 = x226 & n331 ;
  assign n15727 = n15726 ^ n268 ^ 1'b0 ;
  assign n15728 = n15727 ^ n8150 ^ n3945 ;
  assign n15724 = ( n1172 & n1500 ) | ( n1172 & ~n4539 ) | ( n1500 & ~n4539 ) ;
  assign n15725 = ( n419 & n1572 ) | ( n419 & n15724 ) | ( n1572 & n15724 ) ;
  assign n15729 = n15728 ^ n15725 ^ n10409 ;
  assign n15730 = n10056 & ~n15729 ;
  assign n15738 = n15737 ^ n15732 ^ n15730 ;
  assign n15739 = n15738 ^ n8178 ^ 1'b0 ;
  assign n15740 = ~n8820 & n15739 ;
  assign n15741 = n5307 | n6593 ;
  assign n15742 = n7039 ^ n6722 ^ n2544 ;
  assign n15743 = n15742 ^ n11946 ^ 1'b0 ;
  assign n15744 = n15741 | n15743 ;
  assign n15745 = n15744 ^ n9320 ^ 1'b0 ;
  assign n15756 = n3124 ^ n1714 ^ n473 ;
  assign n15750 = n11409 ^ n2336 ^ 1'b0 ;
  assign n15751 = n1485 & n15750 ;
  assign n15752 = x177 & ~n10947 ;
  assign n15753 = n2223 & n15752 ;
  assign n15754 = n3708 & n12980 ;
  assign n15755 = ( ~n15751 & n15753 ) | ( ~n15751 & n15754 ) | ( n15753 & n15754 ) ;
  assign n15746 = n6864 ^ n5525 ^ n1471 ;
  assign n15747 = n11494 ^ n1768 ^ 1'b0 ;
  assign n15748 = ~n15746 & n15747 ;
  assign n15749 = n15748 ^ n8120 ^ x4 ;
  assign n15757 = n15756 ^ n15755 ^ n15749 ;
  assign n15758 = n3497 & ~n9885 ;
  assign n15759 = n7826 & n15758 ;
  assign n15760 = n14159 ^ n2825 ^ n1997 ;
  assign n15761 = ( ~n1242 & n3285 ) | ( ~n1242 & n15760 ) | ( n3285 & n15760 ) ;
  assign n15762 = n15761 ^ n14813 ^ 1'b0 ;
  assign n15763 = n14381 | n15762 ;
  assign n15764 = n15469 ^ n7413 ^ n6943 ;
  assign n15765 = n6820 ^ n6137 ^ n3525 ;
  assign n15766 = ( n14533 & n15764 ) | ( n14533 & n15765 ) | ( n15764 & n15765 ) ;
  assign n15767 = n3278 ^ n2479 ^ 1'b0 ;
  assign n15768 = ( n4375 & n9680 ) | ( n4375 & n15767 ) | ( n9680 & n15767 ) ;
  assign n15769 = n2560 | n11742 ;
  assign n15770 = n15769 ^ n2802 ^ 1'b0 ;
  assign n15771 = ~n3178 & n15770 ;
  assign n15772 = n15771 ^ n9485 ^ 1'b0 ;
  assign n15773 = n15772 ^ n13207 ^ 1'b0 ;
  assign n15774 = ( ~n9249 & n15768 ) | ( ~n9249 & n15773 ) | ( n15768 & n15773 ) ;
  assign n15775 = n15774 ^ n8468 ^ n7295 ;
  assign n15785 = n8468 ^ n4258 ^ 1'b0 ;
  assign n15786 = n15785 ^ n10969 ^ n5355 ;
  assign n15782 = ( n783 & n3588 ) | ( n783 & ~n7447 ) | ( n3588 & ~n7447 ) ;
  assign n15783 = n15782 ^ n3035 ^ 1'b0 ;
  assign n15776 = n12939 ^ n10869 ^ n7493 ;
  assign n15777 = n6775 & ~n8170 ;
  assign n15778 = n2007 & n15777 ;
  assign n15779 = ( n14795 & n15596 ) | ( n14795 & ~n15778 ) | ( n15596 & ~n15778 ) ;
  assign n15780 = n15779 ^ n15744 ^ n9956 ;
  assign n15781 = n15776 & ~n15780 ;
  assign n15784 = n15783 ^ n15781 ^ 1'b0 ;
  assign n15787 = n15786 ^ n15784 ^ n8325 ;
  assign n15788 = n12553 ^ n4818 ^ n273 ;
  assign n15789 = n2570 & n4261 ;
  assign n15790 = ~x66 & n15789 ;
  assign n15791 = n9235 ^ n2859 ^ 1'b0 ;
  assign n15792 = n15790 | n15791 ;
  assign n15793 = n15788 & ~n15792 ;
  assign n15794 = ~n3607 & n3965 ;
  assign n15795 = ~x75 & n15794 ;
  assign n15796 = n6892 & n10060 ;
  assign n15797 = n15796 ^ n1678 ^ 1'b0 ;
  assign n15798 = n3887 & ~n15123 ;
  assign n15799 = n15797 & n15798 ;
  assign n15800 = n818 & ~n15799 ;
  assign n15801 = n15795 & n15800 ;
  assign n15802 = ( x67 & ~n528 ) | ( x67 & n9659 ) | ( ~n528 & n9659 ) ;
  assign n15803 = ( n419 & n2202 ) | ( n419 & n3012 ) | ( n2202 & n3012 ) ;
  assign n15804 = n3247 ^ n874 ^ x141 ;
  assign n15805 = ( n2321 & n3962 ) | ( n2321 & n15804 ) | ( n3962 & n15804 ) ;
  assign n15807 = n3508 ^ n905 ^ 1'b0 ;
  assign n15808 = n10431 & ~n15807 ;
  assign n15809 = n15808 ^ n8413 ^ 1'b0 ;
  assign n15806 = n7214 & n8174 ;
  assign n15810 = n15809 ^ n15806 ^ 1'b0 ;
  assign n15811 = n9639 ^ n927 ^ n542 ;
  assign n15812 = n894 | n15811 ;
  assign n15813 = n6429 & ~n15812 ;
  assign n15814 = n15813 ^ n9940 ^ x207 ;
  assign n15815 = ( n4480 & n12133 ) | ( n4480 & ~n15814 ) | ( n12133 & ~n15814 ) ;
  assign n15816 = ( ~n2402 & n6495 ) | ( ~n2402 & n12226 ) | ( n6495 & n12226 ) ;
  assign n15817 = ( n1436 & n3633 ) | ( n1436 & n9758 ) | ( n3633 & n9758 ) ;
  assign n15818 = n15817 ^ n4805 ^ 1'b0 ;
  assign n15819 = n15378 & n15818 ;
  assign n15820 = ( ~n13382 & n15816 ) | ( ~n13382 & n15819 ) | ( n15816 & n15819 ) ;
  assign n15824 = n11875 ^ n9113 ^ 1'b0 ;
  assign n15825 = n6246 & n15824 ;
  assign n15821 = ( n742 & n2591 ) | ( n742 & ~n4221 ) | ( n2591 & ~n4221 ) ;
  assign n15822 = ( n1074 & n14712 ) | ( n1074 & ~n15821 ) | ( n14712 & ~n15821 ) ;
  assign n15823 = n883 & ~n15822 ;
  assign n15826 = n15825 ^ n15823 ^ 1'b0 ;
  assign n15828 = n507 & n2573 ;
  assign n15829 = n15828 ^ n12012 ^ n3261 ;
  assign n15830 = n7134 | n15829 ;
  assign n15827 = ( ~n847 & n5951 ) | ( ~n847 & n8769 ) | ( n5951 & n8769 ) ;
  assign n15831 = n15830 ^ n15827 ^ n9765 ;
  assign n15832 = n15831 ^ n12561 ^ n8902 ;
  assign n15833 = n356 | n2552 ;
  assign n15834 = n5002 | n9472 ;
  assign n15835 = n15833 | n15834 ;
  assign n15836 = n15835 ^ n6470 ^ 1'b0 ;
  assign n15837 = n9614 ^ n7940 ^ 1'b0 ;
  assign n15838 = n15836 & ~n15837 ;
  assign n15839 = ( n12424 & ~n12502 ) | ( n12424 & n15838 ) | ( ~n12502 & n15838 ) ;
  assign n15840 = ( x54 & n2462 ) | ( x54 & n2561 ) | ( n2462 & n2561 ) ;
  assign n15841 = ( ~n4955 & n14736 ) | ( ~n4955 & n15840 ) | ( n14736 & n15840 ) ;
  assign n15842 = n7603 ^ n2617 ^ n2262 ;
  assign n15843 = n7032 & ~n15842 ;
  assign n15844 = ~n15841 & n15843 ;
  assign n15847 = n15437 ^ n4988 ^ 1'b0 ;
  assign n15845 = n9839 ^ n7251 ^ n4310 ;
  assign n15846 = ( ~n8012 & n13954 ) | ( ~n8012 & n15845 ) | ( n13954 & n15845 ) ;
  assign n15848 = n15847 ^ n15846 ^ n5332 ;
  assign n15858 = ( n290 & ~n5259 ) | ( n290 & n6205 ) | ( ~n5259 & n6205 ) ;
  assign n15859 = n14857 ^ n5443 ^ 1'b0 ;
  assign n15860 = ~n15858 & n15859 ;
  assign n15849 = n1278 ^ n635 ^ n378 ;
  assign n15850 = n15849 ^ n5992 ^ 1'b0 ;
  assign n15851 = ( n8730 & n14016 ) | ( n8730 & n15850 ) | ( n14016 & n15850 ) ;
  assign n15852 = n3639 ^ n2520 ^ 1'b0 ;
  assign n15853 = n3644 ^ n1329 ^ 1'b0 ;
  assign n15854 = n1100 | n15853 ;
  assign n15855 = n15852 | n15854 ;
  assign n15856 = ( n3867 & ~n4405 ) | ( n3867 & n15855 ) | ( ~n4405 & n15855 ) ;
  assign n15857 = ( x217 & n15851 ) | ( x217 & n15856 ) | ( n15851 & n15856 ) ;
  assign n15861 = n15860 ^ n15857 ^ n882 ;
  assign n15862 = n13610 | n15786 ;
  assign n15863 = n4671 & ~n15862 ;
  assign n15864 = ~n1926 & n7253 ;
  assign n15865 = n15864 ^ n10416 ^ 1'b0 ;
  assign n15866 = n5649 ^ n2659 ^ x19 ;
  assign n15868 = ~n11283 & n11724 ;
  assign n15867 = n502 & n2974 ;
  assign n15869 = n15868 ^ n15867 ^ 1'b0 ;
  assign n15870 = ( ~n1104 & n15866 ) | ( ~n1104 & n15869 ) | ( n15866 & n15869 ) ;
  assign n15871 = n15870 ^ n5196 ^ 1'b0 ;
  assign n15874 = n367 & ~n382 ;
  assign n15875 = n15874 ^ n2572 ^ 1'b0 ;
  assign n15876 = ( ~n380 & n1066 ) | ( ~n380 & n15875 ) | ( n1066 & n15875 ) ;
  assign n15877 = n4988 & ~n4999 ;
  assign n15878 = ~n15876 & n15877 ;
  assign n15872 = n2362 & n4247 ;
  assign n15873 = ~n819 & n15872 ;
  assign n15879 = n15878 ^ n15873 ^ n8506 ;
  assign n15880 = ( n1855 & ~n1856 ) | ( n1855 & n4474 ) | ( ~n1856 & n4474 ) ;
  assign n15881 = n15880 ^ n3334 ^ n854 ;
  assign n15882 = n15881 ^ x224 ^ 1'b0 ;
  assign n15883 = ~n9130 & n15882 ;
  assign n15884 = n15883 ^ n12289 ^ n12209 ;
  assign n15885 = ( ~n6132 & n7260 ) | ( ~n6132 & n15884 ) | ( n7260 & n15884 ) ;
  assign n15886 = n3427 | n9616 ;
  assign n15887 = n15411 & n15886 ;
  assign n15888 = n10421 ^ n5054 ^ 1'b0 ;
  assign n15900 = ( n3453 & ~n4810 ) | ( n3453 & n4922 ) | ( ~n4810 & n4922 ) ;
  assign n15901 = n15900 ^ n7319 ^ n7066 ;
  assign n15894 = n825 ^ n486 ^ 1'b0 ;
  assign n15895 = n3617 & ~n15894 ;
  assign n15897 = n6132 ^ n3775 ^ n3524 ;
  assign n15896 = n3844 ^ n3192 ^ x162 ;
  assign n15898 = n15897 ^ n15896 ^ n11401 ;
  assign n15899 = ( n4030 & n15895 ) | ( n4030 & n15898 ) | ( n15895 & n15898 ) ;
  assign n15889 = ( n3617 & ~n4066 ) | ( n3617 & n13338 ) | ( ~n4066 & n13338 ) ;
  assign n15890 = x99 & ~n6142 ;
  assign n15891 = ~n15889 & n15890 ;
  assign n15892 = n7467 | n15891 ;
  assign n15893 = n15892 ^ n6596 ^ 1'b0 ;
  assign n15902 = n15901 ^ n15899 ^ n15893 ;
  assign n15903 = n3245 ^ n1553 ^ n966 ;
  assign n15904 = ( n2321 & n2494 ) | ( n2321 & n15903 ) | ( n2494 & n15903 ) ;
  assign n15905 = n15904 ^ n9332 ^ n4730 ;
  assign n15906 = ( n3534 & n11811 ) | ( n3534 & n15905 ) | ( n11811 & n15905 ) ;
  assign n15907 = n7937 & ~n15553 ;
  assign n15908 = n15313 ^ n8951 ^ n3497 ;
  assign n15909 = ( ~n12985 & n13117 ) | ( ~n12985 & n15908 ) | ( n13117 & n15908 ) ;
  assign n15911 = ~n4673 & n6649 ;
  assign n15912 = n15911 ^ n15173 ^ n5676 ;
  assign n15910 = n749 & ~n3855 ;
  assign n15913 = n15912 ^ n15910 ^ 1'b0 ;
  assign n15914 = n4944 ^ n2062 ^ x156 ;
  assign n15915 = n15914 ^ n8041 ^ 1'b0 ;
  assign n15916 = n15915 ^ n7426 ^ n6214 ;
  assign n15917 = n15913 & ~n15916 ;
  assign n15918 = n15917 ^ n461 ^ 1'b0 ;
  assign n15919 = n15368 ^ n8727 ^ 1'b0 ;
  assign n15920 = n5620 | n6706 ;
  assign n15921 = n7407 & ~n15920 ;
  assign n15922 = n6379 & n9481 ;
  assign n15923 = n15921 & n15922 ;
  assign n15924 = ( n7444 & n15919 ) | ( n7444 & ~n15923 ) | ( n15919 & ~n15923 ) ;
  assign n15925 = n10228 ^ n8666 ^ n5205 ;
  assign n15926 = n7373 ^ n6105 ^ n2575 ;
  assign n15927 = ( n5339 & n10673 ) | ( n5339 & ~n15926 ) | ( n10673 & ~n15926 ) ;
  assign n15928 = n12346 ^ n10268 ^ n800 ;
  assign n15929 = n15928 ^ n11006 ^ 1'b0 ;
  assign n15930 = n6480 | n15929 ;
  assign n15931 = n941 | n12121 ;
  assign n15932 = n15931 ^ n4762 ^ 1'b0 ;
  assign n15933 = n15930 | n15932 ;
  assign n15934 = n15933 ^ n5626 ^ n522 ;
  assign n15935 = n9264 ^ n3569 ^ 1'b0 ;
  assign n15936 = n15935 ^ n11690 ^ n6555 ;
  assign n15937 = n15936 ^ n1290 ^ n599 ;
  assign n15938 = n15937 ^ n481 ^ 1'b0 ;
  assign n15939 = n6246 & ~n15938 ;
  assign n15940 = n665 & n3147 ;
  assign n15941 = n15940 ^ n1927 ^ 1'b0 ;
  assign n15942 = n15941 ^ n952 ^ 1'b0 ;
  assign n15943 = n3449 ^ n665 ^ x53 ;
  assign n15944 = n15943 ^ n5531 ^ n796 ;
  assign n15945 = ( n12656 & ~n13275 ) | ( n12656 & n15944 ) | ( ~n13275 & n15944 ) ;
  assign n15946 = ~n14944 & n15945 ;
  assign n15947 = ( ~n2872 & n3581 ) | ( ~n2872 & n9593 ) | ( n3581 & n9593 ) ;
  assign n15948 = n15947 ^ n10520 ^ 1'b0 ;
  assign n15949 = ( x86 & n1991 ) | ( x86 & ~n2741 ) | ( n1991 & ~n2741 ) ;
  assign n15950 = ( n3285 & n3594 ) | ( n3285 & ~n5121 ) | ( n3594 & ~n5121 ) ;
  assign n15951 = ( n14011 & ~n15949 ) | ( n14011 & n15950 ) | ( ~n15949 & n15950 ) ;
  assign n15954 = n12340 ^ n2910 ^ 1'b0 ;
  assign n15955 = n15954 ^ n2400 ^ n2156 ;
  assign n15952 = n6144 & n9170 ;
  assign n15953 = n15952 ^ n10152 ^ n9673 ;
  assign n15956 = n15955 ^ n15953 ^ n4639 ;
  assign n15957 = ( n4294 & n10727 ) | ( n4294 & ~n12412 ) | ( n10727 & ~n12412 ) ;
  assign n15958 = ( n1041 & ~n13779 ) | ( n1041 & n15957 ) | ( ~n13779 & n15957 ) ;
  assign n15959 = n5092 | n7506 ;
  assign n15960 = ~n15566 & n15959 ;
  assign n15961 = n11322 ^ n8478 ^ n6554 ;
  assign n15962 = n12696 ^ n1920 ^ 1'b0 ;
  assign n15963 = n13441 ^ n3954 ^ 1'b0 ;
  assign n15964 = ~n15962 & n15963 ;
  assign n15965 = n13460 ^ n8055 ^ 1'b0 ;
  assign n15966 = n5444 & n7463 ;
  assign n15967 = n15966 ^ n2168 ^ 1'b0 ;
  assign n15968 = ( n13660 & n15965 ) | ( n13660 & ~n15967 ) | ( n15965 & ~n15967 ) ;
  assign n15969 = n15968 ^ n15331 ^ 1'b0 ;
  assign n15976 = n6708 ^ n5920 ^ 1'b0 ;
  assign n15970 = n6836 ^ n4331 ^ 1'b0 ;
  assign n15971 = n11201 & ~n15970 ;
  assign n15972 = ( n9400 & n10817 ) | ( n9400 & n14099 ) | ( n10817 & n14099 ) ;
  assign n15973 = n15626 & n15972 ;
  assign n15974 = ~n15971 & n15973 ;
  assign n15975 = ( n5298 & ~n5856 ) | ( n5298 & n15974 ) | ( ~n5856 & n15974 ) ;
  assign n15977 = n15976 ^ n15975 ^ 1'b0 ;
  assign n15978 = n7959 & ~n15977 ;
  assign n15980 = n5827 ^ n5670 ^ n537 ;
  assign n15979 = ( n1499 & ~n2265 ) | ( n1499 & n11075 ) | ( ~n2265 & n11075 ) ;
  assign n15981 = n15980 ^ n15979 ^ 1'b0 ;
  assign n15982 = ~n894 & n15981 ;
  assign n15983 = n710 & n4545 ;
  assign n15984 = ~n2472 & n8781 ;
  assign n15985 = n9680 ^ n2088 ^ 1'b0 ;
  assign n15986 = n14767 & n15985 ;
  assign n15987 = ( n2027 & n3173 ) | ( n2027 & n15986 ) | ( n3173 & n15986 ) ;
  assign n15988 = n14645 & ~n15987 ;
  assign n15989 = n15988 ^ n3623 ^ 1'b0 ;
  assign n15990 = n11384 ^ n6482 ^ n3697 ;
  assign n15991 = n7098 & ~n15990 ;
  assign n15992 = n15991 ^ n6339 ^ 1'b0 ;
  assign n15993 = n8777 ^ n3657 ^ n2552 ;
  assign n15994 = ( n2260 & ~n15992 ) | ( n2260 & n15993 ) | ( ~n15992 & n15993 ) ;
  assign n15995 = n13434 ^ n10742 ^ n8102 ;
  assign n15996 = n14010 ^ n13794 ^ 1'b0 ;
  assign n15997 = n13292 & ~n15996 ;
  assign n15998 = n15995 & n15997 ;
  assign n15999 = n15998 ^ n11494 ^ 1'b0 ;
  assign n16000 = ( n11273 & ~n15994 ) | ( n11273 & n15999 ) | ( ~n15994 & n15999 ) ;
  assign n16001 = n3497 ^ n2689 ^ n961 ;
  assign n16002 = ( n2348 & n4023 ) | ( n2348 & n16001 ) | ( n4023 & n16001 ) ;
  assign n16003 = x183 & n4089 ;
  assign n16004 = n670 | n1641 ;
  assign n16005 = ( ~x27 & n12884 ) | ( ~x27 & n16004 ) | ( n12884 & n16004 ) ;
  assign n16006 = n16005 ^ n10082 ^ n9799 ;
  assign n16007 = n3072 & n16006 ;
  assign n16008 = ( ~n16002 & n16003 ) | ( ~n16002 & n16007 ) | ( n16003 & n16007 ) ;
  assign n16009 = x40 & ~n549 ;
  assign n16010 = n5253 & n16009 ;
  assign n16011 = n12068 & ~n16010 ;
  assign n16012 = ( n4999 & n8039 ) | ( n4999 & ~n16011 ) | ( n8039 & ~n16011 ) ;
  assign n16013 = ( n1488 & ~n2401 ) | ( n1488 & n5245 ) | ( ~n2401 & n5245 ) ;
  assign n16014 = n5344 & n16013 ;
  assign n16015 = n16014 ^ n13603 ^ n12826 ;
  assign n16016 = n9078 ^ n3157 ^ 1'b0 ;
  assign n16022 = n4481 ^ n2786 ^ n1580 ;
  assign n16021 = n735 & n9076 ;
  assign n16023 = n16022 ^ n16021 ^ 1'b0 ;
  assign n16017 = n610 | n1712 ;
  assign n16018 = n282 | n16017 ;
  assign n16019 = n16018 ^ n11286 ^ 1'b0 ;
  assign n16020 = ( n7748 & n8253 ) | ( n7748 & n16019 ) | ( n8253 & n16019 ) ;
  assign n16024 = n16023 ^ n16020 ^ n6550 ;
  assign n16025 = ( n328 & n16016 ) | ( n328 & ~n16024 ) | ( n16016 & ~n16024 ) ;
  assign n16026 = ( n12286 & n12731 ) | ( n12286 & ~n15043 ) | ( n12731 & ~n15043 ) ;
  assign n16027 = ~n1057 & n2255 ;
  assign n16028 = ( n8206 & ~n11843 ) | ( n8206 & n16027 ) | ( ~n11843 & n16027 ) ;
  assign n16029 = n16028 ^ n3130 ^ 1'b0 ;
  assign n16030 = n12705 ^ n5531 ^ 1'b0 ;
  assign n16031 = n16029 & ~n16030 ;
  assign n16032 = n6263 ^ n4427 ^ n3973 ;
  assign n16033 = n16032 ^ n14050 ^ 1'b0 ;
  assign n16036 = n3587 ^ n3284 ^ n2417 ;
  assign n16037 = n16036 ^ n13732 ^ n3435 ;
  assign n16034 = n328 & n11614 ;
  assign n16035 = ~n5695 & n16034 ;
  assign n16038 = n16037 ^ n16035 ^ 1'b0 ;
  assign n16039 = n16033 | n16038 ;
  assign n16040 = n4469 & n16039 ;
  assign n16041 = ( n852 & n2680 ) | ( n852 & ~n8640 ) | ( n2680 & ~n8640 ) ;
  assign n16042 = n8674 | n16041 ;
  assign n16043 = n16042 ^ n11422 ^ n2040 ;
  assign n16044 = n16043 ^ n11245 ^ 1'b0 ;
  assign n16045 = ~n12293 & n16044 ;
  assign n16046 = n5275 ^ n4239 ^ n2348 ;
  assign n16047 = ( n2263 & n2433 ) | ( n2263 & n7361 ) | ( n2433 & n7361 ) ;
  assign n16048 = ( n6424 & ~n16046 ) | ( n6424 & n16047 ) | ( ~n16046 & n16047 ) ;
  assign n16049 = n16048 ^ n11475 ^ n1771 ;
  assign n16050 = ( n1288 & ~n5225 ) | ( n1288 & n16049 ) | ( ~n5225 & n16049 ) ;
  assign n16051 = ~n1590 & n16050 ;
  assign n16052 = n595 & n16051 ;
  assign n16055 = ( ~n1225 & n4243 ) | ( ~n1225 & n13205 ) | ( n4243 & n13205 ) ;
  assign n16056 = n16055 ^ n3574 ^ 1'b0 ;
  assign n16057 = n7321 | n16056 ;
  assign n16053 = n9769 & n15699 ;
  assign n16054 = n6919 & n16053 ;
  assign n16058 = n16057 ^ n16054 ^ n759 ;
  assign n16059 = n15160 ^ n6405 ^ 1'b0 ;
  assign n16060 = n559 & n16059 ;
  assign n16061 = n15416 ^ n13900 ^ n9847 ;
  assign n16062 = n1886 ^ n687 ^ 1'b0 ;
  assign n16063 = n4670 & n16062 ;
  assign n16064 = n10947 ^ n2542 ^ 1'b0 ;
  assign n16065 = n4019 ^ n1571 ^ 1'b0 ;
  assign n16066 = n9323 ^ n6245 ^ n6114 ;
  assign n16067 = n2662 ^ n1751 ^ 1'b0 ;
  assign n16068 = n2703 | n16067 ;
  assign n16069 = n6232 | n16068 ;
  assign n16070 = n16069 ^ n5985 ^ n2739 ;
  assign n16071 = ( n16065 & ~n16066 ) | ( n16065 & n16070 ) | ( ~n16066 & n16070 ) ;
  assign n16072 = ( n16063 & ~n16064 ) | ( n16063 & n16071 ) | ( ~n16064 & n16071 ) ;
  assign n16073 = n12272 ^ n6982 ^ 1'b0 ;
  assign n16074 = n16073 ^ n1808 ^ n812 ;
  assign n16075 = ( n3320 & n4072 ) | ( n3320 & n9496 ) | ( n4072 & n9496 ) ;
  assign n16076 = n7007 ^ n6991 ^ n2227 ;
  assign n16077 = n9974 ^ n5396 ^ 1'b0 ;
  assign n16078 = n10930 & ~n16077 ;
  assign n16079 = n364 | n8182 ;
  assign n16080 = n2266 | n16079 ;
  assign n16081 = ~n1820 & n16080 ;
  assign n16082 = n16081 ^ n12479 ^ 1'b0 ;
  assign n16083 = ~n9727 & n16082 ;
  assign n16084 = n10845 | n16083 ;
  assign n16085 = ( n8621 & ~n16078 ) | ( n8621 & n16084 ) | ( ~n16078 & n16084 ) ;
  assign n16086 = n9970 & ~n11536 ;
  assign n16087 = n875 | n9173 ;
  assign n16088 = n16087 ^ n1868 ^ 1'b0 ;
  assign n16089 = n6794 ^ n3155 ^ 1'b0 ;
  assign n16090 = n5984 | n16089 ;
  assign n16091 = ( n4081 & ~n8714 ) | ( n4081 & n16090 ) | ( ~n8714 & n16090 ) ;
  assign n16092 = n16091 ^ n10446 ^ n3542 ;
  assign n16093 = n11271 ^ n9848 ^ n6899 ;
  assign n16094 = n16093 ^ n15853 ^ n6388 ;
  assign n16095 = n16094 ^ n11276 ^ 1'b0 ;
  assign n16096 = ~n1808 & n16095 ;
  assign n16100 = n7972 ^ n7173 ^ 1'b0 ;
  assign n16101 = n7417 | n16100 ;
  assign n16103 = n3629 ^ n2762 ^ 1'b0 ;
  assign n16104 = x157 & n16103 ;
  assign n16102 = ( n2732 & n4698 ) | ( n2732 & ~n5241 ) | ( n4698 & ~n5241 ) ;
  assign n16105 = n16104 ^ n16102 ^ x108 ;
  assign n16106 = ( n6268 & ~n16101 ) | ( n6268 & n16105 ) | ( ~n16101 & n16105 ) ;
  assign n16097 = n3669 & ~n13173 ;
  assign n16098 = n8838 & ~n16097 ;
  assign n16099 = ~n13696 & n16098 ;
  assign n16107 = n16106 ^ n16099 ^ n14077 ;
  assign n16108 = n13996 ^ n13699 ^ 1'b0 ;
  assign n16111 = ( n5018 & n7297 ) | ( n5018 & ~n7329 ) | ( n7297 & ~n7329 ) ;
  assign n16109 = n6529 & ~n10784 ;
  assign n16110 = n10359 & n16109 ;
  assign n16112 = n16111 ^ n16110 ^ n4474 ;
  assign n16113 = ( n2127 & n2356 ) | ( n2127 & n9997 ) | ( n2356 & n9997 ) ;
  assign n16114 = ( ~n399 & n1386 ) | ( ~n399 & n6167 ) | ( n1386 & n6167 ) ;
  assign n16115 = n16113 | n16114 ;
  assign n16116 = n16113 & ~n16115 ;
  assign n16117 = n7603 & ~n11052 ;
  assign n16118 = ( ~n1685 & n6045 ) | ( ~n1685 & n7349 ) | ( n6045 & n7349 ) ;
  assign n16119 = ( n7169 & n13441 ) | ( n7169 & ~n16118 ) | ( n13441 & ~n16118 ) ;
  assign n16120 = ~n16117 & n16119 ;
  assign n16121 = n16120 ^ n1375 ^ 1'b0 ;
  assign n16122 = ( n10400 & n14522 ) | ( n10400 & n16121 ) | ( n14522 & n16121 ) ;
  assign n16124 = ( n4437 & n6333 ) | ( n4437 & n13904 ) | ( n6333 & n13904 ) ;
  assign n16123 = ~n2150 & n8680 ;
  assign n16125 = n16124 ^ n16123 ^ 1'b0 ;
  assign n16126 = n16122 & n16125 ;
  assign n16129 = ~n7798 & n10419 ;
  assign n16127 = n12390 ^ n1317 ^ 1'b0 ;
  assign n16128 = n7451 & n16127 ;
  assign n16130 = n16129 ^ n16128 ^ n10725 ;
  assign n16131 = n16130 ^ n14022 ^ n2962 ;
  assign n16132 = n7434 | n10152 ;
  assign n16133 = n16132 ^ n7871 ^ n3107 ;
  assign n16134 = n8441 ^ n4309 ^ n2245 ;
  assign n16135 = x122 & n6952 ;
  assign n16136 = ~n7466 & n16135 ;
  assign n16137 = ( n3288 & n16134 ) | ( n3288 & n16136 ) | ( n16134 & n16136 ) ;
  assign n16138 = n1777 ^ n690 ^ n490 ;
  assign n16139 = n16138 ^ n4772 ^ x126 ;
  assign n16140 = n16137 & n16139 ;
  assign n16141 = n653 & n3770 ;
  assign n16142 = n5478 | n13717 ;
  assign n16143 = ~n676 & n3287 ;
  assign n16144 = n16143 ^ n15566 ^ 1'b0 ;
  assign n16163 = n14344 ^ n2362 ^ 1'b0 ;
  assign n16164 = ~n570 & n16163 ;
  assign n16159 = ( ~n2449 & n6437 ) | ( ~n2449 & n13130 ) | ( n6437 & n13130 ) ;
  assign n16160 = n16159 ^ n4196 ^ 1'b0 ;
  assign n16161 = n8009 & ~n16160 ;
  assign n16158 = n9314 ^ n2998 ^ n2296 ;
  assign n16162 = n16161 ^ n16158 ^ n2468 ;
  assign n16156 = ( ~n1626 & n4238 ) | ( ~n1626 & n4911 ) | ( n4238 & n4911 ) ;
  assign n16153 = x253 & ~n1272 ;
  assign n16154 = ~n2712 & n16153 ;
  assign n16148 = ( n549 & n943 ) | ( n549 & ~n6143 ) | ( n943 & ~n6143 ) ;
  assign n16149 = n4047 | n16148 ;
  assign n16150 = n16149 ^ n5095 ^ 1'b0 ;
  assign n16151 = n16150 ^ n7209 ^ 1'b0 ;
  assign n16152 = n6985 | n16151 ;
  assign n16155 = n16154 ^ n16152 ^ n5110 ;
  assign n16145 = n10282 ^ n3598 ^ 1'b0 ;
  assign n16146 = n16145 ^ n12070 ^ n3588 ;
  assign n16147 = n16146 ^ n10602 ^ n2786 ;
  assign n16157 = n16156 ^ n16155 ^ n16147 ;
  assign n16165 = n16164 ^ n16162 ^ n16157 ;
  assign n16166 = n3653 ^ n3058 ^ n552 ;
  assign n16167 = n2156 & ~n6946 ;
  assign n16168 = n12028 & n16167 ;
  assign n16169 = n7971 ^ n3786 ^ 1'b0 ;
  assign n16170 = n4616 & ~n16169 ;
  assign n16171 = ( ~n16166 & n16168 ) | ( ~n16166 & n16170 ) | ( n16168 & n16170 ) ;
  assign n16172 = n5556 ^ n795 ^ 1'b0 ;
  assign n16173 = ~n3418 & n9393 ;
  assign n16174 = n16173 ^ n14006 ^ 1'b0 ;
  assign n16175 = ( ~n1181 & n7388 ) | ( ~n1181 & n16174 ) | ( n7388 & n16174 ) ;
  assign n16176 = n16175 ^ n12019 ^ 1'b0 ;
  assign n16177 = n16172 | n16176 ;
  assign n16178 = n16171 & ~n16177 ;
  assign n16179 = n7983 ^ n287 ^ 1'b0 ;
  assign n16180 = n12961 & n16179 ;
  assign n16181 = ( ~n4599 & n5856 ) | ( ~n4599 & n16180 ) | ( n5856 & n16180 ) ;
  assign n16182 = n9790 & n16181 ;
  assign n16183 = n14621 & n16182 ;
  assign n16185 = n9603 ^ x243 ^ 1'b0 ;
  assign n16186 = n11007 & n16185 ;
  assign n16184 = ( n1860 & ~n4139 ) | ( n1860 & n10101 ) | ( ~n4139 & n10101 ) ;
  assign n16187 = n16186 ^ n16184 ^ n2317 ;
  assign n16188 = n16187 ^ n5847 ^ 1'b0 ;
  assign n16189 = n6328 & ~n16188 ;
  assign n16190 = n10722 & n16189 ;
  assign n16191 = n11526 | n14943 ;
  assign n16192 = n6658 | n11172 ;
  assign n16193 = n9591 & ~n16192 ;
  assign n16194 = ( n10220 & n15836 ) | ( n10220 & n16193 ) | ( n15836 & n16193 ) ;
  assign n16195 = n16194 ^ n5420 ^ 1'b0 ;
  assign n16196 = n15921 | n16195 ;
  assign n16197 = n2774 ^ n2268 ^ 1'b0 ;
  assign n16198 = n6839 & n16197 ;
  assign n16199 = n930 | n16198 ;
  assign n16200 = n16199 ^ n958 ^ 1'b0 ;
  assign n16201 = n8703 & ~n16200 ;
  assign n16202 = ( n5313 & n8552 ) | ( n5313 & ~n16201 ) | ( n8552 & ~n16201 ) ;
  assign n16203 = n10060 ^ n9812 ^ n7747 ;
  assign n16204 = n16203 ^ n10090 ^ n7808 ;
  assign n16205 = ~n963 & n8932 ;
  assign n16206 = n16205 ^ n961 ^ 1'b0 ;
  assign n16207 = ( n8023 & ~n11630 ) | ( n8023 & n16206 ) | ( ~n11630 & n16206 ) ;
  assign n16208 = x123 & ~n15438 ;
  assign n16209 = ( ~n4192 & n4658 ) | ( ~n4192 & n8365 ) | ( n4658 & n8365 ) ;
  assign n16210 = n16209 ^ n1227 ^ x241 ;
  assign n16211 = ( n15499 & n16208 ) | ( n15499 & ~n16210 ) | ( n16208 & ~n16210 ) ;
  assign n16212 = n3084 & n7317 ;
  assign n16213 = n16212 ^ n8965 ^ n1713 ;
  assign n16214 = ( n16207 & n16211 ) | ( n16207 & ~n16213 ) | ( n16211 & ~n16213 ) ;
  assign n16215 = n15123 ^ n6420 ^ 1'b0 ;
  assign n16216 = n5965 ^ n5410 ^ n682 ;
  assign n16217 = ( n9766 & n12321 ) | ( n9766 & n16216 ) | ( n12321 & n16216 ) ;
  assign n16218 = n10954 ^ n4657 ^ n1433 ;
  assign n16219 = ( n667 & n5765 ) | ( n667 & n16218 ) | ( n5765 & n16218 ) ;
  assign n16220 = n831 & ~n16219 ;
  assign n16221 = n8456 ^ n4787 ^ 1'b0 ;
  assign n16222 = n16220 | n16221 ;
  assign n16223 = n15633 ^ n3418 ^ n1747 ;
  assign n16224 = n12973 & ~n13198 ;
  assign n16225 = n626 & n16224 ;
  assign n16226 = ( n10041 & n11894 ) | ( n10041 & ~n16225 ) | ( n11894 & ~n16225 ) ;
  assign n16228 = n5173 ^ n2945 ^ n2157 ;
  assign n16227 = n5286 ^ n2455 ^ 1'b0 ;
  assign n16229 = n16228 ^ n16227 ^ n9412 ;
  assign n16230 = ~x246 & n4165 ;
  assign n16231 = n16230 ^ n13986 ^ n10370 ;
  assign n16232 = n10824 ^ n7835 ^ n1873 ;
  assign n16233 = n15310 ^ n10248 ^ n2894 ;
  assign n16234 = ( ~n8560 & n9073 ) | ( ~n8560 & n16233 ) | ( n9073 & n16233 ) ;
  assign n16235 = n14150 ^ n4048 ^ 1'b0 ;
  assign n16236 = ( n6762 & n6767 ) | ( n6762 & ~n12722 ) | ( n6767 & ~n12722 ) ;
  assign n16238 = n6184 & ~n8885 ;
  assign n16237 = ( ~n4640 & n8762 ) | ( ~n4640 & n13989 ) | ( n8762 & n13989 ) ;
  assign n16239 = n16238 ^ n16237 ^ n7828 ;
  assign n16240 = ( x202 & n5251 ) | ( x202 & n6171 ) | ( n5251 & n6171 ) ;
  assign n16241 = ( n4168 & n10733 ) | ( n4168 & n16240 ) | ( n10733 & n16240 ) ;
  assign n16242 = n3727 & n4310 ;
  assign n16243 = ( n922 & n16241 ) | ( n922 & n16242 ) | ( n16241 & n16242 ) ;
  assign n16244 = ~n13795 & n15259 ;
  assign n16245 = n16244 ^ n1491 ^ 1'b0 ;
  assign n16246 = n9571 & ~n14765 ;
  assign n16247 = ( n1096 & n4786 ) | ( n1096 & n11668 ) | ( n4786 & n11668 ) ;
  assign n16248 = n8574 & ~n11682 ;
  assign n16249 = ( n9076 & ~n14868 ) | ( n9076 & n16248 ) | ( ~n14868 & n16248 ) ;
  assign n16252 = n2110 & n6501 ;
  assign n16253 = n16252 ^ n15767 ^ n4792 ;
  assign n16254 = ( ~n2345 & n7649 ) | ( ~n2345 & n11577 ) | ( n7649 & n11577 ) ;
  assign n16255 = ( ~n286 & n16253 ) | ( ~n286 & n16254 ) | ( n16253 & n16254 ) ;
  assign n16256 = n16255 ^ n7103 ^ 1'b0 ;
  assign n16257 = n16027 & n16256 ;
  assign n16250 = n8617 ^ n6039 ^ n5411 ;
  assign n16251 = n16250 ^ n8128 ^ n2632 ;
  assign n16258 = n16257 ^ n16251 ^ 1'b0 ;
  assign n16259 = n16258 ^ n5633 ^ n4467 ;
  assign n16260 = n5943 | n14161 ;
  assign n16261 = ( n9008 & n14096 ) | ( n9008 & n16260 ) | ( n14096 & n16260 ) ;
  assign n16266 = n3617 | n5387 ;
  assign n16264 = n278 & ~n9949 ;
  assign n16265 = n14631 & n16264 ;
  assign n16267 = n16266 ^ n16265 ^ n4311 ;
  assign n16268 = ( n7349 & ~n12272 ) | ( n7349 & n16267 ) | ( ~n12272 & n16267 ) ;
  assign n16262 = n2661 | n4413 ;
  assign n16263 = n16262 ^ n326 ^ 1'b0 ;
  assign n16269 = n16268 ^ n16263 ^ 1'b0 ;
  assign n16270 = n16261 & ~n16269 ;
  assign n16271 = n14946 ^ n1387 ^ 1'b0 ;
  assign n16272 = n6388 | n16271 ;
  assign n16274 = ( x76 & n3538 ) | ( x76 & ~n9974 ) | ( n3538 & ~n9974 ) ;
  assign n16275 = n16274 ^ n11075 ^ n4942 ;
  assign n16273 = ( n4029 & n6845 ) | ( n4029 & ~n11153 ) | ( n6845 & ~n11153 ) ;
  assign n16276 = n16275 ^ n16273 ^ 1'b0 ;
  assign n16277 = ~n16272 & n16276 ;
  assign n16281 = n9763 & n13545 ;
  assign n16278 = n1753 & ~n4774 ;
  assign n16279 = n16278 ^ n6912 ^ 1'b0 ;
  assign n16280 = n6672 | n16279 ;
  assign n16282 = n16281 ^ n16280 ^ n12286 ;
  assign n16283 = n9626 | n11985 ;
  assign n16284 = n8117 ^ n5707 ^ x178 ;
  assign n16285 = ~n5743 & n16284 ;
  assign n16286 = n16283 & n16285 ;
  assign n16287 = ~n2450 & n3361 ;
  assign n16288 = ( ~n1735 & n9538 ) | ( ~n1735 & n10702 ) | ( n9538 & n10702 ) ;
  assign n16289 = n16288 ^ n9879 ^ n4449 ;
  assign n16290 = ( n6454 & n16287 ) | ( n6454 & ~n16289 ) | ( n16287 & ~n16289 ) ;
  assign n16291 = n9109 | n11100 ;
  assign n16292 = n15976 ^ n12247 ^ 1'b0 ;
  assign n16293 = n5976 ^ n3270 ^ x244 ;
  assign n16294 = n12247 ^ n8955 ^ n5621 ;
  assign n16295 = n16293 & n16294 ;
  assign n16296 = n16295 ^ n2290 ^ 1'b0 ;
  assign n16297 = ( n1490 & ~n4679 ) | ( n1490 & n5913 ) | ( ~n4679 & n5913 ) ;
  assign n16298 = ( n777 & n16296 ) | ( n777 & ~n16297 ) | ( n16296 & ~n16297 ) ;
  assign n16299 = n3065 | n3789 ;
  assign n16300 = n16299 ^ n4831 ^ 1'b0 ;
  assign n16301 = ( ~n4687 & n7849 ) | ( ~n4687 & n16300 ) | ( n7849 & n16300 ) ;
  assign n16302 = n10545 ^ n8951 ^ 1'b0 ;
  assign n16303 = n6691 ^ n1573 ^ 1'b0 ;
  assign n16304 = n12666 ^ n6855 ^ n4744 ;
  assign n16305 = n7850 ^ n1894 ^ 1'b0 ;
  assign n16306 = n13782 & ~n16305 ;
  assign n16307 = ( n9969 & ~n11969 ) | ( n9969 & n15327 ) | ( ~n11969 & n15327 ) ;
  assign n16308 = n4330 ^ n2222 ^ 1'b0 ;
  assign n16309 = n10927 & ~n16308 ;
  assign n16310 = n4424 & ~n13545 ;
  assign n16314 = n13892 ^ n5209 ^ n2146 ;
  assign n16311 = ~n9671 & n15424 ;
  assign n16312 = n8173 & n16311 ;
  assign n16313 = n16312 ^ n10372 ^ n7245 ;
  assign n16315 = n16314 ^ n16313 ^ 1'b0 ;
  assign n16316 = ~n11318 & n16315 ;
  assign n16317 = n16316 ^ n9113 ^ 1'b0 ;
  assign n16318 = n16310 & ~n16317 ;
  assign n16319 = ( ~n1452 & n16309 ) | ( ~n1452 & n16318 ) | ( n16309 & n16318 ) ;
  assign n16320 = n12335 ^ n5492 ^ 1'b0 ;
  assign n16321 = n11689 | n16320 ;
  assign n16322 = n2432 | n16321 ;
  assign n16323 = n16322 ^ n5520 ^ 1'b0 ;
  assign n16325 = ( ~n6304 & n7547 ) | ( ~n6304 & n8119 ) | ( n7547 & n8119 ) ;
  assign n16324 = n7992 & n9008 ;
  assign n16326 = n16325 ^ n16324 ^ 1'b0 ;
  assign n16327 = ( n3433 & n11143 ) | ( n3433 & n16326 ) | ( n11143 & n16326 ) ;
  assign n16328 = ~n6538 & n10093 ;
  assign n16329 = n3015 & n16328 ;
  assign n16330 = ~n7440 & n14926 ;
  assign n16331 = n16330 ^ n7192 ^ 1'b0 ;
  assign n16332 = n11493 ^ n7012 ^ n6742 ;
  assign n16333 = n16332 ^ n4812 ^ 1'b0 ;
  assign n16334 = x134 & ~n16333 ;
  assign n16335 = ~n16331 & n16334 ;
  assign n16338 = ( n2127 & n9244 ) | ( n2127 & ~n15384 ) | ( n9244 & ~n15384 ) ;
  assign n16337 = ~n773 & n5625 ;
  assign n16336 = ( ~n5897 & n6723 ) | ( ~n5897 & n10669 ) | ( n6723 & n10669 ) ;
  assign n16339 = n16338 ^ n16337 ^ n16336 ;
  assign n16340 = ( n2017 & ~n16335 ) | ( n2017 & n16339 ) | ( ~n16335 & n16339 ) ;
  assign n16341 = n12006 ^ n3164 ^ 1'b0 ;
  assign n16342 = n1447 & n16341 ;
  assign n16343 = n619 & n10500 ;
  assign n16345 = n2823 ^ n2452 ^ n1793 ;
  assign n16344 = ( n2572 & n6703 ) | ( n2572 & ~n7692 ) | ( n6703 & ~n7692 ) ;
  assign n16346 = n16345 ^ n16344 ^ 1'b0 ;
  assign n16347 = n3439 | n16346 ;
  assign n16348 = ( n1826 & ~n2209 ) | ( n1826 & n2760 ) | ( ~n2209 & n2760 ) ;
  assign n16349 = ( n9105 & n14535 ) | ( n9105 & n16348 ) | ( n14535 & n16348 ) ;
  assign n16350 = n16349 ^ n15583 ^ n9999 ;
  assign n16351 = n340 & n10391 ;
  assign n16352 = ~n11306 & n16351 ;
  assign n16353 = n16352 ^ x216 ^ 1'b0 ;
  assign n16354 = n9489 ^ n3615 ^ n343 ;
  assign n16355 = n3870 ^ n474 ^ 1'b0 ;
  assign n16356 = n16355 ^ n15311 ^ 1'b0 ;
  assign n16357 = ( x89 & ~n16354 ) | ( x89 & n16356 ) | ( ~n16354 & n16356 ) ;
  assign n16359 = ( n400 & ~n2168 ) | ( n400 & n3912 ) | ( ~n2168 & n3912 ) ;
  assign n16358 = n9601 ^ n3620 ^ n3613 ;
  assign n16360 = n16359 ^ n16358 ^ n1497 ;
  assign n16361 = ~n5609 & n16360 ;
  assign n16362 = ~n4379 & n16361 ;
  assign n16363 = n16362 ^ n2749 ^ 1'b0 ;
  assign n16364 = n8102 & n16363 ;
  assign n16365 = ( n925 & n6910 ) | ( n925 & ~n16364 ) | ( n6910 & ~n16364 ) ;
  assign n16366 = ( n5403 & ~n15594 ) | ( n5403 & n16365 ) | ( ~n15594 & n16365 ) ;
  assign n16371 = ( ~n999 & n3424 ) | ( ~n999 & n14145 ) | ( n3424 & n14145 ) ;
  assign n16372 = n16371 ^ n2143 ^ 1'b0 ;
  assign n16373 = ( n2382 & n7401 ) | ( n2382 & n16372 ) | ( n7401 & n16372 ) ;
  assign n16368 = ~n4694 & n12559 ;
  assign n16367 = n5468 ^ n2910 ^ n2290 ;
  assign n16369 = n16368 ^ n16367 ^ 1'b0 ;
  assign n16370 = n6715 & n16369 ;
  assign n16374 = n16373 ^ n16370 ^ 1'b0 ;
  assign n16375 = n4285 & ~n16374 ;
  assign n16376 = ~n3835 & n6437 ;
  assign n16377 = ~n4112 & n16376 ;
  assign n16378 = n16377 ^ n6458 ^ 1'b0 ;
  assign n16382 = ~n7715 & n12985 ;
  assign n16379 = n12806 ^ n8023 ^ n3361 ;
  assign n16380 = n16379 ^ n8817 ^ n5663 ;
  assign n16381 = ( n5616 & n12067 ) | ( n5616 & n16380 ) | ( n12067 & n16380 ) ;
  assign n16383 = n16382 ^ n16381 ^ n5564 ;
  assign n16384 = ( ~n394 & n16378 ) | ( ~n394 & n16383 ) | ( n16378 & n16383 ) ;
  assign n16392 = n1467 | n1873 ;
  assign n16393 = n16392 ^ n2573 ^ 1'b0 ;
  assign n16394 = n1658 | n2523 ;
  assign n16395 = n16393 | n16394 ;
  assign n16396 = n16395 ^ n15024 ^ 1'b0 ;
  assign n16397 = ~n1720 & n16396 ;
  assign n16398 = n9514 ^ n3506 ^ n1582 ;
  assign n16399 = n16397 & n16398 ;
  assign n16400 = n4998 & n16399 ;
  assign n16401 = n16400 ^ n12036 ^ n10762 ;
  assign n16388 = n6081 ^ n2527 ^ 1'b0 ;
  assign n16389 = n4983 & ~n16388 ;
  assign n16390 = n16389 ^ n12050 ^ n4003 ;
  assign n16391 = ( ~n4068 & n4906 ) | ( ~n4068 & n16390 ) | ( n4906 & n16390 ) ;
  assign n16385 = n10492 ^ n8939 ^ n928 ;
  assign n16386 = n3108 & n16385 ;
  assign n16387 = n16386 ^ n1645 ^ 1'b0 ;
  assign n16402 = n16401 ^ n16391 ^ n16387 ;
  assign n16403 = n16402 ^ n3828 ^ n2362 ;
  assign n16405 = n8313 ^ n1066 ^ x128 ;
  assign n16404 = ( n3090 & ~n6976 ) | ( n3090 & n11422 ) | ( ~n6976 & n11422 ) ;
  assign n16406 = n16405 ^ n16404 ^ n556 ;
  assign n16408 = n3034 & ~n6430 ;
  assign n16407 = ~n6895 & n10917 ;
  assign n16409 = n16408 ^ n16407 ^ 1'b0 ;
  assign n16410 = x208 & ~n2963 ;
  assign n16411 = ( n3137 & n12429 ) | ( n3137 & ~n12579 ) | ( n12429 & ~n12579 ) ;
  assign n16412 = n16159 | n16411 ;
  assign n16422 = ( n583 & n1730 ) | ( n583 & ~n5771 ) | ( n1730 & ~n5771 ) ;
  assign n16419 = n1340 & n1977 ;
  assign n16420 = n1898 & n16419 ;
  assign n16418 = ( n1365 & n4279 ) | ( n1365 & ~n8901 ) | ( n4279 & ~n8901 ) ;
  assign n16421 = n16420 ^ n16418 ^ n15102 ;
  assign n16416 = n2324 & ~n4657 ;
  assign n16413 = n8456 & n11373 ;
  assign n16414 = n9451 ^ n3789 ^ 1'b0 ;
  assign n16415 = ( n15845 & n16413 ) | ( n15845 & n16414 ) | ( n16413 & n16414 ) ;
  assign n16417 = n16416 ^ n16415 ^ n9919 ;
  assign n16423 = n16422 ^ n16421 ^ n16417 ;
  assign n16426 = n1661 & n3298 ;
  assign n16424 = n15540 ^ n12554 ^ n12063 ;
  assign n16425 = n16424 ^ n14668 ^ 1'b0 ;
  assign n16427 = n16426 ^ n16425 ^ n8432 ;
  assign n16428 = n16427 ^ n1287 ^ 1'b0 ;
  assign n16429 = n8094 & n16428 ;
  assign n16430 = ( n1548 & ~n6598 ) | ( n1548 & n9151 ) | ( ~n6598 & n9151 ) ;
  assign n16435 = n6114 ^ n4515 ^ n3846 ;
  assign n16436 = n16435 ^ n11071 ^ 1'b0 ;
  assign n16437 = n16436 ^ n7346 ^ 1'b0 ;
  assign n16433 = ( n6246 & n7347 ) | ( n6246 & n11673 ) | ( n7347 & n11673 ) ;
  assign n16432 = ( n511 & ~n5597 ) | ( n511 & n7754 ) | ( ~n5597 & n7754 ) ;
  assign n16434 = n16433 ^ n16432 ^ n13116 ;
  assign n16431 = n11167 & ~n12624 ;
  assign n16438 = n16437 ^ n16434 ^ n16431 ;
  assign n16439 = ( n2550 & ~n11912 ) | ( n2550 & n12570 ) | ( ~n11912 & n12570 ) ;
  assign n16440 = ( ~n456 & n8462 ) | ( ~n456 & n16439 ) | ( n8462 & n16439 ) ;
  assign n16446 = n487 & n5480 ;
  assign n16447 = n7768 ^ n5847 ^ n699 ;
  assign n16448 = ( n7601 & ~n16446 ) | ( n7601 & n16447 ) | ( ~n16446 & n16447 ) ;
  assign n16441 = ( n429 & n7691 ) | ( n429 & ~n10349 ) | ( n7691 & ~n10349 ) ;
  assign n16442 = n16441 ^ n4557 ^ 1'b0 ;
  assign n16443 = ~n11615 & n16442 ;
  assign n16444 = n6558 & ~n8111 ;
  assign n16445 = ( ~n1808 & n16443 ) | ( ~n1808 & n16444 ) | ( n16443 & n16444 ) ;
  assign n16449 = n16448 ^ n16445 ^ n4752 ;
  assign n16450 = n1224 & n7927 ;
  assign n16451 = n4202 & n6208 ;
  assign n16452 = n16451 ^ n8468 ^ n891 ;
  assign n16453 = n11383 ^ n3613 ^ 1'b0 ;
  assign n16454 = ( n550 & ~n5576 ) | ( n550 & n5796 ) | ( ~n5576 & n5796 ) ;
  assign n16455 = ( n3031 & n10617 ) | ( n3031 & n16454 ) | ( n10617 & n16454 ) ;
  assign n16456 = n5930 ^ n3065 ^ 1'b0 ;
  assign n16457 = n4166 & n7536 ;
  assign n16458 = ~n9626 & n16457 ;
  assign n16459 = n16456 & n16458 ;
  assign n16460 = ( n16453 & ~n16455 ) | ( n16453 & n16459 ) | ( ~n16455 & n16459 ) ;
  assign n16461 = n11895 ^ x61 ^ 1'b0 ;
  assign n16462 = n14332 & n16461 ;
  assign n16463 = n16462 ^ n1202 ^ n724 ;
  assign n16465 = ( ~n6474 & n12889 ) | ( ~n6474 & n14879 ) | ( n12889 & n14879 ) ;
  assign n16464 = n11175 & ~n12801 ;
  assign n16466 = n16465 ^ n16464 ^ 1'b0 ;
  assign n16467 = n7937 & ~n9983 ;
  assign n16468 = ( n5182 & n9442 ) | ( n5182 & ~n16467 ) | ( n9442 & ~n16467 ) ;
  assign n16471 = ~n2034 & n10875 ;
  assign n16469 = x191 & ~n3974 ;
  assign n16470 = n10841 & n16469 ;
  assign n16472 = n16471 ^ n16470 ^ 1'b0 ;
  assign n16476 = ( ~n4709 & n6038 ) | ( ~n4709 & n16227 ) | ( n6038 & n16227 ) ;
  assign n16473 = n2997 & ~n4269 ;
  assign n16474 = ~n1605 & n16473 ;
  assign n16475 = n7661 | n16474 ;
  assign n16477 = n16476 ^ n16475 ^ 1'b0 ;
  assign n16478 = n5051 ^ n1152 ^ 1'b0 ;
  assign n16479 = n5696 & n16478 ;
  assign n16480 = ( n3408 & n13434 ) | ( n3408 & n16479 ) | ( n13434 & n16479 ) ;
  assign n16481 = ( ~n2697 & n5255 ) | ( ~n2697 & n7328 ) | ( n5255 & n7328 ) ;
  assign n16482 = ( ~n2580 & n16480 ) | ( ~n2580 & n16481 ) | ( n16480 & n16481 ) ;
  assign n16483 = n3495 ^ n2245 ^ n1604 ;
  assign n16484 = n4503 | n16483 ;
  assign n16485 = n16484 ^ n11017 ^ 1'b0 ;
  assign n16486 = n16485 ^ n10461 ^ x164 ;
  assign n16487 = ( ~x57 & n5664 ) | ( ~x57 & n16486 ) | ( n5664 & n16486 ) ;
  assign n16488 = n16487 ^ n1957 ^ 1'b0 ;
  assign n16489 = ~n16482 & n16488 ;
  assign n16490 = ( n3797 & ~n14277 ) | ( n3797 & n16489 ) | ( ~n14277 & n16489 ) ;
  assign n16491 = ~n7905 & n16490 ;
  assign n16492 = n6210 ^ n5194 ^ n5028 ;
  assign n16493 = n6015 ^ n4728 ^ n2363 ;
  assign n16494 = n7605 ^ n6331 ^ n1466 ;
  assign n16495 = ( n7630 & ~n16493 ) | ( n7630 & n16494 ) | ( ~n16493 & n16494 ) ;
  assign n16496 = n16495 ^ n10877 ^ 1'b0 ;
  assign n16497 = n8852 | n16496 ;
  assign n16498 = x93 & ~n7171 ;
  assign n16499 = ~n9195 & n16498 ;
  assign n16500 = ( n3180 & ~n6769 ) | ( n3180 & n16499 ) | ( ~n6769 & n16499 ) ;
  assign n16501 = ( n16492 & ~n16497 ) | ( n16492 & n16500 ) | ( ~n16497 & n16500 ) ;
  assign n16502 = n16501 ^ n4319 ^ n3646 ;
  assign n16503 = n3030 | n3359 ;
  assign n16504 = n13407 ^ n8846 ^ n4563 ;
  assign n16505 = n4946 | n16504 ;
  assign n16506 = n7331 ^ x111 ^ 1'b0 ;
  assign n16507 = ( n2239 & n15827 ) | ( n2239 & n16506 ) | ( n15827 & n16506 ) ;
  assign n16508 = n16507 ^ n9340 ^ n3245 ;
  assign n16509 = ( n6195 & n16505 ) | ( n6195 & ~n16508 ) | ( n16505 & ~n16508 ) ;
  assign n16510 = ( n2766 & ~n16503 ) | ( n2766 & n16509 ) | ( ~n16503 & n16509 ) ;
  assign n16511 = n7570 ^ x25 ^ 1'b0 ;
  assign n16512 = ( n10655 & ~n14023 ) | ( n10655 & n16511 ) | ( ~n14023 & n16511 ) ;
  assign n16522 = n8474 ^ n2795 ^ 1'b0 ;
  assign n16523 = n16522 ^ n9788 ^ n9646 ;
  assign n16524 = n16523 ^ n8024 ^ 1'b0 ;
  assign n16515 = ( ~x71 & n3178 ) | ( ~x71 & n3936 ) | ( n3178 & n3936 ) ;
  assign n16516 = n4933 & ~n16515 ;
  assign n16517 = n16516 ^ n6257 ^ 1'b0 ;
  assign n16518 = n3685 & ~n12158 ;
  assign n16519 = n16518 ^ n14152 ^ n6018 ;
  assign n16520 = ( ~n9818 & n16517 ) | ( ~n9818 & n16519 ) | ( n16517 & n16519 ) ;
  assign n16521 = n16520 ^ n10700 ^ 1'b0 ;
  assign n16513 = n14302 ^ n8676 ^ n6437 ;
  assign n16514 = n16513 ^ n10135 ^ n8088 ;
  assign n16525 = n16524 ^ n16521 ^ n16514 ;
  assign n16526 = n9150 ^ n6605 ^ n4997 ;
  assign n16527 = n1438 & n1474 ;
  assign n16528 = ( x139 & n16526 ) | ( x139 & n16527 ) | ( n16526 & n16527 ) ;
  assign n16529 = n16528 ^ n1358 ^ 1'b0 ;
  assign n16530 = ( x240 & n1886 ) | ( x240 & n4598 ) | ( n1886 & n4598 ) ;
  assign n16531 = n8180 ^ n3907 ^ n489 ;
  assign n16532 = n16531 ^ n11411 ^ n7684 ;
  assign n16533 = n9439 & n16532 ;
  assign n16538 = ( n5033 & n5739 ) | ( n5033 & n10657 ) | ( n5739 & n10657 ) ;
  assign n16534 = ( ~n1407 & n4499 ) | ( ~n1407 & n6314 ) | ( n4499 & n6314 ) ;
  assign n16535 = ( n594 & ~n4494 ) | ( n594 & n16534 ) | ( ~n4494 & n16534 ) ;
  assign n16536 = n16535 ^ n7984 ^ 1'b0 ;
  assign n16537 = n12485 & n16536 ;
  assign n16539 = n16538 ^ n16537 ^ 1'b0 ;
  assign n16540 = n16539 ^ n8961 ^ n5923 ;
  assign n16541 = ( n16530 & ~n16533 ) | ( n16530 & n16540 ) | ( ~n16533 & n16540 ) ;
  assign n16542 = ( n5176 & n10690 ) | ( n5176 & ~n11238 ) | ( n10690 & ~n11238 ) ;
  assign n16543 = n16542 ^ n5327 ^ 1'b0 ;
  assign n16544 = n1412 | n4808 ;
  assign n16545 = n16544 ^ n605 ^ 1'b0 ;
  assign n16546 = ~n12146 & n16545 ;
  assign n16547 = n5787 ^ n5382 ^ n2011 ;
  assign n16548 = ( n7479 & ~n16546 ) | ( n7479 & n16547 ) | ( ~n16546 & n16547 ) ;
  assign n16549 = n5360 ^ n3901 ^ 1'b0 ;
  assign n16550 = n16548 | n16549 ;
  assign n16551 = ( x129 & n3358 ) | ( x129 & ~n3719 ) | ( n3358 & ~n3719 ) ;
  assign n16552 = n16551 ^ n14504 ^ n11493 ;
  assign n16553 = n4880 & n16552 ;
  assign n16554 = n16553 ^ n3646 ^ 1'b0 ;
  assign n16555 = n16550 & n16554 ;
  assign n16559 = n6167 ^ n3756 ^ 1'b0 ;
  assign n16558 = n5665 & ~n7480 ;
  assign n16560 = n16559 ^ n16558 ^ 1'b0 ;
  assign n16561 = n5050 | n16560 ;
  assign n16556 = n11004 ^ n9878 ^ n7839 ;
  assign n16557 = n16556 ^ n3681 ^ 1'b0 ;
  assign n16562 = n16561 ^ n16557 ^ n13940 ;
  assign n16563 = n13675 ^ n4591 ^ n3251 ;
  assign n16564 = ( n1356 & n6874 ) | ( n1356 & ~n9276 ) | ( n6874 & ~n9276 ) ;
  assign n16565 = n16564 ^ n7995 ^ n2414 ;
  assign n16566 = n752 | n6649 ;
  assign n16567 = n16565 & ~n16566 ;
  assign n16571 = n3971 ^ n1784 ^ n1754 ;
  assign n16572 = ~n7290 & n16571 ;
  assign n16573 = n5884 & n16572 ;
  assign n16568 = n5582 ^ n2161 ^ 1'b0 ;
  assign n16569 = n7024 ^ n1419 ^ 1'b0 ;
  assign n16570 = n16568 & n16569 ;
  assign n16574 = n16573 ^ n16570 ^ 1'b0 ;
  assign n16575 = n16567 & n16574 ;
  assign n16576 = n7247 & ~n10797 ;
  assign n16577 = n16576 ^ n2067 ^ 1'b0 ;
  assign n16578 = ( ~n752 & n4102 ) | ( ~n752 & n16565 ) | ( n4102 & n16565 ) ;
  assign n16579 = n16577 & ~n16578 ;
  assign n16580 = n16579 ^ n4949 ^ 1'b0 ;
  assign n16586 = ( n2151 & n6899 ) | ( n2151 & n9640 ) | ( n6899 & n9640 ) ;
  assign n16585 = n9391 ^ n7378 ^ 1'b0 ;
  assign n16581 = n16111 ^ n2053 ^ n520 ;
  assign n16582 = ( ~n1156 & n6871 ) | ( ~n1156 & n8743 ) | ( n6871 & n8743 ) ;
  assign n16583 = n9283 & n16582 ;
  assign n16584 = ~n16581 & n16583 ;
  assign n16587 = n16586 ^ n16585 ^ n16584 ;
  assign n16588 = n6188 ^ n3225 ^ n395 ;
  assign n16589 = n16588 ^ n2881 ^ n1935 ;
  assign n16590 = n1395 | n11802 ;
  assign n16591 = ( ~n3896 & n5784 ) | ( ~n3896 & n16590 ) | ( n5784 & n16590 ) ;
  assign n16592 = ( ~n2435 & n4466 ) | ( ~n2435 & n9398 ) | ( n4466 & n9398 ) ;
  assign n16597 = ( n1849 & n6403 ) | ( n1849 & ~n12488 ) | ( n6403 & ~n12488 ) ;
  assign n16593 = ( n4529 & ~n6635 ) | ( n4529 & n6943 ) | ( ~n6635 & n6943 ) ;
  assign n16594 = n10349 ^ n6802 ^ n6546 ;
  assign n16595 = ( ~n704 & n2883 ) | ( ~n704 & n16594 ) | ( n2883 & n16594 ) ;
  assign n16596 = n16593 | n16595 ;
  assign n16598 = n16597 ^ n16596 ^ 1'b0 ;
  assign n16599 = n16598 ^ n11410 ^ 1'b0 ;
  assign n16600 = n10091 ^ n1549 ^ n1444 ;
  assign n16601 = ~n11323 & n16600 ;
  assign n16602 = n9480 ^ n4539 ^ 1'b0 ;
  assign n16603 = ~n2355 & n16602 ;
  assign n16604 = ( n9934 & ~n10188 ) | ( n9934 & n16603 ) | ( ~n10188 & n16603 ) ;
  assign n16605 = ( n2765 & n16601 ) | ( n2765 & ~n16604 ) | ( n16601 & ~n16604 ) ;
  assign n16606 = n8692 & ~n12040 ;
  assign n16607 = n16606 ^ n11629 ^ n1698 ;
  assign n16608 = ( ~x94 & n9224 ) | ( ~x94 & n16607 ) | ( n9224 & n16607 ) ;
  assign n16609 = ( n6907 & n6913 ) | ( n6907 & n16608 ) | ( n6913 & n16608 ) ;
  assign n16610 = ( ~n5219 & n5312 ) | ( ~n5219 & n6829 ) | ( n5312 & n6829 ) ;
  assign n16611 = n16610 ^ n11483 ^ n3068 ;
  assign n16612 = ( n3797 & ~n11231 ) | ( n3797 & n16611 ) | ( ~n11231 & n16611 ) ;
  assign n16613 = n16612 ^ n2107 ^ 1'b0 ;
  assign n16614 = n8250 & ~n16613 ;
  assign n16615 = n13858 ^ n4168 ^ n1058 ;
  assign n16616 = ( n15049 & ~n16178 ) | ( n15049 & n16615 ) | ( ~n16178 & n16615 ) ;
  assign n16617 = n6481 ^ n2130 ^ x64 ;
  assign n16618 = ( ~n11428 & n13654 ) | ( ~n11428 & n15595 ) | ( n13654 & n15595 ) ;
  assign n16619 = ~n3504 & n11943 ;
  assign n16620 = n16618 & n16619 ;
  assign n16621 = n4560 ^ n693 ^ 1'b0 ;
  assign n16624 = ~n7227 & n8112 ;
  assign n16622 = n8727 ^ n542 ^ 1'b0 ;
  assign n16623 = n12626 | n16622 ;
  assign n16625 = n16624 ^ n16623 ^ n15054 ;
  assign n16626 = ( n10056 & n16621 ) | ( n10056 & n16625 ) | ( n16621 & n16625 ) ;
  assign n16630 = ( ~n312 & n540 ) | ( ~n312 & n10101 ) | ( n540 & n10101 ) ;
  assign n16628 = n1879 | n3953 ;
  assign n16629 = n12762 & ~n16628 ;
  assign n16631 = n16630 ^ n16629 ^ 1'b0 ;
  assign n16632 = n16631 ^ n7794 ^ x11 ;
  assign n16633 = ( n456 & n10999 ) | ( n456 & n16632 ) | ( n10999 & n16632 ) ;
  assign n16634 = n16633 ^ n5201 ^ n1656 ;
  assign n16627 = n8019 | n14325 ;
  assign n16635 = n16634 ^ n16627 ^ 1'b0 ;
  assign n16636 = n1938 & ~n10976 ;
  assign n16637 = n10965 & n16636 ;
  assign n16638 = ( ~n2981 & n4180 ) | ( ~n2981 & n5080 ) | ( n4180 & n5080 ) ;
  assign n16639 = n5359 ^ n1903 ^ 1'b0 ;
  assign n16640 = n16638 & ~n16639 ;
  assign n16643 = n1553 | n6388 ;
  assign n16644 = n16643 ^ n4152 ^ 1'b0 ;
  assign n16641 = n6414 & ~n15408 ;
  assign n16642 = ~n1849 & n16641 ;
  assign n16645 = n16644 ^ n16642 ^ 1'b0 ;
  assign n16646 = ( n368 & n8434 ) | ( n368 & n16645 ) | ( n8434 & n16645 ) ;
  assign n16647 = n16646 ^ n15132 ^ 1'b0 ;
  assign n16648 = n16640 & ~n16647 ;
  assign n16649 = ( n3151 & n4651 ) | ( n3151 & n16648 ) | ( n4651 & n16648 ) ;
  assign n16650 = ( n509 & ~n7569 ) | ( n509 & n10356 ) | ( ~n7569 & n10356 ) ;
  assign n16651 = n2371 & n16650 ;
  assign n16652 = n16651 ^ n971 ^ 1'b0 ;
  assign n16653 = ( ~n4064 & n4704 ) | ( ~n4064 & n16652 ) | ( n4704 & n16652 ) ;
  assign n16654 = n7004 ^ n4025 ^ 1'b0 ;
  assign n16655 = n16654 ^ n16611 ^ n6956 ;
  assign n16656 = ( n4178 & ~n14160 ) | ( n4178 & n16655 ) | ( ~n14160 & n16655 ) ;
  assign n16657 = n14056 ^ n5089 ^ n2019 ;
  assign n16658 = n15359 ^ n3291 ^ 1'b0 ;
  assign n16659 = n3006 & ~n16658 ;
  assign n16660 = n16659 ^ n15470 ^ n6592 ;
  assign n16661 = n16660 ^ n9714 ^ n3092 ;
  assign n16662 = n7411 & ~n12294 ;
  assign n16663 = n16661 & n16662 ;
  assign n16664 = ( ~n1191 & n5706 ) | ( ~n1191 & n15283 ) | ( n5706 & n15283 ) ;
  assign n16668 = n5234 & n5462 ;
  assign n16669 = n16668 ^ n3732 ^ 1'b0 ;
  assign n16670 = n9339 | n16669 ;
  assign n16671 = n11071 | n16670 ;
  assign n16667 = n3127 ^ n1754 ^ n722 ;
  assign n16665 = ~n5033 & n9293 ;
  assign n16666 = ~n1490 & n16665 ;
  assign n16672 = n16671 ^ n16667 ^ n16666 ;
  assign n16673 = ~n693 & n10366 ;
  assign n16674 = ~n4215 & n14827 ;
  assign n16675 = n16674 ^ n2958 ^ 1'b0 ;
  assign n16676 = ( n4216 & ~n9134 ) | ( n4216 & n16675 ) | ( ~n9134 & n16675 ) ;
  assign n16677 = n14271 ^ n14192 ^ n3901 ;
  assign n16679 = n12497 ^ n12300 ^ 1'b0 ;
  assign n16680 = n1827 & ~n16679 ;
  assign n16681 = n13356 ^ n11076 ^ 1'b0 ;
  assign n16682 = n16681 ^ n15071 ^ 1'b0 ;
  assign n16683 = n16680 & ~n16682 ;
  assign n16678 = n14579 ^ n6493 ^ 1'b0 ;
  assign n16684 = n16683 ^ n16678 ^ n6901 ;
  assign n16685 = x190 & ~n15777 ;
  assign n16686 = n16685 ^ n9472 ^ 1'b0 ;
  assign n16687 = ( ~n537 & n1236 ) | ( ~n537 & n15852 ) | ( n1236 & n15852 ) ;
  assign n16688 = ( n5583 & n13145 ) | ( n5583 & n16687 ) | ( n13145 & n16687 ) ;
  assign n16689 = ( n7220 & n15728 ) | ( n7220 & n16688 ) | ( n15728 & n16688 ) ;
  assign n16690 = ( n1882 & n4911 ) | ( n1882 & n16689 ) | ( n4911 & n16689 ) ;
  assign n16691 = n16690 ^ n13149 ^ n8429 ;
  assign n16692 = n4026 ^ n2771 ^ n2068 ;
  assign n16693 = x149 & ~n16692 ;
  assign n16694 = n16693 ^ n4638 ^ 1'b0 ;
  assign n16695 = n15318 ^ n7924 ^ 1'b0 ;
  assign n16696 = n16695 ^ n10108 ^ 1'b0 ;
  assign n16697 = n12985 & ~n16696 ;
  assign n16698 = n2306 & n16697 ;
  assign n16699 = ~n16694 & n16698 ;
  assign n16700 = n10152 ^ n8310 ^ n1733 ;
  assign n16701 = n16700 ^ n4045 ^ 1'b0 ;
  assign n16702 = n16701 ^ n8208 ^ 1'b0 ;
  assign n16703 = n12673 & n14487 ;
  assign n16704 = ~n12124 & n16703 ;
  assign n16705 = n16704 ^ n9646 ^ n2825 ;
  assign n16706 = ( n4003 & n7184 ) | ( n4003 & ~n10783 ) | ( n7184 & ~n10783 ) ;
  assign n16707 = n16706 ^ n2255 ^ 1'b0 ;
  assign n16708 = n13708 ^ n575 ^ 1'b0 ;
  assign n16709 = ~n16707 & n16708 ;
  assign n16710 = n2570 & ~n3779 ;
  assign n16711 = ~n9418 & n16710 ;
  assign n16712 = n16711 ^ n12570 ^ n520 ;
  assign n16713 = ~n9904 & n16712 ;
  assign n16714 = ~n4589 & n16713 ;
  assign n16715 = ~n7586 & n16714 ;
  assign n16716 = n13945 ^ n7025 ^ n1498 ;
  assign n16717 = n12227 ^ n7609 ^ 1'b0 ;
  assign n16718 = n15489 & ~n16717 ;
  assign n16719 = n16181 & ~n16718 ;
  assign n16720 = ~n4126 & n16719 ;
  assign n16721 = ( n8231 & n12381 ) | ( n8231 & ~n16720 ) | ( n12381 & ~n16720 ) ;
  assign n16722 = n2067 | n5968 ;
  assign n16723 = n16722 ^ n16024 ^ n1077 ;
  assign n16724 = n864 & ~n8337 ;
  assign n16725 = n1218 & n16724 ;
  assign n16726 = ( ~n5245 & n6036 ) | ( ~n5245 & n16725 ) | ( n6036 & n16725 ) ;
  assign n16727 = ( n3285 & n3866 ) | ( n3285 & ~n16726 ) | ( n3866 & ~n16726 ) ;
  assign n16730 = n1475 & n4420 ;
  assign n16731 = ~n3333 & n16730 ;
  assign n16732 = n16731 ^ n14437 ^ n13642 ;
  assign n16729 = n14711 ^ n9791 ^ 1'b0 ;
  assign n16728 = n16362 ^ n5438 ^ n2903 ;
  assign n16733 = n16732 ^ n16729 ^ n16728 ;
  assign n16734 = ~n6243 & n14495 ;
  assign n16735 = n16734 ^ n1125 ^ 1'b0 ;
  assign n16736 = ( ~n1698 & n3754 ) | ( ~n1698 & n5990 ) | ( n3754 & n5990 ) ;
  assign n16737 = n16735 & n16736 ;
  assign n16738 = n16737 ^ n12467 ^ 1'b0 ;
  assign n16739 = ( ~n3986 & n6006 ) | ( ~n3986 & n7180 ) | ( n6006 & n7180 ) ;
  assign n16740 = n16739 ^ n7523 ^ 1'b0 ;
  assign n16741 = n8250 & ~n16740 ;
  assign n16742 = n16741 ^ n8691 ^ n1920 ;
  assign n16743 = n4124 | n5418 ;
  assign n16744 = n16742 & ~n16743 ;
  assign n16745 = n16744 ^ n3498 ^ 1'b0 ;
  assign n16746 = n16745 ^ n12462 ^ 1'b0 ;
  assign n16747 = n16746 ^ n15378 ^ n1718 ;
  assign n16748 = n5672 & n13883 ;
  assign n16749 = ( ~n1361 & n1691 ) | ( ~n1361 & n4072 ) | ( n1691 & n4072 ) ;
  assign n16750 = n16749 ^ n9677 ^ n6019 ;
  assign n16751 = ( n5202 & n9016 ) | ( n5202 & n16750 ) | ( n9016 & n16750 ) ;
  assign n16752 = ( n4563 & n16748 ) | ( n4563 & n16751 ) | ( n16748 & n16751 ) ;
  assign n16753 = n16752 ^ n14952 ^ x164 ;
  assign n16754 = n15140 ^ n13139 ^ 1'b0 ;
  assign n16755 = ( ~n13547 & n16753 ) | ( ~n13547 & n16754 ) | ( n16753 & n16754 ) ;
  assign n16762 = ( n3110 & n7228 ) | ( n3110 & n7262 ) | ( n7228 & n7262 ) ;
  assign n16756 = ( n1359 & ~n1736 ) | ( n1359 & n12365 ) | ( ~n1736 & n12365 ) ;
  assign n16758 = n9712 ^ n7312 ^ n3518 ;
  assign n16757 = n1670 & ~n8405 ;
  assign n16759 = n16758 ^ n16757 ^ 1'b0 ;
  assign n16760 = n16759 ^ n16318 ^ n7981 ;
  assign n16761 = n16756 & ~n16760 ;
  assign n16763 = n16762 ^ n16761 ^ 1'b0 ;
  assign n16765 = n3936 & n4642 ;
  assign n16766 = n16765 ^ n12340 ^ 1'b0 ;
  assign n16764 = n7531 & n11747 ;
  assign n16767 = n16766 ^ n16764 ^ n7603 ;
  assign n16776 = ( n555 & n1251 ) | ( n555 & ~n7668 ) | ( n1251 & ~n7668 ) ;
  assign n16777 = n16776 ^ n3322 ^ n355 ;
  assign n16778 = n13971 ^ n1371 ^ n550 ;
  assign n16779 = ( n15396 & n16777 ) | ( n15396 & ~n16778 ) | ( n16777 & ~n16778 ) ;
  assign n16768 = ( n4978 & n5105 ) | ( n4978 & n11030 ) | ( n5105 & n11030 ) ;
  assign n16769 = ( ~n4027 & n4860 ) | ( ~n4027 & n9816 ) | ( n4860 & n9816 ) ;
  assign n16770 = ( n2646 & ~n16768 ) | ( n2646 & n16769 ) | ( ~n16768 & n16769 ) ;
  assign n16771 = n2224 ^ n308 ^ 1'b0 ;
  assign n16772 = ~n11119 & n16771 ;
  assign n16773 = n16772 ^ n1717 ^ 1'b0 ;
  assign n16774 = x122 & n16773 ;
  assign n16775 = ~n16770 & n16774 ;
  assign n16780 = n16779 ^ n16775 ^ 1'b0 ;
  assign n16781 = n8529 | n16780 ;
  assign n16787 = ( n1990 & n5985 ) | ( n1990 & n12285 ) | ( n5985 & n12285 ) ;
  assign n16788 = ( n14532 & ~n14767 ) | ( n14532 & n16787 ) | ( ~n14767 & n16787 ) ;
  assign n16789 = n9465 & ~n16788 ;
  assign n16782 = ( n3669 & ~n6341 ) | ( n3669 & n15321 ) | ( ~n6341 & n15321 ) ;
  assign n16783 = n16782 ^ n13890 ^ 1'b0 ;
  assign n16784 = n4158 | n16783 ;
  assign n16785 = ~x241 & n11815 ;
  assign n16786 = n16784 | n16785 ;
  assign n16790 = n16789 ^ n16786 ^ 1'b0 ;
  assign n16795 = n15868 ^ n3304 ^ n2205 ;
  assign n16796 = ( n6907 & n14031 ) | ( n6907 & ~n16795 ) | ( n14031 & ~n16795 ) ;
  assign n16791 = ( n1753 & ~n3330 ) | ( n1753 & n7270 ) | ( ~n3330 & n7270 ) ;
  assign n16792 = ( n290 & n7337 ) | ( n290 & n16791 ) | ( n7337 & n16791 ) ;
  assign n16793 = n5285 ^ n1448 ^ x37 ;
  assign n16794 = ( n3242 & ~n16792 ) | ( n3242 & n16793 ) | ( ~n16792 & n16793 ) ;
  assign n16797 = n16796 ^ n16794 ^ n11183 ;
  assign n16798 = n8783 & ~n9958 ;
  assign n16799 = ( ~n8918 & n12533 ) | ( ~n8918 & n16798 ) | ( n12533 & n16798 ) ;
  assign n16800 = n511 & ~n13692 ;
  assign n16801 = n7441 & n16800 ;
  assign n16802 = ( x70 & n4636 ) | ( x70 & ~n13207 ) | ( n4636 & ~n13207 ) ;
  assign n16803 = ( n1257 & n16801 ) | ( n1257 & ~n16802 ) | ( n16801 & ~n16802 ) ;
  assign n16804 = ~n1591 & n16803 ;
  assign n16805 = ~n16803 & n16804 ;
  assign n16806 = ( n2003 & n2823 ) | ( n2003 & ~n9273 ) | ( n2823 & ~n9273 ) ;
  assign n16807 = n16806 ^ n10953 ^ n9385 ;
  assign n16808 = n16807 ^ n2070 ^ 1'b0 ;
  assign n16809 = ~n13325 & n16808 ;
  assign n16810 = n14339 ^ n4545 ^ n2113 ;
  assign n16811 = n6944 ^ n326 ^ x65 ;
  assign n16812 = ( ~n14898 & n16810 ) | ( ~n14898 & n16811 ) | ( n16810 & n16811 ) ;
  assign n16813 = n16812 ^ n14370 ^ 1'b0 ;
  assign n16814 = n3061 ^ n853 ^ 1'b0 ;
  assign n16817 = ~n7749 & n12439 ;
  assign n16815 = n1467 | n1705 ;
  assign n16816 = n2522 | n16815 ;
  assign n16818 = n16817 ^ n16816 ^ 1'b0 ;
  assign n16819 = n3107 & n16818 ;
  assign n16820 = n16819 ^ n4352 ^ n2457 ;
  assign n16821 = ( n2101 & ~n7009 ) | ( n2101 & n12308 ) | ( ~n7009 & n12308 ) ;
  assign n16822 = ( ~n5234 & n14055 ) | ( ~n5234 & n15129 ) | ( n14055 & n15129 ) ;
  assign n16823 = n6403 ^ n4804 ^ n4147 ;
  assign n16824 = n4128 | n16823 ;
  assign n16825 = ~n13826 & n14908 ;
  assign n16826 = ( n3428 & n6888 ) | ( n3428 & ~n11833 ) | ( n6888 & ~n11833 ) ;
  assign n16827 = n16826 ^ n3423 ^ 1'b0 ;
  assign n16828 = n16825 | n16827 ;
  assign n16829 = n3161 & ~n5182 ;
  assign n16833 = n6242 ^ n5246 ^ n669 ;
  assign n16832 = n387 & n10664 ;
  assign n16834 = n16833 ^ n16832 ^ 1'b0 ;
  assign n16835 = ( n1974 & ~n9701 ) | ( n1974 & n16834 ) | ( ~n9701 & n16834 ) ;
  assign n16831 = x18 & n5907 ;
  assign n16830 = ~n8156 & n13355 ;
  assign n16836 = n16835 ^ n16831 ^ n16830 ;
  assign n16839 = n8173 ^ n7571 ^ 1'b0 ;
  assign n16837 = n14031 ^ n11205 ^ n6626 ;
  assign n16838 = n10559 | n16837 ;
  assign n16840 = n16839 ^ n16838 ^ n9600 ;
  assign n16841 = ( n1554 & ~n8073 ) | ( n1554 & n8965 ) | ( ~n8073 & n8965 ) ;
  assign n16842 = ( n4631 & n8603 ) | ( n4631 & ~n16841 ) | ( n8603 & ~n16841 ) ;
  assign n16843 = ( n5996 & ~n16840 ) | ( n5996 & n16842 ) | ( ~n16840 & n16842 ) ;
  assign n16846 = n12697 ^ n9335 ^ 1'b0 ;
  assign n16844 = n15742 ^ n11961 ^ 1'b0 ;
  assign n16845 = n10346 & ~n16844 ;
  assign n16847 = n16846 ^ n16845 ^ 1'b0 ;
  assign n16848 = n1406 & n16847 ;
  assign n16849 = n6754 ^ x42 ^ 1'b0 ;
  assign n16850 = n5257 & n16849 ;
  assign n16851 = ( n4396 & ~n7821 ) | ( n4396 & n16850 ) | ( ~n7821 & n16850 ) ;
  assign n16852 = n1014 | n8672 ;
  assign n16853 = n4796 | n16852 ;
  assign n16854 = n10545 ^ n8869 ^ 1'b0 ;
  assign n16855 = n14405 & n16854 ;
  assign n16856 = ( ~n7104 & n9891 ) | ( ~n7104 & n16855 ) | ( n9891 & n16855 ) ;
  assign n16857 = n16853 & n16856 ;
  assign n16858 = n10845 ^ n7994 ^ n2730 ;
  assign n16861 = n14408 ^ n5546 ^ 1'b0 ;
  assign n16862 = n3791 & n16861 ;
  assign n16863 = n16862 ^ n10604 ^ n5757 ;
  assign n16864 = n16863 ^ n11318 ^ n1966 ;
  assign n16859 = n12673 & n16457 ;
  assign n16860 = n16859 ^ n2820 ^ 1'b0 ;
  assign n16865 = n16864 ^ n16860 ^ n7738 ;
  assign n16866 = n8598 ^ n5896 ^ 1'b0 ;
  assign n16867 = ( n1242 & n4417 ) | ( n1242 & n5402 ) | ( n4417 & n5402 ) ;
  assign n16868 = n16866 & n16867 ;
  assign n16869 = ( n6241 & n12351 ) | ( n6241 & ~n14552 ) | ( n12351 & ~n14552 ) ;
  assign n16870 = ~n284 & n7615 ;
  assign n16871 = n16870 ^ n8733 ^ n3350 ;
  assign n16872 = n6340 & ~n10377 ;
  assign n16873 = n16872 ^ n3034 ^ 1'b0 ;
  assign n16874 = n3004 ^ n1476 ^ n1323 ;
  assign n16875 = n16874 ^ n16659 ^ n9683 ;
  assign n16876 = n4448 & n6341 ;
  assign n16877 = n16876 ^ n13116 ^ 1'b0 ;
  assign n16878 = ( ~n5355 & n9353 ) | ( ~n5355 & n16877 ) | ( n9353 & n16877 ) ;
  assign n16879 = ~n4515 & n7160 ;
  assign n16880 = ~n7636 & n16879 ;
  assign n16881 = ( n662 & ~n4148 ) | ( n662 & n12980 ) | ( ~n4148 & n12980 ) ;
  assign n16882 = n16880 | n16881 ;
  assign n16883 = n16652 ^ n15228 ^ 1'b0 ;
  assign n16884 = n8214 | n16883 ;
  assign n16885 = n7371 & ~n16884 ;
  assign n16886 = n13742 ^ n9931 ^ 1'b0 ;
  assign n16887 = ( n8173 & ~n16745 ) | ( n8173 & n16886 ) | ( ~n16745 & n16886 ) ;
  assign n16888 = ( n1926 & n3619 ) | ( n1926 & ~n4263 ) | ( n3619 & ~n4263 ) ;
  assign n16889 = ( n7100 & ~n13536 ) | ( n7100 & n16888 ) | ( ~n13536 & n16888 ) ;
  assign n16890 = ~n2865 & n16889 ;
  assign n16891 = n16890 ^ n4570 ^ 1'b0 ;
  assign n16892 = n16891 ^ n8551 ^ n4318 ;
  assign n16893 = ( n2158 & ~n5399 ) | ( n2158 & n5703 ) | ( ~n5399 & n5703 ) ;
  assign n16894 = n16893 ^ n16527 ^ n3575 ;
  assign n16895 = n5564 | n16894 ;
  assign n16896 = n16892 | n16895 ;
  assign n16897 = ( n1191 & ~n8378 ) | ( n1191 & n16896 ) | ( ~n8378 & n16896 ) ;
  assign n16898 = n14988 ^ n11699 ^ n814 ;
  assign n16899 = n16898 ^ n11563 ^ 1'b0 ;
  assign n16900 = n14467 ^ n12239 ^ n10399 ;
  assign n16901 = n16900 ^ n9444 ^ 1'b0 ;
  assign n16902 = ~n381 & n10001 ;
  assign n16905 = n10109 ^ n4295 ^ n4250 ;
  assign n16903 = n10001 ^ n4496 ^ n2142 ;
  assign n16904 = ( n3952 & n9597 ) | ( n3952 & ~n16903 ) | ( n9597 & ~n16903 ) ;
  assign n16906 = n16905 ^ n16904 ^ 1'b0 ;
  assign n16907 = n12103 ^ n3260 ^ 1'b0 ;
  assign n16908 = ( n5745 & n9395 ) | ( n5745 & n16907 ) | ( n9395 & n16907 ) ;
  assign n16910 = n9099 ^ n5482 ^ 1'b0 ;
  assign n16911 = n13641 & ~n16910 ;
  assign n16909 = n16530 ^ n4150 ^ 1'b0 ;
  assign n16912 = n16911 ^ n16909 ^ n1327 ;
  assign n16913 = n1298 & n7643 ;
  assign n16914 = ~n10641 & n16913 ;
  assign n16915 = n16914 ^ n3669 ^ n726 ;
  assign n16916 = n5439 & ~n12419 ;
  assign n16917 = ~n363 & n16916 ;
  assign n16918 = n1173 | n16917 ;
  assign n16919 = n16345 ^ n12907 ^ 1'b0 ;
  assign n16920 = n16918 & n16919 ;
  assign n16921 = n16920 ^ n2271 ^ 1'b0 ;
  assign n16922 = ( ~n970 & n15419 ) | ( ~n970 & n16921 ) | ( n15419 & n16921 ) ;
  assign n16928 = n4779 ^ n4245 ^ n2411 ;
  assign n16929 = n10052 | n16928 ;
  assign n16930 = n16929 ^ n16471 ^ 1'b0 ;
  assign n16931 = ( x56 & n10473 ) | ( x56 & n16930 ) | ( n10473 & n16930 ) ;
  assign n16925 = n1524 & n3845 ;
  assign n16923 = ( n3551 & ~n10936 ) | ( n3551 & n11155 ) | ( ~n10936 & n11155 ) ;
  assign n16924 = n6608 & ~n16923 ;
  assign n16926 = n16925 ^ n16924 ^ 1'b0 ;
  assign n16927 = n16926 ^ n13138 ^ 1'b0 ;
  assign n16932 = n16931 ^ n16927 ^ n9357 ;
  assign n16933 = n9624 ^ n7121 ^ n1788 ;
  assign n16934 = n7031 & n10927 ;
  assign n16935 = ~n16933 & n16934 ;
  assign n16936 = n16483 ^ n13554 ^ n821 ;
  assign n16937 = n16936 ^ n5323 ^ x245 ;
  assign n16938 = n4503 | n16937 ;
  assign n16939 = n15189 & ~n16938 ;
  assign n16940 = ( ~n3068 & n16782 ) | ( ~n3068 & n16939 ) | ( n16782 & n16939 ) ;
  assign n16941 = n9391 & ~n12236 ;
  assign n16942 = n16941 ^ n14963 ^ 1'b0 ;
  assign n16943 = ~n16940 & n16942 ;
  assign n16944 = ~n11715 & n16943 ;
  assign n16945 = ( n1139 & n5236 ) | ( n1139 & ~n6817 ) | ( n5236 & ~n6817 ) ;
  assign n16946 = n2181 & n16945 ;
  assign n16947 = ~n8844 & n16946 ;
  assign n16948 = ( n10354 & n10530 ) | ( n10354 & n16220 ) | ( n10530 & n16220 ) ;
  assign n16949 = n2934 ^ n1972 ^ 1'b0 ;
  assign n16950 = ( n2303 & ~n14166 ) | ( n2303 & n16949 ) | ( ~n14166 & n16949 ) ;
  assign n16951 = ( n9164 & ~n9890 ) | ( n9164 & n11642 ) | ( ~n9890 & n11642 ) ;
  assign n16952 = n16951 ^ n1609 ^ 1'b0 ;
  assign n16953 = n2395 | n9794 ;
  assign n16954 = n9979 & ~n16953 ;
  assign n16955 = n16954 ^ n3014 ^ 1'b0 ;
  assign n16956 = ( ~n5294 & n6657 ) | ( ~n5294 & n15545 ) | ( n6657 & n15545 ) ;
  assign n16957 = n16955 & ~n16956 ;
  assign n16958 = n12248 & n12388 ;
  assign n16959 = n13000 ^ n8064 ^ n1970 ;
  assign n16960 = n13948 ^ n8933 ^ n1550 ;
  assign n16961 = ( n1002 & n16959 ) | ( n1002 & n16960 ) | ( n16959 & n16960 ) ;
  assign n16962 = n1332 & ~n10384 ;
  assign n16963 = n12890 & n16962 ;
  assign n16964 = n6523 ^ n5576 ^ x76 ;
  assign n16965 = n16964 ^ n12301 ^ 1'b0 ;
  assign n16966 = n15714 & n16965 ;
  assign n16967 = n16963 & n16966 ;
  assign n16968 = n3822 | n16967 ;
  assign n16969 = n16968 ^ n14755 ^ 1'b0 ;
  assign n16972 = ~n2060 & n15302 ;
  assign n16973 = ~n4154 & n16972 ;
  assign n16970 = ~n9771 & n9808 ;
  assign n16971 = n16970 ^ n9993 ^ n4894 ;
  assign n16974 = n16973 ^ n16971 ^ n8360 ;
  assign n16975 = n3536 & n10538 ;
  assign n16976 = ~n7153 & n16975 ;
  assign n16977 = ( ~x47 & n11409 ) | ( ~x47 & n16976 ) | ( n11409 & n16976 ) ;
  assign n16978 = ~n11389 & n11665 ;
  assign n16979 = n16978 ^ n6249 ^ n3269 ;
  assign n16980 = ( n4135 & n5058 ) | ( n4135 & ~n16979 ) | ( n5058 & ~n16979 ) ;
  assign n16981 = n12229 ^ n4651 ^ 1'b0 ;
  assign n16982 = n3676 & ~n16981 ;
  assign n16983 = n16982 ^ n4867 ^ 1'b0 ;
  assign n16984 = ~n5511 & n16983 ;
  assign n16985 = ( n3965 & ~n4740 ) | ( n3965 & n9483 ) | ( ~n4740 & n9483 ) ;
  assign n16986 = n16985 ^ n5908 ^ n1851 ;
  assign n16987 = n4554 & n11372 ;
  assign n16988 = n15657 & n16987 ;
  assign n16989 = n16988 ^ n14603 ^ n2300 ;
  assign n16990 = n16989 ^ n6365 ^ n4972 ;
  assign n16991 = n16990 ^ n9924 ^ n5178 ;
  assign n17001 = n2080 & ~n6049 ;
  assign n16997 = n3526 | n4120 ;
  assign n16998 = n2530 & ~n16997 ;
  assign n16996 = n3119 | n5549 ;
  assign n16999 = n16998 ^ n16996 ^ n1408 ;
  assign n17000 = n16999 ^ n13631 ^ n5130 ;
  assign n16992 = n7842 ^ n1713 ^ 1'b0 ;
  assign n16993 = n15600 | n16992 ;
  assign n16994 = n16993 ^ n13881 ^ 1'b0 ;
  assign n16995 = n8374 & ~n16994 ;
  assign n17002 = n17001 ^ n17000 ^ n16995 ;
  assign n17003 = n17002 ^ n6550 ^ 1'b0 ;
  assign n17004 = n10967 | n17003 ;
  assign n17008 = ( n4113 & n5442 ) | ( n4113 & ~n6106 ) | ( n5442 & ~n6106 ) ;
  assign n17005 = ( n784 & n3914 ) | ( n784 & ~n4645 ) | ( n3914 & ~n4645 ) ;
  assign n17006 = n17005 ^ n501 ^ 1'b0 ;
  assign n17007 = ( n981 & ~n5976 ) | ( n981 & n17006 ) | ( ~n5976 & n17006 ) ;
  assign n17009 = n17008 ^ n17007 ^ n8607 ;
  assign n17010 = ~x222 & n3528 ;
  assign n17011 = n17010 ^ n6076 ^ 1'b0 ;
  assign n17012 = ( ~n3249 & n3686 ) | ( ~n3249 & n16447 ) | ( n3686 & n16447 ) ;
  assign n17013 = n17011 & n17012 ;
  assign n17014 = ~n14521 & n17013 ;
  assign n17015 = ( n680 & n2643 ) | ( n680 & n3305 ) | ( n2643 & n3305 ) ;
  assign n17016 = n17014 & ~n17015 ;
  assign n17018 = n917 & n3141 ;
  assign n17019 = n11301 & n17018 ;
  assign n17017 = n2886 & ~n5732 ;
  assign n17020 = n17019 ^ n17017 ^ 1'b0 ;
  assign n17021 = n11406 ^ n1284 ^ 1'b0 ;
  assign n17024 = ( ~n2824 & n5449 ) | ( ~n2824 & n9142 ) | ( n5449 & n9142 ) ;
  assign n17025 = n6006 & ~n17024 ;
  assign n17026 = n7661 & n17025 ;
  assign n17027 = n6872 ^ n3255 ^ n2930 ;
  assign n17028 = n817 & n17027 ;
  assign n17029 = n17026 & n17028 ;
  assign n17022 = ( ~n8549 & n9380 ) | ( ~n8549 & n12926 ) | ( n9380 & n12926 ) ;
  assign n17023 = n16836 & ~n17022 ;
  assign n17030 = n17029 ^ n17023 ^ 1'b0 ;
  assign n17031 = n14497 ^ n11483 ^ 1'b0 ;
  assign n17034 = n4772 ^ n541 ^ 1'b0 ;
  assign n17032 = ( n1034 & n3071 ) | ( n1034 & ~n4788 ) | ( n3071 & ~n4788 ) ;
  assign n17033 = n8946 & ~n17032 ;
  assign n17035 = n17034 ^ n17033 ^ 1'b0 ;
  assign n17036 = ( n15345 & ~n17031 ) | ( n15345 & n17035 ) | ( ~n17031 & n17035 ) ;
  assign n17037 = n12707 ^ n5990 ^ x87 ;
  assign n17038 = ( n5298 & n7167 ) | ( n5298 & n11612 ) | ( n7167 & n11612 ) ;
  assign n17039 = ( ~n6148 & n13512 ) | ( ~n6148 & n17038 ) | ( n13512 & n17038 ) ;
  assign n17040 = n17039 ^ n16212 ^ n6971 ;
  assign n17041 = n17037 & ~n17040 ;
  assign n17042 = ( ~n4365 & n15324 ) | ( ~n4365 & n17041 ) | ( n15324 & n17041 ) ;
  assign n17043 = n17042 ^ n9679 ^ 1'b0 ;
  assign n17044 = n17043 ^ n16829 ^ n8410 ;
  assign n17045 = n8466 ^ n1235 ^ 1'b0 ;
  assign n17046 = n8793 ^ n6430 ^ 1'b0 ;
  assign n17047 = n17045 | n17046 ;
  assign n17048 = n17047 ^ n3678 ^ 1'b0 ;
  assign n17049 = n17048 ^ n7401 ^ n1136 ;
  assign n17050 = n5548 ^ n4795 ^ 1'b0 ;
  assign n17051 = n3779 | n17050 ;
  assign n17052 = n918 & ~n17051 ;
  assign n17053 = ~n17049 & n17052 ;
  assign n17054 = n6355 ^ n3191 ^ n1569 ;
  assign n17055 = n17054 ^ n3266 ^ 1'b0 ;
  assign n17056 = n9048 & ~n17055 ;
  assign n17057 = n15425 ^ n6967 ^ 1'b0 ;
  assign n17058 = ( n1601 & n14204 ) | ( n1601 & n17057 ) | ( n14204 & n17057 ) ;
  assign n17059 = ( ~n6045 & n17056 ) | ( ~n6045 & n17058 ) | ( n17056 & n17058 ) ;
  assign n17060 = n4620 & ~n10863 ;
  assign n17061 = n4905 | n17060 ;
  assign n17062 = n17061 ^ n13940 ^ 1'b0 ;
  assign n17063 = ( n2648 & n10402 ) | ( n2648 & ~n17062 ) | ( n10402 & ~n17062 ) ;
  assign n17064 = n13461 ^ n6301 ^ n1764 ;
  assign n17068 = ( n1267 & ~n2565 ) | ( n1267 & n12845 ) | ( ~n2565 & n12845 ) ;
  assign n17065 = n418 | n2678 ;
  assign n17066 = n6242 | n17065 ;
  assign n17067 = n10913 & n17066 ;
  assign n17069 = n17068 ^ n17067 ^ n12075 ;
  assign n17070 = n3901 & n12434 ;
  assign n17071 = ~n2738 & n17070 ;
  assign n17072 = n15731 & ~n17071 ;
  assign n17073 = n3226 ^ n1028 ^ 1'b0 ;
  assign n17074 = ~n1683 & n17073 ;
  assign n17075 = n17074 ^ n1511 ^ 1'b0 ;
  assign n17076 = n8387 ^ n7450 ^ 1'b0 ;
  assign n17077 = n17075 & ~n17076 ;
  assign n17083 = n11383 ^ n634 ^ 1'b0 ;
  assign n17084 = ~n5892 & n17083 ;
  assign n17078 = n8685 ^ n3198 ^ n1612 ;
  assign n17079 = ( ~n6919 & n7114 ) | ( ~n6919 & n11504 ) | ( n7114 & n11504 ) ;
  assign n17080 = n17078 & ~n17079 ;
  assign n17081 = n17080 ^ n14049 ^ 1'b0 ;
  assign n17082 = n17081 ^ n13663 ^ n13023 ;
  assign n17085 = n17084 ^ n17082 ^ 1'b0 ;
  assign n17086 = n17077 & n17085 ;
  assign n17087 = ~n1446 & n11567 ;
  assign n17088 = n5291 ^ n3530 ^ n1768 ;
  assign n17089 = ( n2978 & n5767 ) | ( n2978 & n17088 ) | ( n5767 & n17088 ) ;
  assign n17093 = ( n1315 & ~n1983 ) | ( n1315 & n5612 ) | ( ~n1983 & n5612 ) ;
  assign n17091 = n8472 ^ n2504 ^ 1'b0 ;
  assign n17092 = ( n8891 & n9703 ) | ( n8891 & ~n17091 ) | ( n9703 & ~n17091 ) ;
  assign n17090 = ( n10103 & n10471 ) | ( n10103 & ~n11348 ) | ( n10471 & ~n11348 ) ;
  assign n17094 = n17093 ^ n17092 ^ n17090 ;
  assign n17095 = ( n2738 & n8603 ) | ( n2738 & ~n11483 ) | ( n8603 & ~n11483 ) ;
  assign n17096 = ( n585 & n12280 ) | ( n585 & ~n12689 ) | ( n12280 & ~n12689 ) ;
  assign n17097 = n6988 ^ x58 ^ 1'b0 ;
  assign n17098 = ~n7738 & n17097 ;
  assign n17099 = ( ~n10660 & n11136 ) | ( ~n10660 & n17098 ) | ( n11136 & n17098 ) ;
  assign n17100 = n14871 ^ n2641 ^ x27 ;
  assign n17101 = ( n1496 & ~n8288 ) | ( n1496 & n17100 ) | ( ~n8288 & n17100 ) ;
  assign n17102 = ( n13970 & ~n14856 ) | ( n13970 & n17101 ) | ( ~n14856 & n17101 ) ;
  assign n17103 = n5657 | n17102 ;
  assign n17104 = n13548 & n17103 ;
  assign n17105 = ~n17099 & n17104 ;
  assign n17109 = n11236 ^ n7151 ^ n6834 ;
  assign n17110 = n17109 ^ n7388 ^ 1'b0 ;
  assign n17111 = n17110 ^ n7635 ^ n3027 ;
  assign n17112 = n17111 ^ n16227 ^ n2627 ;
  assign n17106 = ( n1463 & n2738 ) | ( n1463 & n9479 ) | ( n2738 & n9479 ) ;
  assign n17107 = ~n10327 & n17106 ;
  assign n17108 = n17107 ^ n2244 ^ 1'b0 ;
  assign n17113 = n17112 ^ n17108 ^ n382 ;
  assign n17115 = n12438 ^ n3896 ^ 1'b0 ;
  assign n17116 = ~n12236 & n17115 ;
  assign n17117 = ( n1218 & n4476 ) | ( n1218 & n17116 ) | ( n4476 & n17116 ) ;
  assign n17114 = ~n6150 & n7692 ;
  assign n17118 = n17117 ^ n17114 ^ 1'b0 ;
  assign n17119 = n1212 & n7120 ;
  assign n17120 = n17119 ^ n15748 ^ 1'b0 ;
  assign n17128 = ~n2108 & n6164 ;
  assign n17127 = ( n7761 & n12930 ) | ( n7761 & n13109 ) | ( n12930 & n13109 ) ;
  assign n17121 = n16250 ^ n4677 ^ n1243 ;
  assign n17124 = n3287 | n9402 ;
  assign n17122 = n930 | n10411 ;
  assign n17123 = n17122 ^ n9209 ^ n5637 ;
  assign n17125 = n17124 ^ n17123 ^ n3129 ;
  assign n17126 = ( ~n6205 & n17121 ) | ( ~n6205 & n17125 ) | ( n17121 & n17125 ) ;
  assign n17129 = n17128 ^ n17127 ^ n17126 ;
  assign n17130 = n729 & n1913 ;
  assign n17131 = n14045 ^ n3798 ^ 1'b0 ;
  assign n17132 = ~n17130 & n17131 ;
  assign n17133 = n17132 ^ n15786 ^ n10493 ;
  assign n17134 = n14418 ^ n10865 ^ n2029 ;
  assign n17141 = ( n2722 & n3902 ) | ( n2722 & n8738 ) | ( n3902 & n8738 ) ;
  assign n17142 = n12596 ^ n5983 ^ n5443 ;
  assign n17143 = n17141 & ~n17142 ;
  assign n17144 = n17143 ^ n2295 ^ 1'b0 ;
  assign n17140 = n6069 ^ n1108 ^ 1'b0 ;
  assign n17136 = n3378 & ~n6784 ;
  assign n17137 = n6972 & ~n17136 ;
  assign n17138 = n17137 ^ n6528 ^ 1'b0 ;
  assign n17135 = ~n5743 & n9738 ;
  assign n17139 = n17138 ^ n17135 ^ 1'b0 ;
  assign n17145 = n17144 ^ n17140 ^ n17139 ;
  assign n17146 = n10553 | n15533 ;
  assign n17147 = n17146 ^ n5716 ^ 1'b0 ;
  assign n17148 = n17147 ^ n5372 ^ n2053 ;
  assign n17149 = ( n6798 & n10348 ) | ( n6798 & ~n17148 ) | ( n10348 & ~n17148 ) ;
  assign n17150 = n7703 ^ n6930 ^ x150 ;
  assign n17151 = ( x202 & n9466 ) | ( x202 & n9635 ) | ( n9466 & n9635 ) ;
  assign n17152 = n5640 & ~n9251 ;
  assign n17153 = ~n8860 & n17152 ;
  assign n17154 = ( x83 & n17151 ) | ( x83 & ~n17153 ) | ( n17151 & ~n17153 ) ;
  assign n17155 = n13098 ^ n7670 ^ n5335 ;
  assign n17156 = ( n1518 & n12617 ) | ( n1518 & n17155 ) | ( n12617 & n17155 ) ;
  assign n17157 = n17156 ^ n4583 ^ n1996 ;
  assign n17158 = ~n17154 & n17157 ;
  assign n17159 = n11870 & ~n13457 ;
  assign n17160 = n11558 ^ n8844 ^ n7591 ;
  assign n17161 = n17160 ^ n7667 ^ n688 ;
  assign n17162 = ( ~n2755 & n7319 ) | ( ~n2755 & n7597 ) | ( n7319 & n7597 ) ;
  assign n17163 = n17162 ^ n14999 ^ n3561 ;
  assign n17164 = ( n13556 & n17161 ) | ( n13556 & ~n17163 ) | ( n17161 & ~n17163 ) ;
  assign n17165 = ~n5574 & n17164 ;
  assign n17166 = n8749 ^ n332 ^ 1'b0 ;
  assign n17167 = ~n11256 & n17166 ;
  assign n17168 = ( n2255 & n4554 ) | ( n2255 & ~n17167 ) | ( n4554 & ~n17167 ) ;
  assign n17169 = n13875 ^ n4362 ^ 1'b0 ;
  assign n17170 = n17169 ^ n14106 ^ n9033 ;
  assign n17171 = n17170 ^ n14513 ^ n4798 ;
  assign n17172 = n578 | n5363 ;
  assign n17173 = n2432 & ~n6979 ;
  assign n17174 = ~n17172 & n17173 ;
  assign n17175 = ( n669 & n8770 ) | ( n669 & n17174 ) | ( n8770 & n17174 ) ;
  assign n17176 = ~n3142 & n17175 ;
  assign n17177 = n16628 & n17176 ;
  assign n17178 = n17177 ^ n12166 ^ 1'b0 ;
  assign n17179 = ~n11526 & n14842 ;
  assign n17180 = n17179 ^ n6541 ^ 1'b0 ;
  assign n17181 = ~n885 & n4725 ;
  assign n17182 = n17181 ^ n7601 ^ 1'b0 ;
  assign n17183 = ~n4032 & n17182 ;
  assign n17184 = ( n4591 & n17180 ) | ( n4591 & n17183 ) | ( n17180 & n17183 ) ;
  assign n17185 = ( ~n5206 & n5957 ) | ( ~n5206 & n16586 ) | ( n5957 & n16586 ) ;
  assign n17186 = n17185 ^ n10047 ^ n7114 ;
  assign n17187 = n2006 & n3459 ;
  assign n17188 = n15204 ^ n10123 ^ n4008 ;
  assign n17189 = n17188 ^ n6985 ^ n6952 ;
  assign n17190 = ( n7143 & ~n17187 ) | ( n7143 & n17189 ) | ( ~n17187 & n17189 ) ;
  assign n17191 = ( n2481 & n9134 ) | ( n2481 & ~n14945 ) | ( n9134 & ~n14945 ) ;
  assign n17192 = n3258 & ~n17191 ;
  assign n17193 = n11695 ^ n5032 ^ 1'b0 ;
  assign n17194 = ~n17192 & n17193 ;
  assign n17195 = ( ~n17186 & n17190 ) | ( ~n17186 & n17194 ) | ( n17190 & n17194 ) ;
  assign n17196 = n10982 ^ n7202 ^ 1'b0 ;
  assign n17198 = n3456 | n6963 ;
  assign n17199 = n17198 ^ n6465 ^ n3566 ;
  assign n17197 = n7430 & n10232 ;
  assign n17200 = n17199 ^ n17197 ^ 1'b0 ;
  assign n17201 = ( n5935 & ~n12518 ) | ( n5935 & n17200 ) | ( ~n12518 & n17200 ) ;
  assign n17202 = n17201 ^ n13677 ^ 1'b0 ;
  assign n17203 = ~n17196 & n17202 ;
  assign n17204 = n17203 ^ n15906 ^ 1'b0 ;
  assign n17205 = n6987 ^ n3501 ^ n773 ;
  assign n17206 = ( n284 & n3211 ) | ( n284 & ~n17205 ) | ( n3211 & ~n17205 ) ;
  assign n17207 = n17206 ^ n7672 ^ 1'b0 ;
  assign n17208 = ( n5872 & ~n6988 ) | ( n5872 & n16528 ) | ( ~n6988 & n16528 ) ;
  assign n17209 = n553 | n4886 ;
  assign n17210 = n4903 & ~n17209 ;
  assign n17211 = ( n3067 & ~n10384 ) | ( n3067 & n17210 ) | ( ~n10384 & n17210 ) ;
  assign n17212 = ( n4613 & ~n10645 ) | ( n4613 & n12997 ) | ( ~n10645 & n12997 ) ;
  assign n17213 = ( n5384 & ~n6731 ) | ( n5384 & n17212 ) | ( ~n6731 & n17212 ) ;
  assign n17214 = n5402 ^ n1114 ^ 1'b0 ;
  assign n17215 = n7057 | n17214 ;
  assign n17216 = n17215 ^ n6059 ^ 1'b0 ;
  assign n17217 = ( n3669 & n5145 ) | ( n3669 & ~n13103 ) | ( n5145 & ~n13103 ) ;
  assign n17218 = ( ~n10342 & n16631 ) | ( ~n10342 & n17217 ) | ( n16631 & n17217 ) ;
  assign n17219 = n17218 ^ n16375 ^ 1'b0 ;
  assign n17220 = n10245 & n17219 ;
  assign n17221 = n14399 ^ n9609 ^ n6786 ;
  assign n17222 = n10701 ^ n8345 ^ 1'b0 ;
  assign n17223 = n2853 & n17222 ;
  assign n17224 = n2545 ^ n2380 ^ 1'b0 ;
  assign n17225 = n5269 ^ n2462 ^ 1'b0 ;
  assign n17226 = ~n10907 & n17225 ;
  assign n17227 = n7277 ^ n1583 ^ 1'b0 ;
  assign n17228 = n5002 | n17227 ;
  assign n17229 = n9869 & ~n17228 ;
  assign n17230 = n7746 | n17229 ;
  assign n17231 = ( n17224 & ~n17226 ) | ( n17224 & n17230 ) | ( ~n17226 & n17230 ) ;
  assign n17232 = n14094 ^ n2654 ^ 1'b0 ;
  assign n17233 = n4518 ^ n4050 ^ n4036 ;
  assign n17234 = ( n9542 & n11230 ) | ( n9542 & n14600 ) | ( n11230 & n14600 ) ;
  assign n17235 = ( ~n17232 & n17233 ) | ( ~n17232 & n17234 ) | ( n17233 & n17234 ) ;
  assign n17236 = ~n12323 & n16337 ;
  assign n17237 = n14345 ^ n4261 ^ 1'b0 ;
  assign n17238 = n1840 & n17237 ;
  assign n17239 = n17199 ^ n4057 ^ n2130 ;
  assign n17240 = n12878 & n17239 ;
  assign n17241 = n17240 ^ n1678 ^ 1'b0 ;
  assign n17242 = ( ~n6045 & n9773 ) | ( ~n6045 & n17241 ) | ( n9773 & n17241 ) ;
  assign n17243 = n12146 ^ n4285 ^ 1'b0 ;
  assign n17244 = n261 | n17243 ;
  assign n17245 = ( n10903 & n16689 ) | ( n10903 & ~n17244 ) | ( n16689 & ~n17244 ) ;
  assign n17246 = n14436 ^ n3908 ^ 1'b0 ;
  assign n17247 = n17245 & ~n17246 ;
  assign n17251 = ( n673 & n4773 ) | ( n673 & n16250 ) | ( n4773 & n16250 ) ;
  assign n17248 = n9522 ^ n6918 ^ n5328 ;
  assign n17249 = n17248 ^ n16567 ^ n436 ;
  assign n17250 = n3108 & ~n17249 ;
  assign n17252 = n17251 ^ n17250 ^ 1'b0 ;
  assign n17254 = n5961 ^ n4730 ^ n2259 ;
  assign n17255 = n17254 ^ n11665 ^ n6644 ;
  assign n17253 = n11330 | n12523 ;
  assign n17256 = n17255 ^ n17253 ^ 1'b0 ;
  assign n17257 = n17256 ^ n15995 ^ n6761 ;
  assign n17258 = ~n14240 & n16036 ;
  assign n17259 = ~n16036 & n17258 ;
  assign n17260 = n17141 & ~n17259 ;
  assign n17261 = n9431 & n17260 ;
  assign n17262 = n5085 ^ n4217 ^ x71 ;
  assign n17263 = n406 ^ x92 ^ 1'b0 ;
  assign n17264 = x250 & n17263 ;
  assign n17265 = ( n350 & n14106 ) | ( n350 & ~n17264 ) | ( n14106 & ~n17264 ) ;
  assign n17266 = n14783 | n17265 ;
  assign n17267 = ( n17261 & ~n17262 ) | ( n17261 & n17266 ) | ( ~n17262 & n17266 ) ;
  assign n17268 = ~n4935 & n17267 ;
  assign n17269 = ( n3046 & ~n3918 ) | ( n3046 & n15177 ) | ( ~n3918 & n15177 ) ;
  assign n17270 = n6959 ^ n1588 ^ n488 ;
  assign n17271 = n17270 ^ n2710 ^ 1'b0 ;
  assign n17272 = n9831 ^ n5542 ^ 1'b0 ;
  assign n17273 = n5824 ^ n2715 ^ n2210 ;
  assign n17274 = n458 ^ n450 ^ 1'b0 ;
  assign n17275 = n7330 & n17274 ;
  assign n17276 = n7426 & n12922 ;
  assign n17277 = n17276 ^ n12271 ^ n8865 ;
  assign n17279 = n10893 ^ n7051 ^ n1882 ;
  assign n17278 = ( n278 & ~n6978 ) | ( n278 & n13924 ) | ( ~n6978 & n13924 ) ;
  assign n17280 = n17279 ^ n17278 ^ n15891 ;
  assign n17281 = n17277 | n17280 ;
  assign n17282 = n1358 & ~n7566 ;
  assign n17283 = n17281 & n17282 ;
  assign n17284 = n14131 ^ n7279 ^ n1161 ;
  assign n17285 = n2605 | n12930 ;
  assign n17286 = n9304 & n12883 ;
  assign n17287 = n17286 ^ n9408 ^ 1'b0 ;
  assign n17288 = ( ~n1596 & n3007 ) | ( ~n1596 & n4256 ) | ( n3007 & n4256 ) ;
  assign n17289 = n17288 ^ n6690 ^ n2786 ;
  assign n17290 = n4982 & ~n6887 ;
  assign n17291 = ~n5450 & n17290 ;
  assign n17292 = n17291 ^ n7293 ^ 1'b0 ;
  assign n17293 = n17289 & n17292 ;
  assign n17294 = ( n15425 & n17287 ) | ( n15425 & ~n17293 ) | ( n17287 & ~n17293 ) ;
  assign n17295 = n15945 ^ n11424 ^ 1'b0 ;
  assign n17296 = n17294 & n17295 ;
  assign n17297 = ( n5186 & ~n7290 ) | ( n5186 & n11372 ) | ( ~n7290 & n11372 ) ;
  assign n17298 = n3465 | n9775 ;
  assign n17299 = n2442 & ~n17298 ;
  assign n17300 = n15405 & ~n17299 ;
  assign n17301 = n15875 ^ n3729 ^ n1272 ;
  assign n17302 = ( n10254 & ~n15949 ) | ( n10254 & n17301 ) | ( ~n15949 & n17301 ) ;
  assign n17303 = ( n6525 & n17300 ) | ( n6525 & n17302 ) | ( n17300 & n17302 ) ;
  assign n17304 = ( n5302 & n8335 ) | ( n5302 & n8338 ) | ( n8335 & n8338 ) ;
  assign n17305 = ( ~n1077 & n2378 ) | ( ~n1077 & n17304 ) | ( n2378 & n17304 ) ;
  assign n17306 = n9202 ^ n3181 ^ 1'b0 ;
  assign n17307 = n10312 & n17306 ;
  assign n17308 = n12133 ^ n7355 ^ 1'b0 ;
  assign n17309 = n13370 & ~n17308 ;
  assign n17310 = ( ~n1465 & n10557 ) | ( ~n1465 & n10752 ) | ( n10557 & n10752 ) ;
  assign n17312 = ( n1012 & ~n1114 ) | ( n1012 & n5968 ) | ( ~n1114 & n5968 ) ;
  assign n17313 = n17312 ^ n9895 ^ n3988 ;
  assign n17314 = ( ~n4842 & n10992 ) | ( ~n4842 & n17313 ) | ( n10992 & n17313 ) ;
  assign n17311 = ( ~n6719 & n10298 ) | ( ~n6719 & n11384 ) | ( n10298 & n11384 ) ;
  assign n17315 = n17314 ^ n17311 ^ n9312 ;
  assign n17316 = n1805 ^ n1799 ^ n517 ;
  assign n17317 = ( n9123 & n16979 ) | ( n9123 & ~n17316 ) | ( n16979 & ~n17316 ) ;
  assign n17318 = ~n2243 & n4304 ;
  assign n17319 = n17318 ^ n4802 ^ 1'b0 ;
  assign n17320 = n16714 | n17319 ;
  assign n17321 = n6079 ^ n4013 ^ 1'b0 ;
  assign n17322 = ( x132 & n2566 ) | ( x132 & n17321 ) | ( n2566 & n17321 ) ;
  assign n17323 = ( n7569 & n7749 ) | ( n7569 & n9901 ) | ( n7749 & n9901 ) ;
  assign n17324 = n12588 ^ n9902 ^ n1173 ;
  assign n17325 = ( n7503 & n17323 ) | ( n7503 & n17324 ) | ( n17323 & n17324 ) ;
  assign n17326 = ( ~n10398 & n17322 ) | ( ~n10398 & n17325 ) | ( n17322 & n17325 ) ;
  assign n17327 = n17144 ^ n6014 ^ 1'b0 ;
  assign n17336 = ( n2901 & n4566 ) | ( n2901 & n6193 ) | ( n4566 & n6193 ) ;
  assign n17334 = ( n4070 & n6704 ) | ( n4070 & ~n12481 ) | ( n6704 & ~n12481 ) ;
  assign n17328 = ~n1378 & n3542 ;
  assign n17329 = n17328 ^ n2256 ^ 1'b0 ;
  assign n17330 = n3313 ^ n1733 ^ x166 ;
  assign n17331 = n10060 ^ n2646 ^ 1'b0 ;
  assign n17332 = n17330 | n17331 ;
  assign n17333 = ( ~n3158 & n17329 ) | ( ~n3158 & n17332 ) | ( n17329 & n17332 ) ;
  assign n17335 = n17334 ^ n17333 ^ n13665 ;
  assign n17337 = n17336 ^ n17335 ^ n9247 ;
  assign n17338 = n6153 & ~n13813 ;
  assign n17339 = n3670 & n17338 ;
  assign n17340 = n12638 & ~n17339 ;
  assign n17341 = n17340 ^ n16907 ^ 1'b0 ;
  assign n17344 = ( n1710 & n6771 ) | ( n1710 & ~n7452 ) | ( n6771 & ~n7452 ) ;
  assign n17345 = ( n1214 & n13972 ) | ( n1214 & n17344 ) | ( n13972 & n17344 ) ;
  assign n17342 = ( n1061 & ~n3064 ) | ( n1061 & n5997 ) | ( ~n3064 & n5997 ) ;
  assign n17343 = ( ~x142 & n2839 ) | ( ~x142 & n17342 ) | ( n2839 & n17342 ) ;
  assign n17346 = n17345 ^ n17343 ^ 1'b0 ;
  assign n17347 = n16106 & n17346 ;
  assign n17348 = n3051 & n17347 ;
  assign n17349 = ~n3178 & n8112 ;
  assign n17350 = n11143 ^ n6604 ^ n3225 ;
  assign n17351 = n9683 & n9972 ;
  assign n17352 = n4441 & n17351 ;
  assign n17353 = n17350 | n17352 ;
  assign n17354 = n17353 ^ n4322 ^ 1'b0 ;
  assign n17355 = ( n8128 & n17349 ) | ( n8128 & ~n17354 ) | ( n17349 & ~n17354 ) ;
  assign n17360 = ( ~n447 & n1771 ) | ( ~n447 & n10372 ) | ( n1771 & n10372 ) ;
  assign n17356 = n993 | n5488 ;
  assign n17357 = n17356 ^ n9785 ^ 1'b0 ;
  assign n17358 = n17357 ^ n5490 ^ n4306 ;
  assign n17359 = ~n11423 & n17358 ;
  assign n17361 = n17360 ^ n17359 ^ 1'b0 ;
  assign n17362 = ( x194 & ~n2680 ) | ( x194 & n2894 ) | ( ~n2680 & n2894 ) ;
  assign n17363 = n5693 ^ n2315 ^ 1'b0 ;
  assign n17364 = n17363 ^ n9811 ^ 1'b0 ;
  assign n17365 = ( n4275 & n17362 ) | ( n4275 & ~n17364 ) | ( n17362 & ~n17364 ) ;
  assign n17366 = n9991 | n15946 ;
  assign n17367 = n17366 ^ n12418 ^ 1'b0 ;
  assign n17372 = ( n6275 & n10894 ) | ( n6275 & ~n17151 ) | ( n10894 & ~n17151 ) ;
  assign n17373 = n17372 ^ n14314 ^ n2645 ;
  assign n17370 = ( ~n8341 & n11908 ) | ( ~n8341 & n13834 ) | ( n11908 & n13834 ) ;
  assign n17369 = n17054 ^ n3833 ^ 1'b0 ;
  assign n17371 = n17370 ^ n17369 ^ n11360 ;
  assign n17368 = n813 | n3564 ;
  assign n17374 = n17373 ^ n17371 ^ n17368 ;
  assign n17375 = n2218 | n16702 ;
  assign n17376 = x53 & n15814 ;
  assign n17377 = ~n10757 & n17376 ;
  assign n17381 = n17074 ^ n16503 ^ x246 ;
  assign n17378 = n6521 ^ n1048 ^ n642 ;
  assign n17379 = ~n3757 & n17378 ;
  assign n17380 = n9317 & n17379 ;
  assign n17382 = n17381 ^ n17380 ^ n3238 ;
  assign n17383 = ( n2559 & ~n13686 ) | ( n2559 & n16018 ) | ( ~n13686 & n16018 ) ;
  assign n17384 = ( ~n2244 & n8085 ) | ( ~n2244 & n17383 ) | ( n8085 & n17383 ) ;
  assign n17385 = n17060 ^ n3916 ^ 1'b0 ;
  assign n17386 = n811 | n2941 ;
  assign n17387 = ( n1778 & n2402 ) | ( n1778 & n17386 ) | ( n2402 & n17386 ) ;
  assign n17388 = ( ~n280 & n1503 ) | ( ~n280 & n4570 ) | ( n1503 & n4570 ) ;
  assign n17389 = n3543 | n7586 ;
  assign n17390 = n17389 ^ n4224 ^ 1'b0 ;
  assign n17391 = ( n17387 & n17388 ) | ( n17387 & ~n17390 ) | ( n17388 & ~n17390 ) ;
  assign n17392 = ~n1710 & n17391 ;
  assign n17396 = n3768 ^ n3290 ^ 1'b0 ;
  assign n17397 = n3889 & n17396 ;
  assign n17398 = n17397 ^ n2800 ^ n1126 ;
  assign n17395 = n1020 & ~n6681 ;
  assign n17399 = n17398 ^ n17395 ^ n9348 ;
  assign n17393 = ~n6220 & n12226 ;
  assign n17394 = n17393 ^ n7910 ^ n7531 ;
  assign n17400 = n17399 ^ n17394 ^ n8284 ;
  assign n17401 = n2432 & ~n13257 ;
  assign n17402 = ~n5418 & n17401 ;
  assign n17403 = n3166 ^ n3039 ^ 1'b0 ;
  assign n17404 = n9747 ^ n6810 ^ 1'b0 ;
  assign n17405 = ( ~n1386 & n5651 ) | ( ~n1386 & n15294 ) | ( n5651 & n15294 ) ;
  assign n17406 = ( n8110 & n17404 ) | ( n8110 & n17405 ) | ( n17404 & n17405 ) ;
  assign n17407 = ~n13442 & n17349 ;
  assign n17408 = ( n2613 & n4890 ) | ( n2613 & ~n17407 ) | ( n4890 & ~n17407 ) ;
  assign n17409 = ( n1538 & ~n17406 ) | ( n1538 & n17408 ) | ( ~n17406 & n17408 ) ;
  assign n17410 = ( ~n3349 & n8376 ) | ( ~n3349 & n10056 ) | ( n8376 & n10056 ) ;
  assign n17411 = ( ~n5567 & n10291 ) | ( ~n5567 & n17410 ) | ( n10291 & n17410 ) ;
  assign n17412 = ( n11382 & n11730 ) | ( n11382 & ~n15182 ) | ( n11730 & ~n15182 ) ;
  assign n17413 = n927 & n4674 ;
  assign n17414 = ~n12637 & n17413 ;
  assign n17415 = n17414 ^ n12539 ^ n8842 ;
  assign n17416 = n442 | n4620 ;
  assign n17417 = n17416 ^ n13464 ^ 1'b0 ;
  assign n17424 = ( n1889 & n4860 ) | ( n1889 & ~n12632 ) | ( n4860 & ~n12632 ) ;
  assign n17425 = ~n5216 & n17424 ;
  assign n17418 = ~n6442 & n8259 ;
  assign n17419 = ( n1682 & n6817 ) | ( n1682 & ~n17418 ) | ( n6817 & ~n17418 ) ;
  assign n17420 = n10605 ^ n9180 ^ n7357 ;
  assign n17421 = n17420 ^ n9351 ^ 1'b0 ;
  assign n17422 = n14988 & n17421 ;
  assign n17423 = ~n17419 & n17422 ;
  assign n17426 = n17425 ^ n17423 ^ x57 ;
  assign n17427 = ( n3690 & n9755 ) | ( n3690 & n12318 ) | ( n9755 & n12318 ) ;
  assign n17428 = n17427 ^ n13012 ^ n4955 ;
  assign n17430 = ~x70 & n4831 ;
  assign n17431 = n2789 | n17430 ;
  assign n17429 = ( n3506 & n5870 ) | ( n3506 & n8712 ) | ( n5870 & n8712 ) ;
  assign n17432 = n17431 ^ n17429 ^ n2329 ;
  assign n17433 = ( n407 & n4598 ) | ( n407 & ~n7702 ) | ( n4598 & ~n7702 ) ;
  assign n17434 = n6478 & n12219 ;
  assign n17435 = ~n5870 & n15191 ;
  assign n17436 = n4549 ^ n3456 ^ 1'b0 ;
  assign n17437 = x54 & n17436 ;
  assign n17438 = n8614 ^ n5978 ^ 1'b0 ;
  assign n17439 = n17437 | n17438 ;
  assign n17440 = n5547 & n16294 ;
  assign n17441 = n9100 & n17440 ;
  assign n17443 = n2868 & ~n6888 ;
  assign n17444 = n17443 ^ n16542 ^ 1'b0 ;
  assign n17442 = ( ~n4112 & n7110 ) | ( ~n4112 & n10311 ) | ( n7110 & n10311 ) ;
  assign n17445 = n17444 ^ n17442 ^ n14184 ;
  assign n17446 = n12450 & ~n12807 ;
  assign n17447 = ( n6972 & n9336 ) | ( n6972 & n17446 ) | ( n9336 & n17446 ) ;
  assign n17452 = n6725 | n8092 ;
  assign n17448 = ( n587 & n2778 ) | ( n587 & n4670 ) | ( n2778 & n4670 ) ;
  assign n17449 = ~n12728 & n17448 ;
  assign n17450 = n17449 ^ n14761 ^ 1'b0 ;
  assign n17451 = ~n13521 & n17450 ;
  assign n17453 = n17452 ^ n17451 ^ n890 ;
  assign n17462 = n6309 ^ n1009 ^ x221 ;
  assign n17463 = n17462 ^ n9505 ^ 1'b0 ;
  assign n17454 = n2104 & n7267 ;
  assign n17456 = n1942 ^ n1184 ^ 1'b0 ;
  assign n17457 = n2897 | n17456 ;
  assign n17455 = n6204 | n14523 ;
  assign n17458 = n17457 ^ n17455 ^ 1'b0 ;
  assign n17459 = n11951 | n17458 ;
  assign n17460 = n12545 | n17459 ;
  assign n17461 = ~n17454 & n17460 ;
  assign n17464 = n17463 ^ n17461 ^ 1'b0 ;
  assign n17465 = n8874 ^ n1299 ^ 1'b0 ;
  assign n17466 = ( n3857 & ~n12427 ) | ( n3857 & n16717 ) | ( ~n12427 & n16717 ) ;
  assign n17467 = n17026 | n17466 ;
  assign n17468 = n17465 & ~n17467 ;
  assign n17469 = ( n421 & n5975 ) | ( n421 & ~n8097 ) | ( n5975 & ~n8097 ) ;
  assign n17470 = n8836 ^ n2180 ^ n1106 ;
  assign n17471 = n17470 ^ n11318 ^ 1'b0 ;
  assign n17472 = n17469 & ~n17471 ;
  assign n17473 = n17472 ^ n6919 ^ n3059 ;
  assign n17474 = ~n2957 & n13347 ;
  assign n17475 = ~n6767 & n17474 ;
  assign n17476 = n10921 ^ n384 ^ 1'b0 ;
  assign n17477 = n16228 ^ n15483 ^ n3890 ;
  assign n17478 = ( n5021 & ~n5529 ) | ( n5021 & n17477 ) | ( ~n5529 & n17477 ) ;
  assign n17479 = n17478 ^ n7625 ^ 1'b0 ;
  assign n17480 = n17476 & n17479 ;
  assign n17481 = ( n5804 & n17475 ) | ( n5804 & n17480 ) | ( n17475 & n17480 ) ;
  assign n17482 = n4441 & n9316 ;
  assign n17484 = n16454 ^ n9339 ^ n7681 ;
  assign n17483 = n11745 & ~n16480 ;
  assign n17485 = n17484 ^ n17483 ^ 1'b0 ;
  assign n17486 = ( ~n9092 & n17482 ) | ( ~n9092 & n17485 ) | ( n17482 & n17485 ) ;
  assign n17487 = ( n6915 & n7186 ) | ( n6915 & ~n13618 ) | ( n7186 & ~n13618 ) ;
  assign n17490 = n7271 ^ n2206 ^ n1871 ;
  assign n17491 = n6794 ^ n5603 ^ 1'b0 ;
  assign n17492 = n17490 | n17491 ;
  assign n17488 = n10349 ^ x6 ^ 1'b0 ;
  assign n17489 = n17488 ^ n12488 ^ n6499 ;
  assign n17493 = n17492 ^ n17489 ^ n14389 ;
  assign n17499 = ( ~n2679 & n5913 ) | ( ~n2679 & n6127 ) | ( n5913 & n6127 ) ;
  assign n17494 = n15320 ^ n5743 ^ n3856 ;
  assign n17495 = n710 & ~n12257 ;
  assign n17496 = n17495 ^ n2538 ^ 1'b0 ;
  assign n17497 = n17494 | n17496 ;
  assign n17498 = n17497 ^ n4445 ^ 1'b0 ;
  assign n17500 = n17499 ^ n17498 ^ n3659 ;
  assign n17501 = ( n2580 & ~n12035 ) | ( n2580 & n17500 ) | ( ~n12035 & n17500 ) ;
  assign n17502 = n7050 ^ n4642 ^ n2717 ;
  assign n17503 = ( ~n16470 & n17336 ) | ( ~n16470 & n17502 ) | ( n17336 & n17502 ) ;
  assign n17504 = n10723 ^ n742 ^ 1'b0 ;
  assign n17505 = n11719 & ~n17504 ;
  assign n17506 = n15275 & n17505 ;
  assign n17509 = n15278 ^ n5786 ^ 1'b0 ;
  assign n17507 = n15469 ^ n4499 ^ x129 ;
  assign n17508 = n17507 ^ n11798 ^ 1'b0 ;
  assign n17510 = n17509 ^ n17508 ^ n7340 ;
  assign n17511 = n17510 ^ n15628 ^ 1'b0 ;
  assign n17512 = n1449 ^ n1434 ^ 1'b0 ;
  assign n17513 = ~n1221 & n17512 ;
  assign n17514 = ( ~n1600 & n3609 ) | ( ~n1600 & n17513 ) | ( n3609 & n17513 ) ;
  assign n17515 = ( n5918 & n17167 ) | ( n5918 & ~n17514 ) | ( n17167 & ~n17514 ) ;
  assign n17520 = ( n4310 & n5659 ) | ( n4310 & n14809 ) | ( n5659 & n14809 ) ;
  assign n17518 = n1774 & n6217 ;
  assign n17519 = n17518 ^ n6859 ^ 1'b0 ;
  assign n17516 = ( n1618 & ~n5886 ) | ( n1618 & n6200 ) | ( ~n5886 & n6200 ) ;
  assign n17517 = n17516 ^ n16979 ^ n9955 ;
  assign n17521 = n17520 ^ n17519 ^ n17517 ;
  assign n17523 = ~n1953 & n3727 ;
  assign n17522 = x237 & n9332 ;
  assign n17524 = n17523 ^ n17522 ^ 1'b0 ;
  assign n17525 = n9012 ^ n5980 ^ 1'b0 ;
  assign n17526 = n7554 & n17525 ;
  assign n17527 = n17526 ^ n8943 ^ 1'b0 ;
  assign n17528 = n919 | n6651 ;
  assign n17529 = n9883 & ~n17528 ;
  assign n17530 = n12818 ^ n9042 ^ n508 ;
  assign n17531 = ( n2667 & n17529 ) | ( n2667 & ~n17530 ) | ( n17529 & ~n17530 ) ;
  assign n17532 = n800 | n8503 ;
  assign n17533 = n17532 ^ n8363 ^ 1'b0 ;
  assign n17534 = ( ~n6938 & n14799 ) | ( ~n6938 & n17533 ) | ( n14799 & n17533 ) ;
  assign n17535 = n7219 | n17534 ;
  assign n17536 = n9807 ^ n5257 ^ n3538 ;
  assign n17537 = n17536 ^ n16408 ^ x132 ;
  assign n17538 = n10543 ^ n7242 ^ n2536 ;
  assign n17539 = ( n2108 & n2526 ) | ( n2108 & n14266 ) | ( n2526 & n14266 ) ;
  assign n17540 = ( n2406 & n5609 ) | ( n2406 & ~n14600 ) | ( n5609 & ~n14600 ) ;
  assign n17541 = n17540 ^ n11424 ^ n8122 ;
  assign n17542 = ( n1711 & ~n4779 ) | ( n1711 & n17541 ) | ( ~n4779 & n17541 ) ;
  assign n17543 = ( ~n7449 & n16278 ) | ( ~n7449 & n17542 ) | ( n16278 & n17542 ) ;
  assign n17544 = n5937 & ~n17543 ;
  assign n17545 = n10230 ^ n1418 ^ 1'b0 ;
  assign n17546 = n16147 & ~n17545 ;
  assign n17547 = ( n3854 & ~n3911 ) | ( n3854 & n11656 ) | ( ~n3911 & n11656 ) ;
  assign n17548 = ( x27 & ~n10334 ) | ( x27 & n17547 ) | ( ~n10334 & n17547 ) ;
  assign n17553 = n12944 & n17188 ;
  assign n17550 = n4057 ^ n1977 ^ n1833 ;
  assign n17549 = ( ~n865 & n14150 ) | ( ~n865 & n16551 ) | ( n14150 & n16551 ) ;
  assign n17551 = n17550 ^ n17549 ^ n11097 ;
  assign n17552 = ( ~x217 & n8610 ) | ( ~x217 & n17551 ) | ( n8610 & n17551 ) ;
  assign n17554 = n17553 ^ n17552 ^ n2888 ;
  assign n17555 = n8370 & ~n12413 ;
  assign n17556 = n14114 & n17555 ;
  assign n17557 = ( n8595 & ~n12015 ) | ( n8595 & n17556 ) | ( ~n12015 & n17556 ) ;
  assign n17558 = ( n2509 & n4935 ) | ( n2509 & n17557 ) | ( n4935 & n17557 ) ;
  assign n17559 = n7594 & n10211 ;
  assign n17560 = n4529 | n17559 ;
  assign n17561 = n17560 ^ n9346 ^ n8411 ;
  assign n17562 = ( n8064 & n17558 ) | ( n8064 & n17561 ) | ( n17558 & n17561 ) ;
  assign n17563 = ( n5562 & n5668 ) | ( n5562 & ~n13784 ) | ( n5668 & ~n13784 ) ;
  assign n17564 = n10643 ^ n5016 ^ n394 ;
  assign n17565 = n2948 & ~n8161 ;
  assign n17566 = n17565 ^ n8356 ^ 1'b0 ;
  assign n17567 = ( n15850 & n17564 ) | ( n15850 & n17566 ) | ( n17564 & n17566 ) ;
  assign n17568 = ( n3073 & ~n8690 ) | ( n3073 & n12212 ) | ( ~n8690 & n12212 ) ;
  assign n17569 = ( n4931 & n14758 ) | ( n4931 & n17568 ) | ( n14758 & n17568 ) ;
  assign n17570 = ( n17563 & n17567 ) | ( n17563 & ~n17569 ) | ( n17567 & ~n17569 ) ;
  assign n17571 = ( n2074 & n17562 ) | ( n2074 & ~n17570 ) | ( n17562 & ~n17570 ) ;
  assign n17572 = ~x74 & n3859 ;
  assign n17574 = n7017 ^ n2233 ^ n1827 ;
  assign n17573 = n3387 | n7452 ;
  assign n17575 = n17574 ^ n17573 ^ n14426 ;
  assign n17581 = n1745 & ~n7691 ;
  assign n17582 = n17581 ^ n15298 ^ 1'b0 ;
  assign n17583 = ( n7847 & n7854 ) | ( n7847 & n17582 ) | ( n7854 & n17582 ) ;
  assign n17584 = ( n3385 & n8610 ) | ( n3385 & n17583 ) | ( n8610 & n17583 ) ;
  assign n17585 = ( n1210 & n3424 ) | ( n1210 & ~n17584 ) | ( n3424 & ~n17584 ) ;
  assign n17576 = ( ~n2923 & n4836 ) | ( ~n2923 & n8917 ) | ( n4836 & n8917 ) ;
  assign n17577 = n17576 ^ n13611 ^ n3751 ;
  assign n17578 = n8530 | n10007 ;
  assign n17579 = ~n17577 & n17578 ;
  assign n17580 = n17579 ^ n4040 ^ 1'b0 ;
  assign n17586 = n17585 ^ n17580 ^ n4822 ;
  assign n17587 = ( n287 & n380 ) | ( n287 & n834 ) | ( n380 & n834 ) ;
  assign n17588 = n17587 ^ n3180 ^ 1'b0 ;
  assign n17589 = ( n1433 & n13347 ) | ( n1433 & n17588 ) | ( n13347 & n17588 ) ;
  assign n17590 = ~n2880 & n15436 ;
  assign n17591 = ~n10041 & n11842 ;
  assign n17592 = n17590 & ~n17591 ;
  assign n17593 = n10958 ^ n6790 ^ 1'b0 ;
  assign n17594 = ~n648 & n4749 ;
  assign n17595 = n17594 ^ n1673 ^ 1'b0 ;
  assign n17596 = n16908 | n17595 ;
  assign n17597 = n17593 | n17596 ;
  assign n17598 = ( n1077 & n2069 ) | ( n1077 & ~n2096 ) | ( n2069 & ~n2096 ) ;
  assign n17599 = n5009 | n7757 ;
  assign n17600 = n17599 ^ n7814 ^ 1'b0 ;
  assign n17601 = n17600 ^ n9398 ^ 1'b0 ;
  assign n17602 = n17598 & n17601 ;
  assign n17603 = ~n17148 & n17602 ;
  assign n17611 = ( x158 & n636 ) | ( x158 & n14507 ) | ( n636 & n14507 ) ;
  assign n17612 = n4405 | n10486 ;
  assign n17613 = ( n1629 & n4101 ) | ( n1629 & n17612 ) | ( n4101 & n17612 ) ;
  assign n17614 = n17613 ^ n11658 ^ n2047 ;
  assign n17615 = ( n3222 & n17611 ) | ( n3222 & ~n17614 ) | ( n17611 & ~n17614 ) ;
  assign n17604 = n13960 ^ n2918 ^ 1'b0 ;
  assign n17607 = ( n3936 & n4340 ) | ( n3936 & ~n6366 ) | ( n4340 & ~n6366 ) ;
  assign n17605 = n15212 ^ n14628 ^ n8286 ;
  assign n17606 = n17605 ^ n15301 ^ n6184 ;
  assign n17608 = n17607 ^ n17606 ^ n1748 ;
  assign n17609 = ( n4415 & n17604 ) | ( n4415 & ~n17608 ) | ( n17604 & ~n17608 ) ;
  assign n17610 = n13651 & ~n17609 ;
  assign n17616 = n17615 ^ n17610 ^ n10108 ;
  assign n17617 = n16337 ^ n5104 ^ 1'b0 ;
  assign n17618 = n1999 | n17617 ;
  assign n17619 = n8907 ^ x6 ^ 1'b0 ;
  assign n17621 = ( n719 & n1421 ) | ( n719 & n3260 ) | ( n1421 & n3260 ) ;
  assign n17622 = n17621 ^ x147 ^ 1'b0 ;
  assign n17623 = ~n15368 & n17622 ;
  assign n17620 = n12663 ^ n7973 ^ n2515 ;
  assign n17624 = n17623 ^ n17620 ^ n6613 ;
  assign n17625 = ( n7390 & n12798 ) | ( n7390 & ~n17624 ) | ( n12798 & ~n17624 ) ;
  assign n17626 = n7439 ^ n3135 ^ 1'b0 ;
  assign n17627 = ( n3728 & n17324 ) | ( n3728 & ~n17626 ) | ( n17324 & ~n17626 ) ;
  assign n17628 = ~n10262 & n17627 ;
  assign n17629 = n17628 ^ n11509 ^ 1'b0 ;
  assign n17630 = n534 & n14240 ;
  assign n17631 = n17630 ^ n8206 ^ n5162 ;
  assign n17632 = n2160 & n8736 ;
  assign n17633 = ~n17631 & n17632 ;
  assign n17634 = ( n1420 & ~n7426 ) | ( n1420 & n7858 ) | ( ~n7426 & n7858 ) ;
  assign n17635 = n9948 ^ n3892 ^ 1'b0 ;
  assign n17636 = ( n1610 & n14715 ) | ( n1610 & n17635 ) | ( n14715 & n17635 ) ;
  assign n17637 = n5887 & ~n13886 ;
  assign n17638 = ~n5719 & n16709 ;
  assign n17639 = ~n6222 & n17638 ;
  assign n17640 = n8458 ^ n2714 ^ n982 ;
  assign n17641 = n15015 ^ n5279 ^ n777 ;
  assign n17642 = ~n5013 & n12699 ;
  assign n17643 = ~n17641 & n17642 ;
  assign n17644 = n14671 & ~n17643 ;
  assign n17645 = n17644 ^ n1100 ^ 1'b0 ;
  assign n17646 = ( n3360 & n17640 ) | ( n3360 & n17645 ) | ( n17640 & n17645 ) ;
  assign n17647 = ( n2273 & n5189 ) | ( n2273 & ~n9694 ) | ( n5189 & ~n9694 ) ;
  assign n17648 = n6959 & ~n17647 ;
  assign n17649 = ~n3251 & n17648 ;
  assign n17650 = n17649 ^ n13423 ^ 1'b0 ;
  assign n17651 = n15845 ^ n2983 ^ x4 ;
  assign n17652 = n7567 ^ n6130 ^ 1'b0 ;
  assign n17653 = ( n1497 & n17651 ) | ( n1497 & ~n17652 ) | ( n17651 & ~n17652 ) ;
  assign n17654 = n17653 ^ n13663 ^ 1'b0 ;
  assign n17655 = n14449 ^ n4198 ^ 1'b0 ;
  assign n17656 = n9774 & ~n17655 ;
  assign n17657 = n14348 & n17656 ;
  assign n17658 = n10372 | n17657 ;
  assign n17659 = n8186 ^ n5080 ^ 1'b0 ;
  assign n17660 = ( ~n409 & n12264 ) | ( ~n409 & n17659 ) | ( n12264 & n17659 ) ;
  assign n17661 = ( ~n4048 & n12947 ) | ( ~n4048 & n17660 ) | ( n12947 & n17660 ) ;
  assign n17662 = ( ~n830 & n1197 ) | ( ~n830 & n4841 ) | ( n1197 & n4841 ) ;
  assign n17663 = n17662 ^ n16731 ^ n12118 ;
  assign n17665 = ( n747 & ~n4299 ) | ( n747 & n10622 ) | ( ~n4299 & n10622 ) ;
  assign n17666 = n17665 ^ n3536 ^ 1'b0 ;
  assign n17664 = n8187 & ~n16638 ;
  assign n17667 = n17666 ^ n17664 ^ n7640 ;
  assign n17668 = n2733 & ~n6023 ;
  assign n17669 = n1221 & n17668 ;
  assign n17670 = n2406 | n17669 ;
  assign n17671 = n17670 ^ n15378 ^ 1'b0 ;
  assign n17672 = n4844 & ~n5503 ;
  assign n17673 = n5836 ^ n4404 ^ n1029 ;
  assign n17675 = n7855 & ~n15821 ;
  assign n17674 = n5071 & ~n9840 ;
  assign n17676 = n17675 ^ n17674 ^ 1'b0 ;
  assign n17677 = n2802 ^ n494 ^ 1'b0 ;
  assign n17678 = n17677 ^ n13324 ^ n1126 ;
  assign n17679 = ( n5236 & n12628 ) | ( n5236 & ~n17678 ) | ( n12628 & ~n17678 ) ;
  assign n17683 = n15104 ^ n11302 ^ n1401 ;
  assign n17682 = n12183 ^ n8450 ^ n4947 ;
  assign n17680 = n4256 & ~n10966 ;
  assign n17681 = n10877 | n17680 ;
  assign n17684 = n17683 ^ n17682 ^ n17681 ;
  assign n17685 = ( ~n16099 & n16489 ) | ( ~n16099 & n17684 ) | ( n16489 & n17684 ) ;
  assign n17686 = n5484 ^ n3916 ^ n3581 ;
  assign n17687 = ( n2522 & n5080 ) | ( n2522 & ~n17686 ) | ( n5080 & ~n17686 ) ;
  assign n17688 = n16254 ^ n6917 ^ x6 ;
  assign n17689 = n11910 & ~n17688 ;
  assign n17690 = n17689 ^ n9472 ^ 1'b0 ;
  assign n17691 = n17690 ^ n7992 ^ n1971 ;
  assign n17692 = n17691 ^ n2226 ^ 1'b0 ;
  assign n17693 = ~n17687 & n17692 ;
  assign n17694 = ~n2759 & n7764 ;
  assign n17695 = n17694 ^ n5823 ^ n975 ;
  assign n17698 = n17265 ^ n6512 ^ 1'b0 ;
  assign n17699 = x164 & n17698 ;
  assign n17696 = n7905 & ~n14588 ;
  assign n17697 = ~n3303 & n17696 ;
  assign n17700 = n17699 ^ n17697 ^ 1'b0 ;
  assign n17701 = n9670 & ~n17700 ;
  assign n17702 = ( ~n6208 & n17695 ) | ( ~n6208 & n17701 ) | ( n17695 & n17701 ) ;
  assign n17703 = ( n2777 & n17693 ) | ( n2777 & n17702 ) | ( n17693 & n17702 ) ;
  assign n17704 = ( ~n280 & n5915 ) | ( ~n280 & n15352 ) | ( n5915 & n15352 ) ;
  assign n17705 = n17704 ^ n9765 ^ n5392 ;
  assign n17706 = n12128 ^ n4380 ^ 1'b0 ;
  assign n17707 = n12044 ^ n6957 ^ n484 ;
  assign n17708 = ( ~n8102 & n8717 ) | ( ~n8102 & n17707 ) | ( n8717 & n17707 ) ;
  assign n17709 = n17501 ^ n10285 ^ n4665 ;
  assign n17710 = n14203 ^ n13421 ^ n8357 ;
  assign n17711 = n8067 & n17710 ;
  assign n17712 = n17711 ^ n3038 ^ 1'b0 ;
  assign n17713 = n8235 ^ n5187 ^ n1202 ;
  assign n17714 = ~n7069 & n17713 ;
  assign n17715 = ~n13310 & n17714 ;
  assign n17716 = n5833 & ~n6615 ;
  assign n17717 = n2914 & n17716 ;
  assign n17718 = n15888 ^ n15255 ^ n2629 ;
  assign n17719 = n10943 ^ n6643 ^ n667 ;
  assign n17720 = ( n12151 & n12625 ) | ( n12151 & n17707 ) | ( n12625 & n17707 ) ;
  assign n17721 = n16390 ^ n15218 ^ n5690 ;
  assign n17722 = n13425 ^ n5292 ^ n2195 ;
  assign n17723 = n17722 ^ n8175 ^ n707 ;
  assign n17724 = n696 & ~n6525 ;
  assign n17725 = n17490 & n17724 ;
  assign n17726 = n15786 ^ n1307 ^ 1'b0 ;
  assign n17727 = n17726 ^ n12944 ^ n9153 ;
  assign n17728 = n1140 & n8311 ;
  assign n17730 = n3948 ^ n1899 ^ n446 ;
  assign n17731 = n17730 ^ n4257 ^ n1738 ;
  assign n17732 = ( n7728 & ~n10849 ) | ( n7728 & n17731 ) | ( ~n10849 & n17731 ) ;
  assign n17733 = n17732 ^ n1938 ^ 1'b0 ;
  assign n17729 = n5458 | n7817 ;
  assign n17734 = n17733 ^ n17729 ^ 1'b0 ;
  assign n17735 = ~n8532 & n13936 ;
  assign n17736 = n17734 & n17735 ;
  assign n17737 = ( n16171 & ~n17728 ) | ( n16171 & n17736 ) | ( ~n17728 & n17736 ) ;
  assign n17738 = n17727 | n17737 ;
  assign n17739 = ( n5062 & n5743 ) | ( n5062 & ~n8237 ) | ( n5743 & ~n8237 ) ;
  assign n17741 = n9387 ^ n5602 ^ n4275 ;
  assign n17740 = n4017 & n14324 ;
  assign n17742 = n17741 ^ n17740 ^ 1'b0 ;
  assign n17743 = ~n17739 & n17742 ;
  assign n17744 = n17743 ^ n5484 ^ 1'b0 ;
  assign n17745 = n9913 & n17744 ;
  assign n17746 = ( n17725 & ~n17738 ) | ( n17725 & n17745 ) | ( ~n17738 & n17745 ) ;
  assign n17747 = n1124 ^ n708 ^ 1'b0 ;
  assign n17748 = n14174 ^ n7164 ^ n6182 ;
  assign n17749 = ( n13845 & ~n17747 ) | ( n13845 & n17748 ) | ( ~n17747 & n17748 ) ;
  assign n17750 = ( n2517 & ~n13003 ) | ( n2517 & n17749 ) | ( ~n13003 & n17749 ) ;
  assign n17753 = ( ~n3479 & n7118 ) | ( ~n3479 & n10356 ) | ( n7118 & n10356 ) ;
  assign n17754 = ( n2825 & ~n6601 ) | ( n2825 & n17753 ) | ( ~n6601 & n17753 ) ;
  assign n17752 = ( ~n3345 & n4192 ) | ( ~n3345 & n4217 ) | ( n4192 & n4217 ) ;
  assign n17751 = n10914 ^ n7982 ^ n2303 ;
  assign n17755 = n17754 ^ n17752 ^ n17751 ;
  assign n17756 = ( n3976 & n11515 ) | ( n3976 & n17570 ) | ( n11515 & n17570 ) ;
  assign n17757 = n11106 & ~n16181 ;
  assign n17760 = n10140 ^ n500 ^ 1'b0 ;
  assign n17758 = n6317 ^ n4718 ^ n631 ;
  assign n17759 = n17758 ^ n11166 ^ n4372 ;
  assign n17761 = n17760 ^ n17759 ^ 1'b0 ;
  assign n17762 = ~n17757 & n17761 ;
  assign n17771 = n2974 & ~n3227 ;
  assign n17772 = n15406 & n17771 ;
  assign n17773 = n17772 ^ n13015 ^ n3836 ;
  assign n17769 = n16573 ^ n8846 ^ n1614 ;
  assign n17763 = n849 ^ n698 ^ 1'b0 ;
  assign n17764 = n12300 & ~n17763 ;
  assign n17765 = ( x136 & n8459 ) | ( x136 & ~n14007 ) | ( n8459 & ~n14007 ) ;
  assign n17766 = n17765 ^ n12238 ^ 1'b0 ;
  assign n17767 = ( n10473 & n17764 ) | ( n10473 & n17766 ) | ( n17764 & n17766 ) ;
  assign n17768 = n12940 & ~n17767 ;
  assign n17770 = n17769 ^ n17768 ^ 1'b0 ;
  assign n17774 = n17773 ^ n17770 ^ n6693 ;
  assign n17775 = n11106 ^ n7990 ^ n3431 ;
  assign n17776 = n17775 ^ n11769 ^ n5819 ;
  assign n17777 = n5387 | n17776 ;
  assign n17778 = n17777 ^ n17279 ^ n10187 ;
  assign n17779 = n3053 ^ n1534 ^ 1'b0 ;
  assign n17780 = n755 | n12688 ;
  assign n17781 = n11048 | n17780 ;
  assign n17782 = n16542 ^ n15663 ^ 1'b0 ;
  assign n17783 = ( n1408 & n6477 ) | ( n1408 & ~n15049 ) | ( n6477 & ~n15049 ) ;
  assign n17784 = ( ~n2266 & n8056 ) | ( ~n2266 & n12920 ) | ( n8056 & n12920 ) ;
  assign n17785 = ( n11307 & n13292 ) | ( n11307 & n17784 ) | ( n13292 & n17784 ) ;
  assign n17786 = ( n15330 & n17783 ) | ( n15330 & ~n17785 ) | ( n17783 & ~n17785 ) ;
  assign n17787 = n14995 ^ n4202 ^ 1'b0 ;
  assign n17789 = n2060 | n7397 ;
  assign n17790 = n14379 & ~n17789 ;
  assign n17791 = n2760 | n17790 ;
  assign n17792 = n17791 ^ n5988 ^ 1'b0 ;
  assign n17788 = n4169 & n8885 ;
  assign n17793 = n17792 ^ n17788 ^ 1'b0 ;
  assign n17794 = n13892 & ~n17793 ;
  assign n17795 = n17794 ^ n14545 ^ 1'b0 ;
  assign n17796 = n17795 ^ n14369 ^ n8039 ;
  assign n17797 = n12409 ^ n11071 ^ 1'b0 ;
  assign n17798 = ~x108 & n17797 ;
  assign n17799 = ~n10291 & n17798 ;
  assign n17800 = n17799 ^ n5893 ^ 1'b0 ;
  assign n17801 = ( ~n10873 & n11345 ) | ( ~n10873 & n16156 ) | ( n11345 & n16156 ) ;
  assign n17802 = ( n5489 & n7909 ) | ( n5489 & n10787 ) | ( n7909 & n10787 ) ;
  assign n17803 = ( n17800 & n17801 ) | ( n17800 & ~n17802 ) | ( n17801 & ~n17802 ) ;
  assign n17804 = ( ~n3469 & n16632 ) | ( ~n3469 & n17803 ) | ( n16632 & n17803 ) ;
  assign n17805 = ~n3469 & n15381 ;
  assign n17806 = ( ~n898 & n6134 ) | ( ~n898 & n16313 ) | ( n6134 & n16313 ) ;
  assign n17807 = n883 & ~n4327 ;
  assign n17808 = n17807 ^ n6146 ^ 1'b0 ;
  assign n17809 = n793 & n7820 ;
  assign n17810 = ~n10823 & n17809 ;
  assign n17811 = ( n3947 & n5079 ) | ( n3947 & n17810 ) | ( n5079 & n17810 ) ;
  assign n17812 = n8462 ^ n6404 ^ n1477 ;
  assign n17813 = ( n10942 & n13973 ) | ( n10942 & n17812 ) | ( n13973 & n17812 ) ;
  assign n17815 = n7097 | n15575 ;
  assign n17816 = n17815 ^ n7297 ^ 1'b0 ;
  assign n17817 = n17816 ^ n11314 ^ n7765 ;
  assign n17814 = n3149 & n14795 ;
  assign n17818 = n17817 ^ n17814 ^ 1'b0 ;
  assign n17819 = n5844 ^ n5372 ^ n3753 ;
  assign n17820 = n17819 ^ n12027 ^ 1'b0 ;
  assign n17821 = n1185 & n17820 ;
  assign n17822 = n15049 ^ n9534 ^ n5680 ;
  assign n17823 = n17822 ^ n7111 ^ 1'b0 ;
  assign n17826 = ( n3371 & ~n3386 ) | ( n3371 & n12001 ) | ( ~n3386 & n12001 ) ;
  assign n17827 = ( n1793 & n2332 ) | ( n1793 & ~n17826 ) | ( n2332 & ~n17826 ) ;
  assign n17824 = n6408 ^ n2228 ^ n336 ;
  assign n17825 = n12183 & ~n17824 ;
  assign n17828 = n17827 ^ n17825 ^ 1'b0 ;
  assign n17829 = ( ~x61 & n527 ) | ( ~x61 & n5990 ) | ( n527 & n5990 ) ;
  assign n17830 = n17829 ^ n4194 ^ n1925 ;
  assign n17831 = n1688 & n1944 ;
  assign n17832 = ~n5841 & n17831 ;
  assign n17833 = n17830 | n17832 ;
  assign n17834 = n8140 ^ n5737 ^ n2657 ;
  assign n17835 = n17834 ^ n10452 ^ n4417 ;
  assign n17836 = ( ~n6294 & n12883 ) | ( ~n6294 & n17835 ) | ( n12883 & n17835 ) ;
  assign n17840 = ( n2586 & ~n7004 ) | ( n2586 & n7690 ) | ( ~n7004 & n7690 ) ;
  assign n17841 = n17840 ^ n5275 ^ n2714 ;
  assign n17837 = n14581 ^ n6234 ^ n5745 ;
  assign n17838 = n7101 & n17837 ;
  assign n17839 = n17838 ^ n15659 ^ n12669 ;
  assign n17842 = n17841 ^ n17839 ^ n12938 ;
  assign n17845 = n7371 ^ n1753 ^ n1695 ;
  assign n17843 = n7468 ^ n3910 ^ 1'b0 ;
  assign n17844 = n17843 ^ n4537 ^ n1299 ;
  assign n17846 = n17845 ^ n17844 ^ 1'b0 ;
  assign n17847 = n11398 & ~n13796 ;
  assign n17848 = ~n15644 & n17847 ;
  assign n17849 = n9825 | n10841 ;
  assign n17850 = ~n1182 & n17849 ;
  assign n17851 = n14057 ^ n8100 ^ n496 ;
  assign n17852 = n17851 ^ n278 ^ 1'b0 ;
  assign n17853 = ~n10827 & n17852 ;
  assign n17854 = n11718 & n17853 ;
  assign n17858 = n17529 ^ n12262 ^ 1'b0 ;
  assign n17855 = ( ~n3009 & n3387 ) | ( ~n3009 & n9349 ) | ( n3387 & n9349 ) ;
  assign n17856 = n17855 ^ n11312 ^ 1'b0 ;
  assign n17857 = ( ~n3090 & n15711 ) | ( ~n3090 & n17856 ) | ( n15711 & n17856 ) ;
  assign n17859 = n17858 ^ n17857 ^ n1697 ;
  assign n17860 = n16057 ^ n15961 ^ 1'b0 ;
  assign n17861 = n10609 ^ n8760 ^ n5380 ;
  assign n17862 = ( n5750 & ~n7400 ) | ( n5750 & n17861 ) | ( ~n7400 & n17861 ) ;
  assign n17864 = ( n10242 & ~n12614 ) | ( n10242 & n16158 ) | ( ~n12614 & n16158 ) ;
  assign n17863 = x91 & ~n15363 ;
  assign n17865 = n17864 ^ n17863 ^ n4676 ;
  assign n17866 = n3948 & ~n4289 ;
  assign n17871 = n2427 | n7487 ;
  assign n17872 = n17871 ^ n3266 ^ 1'b0 ;
  assign n17869 = ( n4015 & ~n11780 ) | ( n4015 & n16278 ) | ( ~n11780 & n16278 ) ;
  assign n17868 = n15444 ^ n9635 ^ n2366 ;
  assign n17867 = n5552 ^ n3007 ^ 1'b0 ;
  assign n17870 = n17869 ^ n17868 ^ n17867 ;
  assign n17873 = n17872 ^ n17870 ^ n2976 ;
  assign n17874 = ( n16810 & n17734 ) | ( n16810 & ~n17873 ) | ( n17734 & ~n17873 ) ;
  assign n17875 = n4079 | n10519 ;
  assign n17877 = n3063 & n3936 ;
  assign n17878 = n17877 ^ n7089 ^ n6814 ;
  assign n17876 = ~n10665 & n13279 ;
  assign n17879 = n17878 ^ n17876 ^ n11750 ;
  assign n17880 = n8016 ^ n5878 ^ n987 ;
  assign n17881 = ~n1283 & n17880 ;
  assign n17882 = ~n2883 & n2993 ;
  assign n17883 = n2045 & n17882 ;
  assign n17884 = n4850 & n17883 ;
  assign n17885 = n17884 ^ n12111 ^ n7855 ;
  assign n17886 = n17183 ^ n9300 ^ 1'b0 ;
  assign n17887 = ~n10990 & n17886 ;
  assign n17888 = n15104 & n17887 ;
  assign n17889 = n3973 & n17888 ;
  assign n17890 = n8532 | n17108 ;
  assign n17891 = n17889 & ~n17890 ;
  assign n17892 = n3775 ^ n2084 ^ 1'b0 ;
  assign n17893 = n17892 ^ n8300 ^ n5444 ;
  assign n17894 = ( n12152 & n13427 ) | ( n12152 & n15089 ) | ( n13427 & n15089 ) ;
  assign n17895 = ( n9707 & n17893 ) | ( n9707 & ~n17894 ) | ( n17893 & ~n17894 ) ;
  assign n17896 = n7699 ^ n7120 ^ 1'b0 ;
  assign n17897 = ~n15108 & n17896 ;
  assign n17898 = n17897 ^ n16132 ^ n12181 ;
  assign n17899 = ( ~n8031 & n8927 ) | ( ~n8031 & n14275 ) | ( n8927 & n14275 ) ;
  assign n17901 = n4097 & n9829 ;
  assign n17902 = n17901 ^ n1639 ^ 1'b0 ;
  assign n17900 = n15830 ^ n13794 ^ n6068 ;
  assign n17903 = n17902 ^ n17900 ^ 1'b0 ;
  assign n17904 = ~n17899 & n17903 ;
  assign n17905 = n17784 ^ n6466 ^ n2506 ;
  assign n17907 = n7690 ^ n7086 ^ 1'b0 ;
  assign n17908 = n16888 ^ n9413 ^ 1'b0 ;
  assign n17909 = ( n3454 & n17907 ) | ( n3454 & ~n17908 ) | ( n17907 & ~n17908 ) ;
  assign n17910 = n10765 | n17909 ;
  assign n17906 = n5398 ^ n4397 ^ 1'b0 ;
  assign n17911 = n17910 ^ n17906 ^ n12669 ;
  assign n17912 = ~n773 & n2918 ;
  assign n17913 = n17912 ^ n1493 ^ 1'b0 ;
  assign n17914 = n17913 ^ n10601 ^ n1385 ;
  assign n17915 = n11962 & n17914 ;
  assign n17916 = n6936 & ~n17915 ;
  assign n17917 = n17916 ^ n14232 ^ 1'b0 ;
  assign n17918 = x254 & n9162 ;
  assign n17919 = n17918 ^ n11759 ^ n5544 ;
  assign n17920 = ( n9637 & n17917 ) | ( n9637 & n17919 ) | ( n17917 & n17919 ) ;
  assign n17921 = n6925 & n13203 ;
  assign n17922 = ~n4489 & n7227 ;
  assign n17923 = n17922 ^ n12358 ^ n7684 ;
  assign n17924 = n17923 ^ n12248 ^ n8811 ;
  assign n17925 = n14226 ^ n9955 ^ n5216 ;
  assign n17926 = n9104 | n17925 ;
  assign n17927 = n13170 | n17926 ;
  assign n17934 = n6255 ^ n6034 ^ 1'b0 ;
  assign n17935 = n9444 & ~n17934 ;
  assign n17932 = ~n5192 & n16778 ;
  assign n17933 = n17932 ^ n10631 ^ 1'b0 ;
  assign n17936 = n17935 ^ n17933 ^ 1'b0 ;
  assign n17928 = ~n8904 & n14632 ;
  assign n17929 = n17928 ^ n5478 ^ 1'b0 ;
  assign n17930 = n17929 ^ n16152 ^ 1'b0 ;
  assign n17931 = n4328 | n17930 ;
  assign n17937 = n17936 ^ n17931 ^ n13999 ;
  assign n17938 = n2181 & ~n4482 ;
  assign n17939 = ~n3063 & n17938 ;
  assign n17940 = n10387 ^ n6442 ^ n1191 ;
  assign n17941 = n7585 ^ n5136 ^ 1'b0 ;
  assign n17942 = n11982 & n17941 ;
  assign n17943 = n17940 & n17942 ;
  assign n17945 = n1719 | n13303 ;
  assign n17944 = n12793 | n13592 ;
  assign n17946 = n17945 ^ n17944 ^ n11410 ;
  assign n17947 = ( n2104 & n4771 ) | ( n2104 & ~n17946 ) | ( n4771 & ~n17946 ) ;
  assign n17948 = n9855 & ~n17947 ;
  assign n17949 = n17948 ^ n3050 ^ 1'b0 ;
  assign n17950 = ( n1528 & n14243 ) | ( n1528 & n15817 ) | ( n14243 & n15817 ) ;
  assign n17951 = n17950 ^ n16988 ^ n4380 ;
  assign n17952 = n9040 & ~n17270 ;
  assign n17953 = ~n17951 & n17952 ;
  assign n17954 = n8023 ^ n3977 ^ 1'b0 ;
  assign n17955 = n5269 & n17954 ;
  assign n17956 = ~n3538 & n11087 ;
  assign n17957 = n17956 ^ n16400 ^ 1'b0 ;
  assign n17958 = ( ~n1390 & n3841 ) | ( ~n1390 & n17957 ) | ( n3841 & n17957 ) ;
  assign n17959 = ( ~x165 & n17955 ) | ( ~x165 & n17958 ) | ( n17955 & n17958 ) ;
  assign n17960 = n8441 ^ n6488 ^ n2525 ;
  assign n17961 = n11178 ^ n8532 ^ 1'b0 ;
  assign n17962 = n17960 & n17961 ;
  assign n17963 = ( n1236 & n3793 ) | ( n1236 & ~n17962 ) | ( n3793 & ~n17962 ) ;
  assign n17969 = ~n9568 & n13255 ;
  assign n17970 = n17969 ^ n7869 ^ 1'b0 ;
  assign n17967 = ( n1913 & n2610 ) | ( n1913 & ~n3111 ) | ( n2610 & ~n3111 ) ;
  assign n17968 = ( n2542 & ~n5701 ) | ( n2542 & n17967 ) | ( ~n5701 & n17967 ) ;
  assign n17964 = n13413 ^ n12304 ^ n7079 ;
  assign n17965 = ( ~n5626 & n11892 ) | ( ~n5626 & n17964 ) | ( n11892 & n17964 ) ;
  assign n17966 = ~n13380 & n17965 ;
  assign n17971 = n17970 ^ n17968 ^ n17966 ;
  assign n17979 = n2828 ^ n1206 ^ 1'b0 ;
  assign n17977 = n9387 ^ n4503 ^ n3835 ;
  assign n17974 = ( n3085 & n3529 ) | ( n3085 & ~n6309 ) | ( n3529 & ~n6309 ) ;
  assign n17972 = n7066 ^ n5657 ^ 1'b0 ;
  assign n17973 = n17972 ^ n6898 ^ n1598 ;
  assign n17975 = n17974 ^ n17973 ^ n3963 ;
  assign n17976 = n17975 ^ n10172 ^ n1588 ;
  assign n17978 = n17977 ^ n17976 ^ 1'b0 ;
  assign n17980 = n17979 ^ n17978 ^ 1'b0 ;
  assign n17983 = ( n2426 & n7992 ) | ( n2426 & n10238 ) | ( n7992 & n10238 ) ;
  assign n17981 = n11423 ^ n3054 ^ 1'b0 ;
  assign n17982 = ~n15476 & n17981 ;
  assign n17984 = n17983 ^ n17982 ^ n15997 ;
  assign n17986 = n10216 ^ n2547 ^ 1'b0 ;
  assign n17985 = n5326 ^ n4471 ^ x225 ;
  assign n17987 = n17986 ^ n17985 ^ 1'b0 ;
  assign n17988 = n5396 ^ n2352 ^ 1'b0 ;
  assign n17989 = ( n3207 & n6376 ) | ( n3207 & ~n8164 ) | ( n6376 & ~n8164 ) ;
  assign n17990 = n9747 ^ n6095 ^ n353 ;
  assign n17991 = ( n1347 & n8880 ) | ( n1347 & n12355 ) | ( n8880 & n12355 ) ;
  assign n17992 = ( ~n673 & n8630 ) | ( ~n673 & n17991 ) | ( n8630 & n17991 ) ;
  assign n17993 = ( ~n15314 & n15930 ) | ( ~n15314 & n17992 ) | ( n15930 & n17992 ) ;
  assign n17994 = ~n17990 & n17993 ;
  assign n17995 = n10725 ^ n6735 ^ n4858 ;
  assign n17996 = ( n1732 & n5462 ) | ( n1732 & n6246 ) | ( n5462 & n6246 ) ;
  assign n17997 = n13796 ^ n3218 ^ n3161 ;
  assign n17998 = ( n3438 & ~n4720 ) | ( n3438 & n6191 ) | ( ~n4720 & n6191 ) ;
  assign n17999 = ( n6160 & n6670 ) | ( n6160 & n17998 ) | ( n6670 & n17998 ) ;
  assign n18000 = n17999 ^ n5489 ^ n2962 ;
  assign n18001 = ( n3734 & n11680 ) | ( n3734 & ~n13079 ) | ( n11680 & ~n13079 ) ;
  assign n18002 = ( n15822 & n18000 ) | ( n15822 & ~n18001 ) | ( n18000 & ~n18001 ) ;
  assign n18003 = ( n3211 & n11587 ) | ( n3211 & ~n13132 ) | ( n11587 & ~n13132 ) ;
  assign n18004 = ( n1956 & ~n2835 ) | ( n1956 & n2888 ) | ( ~n2835 & n2888 ) ;
  assign n18005 = n18004 ^ n13504 ^ n5505 ;
  assign n18006 = n5603 & ~n18005 ;
  assign n18007 = n15522 ^ n7032 ^ 1'b0 ;
  assign n18008 = n6808 | n18007 ;
  assign n18009 = n6161 & ~n7441 ;
  assign n18010 = ~n6691 & n18009 ;
  assign n18011 = ( n2495 & ~n13894 ) | ( n2495 & n18010 ) | ( ~n13894 & n18010 ) ;
  assign n18012 = n14897 & ~n18011 ;
  assign n18013 = n17824 & n18012 ;
  assign n18014 = ( n4260 & n9083 ) | ( n4260 & n18013 ) | ( n9083 & n18013 ) ;
  assign n18015 = n18014 ^ n3697 ^ 1'b0 ;
  assign n18016 = ~n6210 & n18015 ;
  assign n18017 = n18016 ^ n17107 ^ n12530 ;
  assign n18018 = n3729 & ~n6959 ;
  assign n18019 = n3330 ^ x105 ^ 1'b0 ;
  assign n18020 = ( n2688 & n3407 ) | ( n2688 & n18019 ) | ( n3407 & n18019 ) ;
  assign n18021 = ( n7028 & n7821 ) | ( n7028 & n8371 ) | ( n7821 & n8371 ) ;
  assign n18022 = n14678 ^ n9756 ^ n2674 ;
  assign n18023 = n18022 ^ n10316 ^ 1'b0 ;
  assign n18024 = n18021 & n18023 ;
  assign n18025 = ( ~n759 & n1387 ) | ( ~n759 & n6901 ) | ( n1387 & n6901 ) ;
  assign n18026 = n12069 ^ n8229 ^ n1505 ;
  assign n18027 = ( n4537 & ~n18025 ) | ( n4537 & n18026 ) | ( ~n18025 & n18026 ) ;
  assign n18028 = ( n8014 & ~n17354 ) | ( n8014 & n18027 ) | ( ~n17354 & n18027 ) ;
  assign n18029 = ( n5304 & ~n7265 ) | ( n5304 & n7306 ) | ( ~n7265 & n7306 ) ;
  assign n18030 = n5275 ^ n4151 ^ n1188 ;
  assign n18031 = ( n1042 & ~n4311 ) | ( n1042 & n10022 ) | ( ~n4311 & n10022 ) ;
  assign n18032 = n18030 | n18031 ;
  assign n18033 = n6520 & n17914 ;
  assign n18034 = ( ~n18029 & n18032 ) | ( ~n18029 & n18033 ) | ( n18032 & n18033 ) ;
  assign n18036 = n10727 ^ n7925 ^ 1'b0 ;
  assign n18037 = n18036 ^ n5806 ^ 1'b0 ;
  assign n18038 = n5302 & n12562 ;
  assign n18039 = ( n16907 & n18037 ) | ( n16907 & ~n18038 ) | ( n18037 & ~n18038 ) ;
  assign n18035 = n7504 & ~n12421 ;
  assign n18040 = n18039 ^ n18035 ^ 1'b0 ;
  assign n18041 = ( ~x42 & n4084 ) | ( ~x42 & n8096 ) | ( n4084 & n8096 ) ;
  assign n18042 = n18041 ^ n6034 ^ 1'b0 ;
  assign n18043 = ~n11279 & n18042 ;
  assign n18044 = ~n3645 & n9150 ;
  assign n18045 = n4773 ^ n3799 ^ n1904 ;
  assign n18046 = ( n7751 & n18044 ) | ( n7751 & ~n18045 ) | ( n18044 & ~n18045 ) ;
  assign n18047 = n17902 ^ n6695 ^ n2754 ;
  assign n18054 = ( n8128 & ~n11131 ) | ( n8128 & n15049 ) | ( ~n11131 & n15049 ) ;
  assign n18055 = n15378 & ~n17772 ;
  assign n18056 = n18054 & n18055 ;
  assign n18048 = x171 & ~n2803 ;
  assign n18049 = n18048 ^ n10461 ^ 1'b0 ;
  assign n18050 = n18049 ^ n6508 ^ n4109 ;
  assign n18051 = ( ~n1369 & n14602 ) | ( ~n1369 & n18050 ) | ( n14602 & n18050 ) ;
  assign n18052 = ~n6851 & n18051 ;
  assign n18053 = n18052 ^ n14528 ^ 1'b0 ;
  assign n18057 = n18056 ^ n18053 ^ n14525 ;
  assign n18058 = ( n947 & ~n2964 ) | ( n947 & n8647 ) | ( ~n2964 & n8647 ) ;
  assign n18059 = ( n3414 & n4369 ) | ( n3414 & n18058 ) | ( n4369 & n18058 ) ;
  assign n18060 = n4945 ^ n461 ^ 1'b0 ;
  assign n18061 = ( ~x126 & n5598 ) | ( ~x126 & n11946 ) | ( n5598 & n11946 ) ;
  assign n18062 = ( x24 & ~n18060 ) | ( x24 & n18061 ) | ( ~n18060 & n18061 ) ;
  assign n18065 = n5417 & ~n8167 ;
  assign n18063 = n15456 ^ n15213 ^ 1'b0 ;
  assign n18064 = ~n7878 & n18063 ;
  assign n18066 = n18065 ^ n18064 ^ n9113 ;
  assign n18069 = n13603 ^ n10967 ^ 1'b0 ;
  assign n18067 = ( n6252 & ~n10090 ) | ( n6252 & n15954 ) | ( ~n10090 & n15954 ) ;
  assign n18068 = n15294 | n18067 ;
  assign n18070 = n18069 ^ n18068 ^ n7196 ;
  assign n18071 = n10924 ^ n1722 ^ 1'b0 ;
  assign n18072 = ( n3987 & n4741 ) | ( n3987 & ~n6117 ) | ( n4741 & ~n6117 ) ;
  assign n18073 = n18072 ^ n9908 ^ n8484 ;
  assign n18074 = n1951 | n18073 ;
  assign n18076 = n4415 | n4519 ;
  assign n18077 = n18076 ^ n7012 ^ 1'b0 ;
  assign n18078 = ( ~n5028 & n8403 ) | ( ~n5028 & n18077 ) | ( n8403 & n18077 ) ;
  assign n18079 = n18078 ^ n11617 ^ n1403 ;
  assign n18080 = n18079 ^ n13110 ^ n909 ;
  assign n18075 = ~n10292 & n14341 ;
  assign n18081 = n18080 ^ n18075 ^ n825 ;
  assign n18083 = n13384 ^ n6663 ^ 1'b0 ;
  assign n18084 = n7366 | n18083 ;
  assign n18082 = n16801 ^ n12793 ^ 1'b0 ;
  assign n18085 = n18084 ^ n18082 ^ 1'b0 ;
  assign n18086 = n3101 | n18085 ;
  assign n18087 = n6973 ^ n6938 ^ n2186 ;
  assign n18088 = ~n530 & n14053 ;
  assign n18089 = n18087 & n18088 ;
  assign n18091 = n9197 & ~n11811 ;
  assign n18092 = ~n12134 & n18091 ;
  assign n18090 = ~n4136 & n7954 ;
  assign n18093 = n18092 ^ n18090 ^ 1'b0 ;
  assign n18094 = n4713 ^ x67 ^ 1'b0 ;
  assign n18095 = n18094 ^ n3688 ^ n3083 ;
  assign n18096 = n8660 | n9480 ;
  assign n18097 = ( n4057 & n7153 ) | ( n4057 & ~n13130 ) | ( n7153 & ~n13130 ) ;
  assign n18098 = n2463 & ~n9146 ;
  assign n18099 = n6424 & n18098 ;
  assign n18100 = n1102 & n11722 ;
  assign n18101 = n6803 & n18100 ;
  assign n18102 = n6473 ^ n1058 ^ 1'b0 ;
  assign n18103 = ~n18101 & n18102 ;
  assign n18104 = ~n7444 & n18103 ;
  assign n18105 = ~n11369 & n18104 ;
  assign n18106 = n5582 & ~n6622 ;
  assign n18107 = ( n813 & n993 ) | ( n813 & n6290 ) | ( n993 & n6290 ) ;
  assign n18108 = n2750 & n8454 ;
  assign n18109 = ( ~n2157 & n18107 ) | ( ~n2157 & n18108 ) | ( n18107 & n18108 ) ;
  assign n18110 = n11956 ^ n3633 ^ 1'b0 ;
  assign n18111 = ( n6311 & ~n7282 ) | ( n6311 & n10156 ) | ( ~n7282 & n10156 ) ;
  assign n18112 = n18111 ^ n14597 ^ 1'b0 ;
  assign n18113 = ~n18110 & n18112 ;
  assign n18118 = n762 | n3911 ;
  assign n18119 = n13069 & ~n18118 ;
  assign n18116 = n13361 ^ n8855 ^ 1'b0 ;
  assign n18117 = n18116 ^ n6206 ^ n3622 ;
  assign n18114 = n9030 ^ n5090 ^ n4230 ;
  assign n18115 = n18114 ^ n7301 ^ n3706 ;
  assign n18120 = n18119 ^ n18117 ^ n18115 ;
  assign n18121 = n6908 & ~n18120 ;
  assign n18122 = n18121 ^ n16471 ^ 1'b0 ;
  assign n18125 = ( n2278 & n11794 ) | ( n2278 & n16749 ) | ( n11794 & n16749 ) ;
  assign n18126 = n18125 ^ n4967 ^ n3959 ;
  assign n18127 = ( n4093 & n17475 ) | ( n4093 & n18126 ) | ( n17475 & n18126 ) ;
  assign n18123 = n10232 ^ n9250 ^ 1'b0 ;
  assign n18124 = ~n4363 & n18123 ;
  assign n18128 = n18127 ^ n18124 ^ n4547 ;
  assign n18129 = n12889 ^ n12741 ^ 1'b0 ;
  assign n18130 = n5021 & ~n18129 ;
  assign n18131 = ~n16383 & n17892 ;
  assign n18132 = n9716 & ~n18131 ;
  assign n18133 = ~n18130 & n18132 ;
  assign n18134 = ( n2481 & n9910 ) | ( n2481 & ~n18133 ) | ( n9910 & ~n18133 ) ;
  assign n18135 = n13664 ^ n8099 ^ n982 ;
  assign n18136 = n14892 & n18135 ;
  assign n18137 = ~n4884 & n18136 ;
  assign n18138 = n5234 ^ n2546 ^ 1'b0 ;
  assign n18139 = n18138 ^ n14324 ^ n8484 ;
  assign n18140 = n18139 ^ n14763 ^ n3985 ;
  assign n18141 = ( ~n3311 & n6205 ) | ( ~n3311 & n13291 ) | ( n6205 & n13291 ) ;
  assign n18142 = n18141 ^ n12215 ^ 1'b0 ;
  assign n18143 = n4124 | n12157 ;
  assign n18144 = n18143 ^ n12019 ^ 1'b0 ;
  assign n18145 = n7289 ^ n2668 ^ 1'b0 ;
  assign n18146 = ~x163 & n18145 ;
  assign n18147 = n11379 ^ n5236 ^ x67 ;
  assign n18148 = x226 & ~n6943 ;
  assign n18149 = ~n7609 & n18148 ;
  assign n18150 = ( n8462 & n13465 ) | ( n8462 & ~n18149 ) | ( n13465 & ~n18149 ) ;
  assign n18151 = n18150 ^ n3542 ^ n2300 ;
  assign n18152 = n11757 ^ n10319 ^ n5230 ;
  assign n18153 = n16425 & n18152 ;
  assign n18154 = ( ~n983 & n6698 ) | ( ~n983 & n10342 ) | ( n6698 & n10342 ) ;
  assign n18155 = ( n864 & ~n3728 ) | ( n864 & n15777 ) | ( ~n3728 & n15777 ) ;
  assign n18156 = ( ~n1913 & n4828 ) | ( ~n1913 & n4875 ) | ( n4828 & n4875 ) ;
  assign n18157 = n7139 & ~n18156 ;
  assign n18158 = n18157 ^ n2920 ^ 1'b0 ;
  assign n18159 = n8760 & n18158 ;
  assign n18161 = ~n3399 & n6705 ;
  assign n18162 = n1433 & n18161 ;
  assign n18160 = n6591 | n15552 ;
  assign n18163 = n18162 ^ n18160 ^ 1'b0 ;
  assign n18164 = ( ~n1391 & n18159 ) | ( ~n1391 & n18163 ) | ( n18159 & n18163 ) ;
  assign n18165 = n6454 ^ n5110 ^ 1'b0 ;
  assign n18166 = n5842 & n18165 ;
  assign n18167 = ( n3884 & ~n8001 ) | ( n3884 & n18166 ) | ( ~n8001 & n18166 ) ;
  assign n18168 = n18167 ^ n9005 ^ 1'b0 ;
  assign n18169 = n7907 | n18168 ;
  assign n18170 = n11221 | n17161 ;
  assign n18171 = n10448 ^ n5056 ^ n1929 ;
  assign n18172 = n11817 & n18171 ;
  assign n18173 = ( n11141 & n18170 ) | ( n11141 & ~n18172 ) | ( n18170 & ~n18172 ) ;
  assign n18174 = ( n6535 & ~n18169 ) | ( n6535 & n18173 ) | ( ~n18169 & n18173 ) ;
  assign n18175 = ( n18155 & ~n18164 ) | ( n18155 & n18174 ) | ( ~n18164 & n18174 ) ;
  assign n18176 = n12069 ^ n2011 ^ x191 ;
  assign n18177 = n13161 & n18176 ;
  assign n18178 = n16501 ^ n3895 ^ 1'b0 ;
  assign n18179 = ~n16074 & n18178 ;
  assign n18180 = ( n14576 & ~n18177 ) | ( n14576 & n18179 ) | ( ~n18177 & n18179 ) ;
  assign n18182 = ( n798 & ~n5082 ) | ( n798 & n14899 ) | ( ~n5082 & n14899 ) ;
  assign n18183 = n18182 ^ n13719 ^ n500 ;
  assign n18184 = n18183 ^ n13573 ^ n4810 ;
  assign n18181 = n4143 & n7556 ;
  assign n18185 = n18184 ^ n18181 ^ n14278 ;
  assign n18186 = n12299 ^ n6074 ^ n1956 ;
  assign n18187 = ( n7930 & n11261 ) | ( n7930 & n18186 ) | ( n11261 & n18186 ) ;
  assign n18198 = n9883 ^ n3598 ^ 1'b0 ;
  assign n18199 = n18198 ^ n2166 ^ 1'b0 ;
  assign n18200 = n4924 & ~n18199 ;
  assign n18188 = n5690 ^ n1762 ^ x109 ;
  assign n18189 = ( x248 & ~n1085 ) | ( x248 & n18188 ) | ( ~n1085 & n18188 ) ;
  assign n18190 = n14660 ^ n1323 ^ n1243 ;
  assign n18191 = n16483 ^ n6150 ^ n1099 ;
  assign n18192 = ( n2795 & n18190 ) | ( n2795 & n18191 ) | ( n18190 & n18191 ) ;
  assign n18193 = ~n18189 & n18192 ;
  assign n18194 = n18193 ^ n11683 ^ 1'b0 ;
  assign n18195 = n18194 ^ n4889 ^ 1'b0 ;
  assign n18196 = n7563 & n13944 ;
  assign n18197 = ~n18195 & n18196 ;
  assign n18201 = n18200 ^ n18197 ^ n7783 ;
  assign n18202 = n1280 | n7873 ;
  assign n18203 = n18202 ^ n341 ^ 1'b0 ;
  assign n18204 = n5058 | n18203 ;
  assign n18205 = n5328 ^ n2592 ^ 1'b0 ;
  assign n18206 = n17877 & n18205 ;
  assign n18207 = n18206 ^ n2366 ^ 1'b0 ;
  assign n18208 = n18207 ^ n12247 ^ 1'b0 ;
  assign n18209 = n16454 | n18208 ;
  assign n18210 = ( n991 & n15435 ) | ( n991 & ~n18209 ) | ( n15435 & ~n18209 ) ;
  assign n18211 = ~n15181 & n18210 ;
  assign n18212 = n1558 & n18211 ;
  assign n18213 = n7635 & n18212 ;
  assign n18214 = n332 & n18185 ;
  assign n18215 = ( n7058 & ~n7457 ) | ( n7058 & n7972 ) | ( ~n7457 & n7972 ) ;
  assign n18216 = n18215 ^ n6885 ^ 1'b0 ;
  assign n18217 = n1064 & n18216 ;
  assign n18218 = ( n15015 & n15116 ) | ( n15015 & ~n18217 ) | ( n15116 & ~n18217 ) ;
  assign n18219 = n11208 ^ n9866 ^ n1980 ;
  assign n18222 = n13686 ^ n3151 ^ x23 ;
  assign n18223 = n18222 ^ n11030 ^ n3303 ;
  assign n18220 = n2442 & ~n2566 ;
  assign n18221 = ( n471 & ~n1636 ) | ( n471 & n18220 ) | ( ~n1636 & n18220 ) ;
  assign n18224 = n18223 ^ n18221 ^ n11228 ;
  assign n18225 = ( ~n3858 & n18219 ) | ( ~n3858 & n18224 ) | ( n18219 & n18224 ) ;
  assign n18226 = ~n7785 & n9392 ;
  assign n18227 = n4305 | n7539 ;
  assign n18228 = n5402 | n18227 ;
  assign n18229 = n15555 & n18228 ;
  assign n18230 = n18229 ^ n6064 ^ 1'b0 ;
  assign n18232 = n3884 & ~n11282 ;
  assign n18233 = n18232 ^ n6607 ^ n2816 ;
  assign n18231 = n8838 & n9403 ;
  assign n18234 = n18233 ^ n18231 ^ 1'b0 ;
  assign n18235 = n13009 ^ n12484 ^ 1'b0 ;
  assign n18236 = n5519 | n18235 ;
  assign n18237 = ~n6328 & n6337 ;
  assign n18238 = n18237 ^ n3356 ^ n267 ;
  assign n18239 = n18238 ^ n899 ^ 1'b0 ;
  assign n18245 = n5770 ^ n5395 ^ 1'b0 ;
  assign n18246 = n2140 & n18245 ;
  assign n18240 = n14172 ^ n9754 ^ n4934 ;
  assign n18241 = n3307 | n7089 ;
  assign n18242 = n18241 ^ n14669 ^ n6814 ;
  assign n18243 = ( n4398 & ~n11374 ) | ( n4398 & n18242 ) | ( ~n11374 & n18242 ) ;
  assign n18244 = ~n18240 & n18243 ;
  assign n18247 = n18246 ^ n18244 ^ n5142 ;
  assign n18248 = ( ~n15672 & n18239 ) | ( ~n15672 & n18247 ) | ( n18239 & n18247 ) ;
  assign n18249 = n10150 & ~n13135 ;
  assign n18250 = n18249 ^ n14376 ^ 1'b0 ;
  assign n18251 = n18250 ^ n11511 ^ n10060 ;
  assign n18252 = n18251 ^ n15276 ^ n6669 ;
  assign n18253 = n6614 ^ n3765 ^ n1140 ;
  assign n18254 = n18253 ^ n16225 ^ n10094 ;
  assign n18255 = n9148 ^ n6827 ^ 1'b0 ;
  assign n18256 = ~n4240 & n16001 ;
  assign n18257 = n18256 ^ n494 ^ 1'b0 ;
  assign n18258 = ( ~n387 & n5259 ) | ( ~n387 & n9959 ) | ( n5259 & n9959 ) ;
  assign n18259 = n2871 & ~n13550 ;
  assign n18260 = n18258 & n18259 ;
  assign n18261 = n18257 & ~n18260 ;
  assign n18262 = n10394 ^ n360 ^ 1'b0 ;
  assign n18263 = ( n9344 & n14419 ) | ( n9344 & ~n16813 ) | ( n14419 & ~n16813 ) ;
  assign n18264 = n17183 ^ n6126 ^ n2650 ;
  assign n18265 = ( n929 & n3641 ) | ( n929 & ~n9510 ) | ( n3641 & ~n9510 ) ;
  assign n18266 = n1309 & ~n18265 ;
  assign n18267 = n18266 ^ n15091 ^ 1'b0 ;
  assign n18268 = n15941 ^ n3789 ^ 1'b0 ;
  assign n18269 = ( n633 & n6223 ) | ( n633 & ~n18268 ) | ( n6223 & ~n18268 ) ;
  assign n18270 = ( ~n2643 & n2847 ) | ( ~n2643 & n8482 ) | ( n2847 & n8482 ) ;
  assign n18271 = n11285 ^ n10912 ^ 1'b0 ;
  assign n18272 = ~n18270 & n18271 ;
  assign n18273 = n7029 | n10100 ;
  assign n18274 = ( n5589 & n7004 ) | ( n5589 & ~n17680 ) | ( n7004 & ~n17680 ) ;
  assign n18275 = n18274 ^ n13546 ^ n11688 ;
  assign n18276 = ( n11971 & n18273 ) | ( n11971 & ~n18275 ) | ( n18273 & ~n18275 ) ;
  assign n18277 = n8846 ^ n5192 ^ n2184 ;
  assign n18278 = n18277 ^ n15204 ^ n9530 ;
  assign n18279 = n5937 & n15628 ;
  assign n18280 = n6190 & n18279 ;
  assign n18281 = n18280 ^ n16590 ^ n10085 ;
  assign n18282 = n17397 ^ n10363 ^ 1'b0 ;
  assign n18283 = n18282 ^ n7567 ^ n1106 ;
  assign n18284 = n17339 ^ n13350 ^ 1'b0 ;
  assign n18285 = n18284 ^ n16238 ^ x90 ;
  assign n18286 = n18285 ^ n8093 ^ 1'b0 ;
  assign n18287 = n18283 | n18286 ;
  assign n18289 = n6184 & ~n10310 ;
  assign n18288 = ( n3483 & n11252 ) | ( n3483 & ~n16493 ) | ( n11252 & ~n16493 ) ;
  assign n18290 = n18289 ^ n18288 ^ n497 ;
  assign n18291 = n4468 | n6937 ;
  assign n18292 = ( n1000 & n2036 ) | ( n1000 & n6732 ) | ( n2036 & n6732 ) ;
  assign n18293 = n13121 | n16718 ;
  assign n18294 = ( n18291 & ~n18292 ) | ( n18291 & n18293 ) | ( ~n18292 & n18293 ) ;
  assign n18295 = n721 | n10623 ;
  assign n18296 = ( x180 & ~n6477 ) | ( x180 & n18295 ) | ( ~n6477 & n18295 ) ;
  assign n18297 = n8818 & n18296 ;
  assign n18298 = n1999 | n16405 ;
  assign n18299 = x13 & n18298 ;
  assign n18300 = n18299 ^ n3724 ^ 1'b0 ;
  assign n18301 = n18300 ^ n7875 ^ n5991 ;
  assign n18302 = n16241 ^ n11637 ^ n11012 ;
  assign n18303 = n10640 ^ n8627 ^ n6670 ;
  assign n18304 = ( n4306 & ~n6894 ) | ( n4306 & n18303 ) | ( ~n6894 & n18303 ) ;
  assign n18305 = n11318 ^ n8915 ^ n768 ;
  assign n18306 = n17241 ^ n12476 ^ n6976 ;
  assign n18307 = n5913 | n7249 ;
  assign n18308 = n17300 | n18307 ;
  assign n18309 = n18308 ^ n15359 ^ n5231 ;
  assign n18310 = n18306 & ~n18309 ;
  assign n18311 = n3103 | n12298 ;
  assign n18312 = n5737 & n16530 ;
  assign n18313 = n18312 ^ n5482 ^ 1'b0 ;
  assign n18314 = n18313 ^ n17462 ^ n7753 ;
  assign n18315 = ( ~n1206 & n10817 ) | ( ~n1206 & n11125 ) | ( n10817 & n11125 ) ;
  assign n18316 = n9039 ^ n7749 ^ 1'b0 ;
  assign n18317 = n683 & ~n18316 ;
  assign n18318 = n18315 & n18317 ;
  assign n18319 = n12240 | n18318 ;
  assign n18320 = n5558 | n18319 ;
  assign n18322 = n10021 ^ n9168 ^ n997 ;
  assign n18323 = n18322 ^ n3115 ^ 1'b0 ;
  assign n18324 = n13061 & n18323 ;
  assign n18321 = n4466 & n12219 ;
  assign n18325 = n18324 ^ n18321 ^ n2947 ;
  assign n18326 = n18325 ^ n15677 ^ n3106 ;
  assign n18327 = ( n3037 & n6246 ) | ( n3037 & n8073 ) | ( n6246 & n8073 ) ;
  assign n18328 = n15194 ^ n2621 ^ n2018 ;
  assign n18332 = n11476 ^ n10315 ^ n5552 ;
  assign n18329 = n16354 ^ n6885 ^ 1'b0 ;
  assign n18330 = n7121 & ~n18329 ;
  assign n18331 = ( ~n17737 & n18258 ) | ( ~n17737 & n18330 ) | ( n18258 & n18330 ) ;
  assign n18333 = n18332 ^ n18331 ^ n4963 ;
  assign n18334 = ( ~n6162 & n6572 ) | ( ~n6162 & n18059 ) | ( n6572 & n18059 ) ;
  assign n18335 = n14440 ^ n14175 ^ x196 ;
  assign n18336 = n17655 ^ n5722 ^ 1'b0 ;
  assign n18337 = n18335 & ~n18336 ;
  assign n18340 = x116 & ~n2643 ;
  assign n18341 = n3036 & n18340 ;
  assign n18338 = n1460 & ~n1538 ;
  assign n18339 = n11354 & n18338 ;
  assign n18342 = n18341 ^ n18339 ^ n9412 ;
  assign n18343 = n15273 ^ n14468 ^ n6788 ;
  assign n18344 = n3614 & ~n18343 ;
  assign n18345 = n18344 ^ n17051 ^ 1'b0 ;
  assign n18346 = ( n4156 & n4204 ) | ( n4156 & n18345 ) | ( n4204 & n18345 ) ;
  assign n18347 = n9237 ^ n6905 ^ n2370 ;
  assign n18348 = n18347 ^ n8030 ^ n488 ;
  assign n18349 = ( n3335 & n16197 ) | ( n3335 & ~n18348 ) | ( n16197 & ~n18348 ) ;
  assign n18350 = ~n1933 & n15191 ;
  assign n18351 = n18350 ^ n16018 ^ 1'b0 ;
  assign n18352 = ~n12072 & n13166 ;
  assign n18353 = ~n18351 & n18352 ;
  assign n18354 = n18353 ^ n16170 ^ 1'b0 ;
  assign n18358 = n14865 ^ n7130 ^ 1'b0 ;
  assign n18355 = n1141 & n4472 ;
  assign n18356 = n5525 & n18355 ;
  assign n18357 = ( n525 & ~n11461 ) | ( n525 & n18356 ) | ( ~n11461 & n18356 ) ;
  assign n18359 = n18358 ^ n18357 ^ 1'b0 ;
  assign n18360 = ( n2039 & n3622 ) | ( n2039 & ~n4460 ) | ( n3622 & ~n4460 ) ;
  assign n18361 = n18360 ^ n13513 ^ 1'b0 ;
  assign n18362 = ( ~n496 & n7959 ) | ( ~n496 & n18361 ) | ( n7959 & n18361 ) ;
  assign n18364 = x247 & n5308 ;
  assign n18363 = n2928 | n6970 ;
  assign n18365 = n18364 ^ n18363 ^ 1'b0 ;
  assign n18366 = ( n6919 & ~n9009 ) | ( n6919 & n18365 ) | ( ~n9009 & n18365 ) ;
  assign n18367 = n13200 ^ n12276 ^ 1'b0 ;
  assign n18368 = n7799 ^ n1813 ^ n619 ;
  assign n18371 = n9561 ^ n7473 ^ 1'b0 ;
  assign n18372 = n14237 & n18371 ;
  assign n18369 = n5759 ^ n4780 ^ n786 ;
  assign n18370 = n11076 & ~n18369 ;
  assign n18373 = n18372 ^ n18370 ^ 1'b0 ;
  assign n18374 = ( n4459 & n12102 ) | ( n4459 & n18373 ) | ( n12102 & n18373 ) ;
  assign n18375 = n5212 ^ n1570 ^ 1'b0 ;
  assign n18376 = n9507 & n18375 ;
  assign n18377 = n9335 | n12469 ;
  assign n18378 = ( ~n13908 & n17314 ) | ( ~n13908 & n18377 ) | ( n17314 & n18377 ) ;
  assign n18379 = n18376 & n18378 ;
  assign n18380 = n18374 & n18379 ;
  assign n18381 = n9183 ^ n4792 ^ n1542 ;
  assign n18383 = ~n1032 & n1195 ;
  assign n18384 = n587 & n18383 ;
  assign n18382 = x3 & ~n7310 ;
  assign n18385 = n18384 ^ n18382 ^ 1'b0 ;
  assign n18386 = ( n11667 & ~n12296 ) | ( n11667 & n18385 ) | ( ~n12296 & n18385 ) ;
  assign n18387 = n18381 & n18386 ;
  assign n18388 = n1949 & n5572 ;
  assign n18389 = ( n9347 & n17170 ) | ( n9347 & ~n18388 ) | ( n17170 & ~n18388 ) ;
  assign n18390 = n15574 ^ n6503 ^ n5291 ;
  assign n18391 = n6037 ^ n3909 ^ n2143 ;
  assign n18392 = n6719 & n15499 ;
  assign n18393 = n18391 & n18392 ;
  assign n18394 = n4320 ^ n3532 ^ 1'b0 ;
  assign n18395 = n13285 & n18394 ;
  assign n18396 = n18395 ^ n17255 ^ n13493 ;
  assign n18404 = n13000 ^ n5465 ^ 1'b0 ;
  assign n18401 = n1714 | n1871 ;
  assign n18402 = n18401 ^ n938 ^ 1'b0 ;
  assign n18403 = n18402 ^ n5717 ^ n1351 ;
  assign n18397 = n3766 | n12029 ;
  assign n18398 = n6469 | n10435 ;
  assign n18399 = n11718 | n18398 ;
  assign n18400 = n18397 & n18399 ;
  assign n18405 = n18404 ^ n18403 ^ n18400 ;
  assign n18406 = n18405 ^ n9410 ^ 1'b0 ;
  assign n18407 = ( n2842 & ~n9746 ) | ( n2842 & n10531 ) | ( ~n9746 & n10531 ) ;
  assign n18408 = n4856 & n13441 ;
  assign n18409 = n18408 ^ n706 ^ 1'b0 ;
  assign n18410 = ( n4468 & n16495 ) | ( n4468 & n18409 ) | ( n16495 & n18409 ) ;
  assign n18411 = ( n6187 & n7688 ) | ( n6187 & ~n13910 ) | ( n7688 & ~n13910 ) ;
  assign n18412 = n14235 ^ n5046 ^ 1'b0 ;
  assign n18413 = ( ~n2414 & n8684 ) | ( ~n2414 & n18412 ) | ( n8684 & n18412 ) ;
  assign n18415 = ~n7534 & n17391 ;
  assign n18416 = ~n4652 & n18415 ;
  assign n18414 = ( n4751 & ~n5673 ) | ( n4751 & n8847 ) | ( ~n5673 & n8847 ) ;
  assign n18417 = n18416 ^ n18414 ^ n8269 ;
  assign n18418 = ( n903 & n15379 ) | ( n903 & n18417 ) | ( n15379 & n18417 ) ;
  assign n18419 = n5737 ^ n2044 ^ 1'b0 ;
  assign n18420 = n9285 | n18419 ;
  assign n18421 = n6582 ^ n1958 ^ x112 ;
  assign n18422 = n438 | n18421 ;
  assign n18423 = n18422 ^ n10638 ^ 1'b0 ;
  assign n18424 = n15464 ^ n12955 ^ n7630 ;
  assign n18425 = n18423 | n18424 ;
  assign n18426 = n8922 | n18425 ;
  assign n18430 = n11015 ^ n3865 ^ 1'b0 ;
  assign n18431 = n10283 & n18430 ;
  assign n18432 = n18431 ^ n11056 ^ 1'b0 ;
  assign n18427 = n12065 ^ n11030 ^ n5308 ;
  assign n18428 = ( n6784 & ~n11342 ) | ( n6784 & n18427 ) | ( ~n11342 & n18427 ) ;
  assign n18429 = ~n9983 & n18428 ;
  assign n18433 = n18432 ^ n18429 ^ 1'b0 ;
  assign n18434 = n18433 ^ n9499 ^ 1'b0 ;
  assign n18441 = x75 & ~n3265 ;
  assign n18442 = n4037 & ~n18441 ;
  assign n18443 = n18442 ^ n13749 ^ 1'b0 ;
  assign n18438 = n13234 ^ x31 ^ 1'b0 ;
  assign n18439 = n4684 & ~n18438 ;
  assign n18435 = n1728 ^ n1154 ^ 1'b0 ;
  assign n18436 = n9602 | n18435 ;
  assign n18437 = n2465 & n18436 ;
  assign n18440 = n18439 ^ n18437 ^ 1'b0 ;
  assign n18444 = n18443 ^ n18440 ^ n9711 ;
  assign n18445 = n17123 ^ n16691 ^ x174 ;
  assign n18446 = n4874 | n7192 ;
  assign n18447 = n18446 ^ n17908 ^ 1'b0 ;
  assign n18448 = n11629 ^ n8869 ^ n1804 ;
  assign n18449 = n18448 ^ n13824 ^ n7069 ;
  assign n18450 = n18449 ^ n12358 ^ 1'b0 ;
  assign n18451 = n10914 & ~n13474 ;
  assign n18452 = ~n1741 & n18451 ;
  assign n18453 = n18452 ^ n11891 ^ n2633 ;
  assign n18454 = n1902 & ~n18453 ;
  assign n18455 = n14083 & n18454 ;
  assign n18456 = ( n1790 & n3315 ) | ( n1790 & n16411 ) | ( n3315 & n16411 ) ;
  assign n18457 = n14684 ^ n12216 ^ n12112 ;
  assign n18458 = n4451 & ~n18457 ;
  assign n18459 = n13707 & n18458 ;
  assign n18460 = ~n18456 & n18459 ;
  assign n18461 = n13347 ^ n12176 ^ n1014 ;
  assign n18462 = ( x38 & ~n1438 ) | ( x38 & n1920 ) | ( ~n1438 & n1920 ) ;
  assign n18463 = n18462 ^ n6217 ^ n3991 ;
  assign n18464 = n18417 ^ n9475 ^ 1'b0 ;
  assign n18465 = n18464 ^ n12849 ^ n7994 ;
  assign n18466 = n14304 & n16959 ;
  assign n18467 = n16635 & ~n18466 ;
  assign n18468 = n3918 & ~n9241 ;
  assign n18469 = ~n7856 & n18468 ;
  assign n18470 = x65 & ~n12412 ;
  assign n18471 = ( ~n8058 & n18469 ) | ( ~n8058 & n18470 ) | ( n18469 & n18470 ) ;
  assign n18472 = n16508 & n18471 ;
  assign n18473 = n18472 ^ n17208 ^ n1397 ;
  assign n18474 = n5259 & ~n11283 ;
  assign n18475 = ~n4184 & n7292 ;
  assign n18476 = ~n9205 & n18475 ;
  assign n18477 = n18476 ^ n12596 ^ 1'b0 ;
  assign n18478 = n4069 & n18477 ;
  assign n18479 = n2441 ^ n871 ^ n356 ;
  assign n18480 = ~n1378 & n11603 ;
  assign n18481 = n18480 ^ x128 ^ 1'b0 ;
  assign n18482 = ( n1796 & n18479 ) | ( n1796 & n18481 ) | ( n18479 & n18481 ) ;
  assign n18483 = n18482 ^ n16003 ^ n935 ;
  assign n18484 = n18483 ^ n15375 ^ n1000 ;
  assign n18485 = ( n2190 & n9255 ) | ( n2190 & n18484 ) | ( n9255 & n18484 ) ;
  assign n18487 = n7850 ^ n3053 ^ 1'b0 ;
  assign n18488 = ( n1225 & ~n5340 ) | ( n1225 & n18487 ) | ( ~n5340 & n18487 ) ;
  assign n18486 = n6103 | n11913 ;
  assign n18489 = n18488 ^ n18486 ^ 1'b0 ;
  assign n18490 = n18489 ^ n9506 ^ 1'b0 ;
  assign n18491 = ~n7305 & n18490 ;
  assign n18492 = n18491 ^ n6387 ^ 1'b0 ;
  assign n18493 = ( ~n1596 & n10087 ) | ( ~n1596 & n15204 ) | ( n10087 & n15204 ) ;
  assign n18494 = ( n1408 & n13926 ) | ( n1408 & ~n18493 ) | ( n13926 & ~n18493 ) ;
  assign n18495 = n8255 & ~n15356 ;
  assign n18496 = n16618 & n18495 ;
  assign n18497 = n2319 ^ n1431 ^ 1'b0 ;
  assign n18498 = n18497 ^ n18013 ^ 1'b0 ;
  assign n18499 = n4915 ^ n2411 ^ 1'b0 ;
  assign n18500 = ( ~n6459 & n8932 ) | ( ~n6459 & n12733 ) | ( n8932 & n12733 ) ;
  assign n18501 = n14700 ^ n1497 ^ n1003 ;
  assign n18502 = n18500 & n18501 ;
  assign n18503 = ( ~n17835 & n18499 ) | ( ~n17835 & n18502 ) | ( n18499 & n18502 ) ;
  assign n18504 = ( ~n14398 & n15889 ) | ( ~n14398 & n18280 ) | ( n15889 & n18280 ) ;
  assign n18505 = n7026 & n14348 ;
  assign n18506 = ~n1395 & n9859 ;
  assign n18507 = n15145 & ~n18506 ;
  assign n18508 = n18507 ^ n17121 ^ 1'b0 ;
  assign n18509 = n3267 ^ n2987 ^ n1676 ;
  assign n18510 = n11943 ^ n9344 ^ n5498 ;
  assign n18511 = n18510 ^ n5588 ^ 1'b0 ;
  assign n18512 = ( n4279 & ~n18509 ) | ( n4279 & n18511 ) | ( ~n18509 & n18511 ) ;
  assign n18513 = n5196 ^ n2456 ^ 1'b0 ;
  assign n18514 = n8023 & n18513 ;
  assign n18515 = n3120 & n9338 ;
  assign n18516 = n13194 & n18515 ;
  assign n18518 = ( n2127 & ~n7775 ) | ( n2127 & n10488 ) | ( ~n7775 & n10488 ) ;
  assign n18519 = ( ~n9047 & n12375 ) | ( ~n9047 & n18518 ) | ( n12375 & n18518 ) ;
  assign n18517 = n1880 & ~n3985 ;
  assign n18520 = n18519 ^ n18517 ^ n2619 ;
  assign n18521 = n10431 ^ n8158 ^ n6413 ;
  assign n18522 = n18521 ^ n5830 ^ 1'b0 ;
  assign n18523 = n16447 & ~n18522 ;
  assign n18530 = n3073 | n3146 ;
  assign n18531 = n15392 ^ n12337 ^ n9772 ;
  assign n18532 = ( n1020 & n18530 ) | ( n1020 & n18531 ) | ( n18530 & n18531 ) ;
  assign n18533 = n18532 ^ n14720 ^ n7400 ;
  assign n18524 = n1031 & ~n2198 ;
  assign n18525 = n487 & n18524 ;
  assign n18526 = n919 ^ n279 ^ 1'b0 ;
  assign n18527 = n5192 | n18526 ;
  assign n18528 = n15065 & ~n18527 ;
  assign n18529 = ( n13055 & n18525 ) | ( n13055 & n18528 ) | ( n18525 & n18528 ) ;
  assign n18534 = n18533 ^ n18529 ^ n8769 ;
  assign n18535 = n16432 ^ n16277 ^ 1'b0 ;
  assign n18536 = x28 & n18535 ;
  assign n18537 = n12575 | n16990 ;
  assign n18539 = n13945 ^ n7741 ^ n4585 ;
  assign n18540 = n18539 ^ n9593 ^ n5075 ;
  assign n18538 = ( ~n5019 & n5680 ) | ( ~n5019 & n11724 ) | ( n5680 & n11724 ) ;
  assign n18541 = n18540 ^ n18538 ^ n10279 ;
  assign n18542 = ( n11409 & n16250 ) | ( n11409 & n18541 ) | ( n16250 & n18541 ) ;
  assign n18543 = ~n3022 & n3361 ;
  assign n18544 = ~n470 & n18543 ;
  assign n18545 = n11943 & ~n18544 ;
  assign n18546 = n8163 & n18545 ;
  assign n18547 = n9432 ^ n8393 ^ n1352 ;
  assign n18548 = n7920 & ~n18547 ;
  assign n18549 = n11889 ^ n9214 ^ n1167 ;
  assign n18551 = n12262 ^ n10894 ^ n956 ;
  assign n18550 = n3271 & n6940 ;
  assign n18552 = n18551 ^ n18550 ^ 1'b0 ;
  assign n18553 = ( ~n4057 & n18549 ) | ( ~n4057 & n18552 ) | ( n18549 & n18552 ) ;
  assign n18554 = ( n5024 & n14998 ) | ( n5024 & n15694 ) | ( n14998 & n15694 ) ;
  assign n18555 = ( n7173 & n13770 ) | ( n7173 & n18554 ) | ( n13770 & n18554 ) ;
  assign n18556 = n1152 | n10422 ;
  assign n18557 = n14785 | n18556 ;
  assign n18558 = ( n1407 & n6585 ) | ( n1407 & ~n10771 ) | ( n6585 & ~n10771 ) ;
  assign n18559 = n5262 | n16513 ;
  assign n18560 = n18558 | n18559 ;
  assign n18561 = n2838 | n11766 ;
  assign n18562 = n10124 & ~n18561 ;
  assign n18563 = ( ~n9205 & n11393 ) | ( ~n9205 & n18562 ) | ( n11393 & n18562 ) ;
  assign n18564 = n5502 | n12601 ;
  assign n18565 = n14205 ^ n9830 ^ x6 ;
  assign n18566 = n7536 & ~n18565 ;
  assign n18567 = n18566 ^ n6407 ^ 1'b0 ;
  assign n18569 = n4992 & ~n16001 ;
  assign n18568 = n15817 ^ n13536 ^ n1436 ;
  assign n18570 = n18569 ^ n18568 ^ n3583 ;
  assign n18571 = n5017 | n18570 ;
  assign n18582 = n634 & ~n6370 ;
  assign n18583 = n18582 ^ n2437 ^ 1'b0 ;
  assign n18581 = ( n4433 & ~n5355 ) | ( n4433 & n13028 ) | ( ~n5355 & n13028 ) ;
  assign n18572 = n4880 & ~n18421 ;
  assign n18573 = n18572 ^ n723 ^ 1'b0 ;
  assign n18574 = ( ~n3858 & n4574 ) | ( ~n3858 & n8085 ) | ( n4574 & n8085 ) ;
  assign n18575 = n18574 ^ n12560 ^ n11330 ;
  assign n18576 = ( x142 & n18573 ) | ( x142 & ~n18575 ) | ( n18573 & ~n18575 ) ;
  assign n18577 = ( n4805 & n13055 ) | ( n4805 & ~n18576 ) | ( n13055 & ~n18576 ) ;
  assign n18578 = n18577 ^ n7689 ^ 1'b0 ;
  assign n18579 = ~n7685 & n18578 ;
  assign n18580 = n18579 ^ n8868 ^ 1'b0 ;
  assign n18584 = n18583 ^ n18581 ^ n18580 ;
  assign n18585 = n9117 | n11468 ;
  assign n18586 = n18585 ^ n5456 ^ 1'b0 ;
  assign n18587 = n4109 | n18586 ;
  assign n18588 = n10711 ^ x237 ^ 1'b0 ;
  assign n18589 = n2894 | n18588 ;
  assign n18590 = n2091 & ~n18589 ;
  assign n18591 = n1029 & n5732 ;
  assign n18592 = ( n2408 & n15962 ) | ( n2408 & ~n18591 ) | ( n15962 & ~n18591 ) ;
  assign n18593 = n18592 ^ n16268 ^ n15129 ;
  assign n18594 = n5204 & ~n6392 ;
  assign n18595 = n1074 & n18594 ;
  assign n18596 = n18595 ^ n6361 ^ 1'b0 ;
  assign n18597 = n6855 & ~n18596 ;
  assign n18598 = ( n828 & n1602 ) | ( n828 & ~n7523 ) | ( n1602 & ~n7523 ) ;
  assign n18599 = x121 & n18598 ;
  assign n18600 = n8635 & n18599 ;
  assign n18601 = ( n4397 & ~n5508 ) | ( n4397 & n8979 ) | ( ~n5508 & n8979 ) ;
  assign n18602 = ( n5348 & n9093 ) | ( n5348 & ~n18601 ) | ( n9093 & ~n18601 ) ;
  assign n18603 = x58 & ~n2516 ;
  assign n18604 = n18602 & n18603 ;
  assign n18605 = n8798 & ~n15383 ;
  assign n18606 = n18604 & n18605 ;
  assign n18607 = n3049 & ~n16240 ;
  assign n18608 = ~n8754 & n18607 ;
  assign n18609 = n18240 ^ n16429 ^ 1'b0 ;
  assign n18610 = n18608 | n18609 ;
  assign n18611 = n3801 & n5496 ;
  assign n18612 = n8861 ^ n2455 ^ x19 ;
  assign n18618 = ( n387 & ~n5515 ) | ( n387 & n10040 ) | ( ~n5515 & n10040 ) ;
  assign n18619 = ( n4933 & n7222 ) | ( n4933 & ~n18618 ) | ( n7222 & ~n18618 ) ;
  assign n18615 = ( n10296 & ~n10825 ) | ( n10296 & n15897 ) | ( ~n10825 & n15897 ) ;
  assign n18616 = n18615 ^ n17454 ^ 1'b0 ;
  assign n18617 = n3681 & ~n18616 ;
  assign n18613 = ( ~n1520 & n1578 ) | ( ~n1520 & n8610 ) | ( n1578 & n8610 ) ;
  assign n18614 = n10180 & ~n18613 ;
  assign n18620 = n18619 ^ n18617 ^ n18614 ;
  assign n18621 = ~n13603 & n18620 ;
  assign n18622 = ~n4676 & n18621 ;
  assign n18623 = ( n4066 & n9185 ) | ( n4066 & ~n11178 ) | ( n9185 & ~n11178 ) ;
  assign n18624 = ~n1789 & n2226 ;
  assign n18625 = n18624 ^ n11797 ^ 1'b0 ;
  assign n18626 = n18625 ^ n18449 ^ n15558 ;
  assign n18627 = n18626 ^ n9008 ^ 1'b0 ;
  assign n18628 = ( n10296 & n10874 ) | ( n10296 & n14460 ) | ( n10874 & n14460 ) ;
  assign n18629 = n10084 & ~n10922 ;
  assign n18630 = n11831 & ~n18629 ;
  assign n18631 = n16005 ^ n15056 ^ n2566 ;
  assign n18632 = ( ~n3330 & n18630 ) | ( ~n3330 & n18631 ) | ( n18630 & n18631 ) ;
  assign n18642 = ( n2456 & n6768 ) | ( n2456 & ~n15291 ) | ( n6768 & ~n15291 ) ;
  assign n18643 = ( n5195 & n6906 ) | ( n5195 & n10213 ) | ( n6906 & n10213 ) ;
  assign n18644 = n18643 ^ n9911 ^ n2544 ;
  assign n18645 = ( n1846 & n4645 ) | ( n1846 & ~n18644 ) | ( n4645 & ~n18644 ) ;
  assign n18646 = ~n18642 & n18645 ;
  assign n18639 = n3260 & ~n12366 ;
  assign n18640 = ~x199 & n18639 ;
  assign n18637 = x180 | n1720 ;
  assign n18633 = n6222 & ~n10091 ;
  assign n18634 = ( n3694 & n4026 ) | ( n3694 & ~n18633 ) | ( n4026 & ~n18633 ) ;
  assign n18635 = ~n12298 & n18634 ;
  assign n18636 = n18635 ^ n18036 ^ 1'b0 ;
  assign n18638 = n18637 ^ n18636 ^ n12298 ;
  assign n18641 = n18640 ^ n18638 ^ n11355 ;
  assign n18647 = n18646 ^ n18641 ^ n1384 ;
  assign n18648 = n15809 ^ n4261 ^ n2663 ;
  assign n18660 = n3900 ^ n3766 ^ n2497 ;
  assign n18663 = ( n2070 & n2379 ) | ( n2070 & ~n10701 ) | ( n2379 & ~n10701 ) ;
  assign n18661 = ( n6400 & n9573 ) | ( n6400 & n17840 ) | ( n9573 & n17840 ) ;
  assign n18662 = n8133 & ~n18661 ;
  assign n18664 = n18663 ^ n18662 ^ 1'b0 ;
  assign n18665 = ( n2932 & ~n18660 ) | ( n2932 & n18664 ) | ( ~n18660 & n18664 ) ;
  assign n18657 = n308 | n3103 ;
  assign n18658 = n18657 ^ n1532 ^ 1'b0 ;
  assign n18649 = n9477 ^ n5786 ^ 1'b0 ;
  assign n18650 = ~n827 & n14246 ;
  assign n18651 = n3303 & n18650 ;
  assign n18652 = n18649 | n18651 ;
  assign n18653 = n18652 ^ n13110 ^ 1'b0 ;
  assign n18654 = n2509 | n18653 ;
  assign n18655 = n11726 & n18654 ;
  assign n18656 = n4563 & n18655 ;
  assign n18659 = n18658 ^ n18656 ^ n4068 ;
  assign n18666 = n18665 ^ n18659 ^ n3978 ;
  assign n18667 = ( x35 & n2144 ) | ( x35 & ~n17918 ) | ( n2144 & ~n17918 ) ;
  assign n18668 = n18666 & n18667 ;
  assign n18669 = n18648 & n18668 ;
  assign n18670 = n4322 ^ n3333 ^ 1'b0 ;
  assign n18671 = ( n2592 & ~n3578 ) | ( n2592 & n18670 ) | ( ~n3578 & n18670 ) ;
  assign n18672 = n8954 & ~n13917 ;
  assign n18673 = n18672 ^ n10927 ^ 1'b0 ;
  assign n18674 = n18673 ^ n3372 ^ 1'b0 ;
  assign n18675 = ( n15571 & n18671 ) | ( n15571 & ~n18674 ) | ( n18671 & ~n18674 ) ;
  assign n18676 = ~n6615 & n13652 ;
  assign n18677 = n18676 ^ n14722 ^ n4834 ;
  assign n18678 = n2046 ^ n891 ^ 1'b0 ;
  assign n18679 = n5177 | n18678 ;
  assign n18680 = n18679 ^ n6028 ^ 1'b0 ;
  assign n18681 = ( n14857 & n15727 ) | ( n14857 & n18680 ) | ( n15727 & n18680 ) ;
  assign n18682 = n1297 & ~n18681 ;
  assign n18683 = n18682 ^ n4715 ^ 1'b0 ;
  assign n18684 = ( n6328 & n6693 ) | ( n6328 & n12637 ) | ( n6693 & n12637 ) ;
  assign n18685 = n18684 ^ n1981 ^ 1'b0 ;
  assign n18686 = n18685 ^ n15535 ^ 1'b0 ;
  assign n18687 = ( n2283 & ~n3849 ) | ( n2283 & n10457 ) | ( ~n3849 & n10457 ) ;
  assign n18688 = n6292 | n6381 ;
  assign n18689 = ( n5747 & n8487 ) | ( n5747 & ~n18688 ) | ( n8487 & ~n18688 ) ;
  assign n18690 = n18689 ^ n5880 ^ 1'b0 ;
  assign n18691 = n330 & ~n18690 ;
  assign n18692 = ( ~n8889 & n18687 ) | ( ~n8889 & n18691 ) | ( n18687 & n18691 ) ;
  assign n18693 = n7283 ^ n2332 ^ n1627 ;
  assign n18694 = ( ~n1645 & n5290 ) | ( ~n1645 & n6780 ) | ( n5290 & n6780 ) ;
  assign n18695 = n18694 ^ n12725 ^ 1'b0 ;
  assign n18696 = ( ~n1195 & n2663 ) | ( ~n1195 & n7348 ) | ( n2663 & n7348 ) ;
  assign n18698 = n6644 ^ n2706 ^ 1'b0 ;
  assign n18699 = n1740 | n18698 ;
  assign n18697 = n13079 ^ n549 ^ 1'b0 ;
  assign n18700 = n18699 ^ n18697 ^ 1'b0 ;
  assign n18701 = n13456 ^ n13443 ^ n2969 ;
  assign n18702 = ( n7786 & n17056 ) | ( n7786 & n18701 ) | ( n17056 & n18701 ) ;
  assign n18703 = n5700 | n12286 ;
  assign n18704 = n6363 ^ n1928 ^ n1327 ;
  assign n18705 = n11603 & ~n18704 ;
  assign n18706 = n5249 & n11400 ;
  assign n18707 = ~n5204 & n18706 ;
  assign n18708 = n8148 | n18707 ;
  assign n18709 = ( ~n296 & n4144 ) | ( ~n296 & n12574 ) | ( n4144 & n12574 ) ;
  assign n18710 = ( n5129 & n11724 ) | ( n5129 & n18709 ) | ( n11724 & n18709 ) ;
  assign n18711 = ( n4389 & ~n18708 ) | ( n4389 & n18710 ) | ( ~n18708 & n18710 ) ;
  assign n18712 = n7495 ^ n6857 ^ 1'b0 ;
  assign n18713 = ~n17267 & n18712 ;
  assign n18714 = ( n7512 & n8419 ) | ( n7512 & ~n9597 ) | ( n8419 & ~n9597 ) ;
  assign n18715 = ( n3653 & n10682 ) | ( n3653 & ~n18714 ) | ( n10682 & ~n18714 ) ;
  assign n18716 = n13839 ^ n9546 ^ n7113 ;
  assign n18717 = ~n1116 & n2802 ;
  assign n18718 = ~n7395 & n18717 ;
  assign n18719 = n18718 ^ n15284 ^ n4362 ;
  assign n18720 = ( n7696 & ~n9485 ) | ( n7696 & n13706 ) | ( ~n9485 & n13706 ) ;
  assign n18721 = ( ~n7947 & n11497 ) | ( ~n7947 & n18720 ) | ( n11497 & n18720 ) ;
  assign n18722 = ~n290 & n14500 ;
  assign n18723 = n18722 ^ n17601 ^ 1'b0 ;
  assign n18724 = n9431 | n18723 ;
  assign n18725 = n14766 ^ n12857 ^ n6409 ;
  assign n18726 = ~n11481 & n18725 ;
  assign n18727 = n18726 ^ n14434 ^ 1'b0 ;
  assign n18728 = n18724 | n18727 ;
  assign n18730 = n17300 ^ n1421 ^ 1'b0 ;
  assign n18729 = ( n5566 & n5921 ) | ( n5566 & ~n7728 ) | ( n5921 & ~n7728 ) ;
  assign n18731 = n18730 ^ n18729 ^ n13260 ;
  assign n18732 = n16047 ^ n12688 ^ n9822 ;
  assign n18737 = n9744 & ~n18626 ;
  assign n18738 = n18737 ^ n2395 ^ 1'b0 ;
  assign n18735 = ( ~n798 & n1956 ) | ( ~n798 & n7542 ) | ( n1956 & n7542 ) ;
  assign n18733 = n11155 ^ n7970 ^ n5943 ;
  assign n18734 = n4675 | n18733 ;
  assign n18736 = n18735 ^ n18734 ^ 1'b0 ;
  assign n18739 = n18738 ^ n18736 ^ 1'b0 ;
  assign n18740 = ( n6907 & n7024 ) | ( n6907 & ~n18739 ) | ( n7024 & ~n18739 ) ;
  assign n18741 = ( n16424 & ~n18732 ) | ( n16424 & n18740 ) | ( ~n18732 & n18740 ) ;
  assign n18742 = n5162 ^ x74 ^ 1'b0 ;
  assign n18743 = n18180 ^ n7544 ^ n7056 ;
  assign n18744 = n6363 ^ n5680 ^ 1'b0 ;
  assign n18747 = n2676 & n2928 ;
  assign n18745 = n8264 & n15903 ;
  assign n18746 = n18745 ^ n14628 ^ 1'b0 ;
  assign n18748 = n18747 ^ n18746 ^ n7349 ;
  assign n18749 = ( n735 & n1659 ) | ( n735 & n5849 ) | ( n1659 & n5849 ) ;
  assign n18750 = n351 & n18749 ;
  assign n18751 = n18750 ^ n2797 ^ 1'b0 ;
  assign n18752 = ( n501 & n6869 ) | ( n501 & n10808 ) | ( n6869 & n10808 ) ;
  assign n18753 = n18752 ^ n11675 ^ 1'b0 ;
  assign n18754 = n18751 & ~n18753 ;
  assign n18755 = n18754 ^ n13374 ^ 1'b0 ;
  assign n18756 = n18755 ^ n12630 ^ n7670 ;
  assign n18757 = n3486 ^ n3369 ^ 1'b0 ;
  assign n18758 = n18757 ^ n7365 ^ n422 ;
  assign n18765 = ( n1274 & n3601 ) | ( n1274 & n4294 ) | ( n3601 & n4294 ) ;
  assign n18762 = ( ~n5731 & n7591 ) | ( ~n5731 & n17982 ) | ( n7591 & n17982 ) ;
  assign n18759 = n11810 ^ n4609 ^ 1'b0 ;
  assign n18760 = n1507 | n18759 ;
  assign n18761 = n12069 & ~n18760 ;
  assign n18763 = n18762 ^ n18761 ^ 1'b0 ;
  assign n18764 = n8626 & ~n18763 ;
  assign n18766 = n18765 ^ n18764 ^ n5136 ;
  assign n18767 = ( n2241 & ~n4812 ) | ( n2241 & n12062 ) | ( ~n4812 & n12062 ) ;
  assign n18768 = ( n5419 & n8569 ) | ( n5419 & n18767 ) | ( n8569 & n18767 ) ;
  assign n18769 = ( n3962 & n15900 ) | ( n3962 & ~n18768 ) | ( n15900 & ~n18768 ) ;
  assign n18770 = n11522 | n18769 ;
  assign n18771 = n18766 & ~n18770 ;
  assign n18772 = ( ~x246 & n1466 ) | ( ~x246 & n5270 ) | ( n1466 & n5270 ) ;
  assign n18773 = ( n8315 & n14603 ) | ( n8315 & ~n18772 ) | ( n14603 & ~n18772 ) ;
  assign n18774 = n17793 | n18773 ;
  assign n18775 = n3227 | n5552 ;
  assign n18776 = ( ~n7525 & n16523 ) | ( ~n7525 & n18775 ) | ( n16523 & n18775 ) ;
  assign n18777 = ~n4460 & n8777 ;
  assign n18778 = ~n6493 & n18777 ;
  assign n18779 = ( n1467 & n17974 ) | ( n1467 & ~n18778 ) | ( n17974 & ~n18778 ) ;
  assign n18780 = n8378 & ~n18313 ;
  assign n18781 = ~n18779 & n18780 ;
  assign n18786 = n6331 ^ n4757 ^ n2719 ;
  assign n18784 = n12742 ^ n7928 ^ 1'b0 ;
  assign n18782 = n8924 | n15444 ;
  assign n18783 = n18782 ^ n5389 ^ 1'b0 ;
  assign n18785 = n18784 ^ n18783 ^ n5395 ;
  assign n18787 = n18786 ^ n18785 ^ n4717 ;
  assign n18788 = n17783 ^ n11103 ^ 1'b0 ;
  assign n18789 = ~n2826 & n18788 ;
  assign n18790 = n16586 ^ n7491 ^ n5878 ;
  assign n18791 = n18790 ^ n4729 ^ n3870 ;
  assign n18792 = ( ~n330 & n15371 ) | ( ~n330 & n18791 ) | ( n15371 & n18791 ) ;
  assign n18793 = ( n17147 & ~n18789 ) | ( n17147 & n18792 ) | ( ~n18789 & n18792 ) ;
  assign n18794 = ( n1144 & n1513 ) | ( n1144 & ~n12842 ) | ( n1513 & ~n12842 ) ;
  assign n18795 = n18794 ^ n12542 ^ 1'b0 ;
  assign n18796 = ( n2785 & n3042 ) | ( n2785 & n7259 ) | ( n3042 & n7259 ) ;
  assign n18797 = n3735 & n4399 ;
  assign n18798 = n18797 ^ n7736 ^ 1'b0 ;
  assign n18799 = n18798 ^ n8615 ^ n4447 ;
  assign n18800 = ( n3971 & n6790 ) | ( n3971 & n18131 ) | ( n6790 & n18131 ) ;
  assign n18801 = n8711 ^ n6687 ^ n2764 ;
  assign n18802 = ( n1240 & ~n6798 ) | ( n1240 & n18801 ) | ( ~n6798 & n18801 ) ;
  assign n18803 = n18802 ^ n4709 ^ n834 ;
  assign n18804 = n2430 & n5027 ;
  assign n18805 = n18804 ^ n2633 ^ 1'b0 ;
  assign n18806 = n18805 ^ n10397 ^ n8078 ;
  assign n18807 = n933 & ~n17441 ;
  assign n18808 = ~n11759 & n18807 ;
  assign n18810 = n4454 | n14014 ;
  assign n18811 = n4944 & ~n5138 ;
  assign n18812 = n18575 & n18811 ;
  assign n18813 = n18812 ^ n14871 ^ n5554 ;
  assign n18814 = n18810 & n18813 ;
  assign n18809 = ~n12776 & n15857 ;
  assign n18815 = n18814 ^ n18809 ^ 1'b0 ;
  assign n18816 = ( ~x121 & n2549 ) | ( ~x121 & n18239 ) | ( n2549 & n18239 ) ;
  assign n18817 = n1845 | n15334 ;
  assign n18818 = n13942 ^ n2792 ^ n991 ;
  assign n18819 = ( n1329 & n1791 ) | ( n1329 & ~n5396 ) | ( n1791 & ~n5396 ) ;
  assign n18820 = n3538 | n10306 ;
  assign n18821 = ( ~n5751 & n16694 ) | ( ~n5751 & n18820 ) | ( n16694 & n18820 ) ;
  assign n18822 = n6144 ^ n3131 ^ 1'b0 ;
  assign n18823 = ( n18819 & ~n18821 ) | ( n18819 & n18822 ) | ( ~n18821 & n18822 ) ;
  assign n18824 = n18823 ^ n13009 ^ n3912 ;
  assign n18825 = n10356 ^ n10176 ^ n2666 ;
  assign n18826 = n15459 & n18825 ;
  assign n18827 = n18826 ^ n6668 ^ 1'b0 ;
  assign n18828 = ( n777 & n8714 ) | ( n777 & ~n13981 ) | ( n8714 & ~n13981 ) ;
  assign n18829 = n18828 ^ n2704 ^ 1'b0 ;
  assign n18830 = n7461 ^ n572 ^ 1'b0 ;
  assign n18831 = n18830 ^ n2366 ^ 1'b0 ;
  assign n18832 = n6732 | n18831 ;
  assign n18833 = ( n16945 & ~n17299 ) | ( n16945 & n18832 ) | ( ~n17299 & n18832 ) ;
  assign n18834 = n1392 ^ n837 ^ 1'b0 ;
  assign n18835 = ( n6110 & n8974 ) | ( n6110 & ~n18834 ) | ( n8974 & ~n18834 ) ;
  assign n18836 = n18835 ^ n12221 ^ 1'b0 ;
  assign n18838 = ~n4181 & n10990 ;
  assign n18837 = n6482 ^ n6018 ^ n1685 ;
  assign n18839 = n18838 ^ n18837 ^ 1'b0 ;
  assign n18840 = n17800 | n18839 ;
  assign n18841 = n5540 & ~n7022 ;
  assign n18842 = n18841 ^ n2173 ^ 1'b0 ;
  assign n18843 = ( ~n18836 & n18840 ) | ( ~n18836 & n18842 ) | ( n18840 & n18842 ) ;
  assign n18844 = n6339 ^ n4664 ^ 1'b0 ;
  assign n18845 = n11765 & n18844 ;
  assign n18846 = n4807 ^ n4555 ^ 1'b0 ;
  assign n18847 = ~n3185 & n18846 ;
  assign n18848 = n6855 ^ n3402 ^ 1'b0 ;
  assign n18849 = ( n4283 & n18847 ) | ( n4283 & ~n18848 ) | ( n18847 & ~n18848 ) ;
  assign n18850 = n10958 ^ n7354 ^ n5060 ;
  assign n18851 = n8254 ^ n4201 ^ 1'b0 ;
  assign n18852 = ~n18850 & n18851 ;
  assign n18853 = n15435 ^ n5111 ^ 1'b0 ;
  assign n18854 = ( n4305 & n6164 ) | ( n4305 & n7586 ) | ( n6164 & n7586 ) ;
  assign n18855 = n18854 ^ n13500 ^ n6103 ;
  assign n18860 = ( n393 & ~n10641 ) | ( n393 & n11590 ) | ( ~n10641 & n11590 ) ;
  assign n18857 = ~n4534 & n17582 ;
  assign n18858 = n8205 & n18857 ;
  assign n18859 = ~n447 & n18858 ;
  assign n18861 = n18860 ^ n18859 ^ n11647 ;
  assign n18856 = ( n471 & n3826 ) | ( n471 & n7562 ) | ( n3826 & n7562 ) ;
  assign n18862 = n18861 ^ n18856 ^ n7739 ;
  assign n18863 = ( x4 & ~n4472 ) | ( x4 & n5724 ) | ( ~n4472 & n5724 ) ;
  assign n18864 = n18863 ^ n11093 ^ n282 ;
  assign n18870 = n962 | n2867 ;
  assign n18869 = n13500 ^ n6968 ^ n1146 ;
  assign n18865 = n5777 ^ n2650 ^ 1'b0 ;
  assign n18866 = n18865 ^ n8289 ^ n7730 ;
  assign n18867 = n436 & ~n11025 ;
  assign n18868 = n18866 & n18867 ;
  assign n18871 = n18870 ^ n18869 ^ n18868 ;
  assign n18875 = n17564 ^ n3103 ^ 1'b0 ;
  assign n18872 = ( n3042 & n8784 ) | ( n3042 & ~n11854 ) | ( n8784 & ~n11854 ) ;
  assign n18873 = n13476 & ~n18872 ;
  assign n18874 = n3038 & n18873 ;
  assign n18876 = n18875 ^ n18874 ^ 1'b0 ;
  assign n18877 = n1131 | n15797 ;
  assign n18878 = n18360 & ~n18877 ;
  assign n18879 = ~n7080 & n7663 ;
  assign n18881 = n1701 & ~n5152 ;
  assign n18882 = ~x209 & n18881 ;
  assign n18883 = n18882 ^ n6403 ^ n4525 ;
  assign n18884 = n4139 & ~n18883 ;
  assign n18880 = n15428 ^ n10282 ^ n7120 ;
  assign n18885 = n18884 ^ n18880 ^ n11617 ;
  assign n18886 = n8318 ^ n7294 ^ 1'b0 ;
  assign n18887 = n18886 ^ n14945 ^ n575 ;
  assign n18888 = n3408 ^ n3367 ^ 1'b0 ;
  assign n18889 = n8167 & ~n18888 ;
  assign n18890 = n18889 ^ n13547 ^ n3525 ;
  assign n18891 = n8187 & ~n11766 ;
  assign n18892 = n18890 & n18891 ;
  assign n18893 = n17673 ^ n9927 ^ n2143 ;
  assign n18894 = ~n3571 & n11871 ;
  assign n18895 = ~n3868 & n18894 ;
  assign n18896 = ~n6523 & n9656 ;
  assign n18897 = n500 & n18896 ;
  assign n18898 = n2767 & n18897 ;
  assign n18899 = n18898 ^ n15099 ^ n2240 ;
  assign n18900 = ( n2014 & n18895 ) | ( n2014 & n18899 ) | ( n18895 & n18899 ) ;
  assign n18902 = ( ~n2325 & n4992 ) | ( ~n2325 & n8232 ) | ( n4992 & n8232 ) ;
  assign n18901 = ( n7225 & n8050 ) | ( n7225 & n18658 ) | ( n8050 & n18658 ) ;
  assign n18903 = n18902 ^ n18901 ^ n1365 ;
  assign n18904 = n14448 ^ n9822 ^ n4746 ;
  assign n18905 = n18904 ^ n12827 ^ 1'b0 ;
  assign n18906 = ( n1046 & n4828 ) | ( n1046 & n6016 ) | ( n4828 & n6016 ) ;
  assign n18907 = ( ~n8279 & n18905 ) | ( ~n8279 & n18906 ) | ( n18905 & n18906 ) ;
  assign n18908 = n8664 ^ n8277 ^ 1'b0 ;
  assign n18909 = n11428 | n18908 ;
  assign n18910 = n17189 ^ n16964 ^ n8591 ;
  assign n18911 = n18910 ^ n5256 ^ n2280 ;
  assign n18912 = ~n18909 & n18911 ;
  assign n18913 = n6490 & n18912 ;
  assign n18914 = n17368 ^ n4342 ^ 1'b0 ;
  assign n18915 = ( n5948 & ~n10196 ) | ( n5948 & n12559 ) | ( ~n10196 & n12559 ) ;
  assign n18916 = n5925 ^ n5442 ^ 1'b0 ;
  assign n18917 = ( ~n3906 & n7041 ) | ( ~n3906 & n8044 ) | ( n7041 & n8044 ) ;
  assign n18918 = ( ~n5446 & n12307 ) | ( ~n5446 & n18917 ) | ( n12307 & n18917 ) ;
  assign n18919 = n9857 ^ n2433 ^ n516 ;
  assign n18920 = ( n1594 & ~n4094 ) | ( n1594 & n18919 ) | ( ~n4094 & n18919 ) ;
  assign n18921 = ( x225 & ~n2466 ) | ( x225 & n18920 ) | ( ~n2466 & n18920 ) ;
  assign n18922 = ( ~n5911 & n13072 ) | ( ~n5911 & n18921 ) | ( n13072 & n18921 ) ;
  assign n18923 = n18922 ^ n1649 ^ 1'b0 ;
  assign n18924 = n14151 ^ n6141 ^ n1246 ;
  assign n18925 = n18296 & ~n18924 ;
  assign n18926 = n15438 ^ n15150 ^ 1'b0 ;
  assign n18927 = n8138 & ~n18926 ;
  assign n18928 = n10184 & ~n13462 ;
  assign n18929 = n3190 & n12831 ;
  assign n18930 = n5152 & n18929 ;
  assign n18931 = n18930 ^ n9086 ^ 1'b0 ;
  assign n18932 = n8062 & ~n18931 ;
  assign n18933 = n5901 & ~n18932 ;
  assign n18934 = n320 & n11533 ;
  assign n18935 = n18934 ^ n3294 ^ 1'b0 ;
  assign n18936 = n6963 | n7632 ;
  assign n18937 = n18935 | n18936 ;
  assign n18938 = n3292 ^ n2055 ^ 1'b0 ;
  assign n18939 = n14105 | n18938 ;
  assign n18940 = n12043 | n18939 ;
  assign n18941 = ( n13045 & n18937 ) | ( n13045 & n18940 ) | ( n18937 & n18940 ) ;
  assign n18942 = n4736 & n9020 ;
  assign n18943 = ~n18941 & n18942 ;
  assign n18944 = n2434 & n6073 ;
  assign n18945 = n18944 ^ n11343 ^ n8158 ;
  assign n18946 = n9579 ^ n5048 ^ n2528 ;
  assign n18947 = n18946 ^ n2178 ^ n1344 ;
  assign n18948 = ~n4550 & n11397 ;
  assign n18949 = ~x196 & n18948 ;
  assign n18950 = n18947 & ~n18949 ;
  assign n18951 = ~n18947 & n18950 ;
  assign n18952 = n9656 ^ n7784 ^ n7769 ;
  assign n18953 = ~n3505 & n12398 ;
  assign n18954 = ~n702 & n18953 ;
  assign n18955 = n2870 | n18954 ;
  assign n18956 = n7920 | n18955 ;
  assign n18957 = n2735 | n5424 ;
  assign n18958 = n18957 ^ n825 ^ 1'b0 ;
  assign n18959 = n17333 & n18958 ;
  assign n18960 = n18959 ^ n458 ^ 1'b0 ;
  assign n18961 = n4159 & ~n18960 ;
  assign n18962 = n18961 ^ n16313 ^ 1'b0 ;
  assign n18963 = ( n18952 & n18956 ) | ( n18952 & ~n18962 ) | ( n18956 & ~n18962 ) ;
  assign n18964 = n18951 & n18963 ;
  assign n18967 = ( n7297 & ~n9107 ) | ( n7297 & n13603 ) | ( ~n9107 & n13603 ) ;
  assign n18968 = n18967 ^ n15950 ^ 1'b0 ;
  assign n18969 = n2525 & n18968 ;
  assign n18965 = n17591 ^ n1159 ^ 1'b0 ;
  assign n18966 = ~n12498 & n18965 ;
  assign n18970 = n18969 ^ n18966 ^ 1'b0 ;
  assign n18977 = n4017 & ~n4689 ;
  assign n18978 = n18977 ^ n8295 ^ 1'b0 ;
  assign n18975 = n13270 ^ n8156 ^ n3571 ;
  assign n18971 = ( n784 & n916 ) | ( n784 & ~n3515 ) | ( n916 & ~n3515 ) ;
  assign n18972 = ( n1457 & n13460 ) | ( n1457 & ~n18971 ) | ( n13460 & ~n18971 ) ;
  assign n18973 = n18972 ^ n9405 ^ n8717 ;
  assign n18974 = n18973 ^ n18544 ^ n3254 ;
  assign n18976 = n18975 ^ n18974 ^ n11984 ;
  assign n18979 = n18978 ^ n18976 ^ n18587 ;
  assign n18980 = n10461 ^ n524 ^ 1'b0 ;
  assign n18981 = n1646 | n3973 ;
  assign n18982 = n1546 & ~n18981 ;
  assign n18983 = n18982 ^ n13958 ^ n1455 ;
  assign n18984 = n18983 ^ n8238 ^ n542 ;
  assign n18985 = n765 & n6936 ;
  assign n18986 = n1026 & n18985 ;
  assign n18987 = n18986 ^ n1446 ^ 1'b0 ;
  assign n18988 = n14376 & n18987 ;
  assign n18989 = n12002 ^ n4422 ^ 1'b0 ;
  assign n18990 = n12191 | n18989 ;
  assign n18991 = n360 & ~n11016 ;
  assign n18992 = n9619 | n18991 ;
  assign n18993 = n9157 ^ n5953 ^ 1'b0 ;
  assign n18994 = ~n6834 & n18993 ;
  assign n18995 = n2428 | n4575 ;
  assign n18996 = n18994 | n18995 ;
  assign n18997 = n18996 ^ n7363 ^ n2588 ;
  assign n18998 = ~n18992 & n18997 ;
  assign n18999 = n18990 & n18998 ;
  assign n19000 = n11730 ^ n1996 ^ n1267 ;
  assign n19001 = n7749 | n14966 ;
  assign n19002 = n16511 ^ n12596 ^ n5227 ;
  assign n19003 = ( ~n1763 & n16608 ) | ( ~n1763 & n19002 ) | ( n16608 & n19002 ) ;
  assign n19004 = ( n2889 & n6733 ) | ( n2889 & n7070 ) | ( n6733 & n7070 ) ;
  assign n19005 = ( n3368 & ~n7143 ) | ( n3368 & n19004 ) | ( ~n7143 & n19004 ) ;
  assign n19006 = n19005 ^ n7884 ^ n2492 ;
  assign n19007 = n15332 ^ n5842 ^ n5536 ;
  assign n19008 = ~n9097 & n9993 ;
  assign n19009 = ~n16042 & n19008 ;
  assign n19010 = n9677 & n17513 ;
  assign n19011 = n10163 & n19010 ;
  assign n19012 = n19011 ^ n4883 ^ n3191 ;
  assign n19013 = ( ~n665 & n4477 ) | ( ~n665 & n8274 ) | ( n4477 & n8274 ) ;
  assign n19014 = n18767 ^ n11376 ^ n1325 ;
  assign n19015 = n19014 ^ n10865 ^ 1'b0 ;
  assign n19016 = n834 & ~n19015 ;
  assign n19017 = ~n19013 & n19016 ;
  assign n19018 = n19017 ^ n15517 ^ 1'b0 ;
  assign n19019 = ( x231 & n4640 ) | ( x231 & ~n6330 ) | ( n4640 & ~n6330 ) ;
  assign n19020 = ( n3735 & n14080 ) | ( n3735 & n19019 ) | ( n14080 & n19019 ) ;
  assign n19021 = ( n8668 & ~n10660 ) | ( n8668 & n19020 ) | ( ~n10660 & n19020 ) ;
  assign n19022 = ( ~n1316 & n9285 ) | ( ~n1316 & n14815 ) | ( n9285 & n14815 ) ;
  assign n19023 = ( n548 & ~n6614 ) | ( n548 & n18190 ) | ( ~n6614 & n18190 ) ;
  assign n19024 = n19023 ^ n10151 ^ 1'b0 ;
  assign n19025 = n6060 | n19024 ;
  assign n19026 = n12444 ^ n12326 ^ 1'b0 ;
  assign n19027 = n7393 ^ n5520 ^ n2097 ;
  assign n19028 = n19027 ^ n9346 ^ 1'b0 ;
  assign n19029 = n9486 & n19028 ;
  assign n19030 = ( n12964 & n14887 ) | ( n12964 & ~n19029 ) | ( n14887 & ~n19029 ) ;
  assign n19032 = n7357 & ~n14443 ;
  assign n19033 = n19032 ^ x141 ^ 1'b0 ;
  assign n19031 = n3730 & n5493 ;
  assign n19034 = n19033 ^ n19031 ^ 1'b0 ;
  assign n19035 = ( n10454 & ~n19030 ) | ( n10454 & n19034 ) | ( ~n19030 & n19034 ) ;
  assign n19037 = n1247 & n13584 ;
  assign n19038 = x222 & n19037 ;
  assign n19036 = ( n2820 & ~n9344 ) | ( n2820 & n11021 ) | ( ~n9344 & n11021 ) ;
  assign n19039 = n19038 ^ n19036 ^ n2542 ;
  assign n19047 = n2948 ^ n1279 ^ 1'b0 ;
  assign n19044 = ( ~n764 & n6111 ) | ( ~n764 & n9793 ) | ( n6111 & n9793 ) ;
  assign n19045 = n14628 ^ n11227 ^ n2364 ;
  assign n19046 = n19044 & n19045 ;
  assign n19048 = n19047 ^ n19046 ^ 1'b0 ;
  assign n19049 = n12215 | n19048 ;
  assign n19050 = n2520 & ~n19049 ;
  assign n19040 = n2118 | n4493 ;
  assign n19041 = n14749 ^ n4123 ^ 1'b0 ;
  assign n19042 = n19041 ^ n4909 ^ 1'b0 ;
  assign n19043 = ~n19040 & n19042 ;
  assign n19051 = n19050 ^ n19043 ^ n3853 ;
  assign n19056 = ( n559 & ~n7913 ) | ( n559 & n14600 ) | ( ~n7913 & n14600 ) ;
  assign n19052 = n2720 & ~n9753 ;
  assign n19053 = n19052 ^ n363 ^ x60 ;
  assign n19054 = ~n3230 & n19053 ;
  assign n19055 = ~n10996 & n19054 ;
  assign n19057 = n19056 ^ n19055 ^ n3039 ;
  assign n19058 = n16829 ^ n13284 ^ n11498 ;
  assign n19059 = n11759 ^ n6882 ^ 1'b0 ;
  assign n19060 = n9295 ^ n6797 ^ n2356 ;
  assign n19061 = n3109 ^ n2677 ^ 1'b0 ;
  assign n19062 = n19061 ^ n10169 ^ 1'b0 ;
  assign n19066 = n7788 & n15515 ;
  assign n19067 = n19066 ^ n2922 ^ 1'b0 ;
  assign n19063 = ( n986 & ~n2608 ) | ( n986 & n7318 ) | ( ~n2608 & n7318 ) ;
  assign n19064 = n19063 ^ n18246 ^ n6617 ;
  assign n19065 = n19064 ^ n9467 ^ x120 ;
  assign n19068 = n19067 ^ n19065 ^ n7948 ;
  assign n19069 = ( n5635 & n16645 ) | ( n5635 & ~n19068 ) | ( n16645 & ~n19068 ) ;
  assign n19070 = n17301 ^ n5447 ^ n2818 ;
  assign n19071 = n10762 ^ n4594 ^ n944 ;
  assign n19072 = n12190 & ~n19071 ;
  assign n19073 = n19072 ^ n9341 ^ 1'b0 ;
  assign n19074 = n19073 ^ n7038 ^ 1'b0 ;
  assign n19075 = ~n19070 & n19074 ;
  assign n19076 = ( n1546 & n13145 ) | ( n1546 & n16250 ) | ( n13145 & n16250 ) ;
  assign n19077 = n5662 & ~n19076 ;
  assign n19078 = n19077 ^ n2190 ^ 1'b0 ;
  assign n19079 = n19078 ^ n10189 ^ n890 ;
  assign n19080 = n6774 & n9575 ;
  assign n19081 = n19080 ^ n5663 ^ 1'b0 ;
  assign n19082 = ~n17279 & n19081 ;
  assign n19083 = n19082 ^ n1302 ^ 1'b0 ;
  assign n19084 = n968 & n994 ;
  assign n19085 = ( n353 & n6099 ) | ( n353 & n12025 ) | ( n6099 & n12025 ) ;
  assign n19086 = ( ~n341 & n1926 ) | ( ~n341 & n2100 ) | ( n1926 & n2100 ) ;
  assign n19087 = n4115 & ~n19086 ;
  assign n19088 = n5110 ^ n2633 ^ 1'b0 ;
  assign n19089 = n19088 ^ n16604 ^ 1'b0 ;
  assign n19090 = ( ~n7237 & n17434 ) | ( ~n7237 & n19089 ) | ( n17434 & n19089 ) ;
  assign n19091 = n17605 ^ n8751 ^ n8552 ;
  assign n19092 = n9398 ^ n8976 ^ n8580 ;
  assign n19093 = n18797 & ~n19092 ;
  assign n19094 = ( ~n12330 & n19091 ) | ( ~n12330 & n19093 ) | ( n19091 & n19093 ) ;
  assign n19095 = ( n8478 & n9230 ) | ( n8478 & n19094 ) | ( n9230 & n19094 ) ;
  assign n19096 = n19095 ^ n13355 ^ n6935 ;
  assign n19098 = n19027 ^ n9293 ^ n8161 ;
  assign n19097 = ~n3973 & n14749 ;
  assign n19099 = n19098 ^ n19097 ^ 1'b0 ;
  assign n19100 = n1379 | n15915 ;
  assign n19101 = n19100 ^ n6955 ^ 1'b0 ;
  assign n19102 = n19101 ^ n3519 ^ x227 ;
  assign n19103 = ( ~n8158 & n19099 ) | ( ~n8158 & n19102 ) | ( n19099 & n19102 ) ;
  assign n19104 = ( n8860 & ~n15825 ) | ( n8860 & n19103 ) | ( ~n15825 & n19103 ) ;
  assign n19105 = ( n6733 & n8327 ) | ( n6733 & ~n19104 ) | ( n8327 & ~n19104 ) ;
  assign n19106 = n18589 ^ n10827 ^ n2441 ;
  assign n19107 = n19106 ^ n10936 ^ n6956 ;
  assign n19108 = ~n5592 & n6873 ;
  assign n19109 = ( n578 & n9609 ) | ( n578 & ~n18857 ) | ( n9609 & ~n18857 ) ;
  assign n19110 = ( n819 & ~n17136 ) | ( n819 & n19109 ) | ( ~n17136 & n19109 ) ;
  assign n19111 = ( n19107 & n19108 ) | ( n19107 & n19110 ) | ( n19108 & n19110 ) ;
  assign n19112 = n6985 ^ n5705 ^ n1137 ;
  assign n19122 = n15225 ^ n3441 ^ 1'b0 ;
  assign n19123 = n1865 & n19122 ;
  assign n19121 = n10817 ^ n3615 ^ 1'b0 ;
  assign n19117 = n5117 ^ n1484 ^ 1'b0 ;
  assign n19118 = n2226 & ~n19117 ;
  assign n19119 = ( ~n1407 & n2621 ) | ( ~n1407 & n19118 ) | ( n2621 & n19118 ) ;
  assign n19115 = x119 & ~n4373 ;
  assign n19116 = n19115 ^ n14711 ^ n4870 ;
  assign n19113 = ~n15600 & n19004 ;
  assign n19114 = n11673 & n19113 ;
  assign n19120 = n19119 ^ n19116 ^ n19114 ;
  assign n19124 = n19123 ^ n19121 ^ n19120 ;
  assign n19125 = n1387 & ~n3004 ;
  assign n19126 = n19125 ^ n9305 ^ 1'b0 ;
  assign n19127 = n3523 ^ n603 ^ 1'b0 ;
  assign n19128 = ~n11991 & n19127 ;
  assign n19129 = n19128 ^ n3104 ^ 1'b0 ;
  assign n19130 = ( n2399 & n13666 ) | ( n2399 & n18751 ) | ( n13666 & n18751 ) ;
  assign n19131 = n9376 | n19130 ;
  assign n19132 = ( n4175 & n8694 ) | ( n4175 & ~n19131 ) | ( n8694 & ~n19131 ) ;
  assign n19133 = n2608 | n13971 ;
  assign n19134 = n17773 ^ n3333 ^ n1894 ;
  assign n19135 = ( n10597 & n17936 ) | ( n10597 & n19134 ) | ( n17936 & n19134 ) ;
  assign n19136 = ~n3160 & n6543 ;
  assign n19137 = n19136 ^ n6977 ^ n6083 ;
  assign n19138 = n838 & ~n2169 ;
  assign n19139 = n19138 ^ n5242 ^ 1'b0 ;
  assign n19140 = n817 & ~n19139 ;
  assign n19141 = n19140 ^ n3422 ^ 1'b0 ;
  assign n19142 = n10582 ^ n9995 ^ x33 ;
  assign n19143 = n15804 ^ n2801 ^ n2005 ;
  assign n19144 = n19143 ^ n11457 ^ n5511 ;
  assign n19145 = n9601 & ~n19144 ;
  assign n19146 = ~n3522 & n19145 ;
  assign n19147 = n7182 | n19146 ;
  assign n19148 = n4221 & ~n19147 ;
  assign n19149 = n4865 & ~n19148 ;
  assign n19150 = n19142 & n19149 ;
  assign n19151 = ( n8391 & n19141 ) | ( n8391 & ~n19150 ) | ( n19141 & ~n19150 ) ;
  assign n19152 = n845 & n15314 ;
  assign n19153 = ( n10059 & n19015 ) | ( n10059 & n19152 ) | ( n19015 & n19152 ) ;
  assign n19154 = n18212 ^ n11053 ^ n3059 ;
  assign n19162 = n3561 & n7120 ;
  assign n19163 = n19162 ^ n8494 ^ 1'b0 ;
  assign n19155 = n17054 ^ n9362 ^ n418 ;
  assign n19156 = ( ~n453 & n469 ) | ( ~n453 & n2422 ) | ( n469 & n2422 ) ;
  assign n19157 = n1675 & n2996 ;
  assign n19158 = ( ~n11274 & n19156 ) | ( ~n11274 & n19157 ) | ( n19156 & n19157 ) ;
  assign n19159 = ( ~n2778 & n8050 ) | ( ~n2778 & n19158 ) | ( n8050 & n19158 ) ;
  assign n19160 = n8421 & ~n19159 ;
  assign n19161 = n19155 | n19160 ;
  assign n19164 = n19163 ^ n19161 ^ 1'b0 ;
  assign n19165 = n4017 ^ n3213 ^ 1'b0 ;
  assign n19166 = ~n14319 & n19165 ;
  assign n19167 = n1773 ^ n803 ^ 1'b0 ;
  assign n19168 = ~n3620 & n4072 ;
  assign n19169 = n3620 & n19168 ;
  assign n19170 = n19167 & ~n19169 ;
  assign n19171 = ~n19167 & n19170 ;
  assign n19172 = ( x54 & n370 ) | ( x54 & ~n4154 ) | ( n370 & ~n4154 ) ;
  assign n19173 = ~n6799 & n18664 ;
  assign n19174 = ~n9773 & n19173 ;
  assign n19175 = n19174 ^ n16905 ^ 1'b0 ;
  assign n19176 = ( n2770 & ~n19172 ) | ( n2770 & n19175 ) | ( ~n19172 & n19175 ) ;
  assign n19177 = ( n8644 & ~n19171 ) | ( n8644 & n19176 ) | ( ~n19171 & n19176 ) ;
  assign n19178 = n10111 & ~n10296 ;
  assign n19179 = n16203 ^ n2969 ^ 1'b0 ;
  assign n19180 = n829 | n6139 ;
  assign n19181 = n19179 & ~n19180 ;
  assign n19182 = n2183 | n17889 ;
  assign n19183 = n19182 ^ n2606 ^ 1'b0 ;
  assign n19184 = n17959 ^ n6320 ^ n2323 ;
  assign n19185 = n3216 | n16877 ;
  assign n19187 = n1428 & n7848 ;
  assign n19188 = n948 & n19187 ;
  assign n19186 = n3746 | n6202 ;
  assign n19189 = n19188 ^ n19186 ^ 1'b0 ;
  assign n19190 = n13554 ^ n11208 ^ 1'b0 ;
  assign n19191 = ( n9164 & n11393 ) | ( n9164 & ~n19190 ) | ( n11393 & ~n19190 ) ;
  assign n19192 = n378 & ~n3581 ;
  assign n19193 = n5917 & n19192 ;
  assign n19194 = n5711 | n8067 ;
  assign n19195 = ( n1312 & n19193 ) | ( n1312 & n19194 ) | ( n19193 & n19194 ) ;
  assign n19196 = ( ~n17992 & n19191 ) | ( ~n17992 & n19195 ) | ( n19191 & n19195 ) ;
  assign n19197 = ( n3204 & ~n10504 ) | ( n3204 & n14729 ) | ( ~n10504 & n14729 ) ;
  assign n19198 = ( ~n4807 & n15869 ) | ( ~n4807 & n19197 ) | ( n15869 & n19197 ) ;
  assign n19199 = n6029 ^ n5418 ^ 1'b0 ;
  assign n19200 = n13944 ^ n13052 ^ n4456 ;
  assign n19204 = ~n4331 & n6577 ;
  assign n19205 = ~n7337 & n19204 ;
  assign n19201 = n2125 & ~n6042 ;
  assign n19202 = n19201 ^ n10701 ^ 1'b0 ;
  assign n19203 = n19202 ^ n10617 ^ n4438 ;
  assign n19206 = n19205 ^ n19203 ^ n16365 ;
  assign n19207 = ( n1796 & ~n19200 ) | ( n1796 & n19206 ) | ( ~n19200 & n19206 ) ;
  assign n19208 = n9678 & ~n11534 ;
  assign n19209 = n19207 & n19208 ;
  assign n19211 = n10224 ^ n1326 ^ 1'b0 ;
  assign n19212 = n9870 & ~n19211 ;
  assign n19210 = ( n3769 & n11736 ) | ( n3769 & n15361 ) | ( n11736 & n15361 ) ;
  assign n19213 = n19212 ^ n19210 ^ n3472 ;
  assign n19214 = ( n5214 & ~n17430 ) | ( n5214 & n19213 ) | ( ~n17430 & n19213 ) ;
  assign n19215 = n3970 ^ n3862 ^ n1380 ;
  assign n19216 = ( n1107 & n15395 ) | ( n1107 & n19215 ) | ( n15395 & n19215 ) ;
  assign n19217 = ( n1127 & n2092 ) | ( n1127 & ~n9127 ) | ( n2092 & ~n9127 ) ;
  assign n19218 = n11615 ^ x184 ^ 1'b0 ;
  assign n19219 = n19217 | n19218 ;
  assign n19220 = n19219 ^ n5172 ^ 1'b0 ;
  assign n19221 = n19216 & ~n19220 ;
  assign n19222 = n1970 & ~n13155 ;
  assign n19223 = ( n17264 & n19221 ) | ( n17264 & n19222 ) | ( n19221 & n19222 ) ;
  assign n19224 = ( n2306 & n5492 ) | ( n2306 & ~n9044 ) | ( n5492 & ~n9044 ) ;
  assign n19225 = n19224 ^ n7662 ^ n2295 ;
  assign n19226 = n14246 ^ n2689 ^ n298 ;
  assign n19227 = n10530 ^ n6463 ^ n2634 ;
  assign n19228 = ( ~n7570 & n19226 ) | ( ~n7570 & n19227 ) | ( n19226 & n19227 ) ;
  assign n19229 = ( n6221 & ~n14268 ) | ( n6221 & n19228 ) | ( ~n14268 & n19228 ) ;
  assign n19230 = n7846 ^ n7451 ^ n5565 ;
  assign n19231 = ( n1597 & ~n6037 ) | ( n1597 & n6363 ) | ( ~n6037 & n6363 ) ;
  assign n19232 = ~n11133 & n14892 ;
  assign n19233 = n19232 ^ n8699 ^ 1'b0 ;
  assign n19234 = n10101 | n19233 ;
  assign n19235 = n19231 & ~n19234 ;
  assign n19236 = n19235 ^ n9714 ^ n4249 ;
  assign n19237 = n4156 | n7282 ;
  assign n19238 = n19237 ^ n5874 ^ 1'b0 ;
  assign n19239 = n7977 ^ n2234 ^ 1'b0 ;
  assign n19240 = ( n13620 & n19238 ) | ( n13620 & ~n19239 ) | ( n19238 & ~n19239 ) ;
  assign n19241 = n3997 | n12784 ;
  assign n19242 = n8714 ^ n8026 ^ 1'b0 ;
  assign n19243 = ~n19241 & n19242 ;
  assign n19244 = n2827 ^ n1828 ^ 1'b0 ;
  assign n19245 = n19244 ^ n15544 ^ 1'b0 ;
  assign n19246 = ~n8438 & n19245 ;
  assign n19247 = ( n8356 & ~n9079 ) | ( n8356 & n19246 ) | ( ~n9079 & n19246 ) ;
  assign n19250 = ( n909 & n1457 ) | ( n909 & n7403 ) | ( n1457 & n7403 ) ;
  assign n19248 = ( n2433 & n4418 ) | ( n2433 & n6898 ) | ( n4418 & n6898 ) ;
  assign n19249 = n19248 ^ n7871 ^ n2501 ;
  assign n19251 = n19250 ^ n19249 ^ n12873 ;
  assign n19252 = n4621 | n7952 ;
  assign n19253 = n19252 ^ n9611 ^ n5611 ;
  assign n19259 = n13000 ^ n5790 ^ 1'b0 ;
  assign n19260 = n8036 & ~n19259 ;
  assign n19254 = ~n1657 & n9496 ;
  assign n19255 = ~n2851 & n19254 ;
  assign n19256 = n19255 ^ n10259 ^ 1'b0 ;
  assign n19257 = ( n13978 & n16678 ) | ( n13978 & ~n19256 ) | ( n16678 & ~n19256 ) ;
  assign n19258 = n19257 ^ n10027 ^ n787 ;
  assign n19261 = n19260 ^ n19258 ^ n16633 ;
  assign n19262 = n7068 ^ n4158 ^ n2185 ;
  assign n19263 = n799 | n19262 ;
  assign n19264 = n17174 & ~n19263 ;
  assign n19265 = n2011 & ~n11462 ;
  assign n19266 = n5651 & n19265 ;
  assign n19267 = n11955 ^ n10965 ^ n10239 ;
  assign n19268 = ( n7736 & ~n19266 ) | ( n7736 & n19267 ) | ( ~n19266 & n19267 ) ;
  assign n19269 = ( n895 & ~n16203 ) | ( n895 & n19268 ) | ( ~n16203 & n19268 ) ;
  assign n19270 = ( n3007 & ~n6046 ) | ( n3007 & n19269 ) | ( ~n6046 & n19269 ) ;
  assign n19271 = ( n4339 & n7199 ) | ( n4339 & ~n19231 ) | ( n7199 & ~n19231 ) ;
  assign n19272 = ( ~n11255 & n11640 ) | ( ~n11255 & n19271 ) | ( n11640 & n19271 ) ;
  assign n19273 = ( ~n3185 & n7156 ) | ( ~n3185 & n15900 ) | ( n7156 & n15900 ) ;
  assign n19274 = n19273 ^ n15547 ^ n3845 ;
  assign n19275 = ( n2193 & ~n8069 ) | ( n2193 & n19274 ) | ( ~n8069 & n19274 ) ;
  assign n19276 = ( n4890 & n14703 ) | ( n4890 & n19275 ) | ( n14703 & n19275 ) ;
  assign n19277 = n2818 | n14564 ;
  assign n19278 = x240 & n9444 ;
  assign n19279 = ~n5155 & n19278 ;
  assign n19283 = ( n4547 & n6759 ) | ( n4547 & ~n8097 ) | ( n6759 & ~n8097 ) ;
  assign n19284 = ( n3458 & n9632 ) | ( n3458 & n19283 ) | ( n9632 & n19283 ) ;
  assign n19280 = n6685 & ~n8720 ;
  assign n19281 = ~n9337 & n19280 ;
  assign n19282 = n19281 ^ n8211 ^ x44 ;
  assign n19285 = n19284 ^ n19282 ^ 1'b0 ;
  assign n19286 = ~n19279 & n19285 ;
  assign n19287 = ( n2200 & ~n12101 ) | ( n2200 & n13493 ) | ( ~n12101 & n13493 ) ;
  assign n19292 = n7375 | n12413 ;
  assign n19293 = n14675 | n19292 ;
  assign n19289 = n8372 ^ n7454 ^ n3154 ;
  assign n19290 = ~n14713 & n19289 ;
  assign n19291 = n11567 & n19290 ;
  assign n19294 = n19293 ^ n19291 ^ 1'b0 ;
  assign n19288 = n438 ^ n330 ^ 1'b0 ;
  assign n19295 = n19294 ^ n19288 ^ n2678 ;
  assign n19297 = n1870 & n4261 ;
  assign n19298 = n19297 ^ n12863 ^ n9651 ;
  assign n19299 = ( n3646 & n3887 ) | ( n3646 & ~n19298 ) | ( n3887 & ~n19298 ) ;
  assign n19300 = ( n3082 & ~n16241 ) | ( n3082 & n19299 ) | ( ~n16241 & n19299 ) ;
  assign n19296 = ~n13926 & n17877 ;
  assign n19301 = n19300 ^ n19296 ^ 1'b0 ;
  assign n19302 = n486 & n1376 ;
  assign n19303 = n19302 ^ n10415 ^ 1'b0 ;
  assign n19304 = n10657 ^ n5873 ^ n4822 ;
  assign n19305 = n19303 | n19304 ;
  assign n19306 = ~n441 & n15904 ;
  assign n19307 = n19306 ^ n487 ^ 1'b0 ;
  assign n19308 = ( n932 & n8793 ) | ( n932 & n13719 ) | ( n8793 & n13719 ) ;
  assign n19309 = n15900 ^ n4922 ^ n2306 ;
  assign n19310 = n19309 ^ n12443 ^ 1'b0 ;
  assign n19311 = n7770 | n19310 ;
  assign n19312 = ~n7223 & n13307 ;
  assign n19313 = n19312 ^ n304 ^ 1'b0 ;
  assign n19314 = ( n1023 & n1296 ) | ( n1023 & n2584 ) | ( n1296 & n2584 ) ;
  assign n19315 = ( n989 & n9420 ) | ( n989 & ~n10721 ) | ( n9420 & ~n10721 ) ;
  assign n19316 = n8637 ^ n1933 ^ 1'b0 ;
  assign n19317 = n19315 & ~n19316 ;
  assign n19318 = ( n7996 & n19314 ) | ( n7996 & ~n19317 ) | ( n19314 & ~n19317 ) ;
  assign n19319 = ( n3898 & ~n7152 ) | ( n3898 & n8499 ) | ( ~n7152 & n8499 ) ;
  assign n19320 = n13184 | n19319 ;
  assign n19321 = n10216 | n19320 ;
  assign n19322 = n5374 & ~n7344 ;
  assign n19323 = n15847 & n19322 ;
  assign n19324 = ( ~n1356 & n10034 ) | ( ~n1356 & n17002 ) | ( n10034 & n17002 ) ;
  assign n19325 = n19324 ^ n18126 ^ n6508 ;
  assign n19326 = ( ~n1583 & n6850 ) | ( ~n1583 & n8548 ) | ( n6850 & n8548 ) ;
  assign n19327 = ( n2223 & n3241 ) | ( n2223 & ~n6749 ) | ( n3241 & ~n6749 ) ;
  assign n19328 = ( n8800 & n11955 ) | ( n8800 & n19327 ) | ( n11955 & n19327 ) ;
  assign n19329 = n19328 ^ n10037 ^ n7488 ;
  assign n19330 = n11080 & n19329 ;
  assign n19331 = ~n19326 & n19330 ;
  assign n19332 = x231 & n8450 ;
  assign n19333 = ~n5454 & n19332 ;
  assign n19335 = n3196 ^ n1136 ^ 1'b0 ;
  assign n19336 = x144 & n5110 ;
  assign n19337 = n19336 ^ n3656 ^ 1'b0 ;
  assign n19338 = ( n5000 & n19335 ) | ( n5000 & ~n19337 ) | ( n19335 & ~n19337 ) ;
  assign n19334 = n10543 | n13438 ;
  assign n19339 = n19338 ^ n19334 ^ 1'b0 ;
  assign n19342 = ( n556 & n3371 ) | ( n556 & n9443 ) | ( n3371 & n9443 ) ;
  assign n19340 = n5374 & ~n15026 ;
  assign n19341 = n3811 & n19340 ;
  assign n19343 = n19342 ^ n19341 ^ 1'b0 ;
  assign n19344 = n18038 & ~n19343 ;
  assign n19345 = x2 & ~n6755 ;
  assign n19346 = ( n1119 & n2364 ) | ( n1119 & n19345 ) | ( n2364 & n19345 ) ;
  assign n19347 = n19346 ^ n12572 ^ 1'b0 ;
  assign n19348 = n4312 & n19347 ;
  assign n19359 = n1521 & ~n5175 ;
  assign n19354 = n16455 ^ x212 ^ 1'b0 ;
  assign n19355 = ( n6379 & ~n14941 ) | ( n6379 & n19354 ) | ( ~n14941 & n19354 ) ;
  assign n19356 = n1762 | n4124 ;
  assign n19357 = n19355 | n19356 ;
  assign n19358 = n19357 ^ n9131 ^ n8273 ;
  assign n19352 = n4357 ^ n3137 ^ n1884 ;
  assign n19349 = n4795 ^ n3078 ^ n1072 ;
  assign n19350 = ( n1446 & n11409 ) | ( n1446 & ~n19349 ) | ( n11409 & ~n19349 ) ;
  assign n19351 = n19350 ^ n2020 ^ 1'b0 ;
  assign n19353 = n19352 ^ n19351 ^ n7981 ;
  assign n19360 = n19359 ^ n19358 ^ n19353 ;
  assign n19361 = n536 | n15533 ;
  assign n19362 = n17167 ^ n6408 ^ n6095 ;
  assign n19363 = ( n4692 & ~n7328 ) | ( n4692 & n10316 ) | ( ~n7328 & n10316 ) ;
  assign n19364 = n1426 & n19363 ;
  assign n19365 = n19364 ^ n16453 ^ n11252 ;
  assign n19366 = n2828 & n19365 ;
  assign n19367 = n4228 & n7687 ;
  assign n19368 = n19367 ^ n2132 ^ 1'b0 ;
  assign n19369 = ( n4751 & n14490 ) | ( n4751 & ~n19368 ) | ( n14490 & ~n19368 ) ;
  assign n19370 = ( x62 & n11149 ) | ( x62 & ~n19369 ) | ( n11149 & ~n19369 ) ;
  assign n19371 = n19370 ^ n10326 ^ 1'b0 ;
  assign n19372 = ~n536 & n14217 ;
  assign n19373 = n19372 ^ n541 ^ n393 ;
  assign n19374 = n3146 & ~n16327 ;
  assign n19375 = ~n19373 & n19374 ;
  assign n19376 = ( n6673 & n14736 ) | ( n6673 & ~n16485 ) | ( n14736 & ~n16485 ) ;
  assign n19377 = n606 | n920 ;
  assign n19378 = n13824 & ~n19377 ;
  assign n19379 = n17959 | n19378 ;
  assign n19380 = n3954 & n15699 ;
  assign n19381 = n2847 | n4334 ;
  assign n19382 = n8750 & ~n19381 ;
  assign n19383 = ~n1909 & n13856 ;
  assign n19384 = n19382 & n19383 ;
  assign n19385 = n19384 ^ n13558 ^ n566 ;
  assign n19386 = ( ~n11603 & n12563 ) | ( ~n11603 & n19385 ) | ( n12563 & n19385 ) ;
  assign n19387 = n10152 ^ n9271 ^ n4104 ;
  assign n19389 = n572 & ~n10755 ;
  assign n19390 = n19389 ^ n10557 ^ 1'b0 ;
  assign n19388 = n2884 & ~n14723 ;
  assign n19391 = n19390 ^ n19388 ^ 1'b0 ;
  assign n19392 = ~n19387 & n19391 ;
  assign n19393 = n12346 ^ n1516 ^ 1'b0 ;
  assign n19394 = n9525 ^ n6160 ^ n3465 ;
  assign n19395 = ( n2248 & ~n17935 ) | ( n2248 & n19394 ) | ( ~n17935 & n19394 ) ;
  assign n19396 = ~n11582 & n19395 ;
  assign n19397 = ( n10094 & ~n19393 ) | ( n10094 & n19396 ) | ( ~n19393 & n19396 ) ;
  assign n19406 = n15833 ^ n12952 ^ 1'b0 ;
  assign n19398 = n12188 ^ n10672 ^ 1'b0 ;
  assign n19399 = ( n1214 & ~n9094 ) | ( n1214 & n19398 ) | ( ~n9094 & n19398 ) ;
  assign n19400 = n6817 & n15546 ;
  assign n19401 = n19400 ^ n11295 ^ 1'b0 ;
  assign n19402 = ( n2305 & n6159 ) | ( n2305 & ~n19401 ) | ( n6159 & ~n19401 ) ;
  assign n19403 = n19399 & n19402 ;
  assign n19404 = ~n18619 & n19403 ;
  assign n19405 = n3593 | n19404 ;
  assign n19407 = n19406 ^ n19405 ^ 1'b0 ;
  assign n19410 = ~n5445 & n9575 ;
  assign n19411 = n19410 ^ n6521 ^ 1'b0 ;
  assign n19412 = n19411 ^ n9594 ^ n1750 ;
  assign n19413 = n19412 ^ n17066 ^ n4381 ;
  assign n19408 = n7217 | n13007 ;
  assign n19409 = n2428 & ~n19408 ;
  assign n19414 = n19413 ^ n19409 ^ n8225 ;
  assign n19415 = n12980 ^ n10755 ^ n7766 ;
  assign n19416 = ( n8041 & n12708 ) | ( n8041 & ~n19415 ) | ( n12708 & ~n19415 ) ;
  assign n19417 = n6608 & ~n11923 ;
  assign n19418 = n13610 & n19417 ;
  assign n19419 = ( n838 & n2754 ) | ( n838 & ~n3600 ) | ( n2754 & ~n3600 ) ;
  assign n19420 = ( n845 & ~n10963 ) | ( n845 & n19419 ) | ( ~n10963 & n19419 ) ;
  assign n19421 = n5225 & n19420 ;
  assign n19422 = n19421 ^ n4895 ^ 1'b0 ;
  assign n19423 = ~n14320 & n19422 ;
  assign n19424 = n17945 ^ n7095 ^ 1'b0 ;
  assign n19425 = n19424 ^ n12523 ^ 1'b0 ;
  assign n19426 = ( x232 & ~n13584 ) | ( x232 & n19425 ) | ( ~n13584 & n19425 ) ;
  assign n19427 = ( n4234 & ~n17466 ) | ( n4234 & n19426 ) | ( ~n17466 & n19426 ) ;
  assign n19428 = ( n6705 & n12287 ) | ( n6705 & ~n12848 ) | ( n12287 & ~n12848 ) ;
  assign n19435 = x54 & n751 ;
  assign n19436 = n5554 & n19435 ;
  assign n19437 = n19436 ^ n10574 ^ n2174 ;
  assign n19429 = n7244 ^ n3973 ^ n1971 ;
  assign n19430 = n4492 & n19429 ;
  assign n19431 = ~n10643 & n19430 ;
  assign n19432 = ( n7853 & n14143 ) | ( n7853 & ~n19431 ) | ( n14143 & ~n19431 ) ;
  assign n19433 = n19432 ^ n13809 ^ 1'b0 ;
  assign n19434 = n10802 | n19433 ;
  assign n19438 = n19437 ^ n19434 ^ 1'b0 ;
  assign n19439 = ~n3044 & n19438 ;
  assign n19440 = ( n938 & n4170 ) | ( n938 & ~n15633 ) | ( n4170 & ~n15633 ) ;
  assign n19441 = n4976 & ~n9503 ;
  assign n19442 = n5077 ^ n2221 ^ 1'b0 ;
  assign n19443 = ( n389 & ~n19441 ) | ( n389 & n19442 ) | ( ~n19441 & n19442 ) ;
  assign n19444 = n19443 ^ n17036 ^ 1'b0 ;
  assign n19445 = n18190 ^ n7532 ^ n438 ;
  assign n19446 = ( n1575 & ~n7181 ) | ( n1575 & n16036 ) | ( ~n7181 & n16036 ) ;
  assign n19447 = n17278 & n19446 ;
  assign n19448 = ~n7439 & n19447 ;
  assign n19449 = n19445 | n19448 ;
  assign n19450 = n5661 ^ n2357 ^ n2047 ;
  assign n19451 = ~n1134 & n9853 ;
  assign n19452 = ( n7565 & n19450 ) | ( n7565 & n19451 ) | ( n19450 & n19451 ) ;
  assign n19453 = n19452 ^ n14347 ^ n5809 ;
  assign n19454 = ( n6186 & ~n8790 ) | ( n6186 & n9486 ) | ( ~n8790 & n9486 ) ;
  assign n19455 = ( n1958 & ~n4044 ) | ( n1958 & n19454 ) | ( ~n4044 & n19454 ) ;
  assign n19456 = n7330 & n19455 ;
  assign n19457 = n3319 & n19456 ;
  assign n19458 = ( ~n12308 & n13195 ) | ( ~n12308 & n19457 ) | ( n13195 & n19457 ) ;
  assign n19461 = n4494 & ~n6307 ;
  assign n19459 = n11712 ^ n489 ^ 1'b0 ;
  assign n19460 = ~n1398 & n19459 ;
  assign n19462 = n19461 ^ n19460 ^ 1'b0 ;
  assign n19464 = n17218 ^ n13146 ^ 1'b0 ;
  assign n19465 = n18634 & ~n19464 ;
  assign n19463 = ~n4012 & n13658 ;
  assign n19466 = n19465 ^ n19463 ^ 1'b0 ;
  assign n19467 = n6050 ^ n5042 ^ n2644 ;
  assign n19468 = n5506 ^ n676 ^ 1'b0 ;
  assign n19469 = ~n7415 & n19468 ;
  assign n19470 = ( n9943 & ~n19467 ) | ( n9943 & n19469 ) | ( ~n19467 & n19469 ) ;
  assign n19471 = n18013 ^ n1498 ^ 1'b0 ;
  assign n19472 = ( ~n5740 & n13180 ) | ( ~n5740 & n19471 ) | ( n13180 & n19471 ) ;
  assign n19473 = ( n4269 & n7635 ) | ( n4269 & n13793 ) | ( n7635 & n13793 ) ;
  assign n19474 = ( ~n1237 & n2259 ) | ( ~n1237 & n6079 ) | ( n2259 & n6079 ) ;
  assign n19475 = n19474 ^ n13137 ^ 1'b0 ;
  assign n19476 = n19473 & ~n19475 ;
  assign n19477 = n18489 ^ n3844 ^ n586 ;
  assign n19478 = n19477 ^ n19091 ^ n3800 ;
  assign n19479 = n17553 ^ n15851 ^ n6012 ;
  assign n19480 = ( n19476 & n19478 ) | ( n19476 & n19479 ) | ( n19478 & n19479 ) ;
  assign n19481 = ( n11546 & ~n19472 ) | ( n11546 & n19480 ) | ( ~n19472 & n19480 ) ;
  assign n19482 = n15189 | n17102 ;
  assign n19483 = ( ~n6052 & n6996 ) | ( ~n6052 & n19482 ) | ( n6996 & n19482 ) ;
  assign n19484 = n17879 & n19483 ;
  assign n19485 = ~n3985 & n19484 ;
  assign n19486 = ( ~n4322 & n17564 ) | ( ~n4322 & n17793 ) | ( n17564 & n17793 ) ;
  assign n19487 = ( ~n3609 & n4574 ) | ( ~n3609 & n19486 ) | ( n4574 & n19486 ) ;
  assign n19488 = ( n3426 & n4514 ) | ( n3426 & ~n19487 ) | ( n4514 & ~n19487 ) ;
  assign n19489 = n16018 ^ n9663 ^ n2890 ;
  assign n19490 = n19489 ^ n16495 ^ n2124 ;
  assign n19491 = ( ~n3977 & n6577 ) | ( ~n3977 & n6921 ) | ( n6577 & n6921 ) ;
  assign n19492 = n19491 ^ n13109 ^ n5062 ;
  assign n19493 = n9812 ^ n8867 ^ n7523 ;
  assign n19494 = ( n5177 & n15788 ) | ( n5177 & ~n19493 ) | ( n15788 & ~n19493 ) ;
  assign n19495 = n14215 | n19494 ;
  assign n19496 = n14706 & ~n19495 ;
  assign n19497 = n12553 ^ n6584 ^ n1635 ;
  assign n19498 = ~n14391 & n19497 ;
  assign n19499 = n19496 & n19498 ;
  assign n19500 = n4147 ^ n1028 ^ 1'b0 ;
  assign n19501 = n17369 & n19500 ;
  assign n19502 = ~x22 & n19501 ;
  assign n19503 = n11526 ^ n10082 ^ n5576 ;
  assign n19504 = n6569 ^ n5642 ^ 1'b0 ;
  assign n19505 = n19503 & ~n19504 ;
  assign n19506 = ( n2903 & ~n12250 ) | ( n2903 & n18114 ) | ( ~n12250 & n18114 ) ;
  assign n19507 = ( n19275 & n19505 ) | ( n19275 & n19506 ) | ( n19505 & n19506 ) ;
  assign n19508 = n7169 ^ n4084 ^ 1'b0 ;
  assign n19509 = ( n1116 & n1129 ) | ( n1116 & n19508 ) | ( n1129 & n19508 ) ;
  assign n19510 = n19509 ^ n4017 ^ 1'b0 ;
  assign n19511 = n8133 ^ n5487 ^ n3538 ;
  assign n19512 = ~n13805 & n19511 ;
  assign n19513 = ~n12150 & n19512 ;
  assign n19514 = n17754 & n19513 ;
  assign n19515 = ( x102 & ~n2588 ) | ( x102 & n8602 ) | ( ~n2588 & n8602 ) ;
  assign n19516 = n6763 & ~n9719 ;
  assign n19517 = n19516 ^ n9962 ^ 1'b0 ;
  assign n19518 = ( n786 & n834 ) | ( n786 & ~n2392 ) | ( n834 & ~n2392 ) ;
  assign n19519 = n12940 & ~n19518 ;
  assign n19520 = n19517 & n19519 ;
  assign n19521 = n19520 ^ n5386 ^ 1'b0 ;
  assign n19522 = n19515 | n19521 ;
  assign n19523 = n11296 ^ n10457 ^ n6642 ;
  assign n19524 = ( n9188 & ~n12844 ) | ( n9188 & n13489 ) | ( ~n12844 & n13489 ) ;
  assign n19525 = n2860 ^ x243 ^ 1'b0 ;
  assign n19526 = n717 & ~n19525 ;
  assign n19527 = n1215 & n2185 ;
  assign n19528 = ~x216 & n19527 ;
  assign n19529 = n19528 ^ n14221 ^ n6911 ;
  assign n19530 = ~n3351 & n9222 ;
  assign n19531 = n19530 ^ n10446 ^ 1'b0 ;
  assign n19532 = ( n19526 & n19529 ) | ( n19526 & n19531 ) | ( n19529 & n19531 ) ;
  assign n19533 = n19524 | n19532 ;
  assign n19535 = n16522 ^ n8724 ^ n8273 ;
  assign n19534 = n2443 & ~n17024 ;
  assign n19536 = n19535 ^ n19534 ^ 1'b0 ;
  assign n19537 = ( ~n5102 & n12131 ) | ( ~n5102 & n15283 ) | ( n12131 & n15283 ) ;
  assign n19538 = n9621 | n19537 ;
  assign n19539 = n1461 & ~n19538 ;
  assign n19540 = n19539 ^ n1817 ^ 1'b0 ;
  assign n19541 = n19536 | n19540 ;
  assign n19542 = n7273 ^ n6703 ^ n1741 ;
  assign n19543 = ( n3715 & n4081 ) | ( n3715 & n19542 ) | ( n4081 & n19542 ) ;
  assign n19544 = n12097 ^ n6754 ^ 1'b0 ;
  assign n19545 = n19543 & n19544 ;
  assign n19550 = n13131 ^ n10329 ^ 1'b0 ;
  assign n19548 = ~n1473 & n19157 ;
  assign n19546 = n9413 & ~n11617 ;
  assign n19547 = n19546 ^ n7560 ^ n2866 ;
  assign n19549 = n19548 ^ n19547 ^ 1'b0 ;
  assign n19551 = n19550 ^ n19549 ^ n13512 ;
  assign n19552 = n10414 ^ n6170 ^ n2489 ;
  assign n19553 = n7032 & ~n19552 ;
  assign n19554 = n19553 ^ n18752 ^ 1'b0 ;
  assign n19558 = n7723 ^ n6676 ^ n2522 ;
  assign n19559 = n5196 ^ n3779 ^ 1'b0 ;
  assign n19560 = n19558 | n19559 ;
  assign n19561 = ( n2618 & ~n11213 ) | ( n2618 & n19560 ) | ( ~n11213 & n19560 ) ;
  assign n19555 = ( x60 & ~x135 ) | ( x60 & n9782 ) | ( ~x135 & n9782 ) ;
  assign n19556 = ( n4757 & ~n8150 ) | ( n4757 & n19555 ) | ( ~n8150 & n19555 ) ;
  assign n19557 = ~n10176 & n19556 ;
  assign n19562 = n19561 ^ n19557 ^ 1'b0 ;
  assign n19563 = ( ~n3978 & n8835 ) | ( ~n3978 & n9105 ) | ( n8835 & n9105 ) ;
  assign n19564 = n2586 & n19563 ;
  assign n19565 = ~n3962 & n19564 ;
  assign n19566 = n18806 ^ n4389 ^ 1'b0 ;
  assign n19567 = ~n1346 & n4931 ;
  assign n19568 = n19567 ^ n6604 ^ 1'b0 ;
  assign n19569 = ~n11206 & n19568 ;
  assign n19570 = ~n14414 & n19569 ;
  assign n19571 = ( ~x93 & n15567 ) | ( ~x93 & n19570 ) | ( n15567 & n19570 ) ;
  assign n19572 = ~n10285 & n18094 ;
  assign n19573 = n12131 & ~n14098 ;
  assign n19574 = ( n6223 & n19572 ) | ( n6223 & n19573 ) | ( n19572 & n19573 ) ;
  assign n19575 = ( n2025 & ~n2180 ) | ( n2025 & n6930 ) | ( ~n2180 & n6930 ) ;
  assign n19576 = ( n993 & n8283 ) | ( n993 & ~n19575 ) | ( n8283 & ~n19575 ) ;
  assign n19577 = ( n18892 & n19574 ) | ( n18892 & ~n19576 ) | ( n19574 & ~n19576 ) ;
  assign n19578 = n834 | n1808 ;
  assign n19579 = n6327 & ~n6776 ;
  assign n19580 = n19579 ^ n9851 ^ n576 ;
  assign n19581 = n19092 ^ n5616 ^ 1'b0 ;
  assign n19582 = n19580 & ~n19581 ;
  assign n19583 = ( n13664 & ~n15256 ) | ( n13664 & n19582 ) | ( ~n15256 & n19582 ) ;
  assign n19584 = ( n5189 & n7895 ) | ( n5189 & n16544 ) | ( n7895 & n16544 ) ;
  assign n19585 = n19584 ^ n8231 ^ 1'b0 ;
  assign n19586 = n17362 ^ n4818 ^ n3841 ;
  assign n19587 = n710 & ~n4629 ;
  assign n19588 = n19586 & n19587 ;
  assign n19589 = n1236 & n1917 ;
  assign n19590 = n2545 & n19589 ;
  assign n19591 = n19590 ^ n14040 ^ n5136 ;
  assign n19592 = ( ~n11078 & n19588 ) | ( ~n11078 & n19591 ) | ( n19588 & n19591 ) ;
  assign n19593 = ( n3455 & ~n4404 ) | ( n3455 & n17582 ) | ( ~n4404 & n17582 ) ;
  assign n19594 = n12831 ^ n9668 ^ 1'b0 ;
  assign n19595 = n16145 | n19594 ;
  assign n19596 = ~n4928 & n9456 ;
  assign n19597 = ( n1996 & n11348 ) | ( n1996 & ~n19596 ) | ( n11348 & ~n19596 ) ;
  assign n19598 = n8537 ^ n5832 ^ 1'b0 ;
  assign n19599 = ( n1399 & ~n9924 ) | ( n1399 & n10690 ) | ( ~n9924 & n10690 ) ;
  assign n19600 = n19599 ^ n13867 ^ n1428 ;
  assign n19601 = ~n18276 & n19600 ;
  assign n19602 = n19601 ^ n8478 ^ 1'b0 ;
  assign n19610 = n9890 ^ n3949 ^ 1'b0 ;
  assign n19608 = ( x205 & n4789 ) | ( x205 & n6612 ) | ( n4789 & n6612 ) ;
  assign n19606 = n4865 ^ n4796 ^ n491 ;
  assign n19607 = ( n2203 & n6079 ) | ( n2203 & n19606 ) | ( n6079 & n19606 ) ;
  assign n19609 = n19608 ^ n19607 ^ n5668 ;
  assign n19611 = n19610 ^ n19609 ^ n1219 ;
  assign n19603 = x68 & n1590 ;
  assign n19604 = ( n3115 & n13412 ) | ( n3115 & ~n19603 ) | ( n13412 & ~n19603 ) ;
  assign n19605 = n19604 ^ n11953 ^ 1'b0 ;
  assign n19612 = n19611 ^ n19605 ^ n9144 ;
  assign n19613 = n11870 ^ n2736 ^ n2629 ;
  assign n19614 = n11527 ^ n11468 ^ n8465 ;
  assign n19615 = ( n14065 & ~n19613 ) | ( n14065 & n19614 ) | ( ~n19613 & n19614 ) ;
  assign n19616 = n4846 | n6135 ;
  assign n19617 = n19616 ^ n6042 ^ 1'b0 ;
  assign n19618 = ~n4191 & n9482 ;
  assign n19619 = n10689 & n19618 ;
  assign n19620 = n9637 | n19619 ;
  assign n19621 = n1930 | n19620 ;
  assign n19622 = ( n10219 & n19617 ) | ( n10219 & n19621 ) | ( n19617 & n19621 ) ;
  assign n19623 = ( ~n4615 & n8513 ) | ( ~n4615 & n12346 ) | ( n8513 & n12346 ) ;
  assign n19626 = n2770 & n2997 ;
  assign n19624 = n7830 ^ n3722 ^ n277 ;
  assign n19625 = n19624 ^ n4463 ^ n3595 ;
  assign n19627 = n19626 ^ n19625 ^ 1'b0 ;
  assign n19628 = n8470 ^ n7799 ^ 1'b0 ;
  assign n19632 = n863 & n9535 ;
  assign n19633 = n2373 & n19632 ;
  assign n19634 = n7091 & ~n19633 ;
  assign n19635 = n11781 & n19634 ;
  assign n19636 = n19635 ^ n13674 ^ n10822 ;
  assign n19629 = n7675 ^ n7539 ^ 1'b0 ;
  assign n19630 = n15583 | n19629 ;
  assign n19631 = ( ~n1400 & n11065 ) | ( ~n1400 & n19630 ) | ( n11065 & n19630 ) ;
  assign n19637 = n19636 ^ n19631 ^ 1'b0 ;
  assign n19638 = ~n12236 & n17102 ;
  assign n19639 = ~n6984 & n19638 ;
  assign n19640 = ( n1513 & n19050 ) | ( n1513 & ~n19639 ) | ( n19050 & ~n19639 ) ;
  assign n19641 = n19640 ^ n15694 ^ 1'b0 ;
  assign n19642 = ( n1245 & ~n1843 ) | ( n1245 & n5385 ) | ( ~n1843 & n5385 ) ;
  assign n19643 = n7632 | n19642 ;
  assign n19644 = n19643 ^ n15194 ^ 1'b0 ;
  assign n19645 = n8736 & ~n9177 ;
  assign n19647 = n4723 ^ n2668 ^ 1'b0 ;
  assign n19648 = n4448 & ~n19647 ;
  assign n19646 = ( n13814 & ~n15767 ) | ( n13814 & n16487 ) | ( ~n15767 & n16487 ) ;
  assign n19649 = n19648 ^ n19646 ^ n10825 ;
  assign n19650 = ( x96 & n19645 ) | ( x96 & ~n19649 ) | ( n19645 & ~n19649 ) ;
  assign n19651 = n12898 & ~n14491 ;
  assign n19652 = n19651 ^ n5910 ^ 1'b0 ;
  assign n19654 = n549 & n1351 ;
  assign n19653 = n5877 | n10305 ;
  assign n19655 = n19654 ^ n19653 ^ n2036 ;
  assign n19657 = n3596 ^ n1181 ^ 1'b0 ;
  assign n19658 = n8159 | n19657 ;
  assign n19656 = n3517 ^ n2999 ^ n2025 ;
  assign n19659 = n19658 ^ n19656 ^ 1'b0 ;
  assign n19660 = n5630 ^ n5021 ^ n860 ;
  assign n19661 = n9674 & ~n19660 ;
  assign n19662 = n12213 ^ n1553 ^ 1'b0 ;
  assign n19663 = n19662 ^ n15633 ^ n6131 ;
  assign n19664 = ~n4025 & n11092 ;
  assign n19665 = ~n6617 & n19664 ;
  assign n19676 = n6693 ^ n1585 ^ 1'b0 ;
  assign n19677 = n3914 | n19676 ;
  assign n19666 = ( n640 & n1496 ) | ( n640 & n5086 ) | ( n1496 & n5086 ) ;
  assign n19667 = ( ~n4067 & n10728 ) | ( ~n4067 & n19666 ) | ( n10728 & n19666 ) ;
  assign n19668 = n318 & ~n3022 ;
  assign n19669 = n6389 & n19668 ;
  assign n19670 = n7797 & n15833 ;
  assign n19671 = n19262 ^ n11104 ^ n5491 ;
  assign n19672 = n19671 ^ n18895 ^ n5066 ;
  assign n19673 = n19670 & n19672 ;
  assign n19674 = n19669 & n19673 ;
  assign n19675 = n19667 & ~n19674 ;
  assign n19678 = n19677 ^ n19675 ^ 1'b0 ;
  assign n19679 = ( ~n1048 & n2357 ) | ( ~n1048 & n15897 ) | ( n2357 & n15897 ) ;
  assign n19680 = n19679 ^ n16654 ^ 1'b0 ;
  assign n19681 = n15664 & ~n19680 ;
  assign n19684 = n2477 & n5011 ;
  assign n19685 = ( ~n9915 & n14302 ) | ( ~n9915 & n19684 ) | ( n14302 & n19684 ) ;
  assign n19682 = n2357 ^ n592 ^ 1'b0 ;
  assign n19683 = ~n11230 & n19682 ;
  assign n19686 = n19685 ^ n19683 ^ n2457 ;
  assign n19687 = n2935 & ~n11961 ;
  assign n19688 = ~n3917 & n19687 ;
  assign n19689 = n19688 ^ n14830 ^ 1'b0 ;
  assign n19690 = n14467 ^ n12346 ^ n9264 ;
  assign n19691 = n18773 ^ n2024 ^ x99 ;
  assign n19692 = n17822 ^ n16542 ^ n9012 ;
  assign n19693 = n12893 ^ n6169 ^ n4597 ;
  assign n19694 = n13460 | n16377 ;
  assign n19695 = n19693 & ~n19694 ;
  assign n19696 = ( x145 & n16954 ) | ( x145 & ~n19695 ) | ( n16954 & ~n19695 ) ;
  assign n19703 = n3155 & ~n6028 ;
  assign n19704 = ~n5147 & n19703 ;
  assign n19702 = ~n7713 & n10056 ;
  assign n19705 = n19704 ^ n19702 ^ 1'b0 ;
  assign n19698 = n1037 | n14872 ;
  assign n19699 = n19698 ^ n1499 ^ 1'b0 ;
  assign n19700 = n12390 ^ n8759 ^ 1'b0 ;
  assign n19701 = n19699 | n19700 ;
  assign n19706 = n19705 ^ n19701 ^ n11649 ;
  assign n19697 = n15869 ^ n13489 ^ n12535 ;
  assign n19707 = n19706 ^ n19697 ^ n1295 ;
  assign n19708 = n10918 | n12558 ;
  assign n19709 = n6132 ^ n4769 ^ 1'b0 ;
  assign n19710 = n6921 ^ n4810 ^ 1'b0 ;
  assign n19711 = ~n539 & n19710 ;
  assign n19712 = n19711 ^ n4100 ^ n1431 ;
  assign n19713 = n19712 ^ n4867 ^ 1'b0 ;
  assign n19714 = ( n12267 & ~n19709 ) | ( n12267 & n19713 ) | ( ~n19709 & n19713 ) ;
  assign n19715 = n19684 ^ n9087 ^ n3601 ;
  assign n19716 = ( ~n7698 & n10779 ) | ( ~n7698 & n15169 ) | ( n10779 & n15169 ) ;
  assign n19717 = n8265 & n19716 ;
  assign n19718 = ~n19715 & n19717 ;
  assign n19719 = n1164 & n2042 ;
  assign n19720 = n19718 & n19719 ;
  assign n19721 = n6178 & ~n7286 ;
  assign n19722 = n19721 ^ n8294 ^ 1'b0 ;
  assign n19723 = n11675 ^ n9393 ^ x192 ;
  assign n19724 = n13104 ^ n9666 ^ 1'b0 ;
  assign n19725 = ~n12444 & n19724 ;
  assign n19726 = ( n1520 & ~n19723 ) | ( n1520 & n19725 ) | ( ~n19723 & n19725 ) ;
  assign n19727 = ~n8297 & n14849 ;
  assign n19729 = n8789 ^ n2866 ^ 1'b0 ;
  assign n19730 = n19729 ^ n2484 ^ 1'b0 ;
  assign n19728 = n18025 ^ n5782 ^ n1444 ;
  assign n19731 = n19730 ^ n19728 ^ 1'b0 ;
  assign n19732 = n3230 | n19731 ;
  assign n19733 = n19732 ^ n12007 ^ n10380 ;
  assign n19734 = ~n2705 & n19733 ;
  assign n19735 = n3381 & n19734 ;
  assign n19736 = n3832 ^ n3658 ^ n2523 ;
  assign n19737 = n19736 ^ n12777 ^ n11802 ;
  assign n19741 = n12830 & n15986 ;
  assign n19742 = n19741 ^ n4519 ^ 1'b0 ;
  assign n19738 = n16694 ^ x22 ^ 1'b0 ;
  assign n19739 = ~n4394 & n19738 ;
  assign n19740 = n19739 ^ n12599 ^ n5796 ;
  assign n19743 = n19742 ^ n19740 ^ n3748 ;
  assign n19744 = ~n19737 & n19743 ;
  assign n19746 = ( n2418 & n6348 ) | ( n2418 & ~n7504 ) | ( n6348 & ~n7504 ) ;
  assign n19745 = n12043 ^ n6783 ^ 1'b0 ;
  assign n19747 = n19746 ^ n19745 ^ n6616 ;
  assign n19748 = n15301 ^ n9822 ^ n7058 ;
  assign n19749 = n19748 ^ n19200 ^ n15542 ;
  assign n19750 = n626 | n1242 ;
  assign n19751 = n19750 ^ n5552 ^ 1'b0 ;
  assign n19752 = ( n1343 & ~n3478 ) | ( n1343 & n9953 ) | ( ~n3478 & n9953 ) ;
  assign n19753 = ( n19156 & n19751 ) | ( n19156 & ~n19752 ) | ( n19751 & ~n19752 ) ;
  assign n19754 = n14237 ^ n8845 ^ n7810 ;
  assign n19755 = ~n1979 & n19754 ;
  assign n19756 = n19755 ^ n6113 ^ 1'b0 ;
  assign n19757 = n8258 & n8276 ;
  assign n19758 = n5151 & n19757 ;
  assign n19761 = n3306 | n5066 ;
  assign n19762 = n19761 ^ n5566 ^ 1'b0 ;
  assign n19759 = n8113 ^ n6978 ^ 1'b0 ;
  assign n19760 = n4715 & ~n19759 ;
  assign n19763 = n19762 ^ n19760 ^ 1'b0 ;
  assign n19764 = ~n19758 & n19763 ;
  assign n19765 = n19764 ^ n14109 ^ 1'b0 ;
  assign n19766 = n9915 & n19765 ;
  assign n19767 = n19766 ^ n17489 ^ n2221 ;
  assign n19768 = n19756 | n19767 ;
  assign n19769 = n19768 ^ n13994 ^ 1'b0 ;
  assign n19770 = ~n2762 & n6528 ;
  assign n19771 = n19770 ^ n5604 ^ 1'b0 ;
  assign n19772 = n6912 & n19771 ;
  assign n19773 = n1626 | n19772 ;
  assign n19774 = n19439 ^ n9918 ^ 1'b0 ;
  assign n19775 = ( ~n17588 & n19773 ) | ( ~n17588 & n19774 ) | ( n19773 & n19774 ) ;
  assign n19779 = n15764 ^ n15370 ^ 1'b0 ;
  assign n19780 = n13057 | n19779 ;
  assign n19781 = n19780 ^ n8948 ^ 1'b0 ;
  assign n19782 = n19781 ^ n16564 ^ n11564 ;
  assign n19776 = n582 & ~n7785 ;
  assign n19777 = n13434 ^ n4323 ^ 1'b0 ;
  assign n19778 = n19776 & n19777 ;
  assign n19783 = n19782 ^ n19778 ^ n8264 ;
  assign n19784 = n18516 ^ n9642 ^ 1'b0 ;
  assign n19785 = ( n5830 & n5849 ) | ( n5830 & ~n9223 ) | ( n5849 & ~n9223 ) ;
  assign n19786 = ( ~n9473 & n12367 ) | ( ~n9473 & n19785 ) | ( n12367 & n19785 ) ;
  assign n19787 = ( ~n5195 & n5247 ) | ( ~n5195 & n17766 ) | ( n5247 & n17766 ) ;
  assign n19788 = n19013 ^ n17832 ^ 1'b0 ;
  assign n19789 = n19788 ^ n18922 ^ n4815 ;
  assign n19790 = n7613 ^ n5642 ^ n606 ;
  assign n19791 = n19790 ^ n6497 ^ 1'b0 ;
  assign n19792 = n14789 | n19791 ;
  assign n19793 = n6043 ^ n3351 ^ n696 ;
  assign n19794 = ~n7550 & n19793 ;
  assign n19795 = n19792 & n19794 ;
  assign n19796 = n19795 ^ n7420 ^ 1'b0 ;
  assign n19797 = n17514 & ~n19796 ;
  assign n19798 = n6587 | n8357 ;
  assign n19799 = n19798 ^ n6985 ^ 1'b0 ;
  assign n19800 = ( n7102 & n8842 ) | ( n7102 & ~n13079 ) | ( n8842 & ~n13079 ) ;
  assign n19801 = ( n4431 & ~n6971 ) | ( n4431 & n19800 ) | ( ~n6971 & n19800 ) ;
  assign n19808 = n10305 ^ n6529 ^ n1589 ;
  assign n19809 = n19808 ^ n3352 ^ 1'b0 ;
  assign n19810 = n4165 & ~n19809 ;
  assign n19811 = n19810 ^ n13531 ^ n607 ;
  assign n19805 = n2097 ^ n1638 ^ 1'b0 ;
  assign n19806 = ~n2771 & n19805 ;
  assign n19807 = n19806 ^ n2435 ^ 1'b0 ;
  assign n19802 = ( ~n7260 & n7865 ) | ( ~n7260 & n14862 ) | ( n7865 & n14862 ) ;
  assign n19803 = n19802 ^ n10404 ^ 1'b0 ;
  assign n19804 = n4957 | n19803 ;
  assign n19812 = n19811 ^ n19807 ^ n19804 ;
  assign n19813 = n2147 ^ n1247 ^ 1'b0 ;
  assign n19814 = ( ~n6821 & n6843 ) | ( ~n6821 & n19813 ) | ( n6843 & n19813 ) ;
  assign n19815 = ( n10955 & ~n16493 ) | ( n10955 & n19814 ) | ( ~n16493 & n19814 ) ;
  assign n19816 = n1503 & ~n19815 ;
  assign n19817 = n19816 ^ n18709 ^ 1'b0 ;
  assign n19820 = n7817 ^ n4852 ^ n1689 ;
  assign n19821 = ( n1421 & ~n12455 ) | ( n1421 & n19820 ) | ( ~n12455 & n19820 ) ;
  assign n19818 = n1198 & ~n11302 ;
  assign n19819 = n19818 ^ n8606 ^ 1'b0 ;
  assign n19822 = n19821 ^ n19819 ^ n6035 ;
  assign n19823 = n16927 & n19822 ;
  assign n19824 = ( n17120 & ~n19817 ) | ( n17120 & n19823 ) | ( ~n19817 & n19823 ) ;
  assign n19829 = n6494 | n8261 ;
  assign n19825 = n7426 ^ n1219 ^ 1'b0 ;
  assign n19826 = ~n5549 & n19825 ;
  assign n19827 = ( n1939 & ~n3764 ) | ( n1939 & n19826 ) | ( ~n3764 & n19826 ) ;
  assign n19828 = n19827 ^ n7178 ^ 1'b0 ;
  assign n19830 = n19829 ^ n19828 ^ n13452 ;
  assign n19831 = n11477 ^ x7 ^ 1'b0 ;
  assign n19832 = n6638 | n19831 ;
  assign n19833 = n10109 & ~n19832 ;
  assign n19834 = n19833 ^ n9586 ^ n8109 ;
  assign n19835 = n2722 ^ n1982 ^ n847 ;
  assign n19836 = ( n1804 & ~n2851 ) | ( n1804 & n19835 ) | ( ~n2851 & n19835 ) ;
  assign n19837 = ( n11444 & n19834 ) | ( n11444 & n19836 ) | ( n19834 & n19836 ) ;
  assign n19838 = n5316 ^ n2346 ^ 1'b0 ;
  assign n19839 = ( ~n3817 & n7279 ) | ( ~n3817 & n19838 ) | ( n7279 & n19838 ) ;
  assign n19840 = ( ~n1033 & n1384 ) | ( ~n1033 & n15621 ) | ( n1384 & n15621 ) ;
  assign n19841 = n19840 ^ n10139 ^ 1'b0 ;
  assign n19843 = ( ~n1962 & n3894 ) | ( ~n1962 & n5015 ) | ( n3894 & n5015 ) ;
  assign n19844 = n19843 ^ n6737 ^ n895 ;
  assign n19842 = ( ~n1155 & n5585 ) | ( ~n1155 & n6468 ) | ( n5585 & n6468 ) ;
  assign n19845 = n19844 ^ n19842 ^ 1'b0 ;
  assign n19846 = n7979 & n19845 ;
  assign n19847 = ( ~n7469 & n15774 ) | ( ~n7469 & n19846 ) | ( n15774 & n19846 ) ;
  assign n19848 = ( n6952 & ~n10384 ) | ( n6952 & n14030 ) | ( ~n10384 & n14030 ) ;
  assign n19849 = ( n3176 & n14291 ) | ( n3176 & ~n19848 ) | ( n14291 & ~n19848 ) ;
  assign n19850 = n15491 ^ n3631 ^ x65 ;
  assign n19851 = ( n5144 & ~n8155 ) | ( n5144 & n19850 ) | ( ~n8155 & n19850 ) ;
  assign n19857 = ~n1019 & n7957 ;
  assign n19858 = ~n4616 & n19857 ;
  assign n19852 = n10229 ^ n9057 ^ n6752 ;
  assign n19853 = n6500 ^ n3487 ^ n1330 ;
  assign n19854 = n16435 & ~n19853 ;
  assign n19855 = ( n418 & n12115 ) | ( n418 & ~n19854 ) | ( n12115 & ~n19854 ) ;
  assign n19856 = n19852 & ~n19855 ;
  assign n19859 = n19858 ^ n19856 ^ n10185 ;
  assign n19860 = ~n2899 & n19859 ;
  assign n19861 = n5309 ^ n3663 ^ n2020 ;
  assign n19862 = n5996 & n8154 ;
  assign n19863 = n19862 ^ n14930 ^ 1'b0 ;
  assign n19864 = ( ~x198 & n19861 ) | ( ~x198 & n19863 ) | ( n19861 & n19863 ) ;
  assign n19865 = ( n15583 & n17226 ) | ( n15583 & ~n18720 ) | ( n17226 & ~n18720 ) ;
  assign n19866 = ( n1147 & ~n7209 ) | ( n1147 & n17749 ) | ( ~n7209 & n17749 ) ;
  assign n19867 = ( n1220 & n10594 ) | ( n1220 & ~n19736 ) | ( n10594 & ~n19736 ) ;
  assign n19868 = n9279 & ~n13325 ;
  assign n19869 = n19868 ^ n8046 ^ 1'b0 ;
  assign n19870 = n19869 ^ n2837 ^ n351 ;
  assign n19871 = ~n9114 & n19870 ;
  assign n19872 = ~n10683 & n19871 ;
  assign n19873 = n6144 & ~n18768 ;
  assign n19874 = n19873 ^ n3052 ^ 1'b0 ;
  assign n19875 = n4518 ^ n2156 ^ x45 ;
  assign n19876 = ( n2283 & ~n3391 ) | ( n2283 & n19875 ) | ( ~n3391 & n19875 ) ;
  assign n19877 = n9892 & ~n9976 ;
  assign n19878 = n19877 ^ n880 ^ 1'b0 ;
  assign n19879 = n19878 ^ n6523 ^ n4166 ;
  assign n19880 = n19879 ^ n11942 ^ n10639 ;
  assign n19883 = n12436 ^ n7651 ^ 1'b0 ;
  assign n19881 = ~n6550 & n17564 ;
  assign n19882 = ~n19446 & n19881 ;
  assign n19884 = n19883 ^ n19882 ^ 1'b0 ;
  assign n19885 = ~n6226 & n6994 ;
  assign n19886 = n1712 & n19885 ;
  assign n19887 = ( ~n6724 & n19884 ) | ( ~n6724 & n19886 ) | ( n19884 & n19886 ) ;
  assign n19889 = n19352 ^ n5566 ^ n4349 ;
  assign n19888 = ( n6034 & n7830 ) | ( n6034 & ~n8454 ) | ( n7830 & ~n8454 ) ;
  assign n19890 = n19889 ^ n19888 ^ n2217 ;
  assign n19891 = ( n486 & n14941 ) | ( n486 & n19890 ) | ( n14941 & n19890 ) ;
  assign n19892 = n4330 & ~n9979 ;
  assign n19893 = n19892 ^ n9895 ^ 1'b0 ;
  assign n19894 = n19893 ^ n6171 ^ 1'b0 ;
  assign n19895 = ( n2729 & ~n19891 ) | ( n2729 & n19894 ) | ( ~n19891 & n19894 ) ;
  assign n19896 = ( n4721 & n5594 ) | ( n4721 & n11049 ) | ( n5594 & n11049 ) ;
  assign n19897 = ( ~n809 & n3222 ) | ( ~n809 & n6946 ) | ( n3222 & n6946 ) ;
  assign n19898 = ( ~n4205 & n19896 ) | ( ~n4205 & n19897 ) | ( n19896 & n19897 ) ;
  assign n19899 = ( x242 & n956 ) | ( x242 & n7309 ) | ( n956 & n7309 ) ;
  assign n19900 = ~n3619 & n19899 ;
  assign n19901 = ( ~n5430 & n11507 ) | ( ~n5430 & n15822 ) | ( n11507 & n15822 ) ;
  assign n19902 = n19901 ^ n7667 ^ n7244 ;
  assign n19903 = ( n9014 & n19086 ) | ( n9014 & n19902 ) | ( n19086 & n19902 ) ;
  assign n19904 = ( n8871 & n15571 ) | ( n8871 & n19903 ) | ( n15571 & n19903 ) ;
  assign n19905 = n19904 ^ n14334 ^ n11079 ;
  assign n19906 = n2144 & ~n8061 ;
  assign n19907 = n7784 ^ n6144 ^ 1'b0 ;
  assign n19908 = n4151 & n19907 ;
  assign n19909 = n19906 & n19908 ;
  assign n19910 = ( n2978 & ~n6250 ) | ( n2978 & n8037 ) | ( ~n6250 & n8037 ) ;
  assign n19911 = n5662 ^ n4777 ^ n3206 ;
  assign n19912 = n6540 | n19911 ;
  assign n19913 = n2665 & ~n12092 ;
  assign n19918 = ~n2415 & n3328 ;
  assign n19919 = ~n12746 & n19918 ;
  assign n19920 = ~n8135 & n19919 ;
  assign n19921 = n19920 ^ n12575 ^ n11432 ;
  assign n19922 = n19921 ^ n18975 ^ n7188 ;
  assign n19914 = n16047 ^ n6088 ^ 1'b0 ;
  assign n19915 = n18834 & n19914 ;
  assign n19916 = ( n12180 & n17420 ) | ( n12180 & n19915 ) | ( n17420 & n19915 ) ;
  assign n19917 = n19916 ^ n7168 ^ 1'b0 ;
  assign n19923 = n19922 ^ n19917 ^ n3323 ;
  assign n19924 = ~n6159 & n9494 ;
  assign n19925 = ~n12510 & n13100 ;
  assign n19926 = ~n11966 & n19925 ;
  assign n19927 = n1297 & n14908 ;
  assign n19928 = ~n779 & n19927 ;
  assign n19929 = ( n1940 & n2844 ) | ( n1940 & n5921 ) | ( n2844 & n5921 ) ;
  assign n19930 = n10530 ^ n7871 ^ 1'b0 ;
  assign n19931 = ( n11467 & n19929 ) | ( n11467 & ~n19930 ) | ( n19929 & ~n19930 ) ;
  assign n19936 = ( n438 & n598 ) | ( n438 & n10091 ) | ( n598 & n10091 ) ;
  assign n19937 = ( n4555 & ~n8082 ) | ( n4555 & n19936 ) | ( ~n8082 & n19936 ) ;
  assign n19938 = n19937 ^ n19071 ^ n13500 ;
  assign n19939 = n19938 ^ n16564 ^ n5511 ;
  assign n19933 = n455 | n828 ;
  assign n19934 = n14610 | n19933 ;
  assign n19932 = x98 & ~n3268 ;
  assign n19935 = n19934 ^ n19932 ^ 1'b0 ;
  assign n19940 = n19939 ^ n19935 ^ 1'b0 ;
  assign n19959 = n9047 ^ n7318 ^ 1'b0 ;
  assign n19960 = n11800 & n19959 ;
  assign n19961 = n1200 & n19960 ;
  assign n19953 = n2128 ^ n1323 ^ x141 ;
  assign n19952 = n4712 ^ n4492 ^ n3502 ;
  assign n19954 = n19953 ^ n19952 ^ 1'b0 ;
  assign n19955 = n5232 & n19954 ;
  assign n19956 = n15042 ^ n579 ^ 1'b0 ;
  assign n19957 = n19955 & ~n19956 ;
  assign n19958 = ~n11231 & n19957 ;
  assign n19962 = n19961 ^ n19958 ^ 1'b0 ;
  assign n19963 = n19962 ^ n10074 ^ 1'b0 ;
  assign n19964 = n16561 | n19963 ;
  assign n19941 = ( n5841 & n6963 ) | ( n5841 & n11907 ) | ( n6963 & n11907 ) ;
  assign n19942 = ~n3966 & n19941 ;
  assign n19943 = n19942 ^ n7361 ^ 1'b0 ;
  assign n19946 = n1220 & ~n10038 ;
  assign n19944 = n7699 ^ n4784 ^ n2566 ;
  assign n19945 = ( n9576 & n14195 ) | ( n9576 & ~n19944 ) | ( n14195 & ~n19944 ) ;
  assign n19947 = n19946 ^ n19945 ^ n7442 ;
  assign n19948 = n19947 ^ n19604 ^ 1'b0 ;
  assign n19949 = ~n3723 & n19948 ;
  assign n19950 = ( n3663 & n19943 ) | ( n3663 & ~n19949 ) | ( n19943 & ~n19949 ) ;
  assign n19951 = n2310 & n19950 ;
  assign n19965 = n19964 ^ n19951 ^ 1'b0 ;
  assign n19969 = n10336 ^ n7884 ^ n3832 ;
  assign n19970 = ( ~n1082 & n5089 ) | ( ~n1082 & n19969 ) | ( n5089 & n19969 ) ;
  assign n19966 = n2254 & ~n13455 ;
  assign n19967 = ~n8740 & n19966 ;
  assign n19968 = n6188 | n19967 ;
  assign n19971 = n19970 ^ n19968 ^ 1'b0 ;
  assign n19972 = n424 & n19971 ;
  assign n19973 = n19302 & n19972 ;
  assign n19974 = n12004 ^ n2964 ^ x183 ;
  assign n19975 = n2549 ^ n2100 ^ 1'b0 ;
  assign n19976 = n19957 & n19975 ;
  assign n19980 = n2689 & ~n7152 ;
  assign n19981 = n19980 ^ n7072 ^ 1'b0 ;
  assign n19977 = n12725 ^ n4232 ^ 1'b0 ;
  assign n19978 = n8552 | n19977 ;
  assign n19979 = ( ~n2877 & n6851 ) | ( ~n2877 & n19978 ) | ( n6851 & n19978 ) ;
  assign n19982 = n19981 ^ n19979 ^ 1'b0 ;
  assign n19983 = n553 ^ n522 ^ x101 ;
  assign n19984 = n13031 | n19983 ;
  assign n19985 = n4908 | n11435 ;
  assign n19986 = n19985 ^ n3245 ^ 1'b0 ;
  assign n19987 = ( ~n3794 & n6633 ) | ( ~n3794 & n19986 ) | ( n6633 & n19986 ) ;
  assign n19988 = n19984 & ~n19987 ;
  assign n19989 = n19988 ^ n18653 ^ 1'b0 ;
  assign n19990 = n16814 ^ x173 ^ 1'b0 ;
  assign n19991 = n17301 & ~n19990 ;
  assign n19992 = n6111 ^ n2132 ^ 1'b0 ;
  assign n19993 = ~n6259 & n19992 ;
  assign n19994 = n19993 ^ n15782 ^ 1'b0 ;
  assign n19995 = n13928 ^ n9477 ^ 1'b0 ;
  assign n19996 = n19995 ^ n5963 ^ n5714 ;
  assign n19997 = n11491 | n16637 ;
  assign n19998 = n19997 ^ n11639 ^ 1'b0 ;
  assign n19999 = ( ~x166 & n1116 ) | ( ~x166 & n8325 ) | ( n1116 & n8325 ) ;
  assign n20000 = n19999 ^ n18875 ^ 1'b0 ;
  assign n20001 = ~n19998 & n20000 ;
  assign n20002 = n19827 ^ n2475 ^ 1'b0 ;
  assign n20003 = ~n5884 & n8200 ;
  assign n20004 = n20003 ^ n19608 ^ 1'b0 ;
  assign n20005 = ( n9811 & n20002 ) | ( n9811 & n20004 ) | ( n20002 & n20004 ) ;
  assign n20006 = ( n3024 & ~n4667 ) | ( n3024 & n15284 ) | ( ~n4667 & n15284 ) ;
  assign n20007 = n5787 & ~n20006 ;
  assign n20008 = n7464 & n20007 ;
  assign n20012 = ( ~n391 & n2164 ) | ( ~n391 & n14175 ) | ( n2164 & n14175 ) ;
  assign n20013 = n20012 ^ n2913 ^ 1'b0 ;
  assign n20009 = ~n3315 & n11934 ;
  assign n20010 = n20009 ^ n19053 ^ 1'b0 ;
  assign n20011 = ~n11999 & n20010 ;
  assign n20014 = n20013 ^ n20011 ^ 1'b0 ;
  assign n20015 = ( n640 & n6788 ) | ( n640 & n16802 ) | ( n6788 & n16802 ) ;
  assign n20016 = n19879 ^ n4101 ^ n2610 ;
  assign n20017 = n20015 & ~n20016 ;
  assign n20018 = ~n20014 & n20017 ;
  assign n20019 = n710 & ~n2994 ;
  assign n20020 = n20019 ^ n18575 ^ 1'b0 ;
  assign n20021 = n669 & n18281 ;
  assign n20022 = n1691 & ~n9820 ;
  assign n20023 = n20022 ^ n6595 ^ 1'b0 ;
  assign n20024 = n4916 & ~n20023 ;
  assign n20025 = n4100 ^ n1876 ^ 1'b0 ;
  assign n20026 = n15157 & n16105 ;
  assign n20027 = ( n15376 & n20025 ) | ( n15376 & ~n20026 ) | ( n20025 & ~n20026 ) ;
  assign n20033 = n3641 ^ n2150 ^ n1394 ;
  assign n20032 = n13940 ^ n4232 ^ 1'b0 ;
  assign n20028 = n7327 | n10966 ;
  assign n20029 = n20028 ^ n14883 ^ 1'b0 ;
  assign n20030 = n20029 ^ n12886 ^ n9974 ;
  assign n20031 = n20030 ^ n8152 ^ n2699 ;
  assign n20034 = n20033 ^ n20032 ^ n20031 ;
  assign n20035 = n7943 ^ n1965 ^ n633 ;
  assign n20036 = n20035 ^ n15073 ^ 1'b0 ;
  assign n20037 = n20036 ^ n18284 ^ n12414 ;
  assign n20038 = ( ~n2186 & n2747 ) | ( ~n2186 & n10982 ) | ( n2747 & n10982 ) ;
  assign n20039 = n20038 ^ n3910 ^ n981 ;
  assign n20052 = n693 & n19893 ;
  assign n20057 = n1217 | n4147 ;
  assign n20058 = n1842 | n20057 ;
  assign n20053 = ~n7615 & n8037 ;
  assign n20054 = ~n8213 & n20053 ;
  assign n20055 = n6940 & ~n20054 ;
  assign n20056 = n13531 & n20055 ;
  assign n20059 = n20058 ^ n20056 ^ n10260 ;
  assign n20060 = ( n4896 & ~n20052 ) | ( n4896 & n20059 ) | ( ~n20052 & n20059 ) ;
  assign n20040 = n6417 | n8203 ;
  assign n20041 = ~n4874 & n20040 ;
  assign n20042 = n20041 ^ n5672 ^ 1'b0 ;
  assign n20043 = n20042 ^ n14465 ^ n2286 ;
  assign n20049 = ( n861 & ~n5578 ) | ( n861 & n15010 ) | ( ~n5578 & n15010 ) ;
  assign n20046 = n5122 & n17509 ;
  assign n20047 = n20046 ^ n9843 ^ 1'b0 ;
  assign n20048 = ( n5062 & n15412 ) | ( n5062 & ~n20047 ) | ( n15412 & ~n20047 ) ;
  assign n20044 = n8108 ^ n1408 ^ 1'b0 ;
  assign n20045 = n20044 ^ n13020 ^ n8447 ;
  assign n20050 = n20049 ^ n20048 ^ n20045 ;
  assign n20051 = n20043 | n20050 ;
  assign n20061 = n20060 ^ n20051 ^ 1'b0 ;
  assign n20062 = n3514 ^ n2430 ^ n431 ;
  assign n20063 = n10001 & n13324 ;
  assign n20064 = ~n1326 & n20063 ;
  assign n20065 = ( ~n10359 & n20062 ) | ( ~n10359 & n20064 ) | ( n20062 & n20064 ) ;
  assign n20068 = n3803 | n11304 ;
  assign n20069 = n340 | n20068 ;
  assign n20066 = ~n5485 & n19355 ;
  assign n20067 = ~n10702 & n20066 ;
  assign n20070 = n20069 ^ n20067 ^ n3569 ;
  assign n20071 = n4225 ^ n2224 ^ n296 ;
  assign n20072 = ( n2319 & n12346 ) | ( n2319 & ~n20071 ) | ( n12346 & ~n20071 ) ;
  assign n20073 = ( n3158 & n8137 ) | ( n3158 & n18194 ) | ( n8137 & n18194 ) ;
  assign n20074 = ( ~n2745 & n6336 ) | ( ~n2745 & n6705 ) | ( n6336 & n6705 ) ;
  assign n20075 = n20074 ^ n10466 ^ n1897 ;
  assign n20076 = ( x236 & n2189 ) | ( x236 & n9635 ) | ( n2189 & n9635 ) ;
  assign n20077 = ( n1025 & n5915 ) | ( n1025 & n9614 ) | ( n5915 & n9614 ) ;
  assign n20078 = n808 & n20077 ;
  assign n20079 = n20076 & n20078 ;
  assign n20080 = n5401 ^ n1365 ^ 1'b0 ;
  assign n20081 = n7148 | n20080 ;
  assign n20082 = n20081 ^ n19364 ^ 1'b0 ;
  assign n20083 = ( ~n20075 & n20079 ) | ( ~n20075 & n20082 ) | ( n20079 & n20082 ) ;
  assign n20084 = n925 & n17265 ;
  assign n20085 = n20083 & n20084 ;
  assign n20086 = n8881 & n11244 ;
  assign n20087 = n18767 ^ n13141 ^ 1'b0 ;
  assign n20088 = n20086 | n20087 ;
  assign n20089 = n15619 ^ n14211 ^ 1'b0 ;
  assign n20090 = ( ~n348 & n3281 ) | ( ~n348 & n4590 ) | ( n3281 & n4590 ) ;
  assign n20091 = n20090 ^ n17154 ^ n6654 ;
  assign n20092 = n1002 & ~n20091 ;
  assign n20093 = n10490 & n20092 ;
  assign n20094 = n2317 ^ n2288 ^ 1'b0 ;
  assign n20095 = n20094 ^ n17166 ^ 1'b0 ;
  assign n20096 = n3226 & ~n20095 ;
  assign n20097 = n20096 ^ n5778 ^ 1'b0 ;
  assign n20098 = n20097 ^ n4921 ^ 1'b0 ;
  assign n20099 = n3568 ^ n2914 ^ n984 ;
  assign n20100 = ( ~n8369 & n16684 ) | ( ~n8369 & n20099 ) | ( n16684 & n20099 ) ;
  assign n20106 = n16111 ^ n3163 ^ 1'b0 ;
  assign n20104 = n1809 ^ n1490 ^ 1'b0 ;
  assign n20102 = ( n2773 & ~n4339 ) | ( n2773 & n8158 ) | ( ~n4339 & n8158 ) ;
  assign n20103 = n20102 ^ n3082 ^ 1'b0 ;
  assign n20101 = ( ~x86 & n7682 ) | ( ~x86 & n14017 ) | ( n7682 & n14017 ) ;
  assign n20105 = n20104 ^ n20103 ^ n20101 ;
  assign n20107 = n20106 ^ n20105 ^ n10612 ;
  assign n20111 = n4314 & ~n5258 ;
  assign n20112 = n20111 ^ n17166 ^ 1'b0 ;
  assign n20113 = n20112 ^ n14742 ^ n4299 ;
  assign n20114 = n7843 & n14250 ;
  assign n20115 = ~n20113 & n20114 ;
  assign n20116 = n8097 & n20115 ;
  assign n20108 = ~n4547 & n17265 ;
  assign n20109 = n20108 ^ n10267 ^ 1'b0 ;
  assign n20110 = n16751 & ~n20109 ;
  assign n20117 = n20116 ^ n20110 ^ 1'b0 ;
  assign n20118 = ~n5017 & n8170 ;
  assign n20119 = n6377 ^ n1791 ^ 1'b0 ;
  assign n20120 = n20119 ^ n13641 ^ n13583 ;
  assign n20121 = n3097 & n20120 ;
  assign n20122 = n10737 & n15546 ;
  assign n20123 = n20122 ^ n3517 ^ 1'b0 ;
  assign n20124 = ~n11522 & n20123 ;
  assign n20125 = n20124 ^ n19349 ^ n257 ;
  assign n20126 = n3074 ^ n2168 ^ n1313 ;
  assign n20127 = ( n12325 & n12813 ) | ( n12325 & n20126 ) | ( n12813 & n20126 ) ;
  assign n20128 = n20127 ^ n20040 ^ n16010 ;
  assign n20129 = n12418 | n20128 ;
  assign n20130 = n5694 ^ n3309 ^ n2583 ;
  assign n20131 = ( n2987 & n8567 ) | ( n2987 & ~n15071 ) | ( n8567 & ~n15071 ) ;
  assign n20132 = ~n7207 & n20131 ;
  assign n20133 = ( ~n3219 & n20130 ) | ( ~n3219 & n20132 ) | ( n20130 & n20132 ) ;
  assign n20134 = n10111 & ~n19236 ;
  assign n20135 = n20134 ^ n14871 ^ 1'b0 ;
  assign n20136 = ( n7799 & ~n11147 ) | ( n7799 & n19644 ) | ( ~n11147 & n19644 ) ;
  assign n20137 = n971 & ~n18958 ;
  assign n20138 = ( ~n2491 & n6268 ) | ( ~n2491 & n6622 ) | ( n6268 & n6622 ) ;
  assign n20139 = n2614 & n20138 ;
  assign n20140 = ~n4627 & n20139 ;
  assign n20141 = ( x212 & n16441 ) | ( x212 & ~n20140 ) | ( n16441 & ~n20140 ) ;
  assign n20142 = ~n4547 & n5093 ;
  assign n20143 = n8087 & n16511 ;
  assign n20144 = ~n979 & n2179 ;
  assign n20145 = n20144 ^ n2052 ^ 1'b0 ;
  assign n20146 = n20145 ^ n13556 ^ n7870 ;
  assign n20147 = x57 & ~n2555 ;
  assign n20148 = n20147 ^ n3707 ^ 1'b0 ;
  assign n20149 = ~n6205 & n20148 ;
  assign n20150 = n13234 & n20149 ;
  assign n20151 = ( n5481 & ~n13944 ) | ( n5481 & n20150 ) | ( ~n13944 & n20150 ) ;
  assign n20153 = n8498 & n9716 ;
  assign n20154 = n4452 & n20153 ;
  assign n20152 = n19216 ^ n13932 ^ n9728 ;
  assign n20155 = n20154 ^ n20152 ^ 1'b0 ;
  assign n20157 = ~n5300 & n12708 ;
  assign n20158 = n20157 ^ n15778 ^ n9787 ;
  assign n20159 = n10486 ^ n3052 ^ 1'b0 ;
  assign n20160 = n20158 & ~n20159 ;
  assign n20156 = ( n628 & n5448 ) | ( n628 & n17092 ) | ( n5448 & n17092 ) ;
  assign n20161 = n20160 ^ n20156 ^ 1'b0 ;
  assign n20164 = n8342 ^ n3263 ^ n2608 ;
  assign n20162 = ( n1139 & ~n3633 ) | ( n1139 & n3803 ) | ( ~n3633 & n3803 ) ;
  assign n20163 = ( n3601 & n7600 ) | ( n3601 & ~n20162 ) | ( n7600 & ~n20162 ) ;
  assign n20165 = n20164 ^ n20163 ^ n8480 ;
  assign n20166 = ( n3358 & ~n11962 ) | ( n3358 & n20165 ) | ( ~n11962 & n20165 ) ;
  assign n20167 = n18822 & ~n19473 ;
  assign n20168 = ( n2162 & n6759 ) | ( n2162 & n20167 ) | ( n6759 & n20167 ) ;
  assign n20175 = ( n4097 & ~n8171 ) | ( n4097 & n17773 ) | ( ~n8171 & n17773 ) ;
  assign n20172 = n1387 & ~n7136 ;
  assign n20173 = ~n9358 & n20172 ;
  assign n20169 = ( ~n1452 & n4130 ) | ( ~n1452 & n12606 ) | ( n4130 & n12606 ) ;
  assign n20170 = n3208 | n20169 ;
  assign n20171 = ( n8254 & n12863 ) | ( n8254 & ~n20170 ) | ( n12863 & ~n20170 ) ;
  assign n20174 = n20173 ^ n20171 ^ n781 ;
  assign n20176 = n20175 ^ n20174 ^ 1'b0 ;
  assign n20178 = n6310 & n9896 ;
  assign n20177 = n6230 & n7837 ;
  assign n20179 = n20178 ^ n20177 ^ 1'b0 ;
  assign n20180 = n6143 ^ n1212 ^ 1'b0 ;
  assign n20181 = n20180 ^ n10202 ^ n3613 ;
  assign n20182 = n20181 ^ n10443 ^ 1'b0 ;
  assign n20183 = ( n4570 & n16907 ) | ( n4570 & ~n19452 ) | ( n16907 & ~n19452 ) ;
  assign n20184 = n2989 | n20183 ;
  assign n20185 = ( n1991 & n8847 ) | ( n1991 & n20184 ) | ( n8847 & n20184 ) ;
  assign n20186 = n5028 & ~n9130 ;
  assign n20187 = n20186 ^ n5015 ^ 1'b0 ;
  assign n20188 = n1413 & ~n7116 ;
  assign n20189 = n20188 ^ n2941 ^ 1'b0 ;
  assign n20191 = n9109 ^ n278 ^ 1'b0 ;
  assign n20192 = n4444 & ~n20191 ;
  assign n20190 = ( ~n2442 & n4351 ) | ( ~n2442 & n7123 ) | ( n4351 & n7123 ) ;
  assign n20193 = n20192 ^ n20190 ^ n2258 ;
  assign n20194 = ( n20187 & n20189 ) | ( n20187 & n20193 ) | ( n20189 & n20193 ) ;
  assign n20195 = n6029 | n12479 ;
  assign n20196 = n20195 ^ n16714 ^ 1'b0 ;
  assign n20197 = n7227 & ~n17983 ;
  assign n20198 = n13929 ^ n2852 ^ 1'b0 ;
  assign n20199 = n11543 | n13531 ;
  assign n20200 = n20198 | n20199 ;
  assign n20201 = n12358 ^ n6992 ^ 1'b0 ;
  assign n20202 = n20200 & n20201 ;
  assign n20203 = n20202 ^ n16598 ^ n11455 ;
  assign n20204 = ( n4192 & ~n15669 ) | ( n4192 & n16423 ) | ( ~n15669 & n16423 ) ;
  assign n20211 = n6533 ^ n1983 ^ 1'b0 ;
  assign n20212 = n19047 & ~n20211 ;
  assign n20205 = ( n2098 & n4381 ) | ( n2098 & ~n9979 ) | ( n4381 & ~n9979 ) ;
  assign n20206 = n1554 & n4668 ;
  assign n20207 = ( ~n1087 & n13127 ) | ( ~n1087 & n20206 ) | ( n13127 & n20206 ) ;
  assign n20208 = ( n476 & ~n20205 ) | ( n476 & n20207 ) | ( ~n20205 & n20207 ) ;
  assign n20209 = ( ~n6710 & n14783 ) | ( ~n6710 & n20208 ) | ( n14783 & n20208 ) ;
  assign n20210 = ~n16637 & n20209 ;
  assign n20213 = n20212 ^ n20210 ^ 1'b0 ;
  assign n20216 = n11149 ^ n5481 ^ 1'b0 ;
  assign n20214 = n17075 ^ n5256 ^ 1'b0 ;
  assign n20215 = n13266 | n20214 ;
  assign n20217 = n20216 ^ n20215 ^ n5392 ;
  assign n20218 = n793 & ~n16697 ;
  assign n20219 = ( n5857 & ~n11584 ) | ( n5857 & n20218 ) | ( ~n11584 & n20218 ) ;
  assign n20220 = x15 & ~n1398 ;
  assign n20221 = ~x93 & n20220 ;
  assign n20222 = ( n5974 & ~n11397 ) | ( n5974 & n20221 ) | ( ~n11397 & n20221 ) ;
  assign n20223 = ( ~n3106 & n12054 ) | ( ~n3106 & n20222 ) | ( n12054 & n20222 ) ;
  assign n20224 = ( n14153 & n17762 ) | ( n14153 & n20223 ) | ( n17762 & n20223 ) ;
  assign n20225 = ~n1125 & n12255 ;
  assign n20226 = n12419 ^ n4842 ^ 1'b0 ;
  assign n20227 = n13531 ^ n931 ^ 1'b0 ;
  assign n20228 = n8269 & ~n20227 ;
  assign n20229 = n20228 ^ n13923 ^ 1'b0 ;
  assign n20230 = ( n5904 & n20226 ) | ( n5904 & n20229 ) | ( n20226 & n20229 ) ;
  assign n20234 = n4358 | n16385 ;
  assign n20232 = ( n8810 & n12560 ) | ( n8810 & n14527 ) | ( n12560 & n14527 ) ;
  assign n20233 = ( ~n8352 & n18660 ) | ( ~n8352 & n20232 ) | ( n18660 & n20232 ) ;
  assign n20231 = n3734 | n6006 ;
  assign n20235 = n20234 ^ n20233 ^ n20231 ;
  assign n20236 = n13798 ^ n2235 ^ 1'b0 ;
  assign n20237 = n13405 ^ n3869 ^ n3554 ;
  assign n20238 = n1122 & ~n20237 ;
  assign n20239 = n20238 ^ x77 ^ 1'b0 ;
  assign n20240 = ( n2905 & n20236 ) | ( n2905 & ~n20239 ) | ( n20236 & ~n20239 ) ;
  assign n20241 = n8864 ^ n375 ^ 1'b0 ;
  assign n20243 = n10722 & n11008 ;
  assign n20244 = n20243 ^ n12857 ^ 1'b0 ;
  assign n20245 = n10430 ^ x75 ^ 1'b0 ;
  assign n20246 = n20244 | n20245 ;
  assign n20242 = n525 & ~n4493 ;
  assign n20247 = n20246 ^ n20242 ^ 1'b0 ;
  assign n20248 = ~n8397 & n10335 ;
  assign n20249 = n5978 & n20248 ;
  assign n20250 = n20249 ^ n19474 ^ n5442 ;
  assign n20251 = n4592 & n12763 ;
  assign n20252 = ~n8875 & n20251 ;
  assign n20259 = n3244 | n3588 ;
  assign n20260 = n20259 ^ n6978 ^ 1'b0 ;
  assign n20261 = n8607 & ~n20260 ;
  assign n20262 = ( n6583 & n7661 ) | ( n6583 & n20261 ) | ( n7661 & n20261 ) ;
  assign n20253 = n13756 ^ n797 ^ 1'b0 ;
  assign n20254 = n3853 & ~n20253 ;
  assign n20255 = n8180 ^ n5067 ^ n3280 ;
  assign n20256 = n20255 ^ n13700 ^ n3130 ;
  assign n20257 = ( n5531 & n20254 ) | ( n5531 & ~n20256 ) | ( n20254 & ~n20256 ) ;
  assign n20258 = ~n2985 & n20257 ;
  assign n20263 = n20262 ^ n20258 ^ 1'b0 ;
  assign n20264 = n4922 | n16865 ;
  assign n20265 = n1079 | n4273 ;
  assign n20266 = n20265 ^ n10733 ^ 1'b0 ;
  assign n20267 = n9999 & ~n13746 ;
  assign n20268 = ~n8887 & n20267 ;
  assign n20269 = n7112 ^ n4640 ^ n4570 ;
  assign n20270 = ~n2881 & n3219 ;
  assign n20271 = n20270 ^ n19508 ^ 1'b0 ;
  assign n20272 = n20271 ^ n12170 ^ 1'b0 ;
  assign n20273 = n7720 & n20272 ;
  assign n20274 = ( n8770 & n20269 ) | ( n8770 & ~n20273 ) | ( n20269 & ~n20273 ) ;
  assign n20275 = ( n20266 & n20268 ) | ( n20266 & ~n20274 ) | ( n20268 & ~n20274 ) ;
  assign n20276 = n3310 & n3472 ;
  assign n20277 = ( n4067 & n12099 ) | ( n4067 & ~n20276 ) | ( n12099 & ~n20276 ) ;
  assign n20278 = n20277 ^ n12977 ^ n12458 ;
  assign n20279 = ( x9 & n4935 ) | ( x9 & n12034 ) | ( n4935 & n12034 ) ;
  assign n20280 = ( ~n5799 & n8528 ) | ( ~n5799 & n20279 ) | ( n8528 & n20279 ) ;
  assign n20281 = ~n2668 & n13759 ;
  assign n20282 = n20281 ^ n1240 ^ 1'b0 ;
  assign n20284 = n1591 | n7889 ;
  assign n20285 = n480 | n20284 ;
  assign n20283 = ( ~n1481 & n1590 ) | ( ~n1481 & n7047 ) | ( n1590 & n7047 ) ;
  assign n20286 = n20285 ^ n20283 ^ n487 ;
  assign n20287 = n20286 ^ n17710 ^ 1'b0 ;
  assign n20288 = n11658 ^ n8391 ^ n323 ;
  assign n20289 = n10647 & ~n13573 ;
  assign n20290 = n20289 ^ n3672 ^ 1'b0 ;
  assign n20291 = n20290 ^ n6268 ^ x245 ;
  assign n20293 = n11520 ^ n570 ^ 1'b0 ;
  assign n20292 = ( n3564 & n6345 ) | ( n3564 & ~n8405 ) | ( n6345 & ~n8405 ) ;
  assign n20294 = n20293 ^ n20292 ^ n3101 ;
  assign n20295 = n5633 | n20294 ;
  assign n20296 = n20295 ^ n19570 ^ 1'b0 ;
  assign n20297 = ( n20288 & n20291 ) | ( n20288 & ~n20296 ) | ( n20291 & ~n20296 ) ;
  assign n20298 = ( n3752 & ~n9805 ) | ( n3752 & n15899 ) | ( ~n9805 & n15899 ) ;
  assign n20299 = ( n1093 & ~n8067 ) | ( n1093 & n20298 ) | ( ~n8067 & n20298 ) ;
  assign n20300 = ( n4334 & n5009 ) | ( n4334 & n8067 ) | ( n5009 & n8067 ) ;
  assign n20301 = n20300 ^ n6937 ^ n6336 ;
  assign n20302 = ( n3441 & n7664 ) | ( n3441 & ~n11692 ) | ( n7664 & ~n11692 ) ;
  assign n20303 = n15313 ^ n11992 ^ n7884 ;
  assign n20307 = ( ~n6267 & n6716 ) | ( ~n6267 & n9992 ) | ( n6716 & n9992 ) ;
  assign n20308 = n20307 ^ n10448 ^ n9927 ;
  assign n20309 = ( x33 & n7322 ) | ( x33 & n11706 ) | ( n7322 & n11706 ) ;
  assign n20310 = ( ~n14277 & n20308 ) | ( ~n14277 & n20309 ) | ( n20308 & n20309 ) ;
  assign n20304 = n16385 ^ n8499 ^ 1'b0 ;
  assign n20305 = n8174 & ~n20304 ;
  assign n20306 = n20305 ^ n4671 ^ 1'b0 ;
  assign n20311 = n20310 ^ n20306 ^ 1'b0 ;
  assign n20312 = n3961 ^ n3415 ^ 1'b0 ;
  assign n20313 = ( ~n2520 & n4890 ) | ( ~n2520 & n20312 ) | ( n4890 & n20312 ) ;
  assign n20314 = ~n2066 & n17624 ;
  assign n20315 = ( ~n489 & n4112 ) | ( ~n489 & n20314 ) | ( n4112 & n20314 ) ;
  assign n20316 = n13098 ^ n1851 ^ n829 ;
  assign n20324 = n16371 ^ n4022 ^ n534 ;
  assign n20317 = n11772 ^ n9582 ^ n6379 ;
  assign n20320 = n18530 ^ n7102 ^ n7029 ;
  assign n20318 = x115 & ~n9047 ;
  assign n20319 = ~n6158 & n20318 ;
  assign n20321 = n20320 ^ n20319 ^ 1'b0 ;
  assign n20322 = ( ~n1844 & n20317 ) | ( ~n1844 & n20321 ) | ( n20317 & n20321 ) ;
  assign n20323 = n2822 | n20322 ;
  assign n20325 = n20324 ^ n20323 ^ 1'b0 ;
  assign n20326 = n20325 ^ n8480 ^ n1154 ;
  assign n20330 = n10963 ^ n4170 ^ 1'b0 ;
  assign n20331 = n20330 ^ n10154 ^ 1'b0 ;
  assign n20332 = n20331 ^ n14544 ^ 1'b0 ;
  assign n20333 = n5546 | n20332 ;
  assign n20327 = ( n2988 & n10448 ) | ( n2988 & ~n13170 ) | ( n10448 & ~n13170 ) ;
  assign n20328 = ( n1251 & n3043 ) | ( n1251 & n20327 ) | ( n3043 & n20327 ) ;
  assign n20329 = n20328 ^ n18427 ^ n16846 ;
  assign n20334 = n20333 ^ n20329 ^ n14765 ;
  assign n20335 = n14524 & n20334 ;
  assign n20336 = ( n6026 & n6491 ) | ( n6026 & ~n14712 ) | ( n6491 & ~n14712 ) ;
  assign n20337 = ( n1720 & n14533 ) | ( n1720 & ~n20336 ) | ( n14533 & ~n20336 ) ;
  assign n20338 = ( n548 & n5572 ) | ( n548 & ~n11140 ) | ( n5572 & ~n11140 ) ;
  assign n20339 = ( n3593 & ~n3975 ) | ( n3593 & n9810 ) | ( ~n3975 & n9810 ) ;
  assign n20340 = ( n2075 & n3657 ) | ( n2075 & n20339 ) | ( n3657 & n20339 ) ;
  assign n20341 = n20340 ^ n18949 ^ 1'b0 ;
  assign n20342 = ( n2819 & n20338 ) | ( n2819 & ~n20341 ) | ( n20338 & ~n20341 ) ;
  assign n20343 = n20342 ^ n16058 ^ n12277 ;
  assign n20344 = ( ~n4520 & n20337 ) | ( ~n4520 & n20343 ) | ( n20337 & n20343 ) ;
  assign n20345 = n12907 ^ n9796 ^ n9737 ;
  assign n20346 = n20345 ^ n6882 ^ n987 ;
  assign n20347 = n461 & ~n12507 ;
  assign n20348 = n6139 & n20347 ;
  assign n20349 = n12023 & ~n20348 ;
  assign n20350 = n1009 & n20349 ;
  assign n20351 = n8267 ^ n6560 ^ n2955 ;
  assign n20352 = n4997 | n10734 ;
  assign n20353 = n20352 ^ n19889 ^ 1'b0 ;
  assign n20354 = n3997 | n7643 ;
  assign n20355 = ( n3541 & ~n18847 ) | ( n3541 & n20354 ) | ( ~n18847 & n20354 ) ;
  assign n20356 = n20355 ^ n16036 ^ 1'b0 ;
  assign n20357 = n6745 ^ n3462 ^ 1'b0 ;
  assign n20358 = n3239 & n20357 ;
  assign n20359 = n3740 & ~n20358 ;
  assign n20360 = n4593 & ~n20359 ;
  assign n20361 = n20360 ^ n4603 ^ 1'b0 ;
  assign n20362 = n20356 | n20361 ;
  assign n20363 = ( n20351 & ~n20353 ) | ( n20351 & n20362 ) | ( ~n20353 & n20362 ) ;
  assign n20364 = n1169 & n17893 ;
  assign n20365 = n20364 ^ n7859 ^ 1'b0 ;
  assign n20366 = n20365 ^ n13560 ^ n333 ;
  assign n20367 = n5071 & ~n19156 ;
  assign n20368 = n20367 ^ n11961 ^ 1'b0 ;
  assign n20369 = ( n1048 & n9773 ) | ( n1048 & ~n20368 ) | ( n9773 & ~n20368 ) ;
  assign n20370 = ( n7757 & ~n11063 ) | ( n7757 & n16771 ) | ( ~n11063 & n16771 ) ;
  assign n20371 = ( n8316 & n20369 ) | ( n8316 & ~n20370 ) | ( n20369 & ~n20370 ) ;
  assign n20372 = n20371 ^ n11878 ^ 1'b0 ;
  assign n20380 = ( n4525 & n7171 ) | ( n4525 & ~n15965 ) | ( n7171 & ~n15965 ) ;
  assign n20378 = n13459 ^ n2139 ^ 1'b0 ;
  assign n20376 = n9078 | n13691 ;
  assign n20377 = n20376 ^ n1845 ^ 1'b0 ;
  assign n20379 = n20378 ^ n20377 ^ n13190 ;
  assign n20373 = ( ~n8064 & n14934 ) | ( ~n8064 & n15622 ) | ( n14934 & n15622 ) ;
  assign n20374 = n18452 ^ n12315 ^ 1'b0 ;
  assign n20375 = n20373 & n20374 ;
  assign n20381 = n20380 ^ n20379 ^ n20375 ;
  assign n20382 = n12208 ^ n8802 ^ n1791 ;
  assign n20383 = n919 | n11238 ;
  assign n20384 = n9709 | n20383 ;
  assign n20385 = n20384 ^ n9169 ^ n1465 ;
  assign n20386 = n18337 ^ n12039 ^ 1'b0 ;
  assign n20387 = n20385 & n20386 ;
  assign n20388 = ( n4448 & ~n11426 ) | ( n4448 & n12883 ) | ( ~n11426 & n12883 ) ;
  assign n20392 = ( ~n789 & n4558 ) | ( ~n789 & n9245 ) | ( n4558 & n9245 ) ;
  assign n20389 = n14270 & n17169 ;
  assign n20390 = n20389 ^ n7310 ^ n5856 ;
  assign n20391 = n20390 ^ n6255 ^ 1'b0 ;
  assign n20393 = n20392 ^ n20391 ^ 1'b0 ;
  assign n20394 = n20393 ^ n14157 ^ n14123 ;
  assign n20400 = n12906 ^ n3493 ^ n571 ;
  assign n20395 = n14334 ^ n1565 ^ 1'b0 ;
  assign n20396 = n8512 ^ n5402 ^ n4219 ;
  assign n20397 = n20396 ^ n8267 ^ 1'b0 ;
  assign n20398 = n20395 & n20397 ;
  assign n20399 = n20398 ^ n11356 ^ 1'b0 ;
  assign n20401 = n20400 ^ n20399 ^ n6975 ;
  assign n20402 = ( ~n5811 & n11427 ) | ( ~n5811 & n20385 ) | ( n11427 & n20385 ) ;
  assign n20403 = ( n4110 & n4902 ) | ( n4110 & n11065 ) | ( n4902 & n11065 ) ;
  assign n20414 = ( ~n2392 & n8115 ) | ( ~n2392 & n14825 ) | ( n8115 & n14825 ) ;
  assign n20415 = ( ~n8806 & n13497 ) | ( ~n8806 & n20414 ) | ( n13497 & n20414 ) ;
  assign n20413 = n868 & n11191 ;
  assign n20416 = n20415 ^ n20413 ^ 1'b0 ;
  assign n20404 = n8718 ^ n849 ^ 1'b0 ;
  assign n20405 = n4631 & ~n20404 ;
  assign n20406 = n4590 | n11241 ;
  assign n20407 = n2724 | n20406 ;
  assign n20408 = n20407 ^ n11609 ^ n1106 ;
  assign n20409 = ( n11781 & n20395 ) | ( n11781 & n20408 ) | ( n20395 & n20408 ) ;
  assign n20410 = n20409 ^ n633 ^ 1'b0 ;
  assign n20411 = n20405 & ~n20410 ;
  assign n20412 = n20411 ^ n19335 ^ n14192 ;
  assign n20417 = n20416 ^ n20412 ^ 1'b0 ;
  assign n20418 = n9420 & ~n20417 ;
  assign n20419 = n20403 & n20418 ;
  assign n20420 = n11826 & n20419 ;
  assign n20423 = ( x191 & n7944 ) | ( x191 & n19941 ) | ( n7944 & n19941 ) ;
  assign n20422 = n10356 & n14181 ;
  assign n20421 = n7739 ^ n4599 ^ n1814 ;
  assign n20424 = n20423 ^ n20422 ^ n20421 ;
  assign n20425 = n20033 ^ n11971 ^ n8774 ;
  assign n20426 = n12238 ^ n1827 ^ 1'b0 ;
  assign n20427 = n270 | n20426 ;
  assign n20428 = n14825 ^ n12013 ^ 1'b0 ;
  assign n20429 = ( n20425 & ~n20427 ) | ( n20425 & n20428 ) | ( ~n20427 & n20428 ) ;
  assign n20430 = ( ~n5656 & n9722 ) | ( ~n5656 & n15186 ) | ( n9722 & n15186 ) ;
  assign n20431 = n8760 ^ n1463 ^ 1'b0 ;
  assign n20432 = n6694 ^ n5138 ^ 1'b0 ;
  assign n20433 = n20432 ^ n6927 ^ n1179 ;
  assign n20434 = n20433 ^ n8337 ^ n4307 ;
  assign n20435 = ( ~n3806 & n6300 ) | ( ~n3806 & n20434 ) | ( n6300 & n20434 ) ;
  assign n20436 = n8866 ^ n1226 ^ 1'b0 ;
  assign n20437 = ( x3 & ~n5481 ) | ( x3 & n14202 ) | ( ~n5481 & n14202 ) ;
  assign n20438 = n6827 ^ n2660 ^ 1'b0 ;
  assign n20439 = ( n5083 & n15227 ) | ( n5083 & n20438 ) | ( n15227 & n20438 ) ;
  assign n20440 = n20266 & n20439 ;
  assign n20441 = n20440 ^ n2509 ^ 1'b0 ;
  assign n20442 = n20441 ^ n13012 ^ 1'b0 ;
  assign n20443 = n16414 | n20442 ;
  assign n20444 = n20443 ^ n1486 ^ 1'b0 ;
  assign n20445 = n20444 ^ n3859 ^ 1'b0 ;
  assign n20446 = n10174 & ~n20445 ;
  assign n20447 = n8080 & n20446 ;
  assign n20448 = ~n20437 & n20447 ;
  assign n20449 = n2960 & ~n20448 ;
  assign n20450 = ( n12019 & n20436 ) | ( n12019 & n20449 ) | ( n20436 & n20449 ) ;
  assign n20451 = ( ~n19806 & n20435 ) | ( ~n19806 & n20450 ) | ( n20435 & n20450 ) ;
  assign n20452 = n8688 ^ n7717 ^ 1'b0 ;
  assign n20453 = n20451 | n20452 ;
  assign n20454 = n18065 ^ n17378 ^ n16398 ;
  assign n20455 = ( ~n11712 & n19281 ) | ( ~n11712 & n20454 ) | ( n19281 & n20454 ) ;
  assign n20456 = ~n3483 & n20328 ;
  assign n20457 = ~n18201 & n20456 ;
  assign n20458 = ( n921 & n5248 ) | ( n921 & n16748 ) | ( n5248 & n16748 ) ;
  assign n20459 = n20458 ^ n1944 ^ 1'b0 ;
  assign n20460 = n5169 | n20459 ;
  assign n20461 = n6632 | n16565 ;
  assign n20462 = n13070 & ~n20461 ;
  assign n20463 = ( n4215 & n12176 ) | ( n4215 & n20462 ) | ( n12176 & n20462 ) ;
  assign n20464 = ~n18736 & n20463 ;
  assign n20465 = n6430 & ~n19686 ;
  assign n20466 = n12678 ^ n6330 ^ n2461 ;
  assign n20467 = n8838 ^ n8311 ^ 1'b0 ;
  assign n20468 = ( n11998 & ~n20466 ) | ( n11998 & n20467 ) | ( ~n20466 & n20467 ) ;
  assign n20469 = ( n1520 & ~n4930 ) | ( n1520 & n10552 ) | ( ~n4930 & n10552 ) ;
  assign n20470 = n10950 ^ n3525 ^ 1'b0 ;
  assign n20471 = n327 & ~n20470 ;
  assign n20472 = n20469 & n20471 ;
  assign n20473 = n20472 ^ n15772 ^ 1'b0 ;
  assign n20474 = n14198 ^ n11509 ^ 1'b0 ;
  assign n20476 = ( n5866 & n7220 ) | ( n5866 & n14030 ) | ( n7220 & n14030 ) ;
  assign n20475 = ( n1309 & n1982 ) | ( n1309 & n5319 ) | ( n1982 & n5319 ) ;
  assign n20477 = n20476 ^ n20475 ^ 1'b0 ;
  assign n20478 = ( ~n15026 & n19889 ) | ( ~n15026 & n20477 ) | ( n19889 & n20477 ) ;
  assign n20479 = n2685 | n10291 ;
  assign n20480 = n14000 & ~n20479 ;
  assign n20481 = n20480 ^ n3593 ^ 1'b0 ;
  assign n20482 = n9506 ^ n7009 ^ 1'b0 ;
  assign n20483 = n1400 & ~n20482 ;
  assign n20490 = n20025 ^ n16530 ^ n1079 ;
  assign n20487 = n17116 ^ n5574 ^ 1'b0 ;
  assign n20488 = n19729 | n20487 ;
  assign n20489 = n595 | n20488 ;
  assign n20491 = n20490 ^ n20489 ^ 1'b0 ;
  assign n20484 = n5918 ^ n5682 ^ 1'b0 ;
  assign n20485 = n13874 & ~n20484 ;
  assign n20486 = n20485 ^ n13294 ^ n3500 ;
  assign n20492 = n20491 ^ n20486 ^ n5911 ;
  assign n20493 = ( n2150 & ~n6221 ) | ( n2150 & n18176 ) | ( ~n6221 & n18176 ) ;
  assign n20494 = ( n9068 & n16146 ) | ( n9068 & ~n20493 ) | ( n16146 & ~n20493 ) ;
  assign n20495 = n13442 & ~n14045 ;
  assign n20496 = n12402 & n20495 ;
  assign n20497 = n20496 ^ n2922 ^ 1'b0 ;
  assign n20498 = n12624 ^ n12602 ^ n5412 ;
  assign n20499 = n2535 | n20498 ;
  assign n20500 = n20497 & ~n20499 ;
  assign n20501 = n3959 & n8111 ;
  assign n20502 = n11657 & n17244 ;
  assign n20503 = n16601 ^ n7835 ^ n6520 ;
  assign n20504 = ( ~n16037 & n20502 ) | ( ~n16037 & n20503 ) | ( n20502 & n20503 ) ;
  assign n20505 = ( ~n4113 & n19271 ) | ( ~n4113 & n20504 ) | ( n19271 & n20504 ) ;
  assign n20506 = ( x23 & ~n971 ) | ( x23 & n5624 ) | ( ~n971 & n5624 ) ;
  assign n20507 = n20506 ^ n11720 ^ 1'b0 ;
  assign n20508 = ( ~n911 & n5761 ) | ( ~n911 & n13891 ) | ( n5761 & n13891 ) ;
  assign n20509 = n20508 ^ n14383 ^ n565 ;
  assign n20510 = n2913 ^ n819 ^ x245 ;
  assign n20511 = n14285 & n20510 ;
  assign n20512 = n10212 ^ n7463 ^ n3251 ;
  assign n20514 = n6642 | n9597 ;
  assign n20515 = n3554 & ~n20514 ;
  assign n20516 = n20515 ^ n4017 ^ 1'b0 ;
  assign n20513 = ( n289 & n10935 ) | ( n289 & ~n16111 ) | ( n10935 & ~n16111 ) ;
  assign n20517 = n20516 ^ n20513 ^ 1'b0 ;
  assign n20518 = n20512 & ~n20517 ;
  assign n20519 = n14309 & n20518 ;
  assign n20520 = ~n20511 & n20519 ;
  assign n20521 = n9450 ^ n7225 ^ n3405 ;
  assign n20522 = n20521 ^ n8615 ^ n3636 ;
  assign n20523 = n3690 & ~n4165 ;
  assign n20524 = ( n1532 & ~n13674 ) | ( n1532 & n20523 ) | ( ~n13674 & n20523 ) ;
  assign n20525 = n18975 ^ n11384 ^ n3035 ;
  assign n20526 = ( n2974 & ~n3286 ) | ( n2974 & n20525 ) | ( ~n3286 & n20525 ) ;
  assign n20527 = n20526 ^ n10326 ^ n5534 ;
  assign n20528 = n16118 ^ n5350 ^ 1'b0 ;
  assign n20529 = ( ~n20524 & n20527 ) | ( ~n20524 & n20528 ) | ( n20527 & n20528 ) ;
  assign n20530 = n13999 | n15475 ;
  assign n20531 = n3546 ^ n1491 ^ 1'b0 ;
  assign n20532 = n18388 & ~n20531 ;
  assign n20533 = n20532 ^ n13371 ^ n10565 ;
  assign n20534 = n578 & ~n20533 ;
  assign n20535 = n16522 & ~n19193 ;
  assign n20536 = n20535 ^ n1622 ^ n1046 ;
  assign n20537 = ~n2257 & n18000 ;
  assign n20538 = ( n20534 & n20536 ) | ( n20534 & n20537 ) | ( n20536 & n20537 ) ;
  assign n20543 = ( n7217 & n8332 ) | ( n7217 & ~n14122 ) | ( n8332 & ~n14122 ) ;
  assign n20539 = ~n979 & n8193 ;
  assign n20540 = n13671 ^ n1336 ^ 1'b0 ;
  assign n20541 = n20539 & ~n20540 ;
  assign n20542 = n20541 ^ n3389 ^ 1'b0 ;
  assign n20544 = n20543 ^ n20542 ^ n3989 ;
  assign n20546 = ( n915 & n17141 ) | ( n915 & ~n18125 ) | ( n17141 & ~n18125 ) ;
  assign n20545 = n1572 & n12762 ;
  assign n20547 = n20546 ^ n20545 ^ n1751 ;
  assign n20548 = n5044 ^ n1431 ^ n263 ;
  assign n20549 = ( ~n4625 & n8120 ) | ( ~n4625 & n15218 ) | ( n8120 & n15218 ) ;
  assign n20550 = ( n3129 & n8270 ) | ( n3129 & n8332 ) | ( n8270 & n8332 ) ;
  assign n20551 = ( ~n2865 & n10790 ) | ( ~n2865 & n20550 ) | ( n10790 & n20550 ) ;
  assign n20552 = n1921 & n3701 ;
  assign n20553 = ( n2430 & n6923 ) | ( n2430 & n11577 ) | ( n6923 & n11577 ) ;
  assign n20554 = ( n18244 & n20552 ) | ( n18244 & ~n20553 ) | ( n20552 & ~n20553 ) ;
  assign n20555 = n7153 | n14275 ;
  assign n20556 = n3832 | n20555 ;
  assign n20557 = n20556 ^ n8075 ^ 1'b0 ;
  assign n20558 = n20557 ^ n12121 ^ n974 ;
  assign n20559 = n11791 ^ n11483 ^ 1'b0 ;
  assign n20560 = n20558 & ~n20559 ;
  assign n20561 = n9917 & n13792 ;
  assign n20562 = n20561 ^ n10832 ^ 1'b0 ;
  assign n20563 = ( n20554 & n20560 ) | ( n20554 & ~n20562 ) | ( n20560 & ~n20562 ) ;
  assign n20564 = n14643 ^ n6060 ^ n3260 ;
  assign n20565 = ( n1650 & ~n4192 ) | ( n1650 & n4240 ) | ( ~n4192 & n4240 ) ;
  assign n20566 = ( n7450 & n20564 ) | ( n7450 & ~n20565 ) | ( n20564 & ~n20565 ) ;
  assign n20567 = n20566 ^ n4124 ^ 1'b0 ;
  assign n20568 = ( n6039 & n16097 ) | ( n6039 & n20567 ) | ( n16097 & n20567 ) ;
  assign n20569 = n478 & n20568 ;
  assign n20570 = n3501 ^ n3288 ^ n1482 ;
  assign n20571 = n20570 ^ n3927 ^ 1'b0 ;
  assign n20572 = n2590 & ~n14519 ;
  assign n20573 = n20571 & ~n20572 ;
  assign n20574 = n20569 & n20573 ;
  assign n20577 = n4444 ^ n3271 ^ 1'b0 ;
  assign n20578 = ~n2476 & n20577 ;
  assign n20575 = n17551 ^ n8866 ^ 1'b0 ;
  assign n20576 = n20575 ^ n3044 ^ n440 ;
  assign n20579 = n20578 ^ n20576 ^ n12211 ;
  assign n20580 = n13470 ^ n8255 ^ 1'b0 ;
  assign n20581 = ( n3185 & n11894 ) | ( n3185 & n12847 ) | ( n11894 & n12847 ) ;
  assign n20582 = n20581 ^ n9479 ^ 1'b0 ;
  assign n20583 = n20580 | n20582 ;
  assign n20585 = n6788 ^ n1595 ^ 1'b0 ;
  assign n20584 = n5033 ^ n4486 ^ n2029 ;
  assign n20586 = n20585 ^ n20584 ^ 1'b0 ;
  assign n20587 = n17783 & n20586 ;
  assign n20588 = n7862 ^ n5416 ^ n3483 ;
  assign n20589 = n15320 ^ n10294 ^ n5037 ;
  assign n20590 = n20589 ^ n14146 ^ n12077 ;
  assign n20591 = ( n20587 & ~n20588 ) | ( n20587 & n20590 ) | ( ~n20588 & n20590 ) ;
  assign n20592 = n20591 ^ n19083 ^ 1'b0 ;
  assign n20593 = n700 & ~n3488 ;
  assign n20594 = n10124 & n20593 ;
  assign n20595 = ( n798 & ~n864 ) | ( n798 & n7982 ) | ( ~n864 & n7982 ) ;
  assign n20596 = n5746 ^ n1591 ^ 1'b0 ;
  assign n20597 = n4691 | n13779 ;
  assign n20598 = ( n7035 & ~n20596 ) | ( n7035 & n20597 ) | ( ~n20596 & n20597 ) ;
  assign n20599 = ( n2738 & n20595 ) | ( n2738 & ~n20598 ) | ( n20595 & ~n20598 ) ;
  assign n20600 = n16180 ^ n15853 ^ n4960 ;
  assign n20601 = ( n11584 & n20599 ) | ( n11584 & ~n20600 ) | ( n20599 & ~n20600 ) ;
  assign n20602 = ~n20594 & n20601 ;
  assign n20603 = ( ~n1317 & n4557 ) | ( ~n1317 & n6579 ) | ( n4557 & n6579 ) ;
  assign n20604 = n20603 ^ n17829 ^ n14575 ;
  assign n20605 = n17657 ^ n716 ^ 1'b0 ;
  assign n20606 = n704 & n3916 ;
  assign n20607 = n19002 | n20606 ;
  assign n20608 = n16137 & ~n20607 ;
  assign n20609 = n5249 ^ n1037 ^ x196 ;
  assign n20611 = n14674 ^ n10010 ^ 1'b0 ;
  assign n20612 = n6338 | n20611 ;
  assign n20610 = n11712 & n15059 ;
  assign n20613 = n20612 ^ n20610 ^ 1'b0 ;
  assign n20614 = ~n7995 & n17084 ;
  assign n20615 = ~n20613 & n20614 ;
  assign n20616 = n4509 | n11923 ;
  assign n20617 = ( ~n5221 & n8738 ) | ( ~n5221 & n20616 ) | ( n8738 & n20616 ) ;
  assign n20618 = n11811 ^ n10253 ^ n5811 ;
  assign n20619 = n13162 ^ n7890 ^ n5456 ;
  assign n20620 = n11126 ^ n9769 ^ n1652 ;
  assign n20621 = n20619 & ~n20620 ;
  assign n20622 = n3532 & n6329 ;
  assign n20623 = ~n4358 & n13403 ;
  assign n20624 = n504 & ~n20623 ;
  assign n20625 = n20624 ^ n9087 ^ 1'b0 ;
  assign n20627 = ( n1693 & n10356 ) | ( n1693 & n14246 ) | ( n10356 & n14246 ) ;
  assign n20626 = n8083 | n11984 ;
  assign n20628 = n20627 ^ n20626 ^ 1'b0 ;
  assign n20629 = n3135 | n5981 ;
  assign n20630 = n20629 ^ n3158 ^ 1'b0 ;
  assign n20631 = ( n14060 & n18171 ) | ( n14060 & n20630 ) | ( n18171 & n20630 ) ;
  assign n20632 = ( ~n3916 & n19017 ) | ( ~n3916 & n20631 ) | ( n19017 & n20631 ) ;
  assign n20633 = n7723 ^ n4733 ^ x169 ;
  assign n20634 = n8443 & n20633 ;
  assign n20635 = n14112 ^ n6587 ^ n5020 ;
  assign n20636 = n20635 ^ n14933 ^ n5929 ;
  assign n20637 = n20636 ^ n11588 ^ 1'b0 ;
  assign n20638 = n2275 | n20637 ;
  assign n20639 = n20638 ^ n3874 ^ 1'b0 ;
  assign n20640 = n2181 | n18414 ;
  assign n20641 = n18784 ^ n7174 ^ n2182 ;
  assign n20642 = n2035 & ~n15166 ;
  assign n20643 = ( ~n11924 & n20641 ) | ( ~n11924 & n20642 ) | ( n20641 & n20642 ) ;
  assign n20644 = n15582 ^ n13999 ^ 1'b0 ;
  assign n20645 = n2680 & n20644 ;
  assign n20649 = n20307 ^ n5725 ^ 1'b0 ;
  assign n20646 = ~n12603 & n18149 ;
  assign n20647 = n9267 & n20646 ;
  assign n20648 = n20647 ^ n18155 ^ 1'b0 ;
  assign n20650 = n20649 ^ n20648 ^ n5797 ;
  assign n20651 = ( n4328 & ~n12890 ) | ( n4328 & n20650 ) | ( ~n12890 & n20650 ) ;
  assign n20652 = ( n14190 & ~n20645 ) | ( n14190 & n20651 ) | ( ~n20645 & n20651 ) ;
  assign n20653 = n18175 ^ n15118 ^ 1'b0 ;
  assign n20654 = n20652 | n20653 ;
  assign n20655 = n6199 & ~n6500 ;
  assign n20656 = n11845 & n20655 ;
  assign n20657 = n20656 ^ n16493 ^ n2081 ;
  assign n20658 = ( ~n2923 & n7294 ) | ( ~n2923 & n7870 ) | ( n7294 & n7870 ) ;
  assign n20659 = ( ~n5666 & n20657 ) | ( ~n5666 & n20658 ) | ( n20657 & n20658 ) ;
  assign n20660 = n1312 & ~n11164 ;
  assign n20661 = n2001 & n20660 ;
  assign n20662 = n20661 ^ n10150 ^ 1'b0 ;
  assign n20663 = n7225 ^ n5596 ^ 1'b0 ;
  assign n20664 = ( n10881 & n11803 ) | ( n10881 & ~n20663 ) | ( n11803 & ~n20663 ) ;
  assign n20665 = n20664 ^ n5838 ^ 1'b0 ;
  assign n20666 = x61 & n5585 ;
  assign n20667 = n20666 ^ n18921 ^ n12109 ;
  assign n20668 = n8679 | n14097 ;
  assign n20669 = n20668 ^ n9071 ^ 1'b0 ;
  assign n20670 = n10870 & n20669 ;
  assign n20671 = n7315 ^ n6029 ^ n4713 ;
  assign n20672 = n20671 ^ n8173 ^ 1'b0 ;
  assign n20673 = n13016 ^ n7542 ^ n501 ;
  assign n20674 = n20673 ^ n15804 ^ n8680 ;
  assign n20675 = n5053 ^ n2981 ^ n2664 ;
  assign n20676 = n20675 ^ n10570 ^ n287 ;
  assign n20677 = ( n4527 & ~n14236 ) | ( n4527 & n20676 ) | ( ~n14236 & n20676 ) ;
  assign n20678 = ( ~n11250 & n12634 ) | ( ~n11250 & n20677 ) | ( n12634 & n20677 ) ;
  assign n20679 = ( ~x215 & n14186 ) | ( ~x215 & n20678 ) | ( n14186 & n20678 ) ;
  assign n20680 = n20679 ^ n6244 ^ 1'b0 ;
  assign n20681 = n20674 | n20680 ;
  assign n20682 = ~n9479 & n16762 ;
  assign n20683 = ~n6223 & n20682 ;
  assign n20684 = n7027 ^ n5024 ^ n5006 ;
  assign n20685 = n3147 & ~n6223 ;
  assign n20686 = ( n2367 & ~n2766 ) | ( n2367 & n10627 ) | ( ~n2766 & n10627 ) ;
  assign n20687 = ( ~n5158 & n5756 ) | ( ~n5158 & n13063 ) | ( n5756 & n13063 ) ;
  assign n20688 = ( n20685 & ~n20686 ) | ( n20685 & n20687 ) | ( ~n20686 & n20687 ) ;
  assign n20689 = n20688 ^ n17045 ^ n9903 ;
  assign n20690 = ~n3021 & n14736 ;
  assign n20691 = n20690 ^ n4798 ^ n4726 ;
  assign n20692 = n8166 & n15236 ;
  assign n20693 = ~n17972 & n20692 ;
  assign n20694 = ( n7996 & ~n13341 ) | ( n7996 & n20693 ) | ( ~n13341 & n20693 ) ;
  assign n20696 = ( n4097 & n9185 ) | ( n4097 & ~n13578 ) | ( n9185 & ~n13578 ) ;
  assign n20697 = n20696 ^ n4371 ^ n808 ;
  assign n20695 = ~n4910 & n12749 ;
  assign n20698 = n20697 ^ n20695 ^ 1'b0 ;
  assign n20699 = n20698 ^ n9239 ^ 1'b0 ;
  assign n20700 = n8668 | n15611 ;
  assign n20701 = n4841 | n20700 ;
  assign n20704 = n20462 ^ n13629 ^ 1'b0 ;
  assign n20702 = n16065 ^ n12004 ^ n9602 ;
  assign n20703 = ~n2265 & n20702 ;
  assign n20705 = n20704 ^ n20703 ^ 1'b0 ;
  assign n20706 = ( n3412 & ~n11393 ) | ( n3412 & n12708 ) | ( ~n11393 & n12708 ) ;
  assign n20707 = n20706 ^ n3509 ^ n1578 ;
  assign n20708 = n13042 ^ n10446 ^ n1665 ;
  assign n20709 = n19259 ^ n6955 ^ 1'b0 ;
  assign n20710 = ~n20708 & n20709 ;
  assign n20711 = n20710 ^ n11972 ^ n6571 ;
  assign n20712 = ~n20707 & n20711 ;
  assign n20713 = ~n19916 & n20712 ;
  assign n20714 = n9464 ^ n5447 ^ n2217 ;
  assign n20715 = ( ~n3053 & n6186 ) | ( ~n3053 & n6223 ) | ( n6186 & n6223 ) ;
  assign n20716 = ( x93 & n19349 ) | ( x93 & ~n20715 ) | ( n19349 & ~n20715 ) ;
  assign n20717 = n12452 ^ n9721 ^ n1805 ;
  assign n20718 = n12109 ^ n10764 ^ 1'b0 ;
  assign n20719 = n20717 | n20718 ;
  assign n20720 = n20719 ^ n11260 ^ x27 ;
  assign n20721 = n7952 & n14053 ;
  assign n20722 = ~x224 & n20721 ;
  assign n20723 = ( n6480 & ~n14227 ) | ( n6480 & n17892 ) | ( ~n14227 & n17892 ) ;
  assign n20724 = n10983 ^ n10418 ^ n7176 ;
  assign n20725 = ~n5735 & n20724 ;
  assign n20726 = ~n7141 & n20725 ;
  assign n20727 = ( x227 & ~n1587 ) | ( x227 & n3326 ) | ( ~n1587 & n3326 ) ;
  assign n20728 = ( n8024 & ~n8866 ) | ( n8024 & n20727 ) | ( ~n8866 & n20727 ) ;
  assign n20729 = n20728 ^ n14232 ^ n3543 ;
  assign n20730 = n7907 ^ n3713 ^ 1'b0 ;
  assign n20731 = ~n13091 & n20730 ;
  assign n20732 = ( ~n13651 & n20729 ) | ( ~n13651 & n20731 ) | ( n20729 & n20731 ) ;
  assign n20733 = ( n18896 & n20726 ) | ( n18896 & ~n20732 ) | ( n20726 & ~n20732 ) ;
  assign n20734 = n19478 ^ n9712 ^ n6861 ;
  assign n20735 = n6039 ^ n5237 ^ n2883 ;
  assign n20736 = n20735 ^ n13513 ^ n7348 ;
  assign n20737 = n20736 ^ n18547 ^ n8946 ;
  assign n20738 = ( ~n11913 & n13079 ) | ( ~n11913 & n20737 ) | ( n13079 & n20737 ) ;
  assign n20740 = n4713 & ~n12229 ;
  assign n20741 = n20740 ^ n14455 ^ 1'b0 ;
  assign n20739 = n4917 ^ n4015 ^ n790 ;
  assign n20742 = n20741 ^ n20739 ^ 1'b0 ;
  assign n20743 = n19781 & n20742 ;
  assign n20744 = ( ~n639 & n5896 ) | ( ~n639 & n7764 ) | ( n5896 & n7764 ) ;
  assign n20745 = ( n3027 & n3126 ) | ( n3027 & n20744 ) | ( n3126 & n20744 ) ;
  assign n20746 = n1827 & n6865 ;
  assign n20747 = n20746 ^ n9535 ^ n9382 ;
  assign n20748 = ( n7863 & ~n13403 ) | ( n7863 & n20747 ) | ( ~n13403 & n20747 ) ;
  assign n20749 = n20748 ^ n20606 ^ n1304 ;
  assign n20751 = n16923 ^ n11533 ^ n10061 ;
  assign n20752 = ( n1795 & n7176 ) | ( n1795 & n20751 ) | ( n7176 & n20751 ) ;
  assign n20750 = n12760 & ~n15471 ;
  assign n20753 = n20752 ^ n20750 ^ n12571 ;
  assign n20757 = n9736 & ~n11155 ;
  assign n20758 = n20757 ^ n19450 ^ 1'b0 ;
  assign n20759 = n20758 ^ n7398 ^ n6737 ;
  assign n20754 = n13792 ^ n12182 ^ 1'b0 ;
  assign n20755 = n9127 ^ n259 ^ 1'b0 ;
  assign n20756 = n20754 & n20755 ;
  assign n20760 = n20759 ^ n20756 ^ n1603 ;
  assign n20761 = n10808 ^ x237 ^ 1'b0 ;
  assign n20762 = n599 | n20761 ;
  assign n20763 = ( n4998 & n5592 ) | ( n4998 & ~n15166 ) | ( n5592 & ~n15166 ) ;
  assign n20764 = ( n7260 & n20762 ) | ( n7260 & n20763 ) | ( n20762 & n20763 ) ;
  assign n20765 = n8659 ^ n3844 ^ n2275 ;
  assign n20766 = ( ~n12239 & n14726 ) | ( ~n12239 & n20765 ) | ( n14726 & n20765 ) ;
  assign n20767 = n4440 | n20766 ;
  assign n20768 = n20767 ^ n11240 ^ 1'b0 ;
  assign n20769 = n11730 ^ n5368 ^ n4524 ;
  assign n20770 = n15022 ^ n12930 ^ 1'b0 ;
  assign n20771 = n15167 & n20770 ;
  assign n20772 = n1135 & n1930 ;
  assign n20773 = n20772 ^ n5250 ^ 1'b0 ;
  assign n20774 = n11338 ^ n10314 ^ 1'b0 ;
  assign n20775 = ( n7880 & ~n12907 ) | ( n7880 & n20774 ) | ( ~n12907 & n20774 ) ;
  assign n20776 = n19106 ^ n18645 ^ n9303 ;
  assign n20782 = n8026 ^ n2770 ^ n721 ;
  assign n20783 = n20782 ^ n4672 ^ 1'b0 ;
  assign n20784 = n7661 | n20783 ;
  assign n20777 = ( ~n4860 & n6994 ) | ( ~n4860 & n10699 ) | ( n6994 & n10699 ) ;
  assign n20778 = n20777 ^ n13001 ^ 1'b0 ;
  assign n20779 = n2067 | n20778 ;
  assign n20780 = n18842 | n20779 ;
  assign n20781 = n20780 ^ n20437 ^ 1'b0 ;
  assign n20785 = n20784 ^ n20781 ^ 1'b0 ;
  assign n20786 = n20776 | n20785 ;
  assign n20787 = n12975 ^ n9747 ^ 1'b0 ;
  assign n20788 = ( n7667 & n12519 ) | ( n7667 & ~n19539 ) | ( n12519 & ~n19539 ) ;
  assign n20789 = ~x151 & n20788 ;
  assign n20790 = n20787 | n20789 ;
  assign n20791 = n14079 & ~n20790 ;
  assign n20794 = n9167 ^ n6824 ^ 1'b0 ;
  assign n20795 = n17765 & n20794 ;
  assign n20796 = n20795 ^ n933 ^ 1'b0 ;
  assign n20793 = ( n1955 & ~n3668 ) | ( n1955 & n14826 ) | ( ~n3668 & n14826 ) ;
  assign n20792 = n10383 ^ n10358 ^ n10334 ;
  assign n20797 = n20796 ^ n20793 ^ n20792 ;
  assign n20798 = n16252 ^ n1590 ^ 1'b0 ;
  assign n20799 = n20798 ^ n10150 ^ n4067 ;
  assign n20800 = ( n2100 & n3163 ) | ( n2100 & n3431 ) | ( n3163 & n3431 ) ;
  assign n20801 = n3360 & ~n14444 ;
  assign n20802 = n20800 & ~n20801 ;
  assign n20803 = ~n8197 & n20802 ;
  assign n20804 = ( n3410 & ~n7483 ) | ( n3410 & n9014 ) | ( ~n7483 & n9014 ) ;
  assign n20805 = n20804 ^ n16455 ^ n15932 ;
  assign n20806 = n3336 | n15421 ;
  assign n20807 = x42 | n20806 ;
  assign n20808 = ~n12102 & n16166 ;
  assign n20809 = ( n4641 & n6046 ) | ( n4641 & ~n20808 ) | ( n6046 & ~n20808 ) ;
  assign n20810 = ( ~n5996 & n20807 ) | ( ~n5996 & n20809 ) | ( n20807 & n20809 ) ;
  assign n20811 = n6672 ^ n3102 ^ n2092 ;
  assign n20812 = ( ~n2598 & n9956 ) | ( ~n2598 & n20811 ) | ( n9956 & n20811 ) ;
  assign n20813 = n11238 ^ n7805 ^ 1'b0 ;
  assign n20814 = n20600 & n20813 ;
  assign n20815 = n17990 ^ n8990 ^ 1'b0 ;
  assign n20816 = n8339 & n20815 ;
  assign n20817 = ( n1366 & n2956 ) | ( n1366 & ~n17088 ) | ( n2956 & ~n17088 ) ;
  assign n20818 = ( ~n1875 & n17592 ) | ( ~n1875 & n20817 ) | ( n17592 & n20817 ) ;
  assign n20822 = n2800 | n10826 ;
  assign n20823 = n3138 & ~n20822 ;
  assign n20824 = n20823 ^ n914 ^ 1'b0 ;
  assign n20819 = n10943 ^ n5572 ^ 1'b0 ;
  assign n20820 = n6486 | n20819 ;
  assign n20821 = n12947 & ~n20820 ;
  assign n20825 = n20824 ^ n20821 ^ 1'b0 ;
  assign n20826 = n1664 & n5469 ;
  assign n20827 = ( n4023 & ~n12405 ) | ( n4023 & n20826 ) | ( ~n12405 & n20826 ) ;
  assign n20828 = n14857 ^ n4656 ^ 1'b0 ;
  assign n20829 = n6671 & n20828 ;
  assign n20830 = n19258 & n20829 ;
  assign n20831 = ~n20827 & n20830 ;
  assign n20832 = n7467 | n11971 ;
  assign n20833 = n5941 | n20832 ;
  assign n20834 = n20833 ^ n3803 ^ n2168 ;
  assign n20835 = ~n4238 & n18982 ;
  assign n20836 = n20834 & ~n20835 ;
  assign n20837 = n16742 ^ n5423 ^ n5381 ;
  assign n20838 = ( n1602 & ~n9039 ) | ( n1602 & n13205 ) | ( ~n9039 & n13205 ) ;
  assign n20839 = n20838 ^ n12630 ^ n983 ;
  assign n20840 = ( n12936 & n16785 ) | ( n12936 & ~n20839 ) | ( n16785 & ~n20839 ) ;
  assign n20841 = n2807 | n2994 ;
  assign n20842 = n20840 & ~n20841 ;
  assign n20843 = ( n5471 & n5538 ) | ( n5471 & ~n20842 ) | ( n5538 & ~n20842 ) ;
  assign n20845 = ( ~n4273 & n4427 ) | ( ~n4273 & n7709 ) | ( n4427 & n7709 ) ;
  assign n20844 = ( n4427 & n6898 ) | ( n4427 & ~n7341 ) | ( n6898 & ~n7341 ) ;
  assign n20846 = n20845 ^ n20844 ^ n9872 ;
  assign n20847 = n20846 ^ n14073 ^ 1'b0 ;
  assign n20848 = ( n16145 & n17387 ) | ( n16145 & ~n20847 ) | ( n17387 & ~n20847 ) ;
  assign n20849 = n20848 ^ n2966 ^ 1'b0 ;
  assign n20850 = n2757 & n20849 ;
  assign n20853 = ( n3695 & n7975 ) | ( n3695 & n11476 ) | ( n7975 & n11476 ) ;
  assign n20851 = n15921 ^ n2911 ^ n2885 ;
  assign n20852 = n20851 ^ n13913 ^ n7842 ;
  assign n20854 = n20853 ^ n20852 ^ n8599 ;
  assign n20855 = n13413 ^ n5086 ^ 1'b0 ;
  assign n20856 = ( n3492 & n5929 ) | ( n3492 & ~n7708 ) | ( n5929 & ~n7708 ) ;
  assign n20857 = n17519 ^ n5814 ^ 1'b0 ;
  assign n20858 = ~n20856 & n20857 ;
  assign n20859 = ( n20132 & ~n20855 ) | ( n20132 & n20858 ) | ( ~n20855 & n20858 ) ;
  assign n20860 = n17875 ^ n2427 ^ 1'b0 ;
  assign n20861 = n2021 & n20860 ;
  assign n20862 = ( n8577 & n20377 ) | ( n8577 & n20861 ) | ( n20377 & n20861 ) ;
  assign n20863 = ( n2985 & n3710 ) | ( n2985 & n11914 ) | ( n3710 & n11914 ) ;
  assign n20864 = ( n4999 & n8903 ) | ( n4999 & n18283 ) | ( n8903 & n18283 ) ;
  assign n20865 = n14879 ^ n9471 ^ n2397 ;
  assign n20866 = n20865 ^ n6833 ^ 1'b0 ;
  assign n20867 = ~n20864 & n20866 ;
  assign n20868 = ( x87 & n828 ) | ( x87 & n1125 ) | ( n828 & n1125 ) ;
  assign n20869 = x243 & ~n13659 ;
  assign n20870 = n20869 ^ n661 ^ 1'b0 ;
  assign n20871 = n20868 | n20870 ;
  assign n20878 = n17946 ^ n5942 ^ n3846 ;
  assign n20875 = n10849 ^ n7585 ^ n1041 ;
  assign n20872 = ( ~n3703 & n10363 ) | ( ~n3703 & n14444 ) | ( n10363 & n14444 ) ;
  assign n20873 = ( n5002 & ~n8197 ) | ( n5002 & n20872 ) | ( ~n8197 & n20872 ) ;
  assign n20874 = n1001 & ~n20873 ;
  assign n20876 = n20875 ^ n20874 ^ 1'b0 ;
  assign n20877 = n20876 ^ n19227 ^ 1'b0 ;
  assign n20879 = n20878 ^ n20877 ^ 1'b0 ;
  assign n20880 = n2650 & n14631 ;
  assign n20881 = n20880 ^ n887 ^ 1'b0 ;
  assign n20882 = n20881 ^ n7057 ^ n1428 ;
  assign n20883 = ( n515 & n4760 ) | ( n515 & n10329 ) | ( n4760 & n10329 ) ;
  assign n20884 = n2562 & ~n4438 ;
  assign n20885 = n9346 ^ n825 ^ 1'b0 ;
  assign n20886 = n20884 | n20885 ;
  assign n20887 = x60 & ~n8263 ;
  assign n20888 = ( n662 & n17435 ) | ( n662 & ~n20887 ) | ( n17435 & ~n20887 ) ;
  assign n20889 = n5340 ^ n3397 ^ n3379 ;
  assign n20890 = n20889 ^ n3967 ^ 1'b0 ;
  assign n20891 = n20890 ^ n6984 ^ 1'b0 ;
  assign n20892 = n20891 ^ n1676 ^ 1'b0 ;
  assign n20896 = n11503 & ~n18794 ;
  assign n20893 = n552 & n1165 ;
  assign n20894 = n20893 ^ n8731 ^ 1'b0 ;
  assign n20895 = n7586 | n20894 ;
  assign n20897 = n20896 ^ n20895 ^ 1'b0 ;
  assign n20898 = n19573 ^ n12562 ^ n3270 ;
  assign n20899 = ( n1098 & n6204 ) | ( n1098 & ~n17998 ) | ( n6204 & ~n17998 ) ;
  assign n20900 = n20899 ^ n15471 ^ 1'b0 ;
  assign n20901 = ( ~n1066 & n2622 ) | ( ~n1066 & n11742 ) | ( n2622 & n11742 ) ;
  assign n20902 = ( n4239 & n9061 ) | ( n4239 & ~n10584 ) | ( n9061 & ~n10584 ) ;
  assign n20903 = n14842 ^ n13339 ^ n1072 ;
  assign n20904 = ( n7025 & n11450 ) | ( n7025 & ~n20903 ) | ( n11450 & ~n20903 ) ;
  assign n20905 = n20904 ^ n2520 ^ 1'b0 ;
  assign n20906 = ~n20902 & n20905 ;
  assign n20907 = n1760 & ~n4047 ;
  assign n20908 = ~n17683 & n20907 ;
  assign n20909 = ( n1901 & n18598 ) | ( n1901 & ~n20908 ) | ( n18598 & ~n20908 ) ;
  assign n20910 = ( n2998 & n7905 ) | ( n2998 & ~n8967 ) | ( n7905 & ~n8967 ) ;
  assign n20911 = ( n5381 & n7415 ) | ( n5381 & ~n20910 ) | ( n7415 & ~n20910 ) ;
  assign n20912 = ( ~n8357 & n13470 ) | ( ~n8357 & n20911 ) | ( n13470 & n20911 ) ;
  assign n20913 = n12248 ^ n11940 ^ 1'b0 ;
  assign n20914 = ( n3794 & ~n20912 ) | ( n3794 & n20913 ) | ( ~n20912 & n20913 ) ;
  assign n20915 = n9486 ^ n5864 ^ 1'b0 ;
  assign n20916 = ( n9744 & ~n10845 ) | ( n9744 & n20056 ) | ( ~n10845 & n20056 ) ;
  assign n20917 = ( n563 & n20915 ) | ( n563 & n20916 ) | ( n20915 & n20916 ) ;
  assign n20918 = n20917 ^ n9446 ^ 1'b0 ;
  assign n20919 = n1020 & ~n20918 ;
  assign n20920 = n3932 & ~n13001 ;
  assign n20921 = n18060 ^ n3128 ^ 1'b0 ;
  assign n20922 = n15452 | n20921 ;
  assign n20923 = n6010 & n20922 ;
  assign n20924 = n3878 ^ n3713 ^ n691 ;
  assign n20925 = ( n6383 & n17458 ) | ( n6383 & ~n20924 ) | ( n17458 & ~n20924 ) ;
  assign n20926 = ( n1141 & ~n4673 ) | ( n1141 & n20925 ) | ( ~n4673 & n20925 ) ;
  assign n20928 = n355 | n4323 ;
  assign n20929 = n20928 ^ n13306 ^ 1'b0 ;
  assign n20927 = n16333 ^ n4250 ^ n418 ;
  assign n20930 = n20929 ^ n20927 ^ 1'b0 ;
  assign n20931 = ( n2737 & n5774 ) | ( n2737 & ~n9477 ) | ( n5774 & ~n9477 ) ;
  assign n20932 = ( n2512 & n5257 ) | ( n2512 & n8187 ) | ( n5257 & n8187 ) ;
  assign n20933 = n2224 & n20932 ;
  assign n20934 = ( n7423 & n20931 ) | ( n7423 & ~n20933 ) | ( n20931 & ~n20933 ) ;
  assign n20935 = ( ~n1201 & n8142 ) | ( ~n1201 & n20934 ) | ( n8142 & n20934 ) ;
  assign n20936 = ~n11839 & n20935 ;
  assign n20937 = n10272 ^ n6049 ^ n4207 ;
  assign n20938 = n10300 & ~n15825 ;
  assign n20939 = ( n4851 & n9482 ) | ( n4851 & n10708 ) | ( n9482 & n10708 ) ;
  assign n20940 = ( n4320 & n5611 ) | ( n4320 & n17431 ) | ( n5611 & n17431 ) ;
  assign n20941 = n12012 ^ n7807 ^ n2440 ;
  assign n20942 = ( ~n968 & n20940 ) | ( ~n968 & n20941 ) | ( n20940 & n20941 ) ;
  assign n20943 = n20942 ^ n9946 ^ n1806 ;
  assign n20944 = n20943 ^ n18753 ^ 1'b0 ;
  assign n20945 = n20939 & ~n20944 ;
  assign n20946 = n6573 ^ n5916 ^ 1'b0 ;
  assign n20947 = ( ~n15089 & n15827 ) | ( ~n15089 & n20946 ) | ( n15827 & n20946 ) ;
  assign n20948 = ( n12814 & n20945 ) | ( n12814 & ~n20947 ) | ( n20945 & ~n20947 ) ;
  assign n20949 = n6170 ^ n1047 ^ x129 ;
  assign n20950 = ( n4586 & n9124 ) | ( n4586 & n20949 ) | ( n9124 & n20949 ) ;
  assign n20951 = n20950 ^ n13894 ^ n2137 ;
  assign n20952 = n11274 ^ n6913 ^ n2806 ;
  assign n20953 = ~n5637 & n20952 ;
  assign n20954 = n12901 & n20953 ;
  assign n20959 = n2781 ^ n2765 ^ 1'b0 ;
  assign n20960 = ~n5133 & n20959 ;
  assign n20955 = ~n3995 & n17012 ;
  assign n20956 = ~n12365 & n20955 ;
  assign n20957 = n7467 | n20956 ;
  assign n20958 = n4257 & ~n20957 ;
  assign n20961 = n20960 ^ n20958 ^ 1'b0 ;
  assign n20962 = n20954 | n20961 ;
  assign n20963 = n16397 & n20962 ;
  assign n20964 = n4672 & ~n18649 ;
  assign n20965 = n20964 ^ n3881 ^ 1'b0 ;
  assign n20966 = n20965 ^ n13066 ^ 1'b0 ;
  assign n20967 = n3350 & ~n20966 ;
  assign n20968 = n5737 & n7970 ;
  assign n20969 = ~n3840 & n20968 ;
  assign n20970 = n20969 ^ n1361 ^ 1'b0 ;
  assign n20971 = n20970 ^ n13909 ^ n12282 ;
  assign n20972 = n899 | n3490 ;
  assign n20973 = ~n10922 & n15835 ;
  assign n20974 = n20972 & ~n20973 ;
  assign n20975 = n20974 ^ n17705 ^ n507 ;
  assign n20976 = ( n12858 & n15660 ) | ( n12858 & ~n15918 ) | ( n15660 & ~n15918 ) ;
  assign n20977 = ~n1106 & n2290 ;
  assign n20978 = n8614 ^ n5620 ^ n2581 ;
  assign n20979 = ( n447 & n7015 ) | ( n447 & ~n20978 ) | ( n7015 & ~n20978 ) ;
  assign n20980 = n20979 ^ n9208 ^ 1'b0 ;
  assign n20981 = n16542 & ~n19082 ;
  assign n20982 = ( n9777 & n17600 ) | ( n9777 & ~n20981 ) | ( n17600 & ~n20981 ) ;
  assign n20987 = n12247 ^ n9270 ^ 1'b0 ;
  assign n20984 = n350 & ~n469 ;
  assign n20985 = n20984 ^ n6039 ^ 1'b0 ;
  assign n20983 = n5592 & ~n11256 ;
  assign n20986 = n20985 ^ n20983 ^ n2198 ;
  assign n20988 = n20987 ^ n20986 ^ n11313 ;
  assign n20989 = n9745 ^ n3519 ^ n1152 ;
  assign n20990 = n13094 ^ n7649 ^ n398 ;
  assign n20991 = n1561 | n20990 ;
  assign n20992 = n6622 | n20991 ;
  assign n20993 = n20989 & n20992 ;
  assign n20995 = n3200 | n3799 ;
  assign n20996 = n20995 ^ n8749 ^ n1490 ;
  assign n20997 = n20996 ^ n5034 ^ 1'b0 ;
  assign n20998 = n20997 ^ n9452 ^ 1'b0 ;
  assign n20999 = n20998 ^ n12905 ^ n6357 ;
  assign n20994 = n8248 | n15654 ;
  assign n21000 = n20999 ^ n20994 ^ 1'b0 ;
  assign n21002 = ( ~n331 & n5329 ) | ( ~n331 & n12468 ) | ( n5329 & n12468 ) ;
  assign n21003 = n4498 | n21002 ;
  assign n21004 = n21003 ^ n13062 ^ 1'b0 ;
  assign n21005 = ~n3800 & n21004 ;
  assign n21006 = n21005 ^ n20998 ^ n5525 ;
  assign n21001 = n324 & ~n3340 ;
  assign n21007 = n21006 ^ n21001 ^ 1'b0 ;
  assign n21008 = n9193 ^ n2083 ^ 1'b0 ;
  assign n21009 = n21008 ^ n8083 ^ n2043 ;
  assign n21010 = n13161 ^ n2851 ^ 1'b0 ;
  assign n21011 = ( n1625 & ~n15453 ) | ( n1625 & n21010 ) | ( ~n15453 & n21010 ) ;
  assign n21012 = n21011 ^ n19497 ^ n7514 ;
  assign n21013 = n4397 | n7054 ;
  assign n21014 = n15697 ^ n13503 ^ 1'b0 ;
  assign n21015 = ( n6630 & n8030 ) | ( n6630 & n16042 ) | ( n8030 & n16042 ) ;
  assign n21016 = ~n2965 & n21015 ;
  assign n21017 = ( n4670 & ~n9930 ) | ( n4670 & n19808 ) | ( ~n9930 & n19808 ) ;
  assign n21018 = ( ~n875 & n5098 ) | ( ~n875 & n6523 ) | ( n5098 & n6523 ) ;
  assign n21019 = ( ~n8842 & n16319 ) | ( ~n8842 & n21018 ) | ( n16319 & n21018 ) ;
  assign n21020 = n15939 & n18551 ;
  assign n21021 = n21020 ^ n17645 ^ 1'b0 ;
  assign n21022 = n13504 ^ n8967 ^ n4725 ;
  assign n21023 = x222 & ~n21022 ;
  assign n21024 = n21023 ^ n2603 ^ n1953 ;
  assign n21025 = ( n8430 & ~n14741 ) | ( n8430 & n21024 ) | ( ~n14741 & n21024 ) ;
  assign n21026 = n3311 | n21025 ;
  assign n21027 = n21026 ^ n19579 ^ 1'b0 ;
  assign n21028 = n10893 ^ n6613 ^ n6062 ;
  assign n21031 = n12442 ^ n7761 ^ n7560 ;
  assign n21029 = n378 & ~n2488 ;
  assign n21030 = n21029 ^ n10892 ^ 1'b0 ;
  assign n21032 = n21031 ^ n21030 ^ x125 ;
  assign n21033 = n21032 ^ n3176 ^ 1'b0 ;
  assign n21034 = n5237 & n21033 ;
  assign n21035 = ( n1365 & ~n5818 ) | ( n1365 & n21034 ) | ( ~n5818 & n21034 ) ;
  assign n21036 = n8422 & ~n20777 ;
  assign n21037 = n21036 ^ n12742 ^ 1'b0 ;
  assign n21038 = n3962 | n20690 ;
  assign n21039 = n14874 ^ n12582 ^ 1'b0 ;
  assign n21040 = ( n6327 & n21038 ) | ( n6327 & ~n21039 ) | ( n21038 & ~n21039 ) ;
  assign n21041 = ~n4124 & n12953 ;
  assign n21042 = n21041 ^ x133 ^ 1'b0 ;
  assign n21043 = n21040 & ~n21042 ;
  assign n21044 = n21043 ^ n10781 ^ 1'b0 ;
  assign n21046 = n7585 ^ n5468 ^ n1390 ;
  assign n21045 = n16729 ^ n13935 ^ n5066 ;
  assign n21047 = n21046 ^ n21045 ^ n17404 ;
  assign n21048 = ( n678 & n1484 ) | ( n678 & n7017 ) | ( n1484 & n7017 ) ;
  assign n21049 = n9562 | n21048 ;
  assign n21050 = ( n2509 & ~n11389 ) | ( n2509 & n12526 ) | ( ~n11389 & n12526 ) ;
  assign n21051 = ~n3118 & n21050 ;
  assign n21061 = n315 & n5580 ;
  assign n21060 = n18388 ^ n5751 ^ n1436 ;
  assign n21052 = n1425 & ~n4784 ;
  assign n21053 = n21052 ^ n704 ^ 1'b0 ;
  assign n21054 = n2185 | n8780 ;
  assign n21055 = n21054 ^ n12720 ^ n8540 ;
  assign n21056 = n7124 | n10969 ;
  assign n21057 = n7337 & n21056 ;
  assign n21058 = n21057 ^ n8438 ^ n2232 ;
  assign n21059 = ( ~n21053 & n21055 ) | ( ~n21053 & n21058 ) | ( n21055 & n21058 ) ;
  assign n21062 = n21061 ^ n21060 ^ n21059 ;
  assign n21063 = x249 & ~n15317 ;
  assign n21064 = ~n2981 & n21063 ;
  assign n21065 = n15873 | n17232 ;
  assign n21066 = ~n20915 & n21065 ;
  assign n21067 = ~n11175 & n21066 ;
  assign n21071 = ( n2804 & n5637 ) | ( n2804 & n14007 ) | ( n5637 & n14007 ) ;
  assign n21068 = n13657 ^ n3707 ^ 1'b0 ;
  assign n21069 = n13412 & n21068 ;
  assign n21070 = ( n4165 & n10119 ) | ( n4165 & ~n21069 ) | ( n10119 & ~n21069 ) ;
  assign n21072 = n21071 ^ n21070 ^ n13195 ;
  assign n21076 = ( n1539 & n3064 ) | ( n1539 & n9387 ) | ( n3064 & n9387 ) ;
  assign n21073 = n7030 ^ n864 ^ 1'b0 ;
  assign n21074 = ~n1571 & n21073 ;
  assign n21075 = ( ~n2517 & n9004 ) | ( ~n2517 & n21074 ) | ( n9004 & n21074 ) ;
  assign n21077 = n21076 ^ n21075 ^ n8978 ;
  assign n21078 = n21077 ^ n5591 ^ n2059 ;
  assign n21079 = ( n4192 & ~n8882 ) | ( n4192 & n12361 ) | ( ~n8882 & n12361 ) ;
  assign n21080 = ( n4170 & n6827 ) | ( n4170 & ~n21079 ) | ( n6827 & ~n21079 ) ;
  assign n21081 = ( n793 & ~n12387 ) | ( n793 & n21080 ) | ( ~n12387 & n21080 ) ;
  assign n21082 = n8771 ^ n7182 ^ n5108 ;
  assign n21083 = n3471 & ~n10998 ;
  assign n21084 = n5186 & n13577 ;
  assign n21085 = n8928 & n21084 ;
  assign n21086 = ( ~n604 & n6151 ) | ( ~n604 & n21085 ) | ( n6151 & n21085 ) ;
  assign n21087 = ~x42 & n21086 ;
  assign n21088 = n10201 & ~n11690 ;
  assign n21089 = ( n21083 & n21087 ) | ( n21083 & n21088 ) | ( n21087 & n21088 ) ;
  assign n21090 = ~n2309 & n9264 ;
  assign n21091 = n21090 ^ x208 ^ 1'b0 ;
  assign n21092 = ~n13543 & n21091 ;
  assign n21093 = n20672 ^ n8195 ^ 1'b0 ;
  assign n21094 = n19462 & n21093 ;
  assign n21095 = n6509 & n7735 ;
  assign n21096 = n18094 & n21095 ;
  assign n21097 = n21096 ^ n10547 ^ n4050 ;
  assign n21098 = ( n2615 & ~n18820 ) | ( n2615 & n20762 ) | ( ~n18820 & n20762 ) ;
  assign n21099 = n1412 & n3161 ;
  assign n21100 = n21099 ^ n14089 ^ n3920 ;
  assign n21101 = n3397 ^ n456 ^ 1'b0 ;
  assign n21102 = ~n9892 & n17641 ;
  assign n21103 = ~n21101 & n21102 ;
  assign n21109 = n14120 ^ n3368 ^ n858 ;
  assign n21110 = ( n10333 & n14037 ) | ( n10333 & n15421 ) | ( n14037 & n15421 ) ;
  assign n21111 = ( n7898 & n21109 ) | ( n7898 & n21110 ) | ( n21109 & n21110 ) ;
  assign n21112 = n11171 & n16397 ;
  assign n21113 = n21112 ^ n5445 ^ 1'b0 ;
  assign n21114 = n883 & n1814 ;
  assign n21115 = n3167 & n21114 ;
  assign n21116 = ( n6397 & ~n6915 ) | ( n6397 & n21115 ) | ( ~n6915 & n21115 ) ;
  assign n21117 = ( n21111 & n21113 ) | ( n21111 & n21116 ) | ( n21113 & n21116 ) ;
  assign n21104 = ( n2003 & ~n12746 ) | ( n2003 & n20294 ) | ( ~n12746 & n20294 ) ;
  assign n21105 = x159 | n15102 ;
  assign n21106 = n21105 ^ n8981 ^ n4677 ;
  assign n21107 = n8769 | n21106 ;
  assign n21108 = ( n15545 & ~n21104 ) | ( n15545 & n21107 ) | ( ~n21104 & n21107 ) ;
  assign n21118 = n21117 ^ n21108 ^ 1'b0 ;
  assign n21119 = ~n2202 & n9039 ;
  assign n21120 = ( n13279 & n16885 ) | ( n13279 & ~n21119 ) | ( n16885 & ~n21119 ) ;
  assign n21121 = n21120 ^ n3539 ^ 1'b0 ;
  assign n21122 = n21118 | n21121 ;
  assign n21123 = n11379 ^ n6783 ^ 1'b0 ;
  assign n21124 = ( ~n15694 & n17821 ) | ( ~n15694 & n21123 ) | ( n17821 & n21123 ) ;
  assign n21125 = n14252 ^ n7671 ^ 1'b0 ;
  assign n21126 = ( ~n9019 & n11948 ) | ( ~n9019 & n15047 ) | ( n11948 & n15047 ) ;
  assign n21127 = ( x65 & n20679 ) | ( x65 & n21126 ) | ( n20679 & n21126 ) ;
  assign n21128 = n17458 ^ n3921 ^ n666 ;
  assign n21129 = n21128 ^ n18602 ^ 1'b0 ;
  assign n21130 = n15030 | n21129 ;
  assign n21131 = n21130 ^ n16669 ^ 1'b0 ;
  assign n21132 = ( n5362 & n14881 ) | ( n5362 & n16728 ) | ( n14881 & n16728 ) ;
  assign n21133 = ~n3505 & n16209 ;
  assign n21134 = ~n4110 & n21133 ;
  assign n21135 = n14003 & ~n21134 ;
  assign n21136 = ~n15976 & n21135 ;
  assign n21137 = n18895 ^ n9340 ^ n5583 ;
  assign n21138 = n10725 ^ n7101 ^ 1'b0 ;
  assign n21139 = n15311 & ~n21138 ;
  assign n21143 = n21002 ^ n2333 ^ n1472 ;
  assign n21140 = n7508 & n17045 ;
  assign n21141 = ~n16491 & n21140 ;
  assign n21142 = ~n7699 & n21141 ;
  assign n21144 = n21143 ^ n21142 ^ 1'b0 ;
  assign n21145 = n21139 & n21144 ;
  assign n21146 = ~n21137 & n21145 ;
  assign n21147 = n21146 ^ n8844 ^ 1'b0 ;
  assign n21150 = n6294 & ~n12563 ;
  assign n21151 = ( n13836 & n16355 ) | ( n13836 & ~n21150 ) | ( n16355 & ~n21150 ) ;
  assign n21148 = n11526 ^ n10302 ^ 1'b0 ;
  assign n21149 = ( n5532 & n14485 ) | ( n5532 & n21148 ) | ( n14485 & n21148 ) ;
  assign n21152 = n21151 ^ n21149 ^ n10457 ;
  assign n21153 = n11548 ^ n8720 ^ n6200 ;
  assign n21154 = ( n5804 & ~n13066 ) | ( n5804 & n15347 ) | ( ~n13066 & n15347 ) ;
  assign n21155 = n21154 ^ n5152 ^ 1'b0 ;
  assign n21158 = n11760 ^ n5904 ^ n5529 ;
  assign n21156 = n8421 | n10397 ;
  assign n21157 = n21156 ^ n13298 ^ 1'b0 ;
  assign n21159 = n21158 ^ n21157 ^ n12202 ;
  assign n21172 = ( ~x88 & n798 ) | ( ~x88 & n5199 ) | ( n798 & n5199 ) ;
  assign n21173 = n4485 | n21172 ;
  assign n21174 = n21173 ^ n14594 ^ 1'b0 ;
  assign n21162 = n3659 ^ n1237 ^ 1'b0 ;
  assign n21163 = n6911 & n21162 ;
  assign n21160 = n17733 ^ n14473 ^ n9439 ;
  assign n21161 = n3719 & ~n21160 ;
  assign n21164 = n21163 ^ n21161 ^ 1'b0 ;
  assign n21165 = n17968 ^ n9179 ^ n1953 ;
  assign n21168 = n10550 ^ n5227 ^ n357 ;
  assign n21166 = n5797 ^ n3255 ^ 1'b0 ;
  assign n21167 = ~x227 & n21166 ;
  assign n21169 = n21168 ^ n21167 ^ n4197 ;
  assign n21170 = n9093 & n21169 ;
  assign n21171 = ( n21164 & ~n21165 ) | ( n21164 & n21170 ) | ( ~n21165 & n21170 ) ;
  assign n21175 = n21174 ^ n21171 ^ 1'b0 ;
  assign n21176 = ( ~n17458 & n21159 ) | ( ~n17458 & n21175 ) | ( n21159 & n21175 ) ;
  assign n21177 = n5067 | n11236 ;
  assign n21178 = ( n13228 & n14929 ) | ( n13228 & n21177 ) | ( n14929 & n21177 ) ;
  assign n21179 = n21178 ^ n18793 ^ n15902 ;
  assign n21180 = n13426 ^ n6524 ^ n1719 ;
  assign n21181 = ( ~n9174 & n12689 ) | ( ~n9174 & n16646 ) | ( n12689 & n16646 ) ;
  assign n21182 = ( n903 & n11332 ) | ( n903 & ~n21181 ) | ( n11332 & ~n21181 ) ;
  assign n21183 = n14284 ^ n8104 ^ n1753 ;
  assign n21184 = n21183 ^ n15007 ^ x164 ;
  assign n21185 = n15660 ^ n2116 ^ n1238 ;
  assign n21186 = ( n14699 & ~n19552 ) | ( n14699 & n21185 ) | ( ~n19552 & n21185 ) ;
  assign n21187 = ( ~n7488 & n16592 ) | ( ~n7488 & n21186 ) | ( n16592 & n21186 ) ;
  assign n21188 = ( ~n21025 & n21184 ) | ( ~n21025 & n21187 ) | ( n21184 & n21187 ) ;
  assign n21189 = ( x40 & n3727 ) | ( x40 & ~n5942 ) | ( n3727 & ~n5942 ) ;
  assign n21190 = n19573 ^ n5307 ^ 1'b0 ;
  assign n21191 = ( n18778 & n21189 ) | ( n18778 & n21190 ) | ( n21189 & n21190 ) ;
  assign n21192 = ( n12300 & n21188 ) | ( n12300 & n21191 ) | ( n21188 & n21191 ) ;
  assign n21193 = n6736 ^ n1285 ^ n328 ;
  assign n21196 = ( n15071 & n20355 ) | ( n15071 & n20669 ) | ( n20355 & n20669 ) ;
  assign n21194 = n16326 ^ n6760 ^ n6047 ;
  assign n21195 = n5515 & ~n21194 ;
  assign n21197 = n21196 ^ n21195 ^ 1'b0 ;
  assign n21198 = n644 & n6585 ;
  assign n21199 = ( x13 & ~n14246 ) | ( x13 & n19216 ) | ( ~n14246 & n19216 ) ;
  assign n21200 = ( n3878 & n4362 ) | ( n3878 & ~n4922 ) | ( n4362 & ~n4922 ) ;
  assign n21201 = ( n10875 & n21199 ) | ( n10875 & ~n21200 ) | ( n21199 & ~n21200 ) ;
  assign n21202 = ( n4514 & ~n21198 ) | ( n4514 & n21201 ) | ( ~n21198 & n21201 ) ;
  assign n21203 = n3641 & ~n17801 ;
  assign n21204 = n21203 ^ n1576 ^ 1'b0 ;
  assign n21205 = n17950 & ~n21204 ;
  assign n21206 = n21205 ^ n18188 ^ 1'b0 ;
  assign n21207 = ~n12519 & n21206 ;
  assign n21211 = n17481 ^ n11837 ^ 1'b0 ;
  assign n21212 = n16898 | n21211 ;
  assign n21208 = n20231 ^ n12570 ^ n8997 ;
  assign n21209 = ( n5877 & n18751 ) | ( n5877 & n21208 ) | ( n18751 & n21208 ) ;
  assign n21210 = ~n325 & n21209 ;
  assign n21213 = n21212 ^ n21210 ^ 1'b0 ;
  assign n21214 = n5664 & n12264 ;
  assign n21215 = n15341 & n21214 ;
  assign n21216 = n10766 ^ n8261 ^ n636 ;
  assign n21217 = ( n2331 & ~n7662 ) | ( n2331 & n21216 ) | ( ~n7662 & n21216 ) ;
  assign n21218 = n1875 | n2186 ;
  assign n21219 = n7534 & ~n21218 ;
  assign n21220 = ( n12560 & n17520 ) | ( n12560 & ~n21219 ) | ( n17520 & ~n21219 ) ;
  assign n21221 = ( ~n14883 & n21217 ) | ( ~n14883 & n21220 ) | ( n21217 & n21220 ) ;
  assign n21222 = n5293 | n7601 ;
  assign n21223 = x92 | n21222 ;
  assign n21224 = n21223 ^ n12368 ^ n11707 ;
  assign n21231 = n11479 & n19446 ;
  assign n21232 = n21231 ^ n20466 ^ 1'b0 ;
  assign n21233 = n17127 & n21232 ;
  assign n21225 = n12249 ^ n7349 ^ n6935 ;
  assign n21226 = n21225 ^ n7443 ^ n4247 ;
  assign n21227 = ( n2953 & ~n3908 ) | ( n2953 & n16486 ) | ( ~n3908 & n16486 ) ;
  assign n21228 = n21227 ^ n17946 ^ n4124 ;
  assign n21229 = n21226 & n21228 ;
  assign n21230 = n15028 & ~n21229 ;
  assign n21234 = n21233 ^ n21230 ^ 1'b0 ;
  assign n21236 = n7738 ^ n4689 ^ x67 ;
  assign n21235 = ( n3016 & n4299 ) | ( n3016 & ~n19109 ) | ( n4299 & ~n19109 ) ;
  assign n21237 = n21236 ^ n21235 ^ n440 ;
  assign n21238 = ( ~n2943 & n3509 ) | ( ~n2943 & n5834 ) | ( n3509 & n5834 ) ;
  assign n21239 = ( ~n2319 & n11678 ) | ( ~n2319 & n21238 ) | ( n11678 & n21238 ) ;
  assign n21240 = n16284 & ~n21239 ;
  assign n21241 = ~n21237 & n21240 ;
  assign n21242 = ( n1875 & ~n2442 ) | ( n1875 & n10439 ) | ( ~n2442 & n10439 ) ;
  assign n21243 = ( ~n8110 & n14328 ) | ( ~n8110 & n21242 ) | ( n14328 & n21242 ) ;
  assign n21244 = ( n4570 & n10775 ) | ( n4570 & ~n21243 ) | ( n10775 & ~n21243 ) ;
  assign n21255 = n19953 ^ n17430 ^ n2357 ;
  assign n21252 = n11564 ^ n4026 ^ n1499 ;
  assign n21253 = ( n15067 & n16028 ) | ( n15067 & n21252 ) | ( n16028 & n21252 ) ;
  assign n21254 = ( ~n5740 & n15109 ) | ( ~n5740 & n21253 ) | ( n15109 & n21253 ) ;
  assign n21256 = n21255 ^ n21254 ^ 1'b0 ;
  assign n21257 = n19108 | n21256 ;
  assign n21248 = ( x128 & n3009 ) | ( x128 & ~n6200 ) | ( n3009 & ~n6200 ) ;
  assign n21249 = ( n10722 & n19511 ) | ( n10722 & ~n21248 ) | ( n19511 & ~n21248 ) ;
  assign n21245 = n13564 ^ n4815 ^ 1'b0 ;
  assign n21246 = n21245 ^ n12564 ^ 1'b0 ;
  assign n21247 = n21246 ^ n15047 ^ n5017 ;
  assign n21250 = n21249 ^ n21247 ^ 1'b0 ;
  assign n21251 = n19921 & ~n21250 ;
  assign n21258 = n21257 ^ n21251 ^ n6345 ;
  assign n21263 = n3690 ^ n2961 ^ n321 ;
  assign n21264 = n6567 & n15071 ;
  assign n21265 = ( n503 & ~n21263 ) | ( n503 & n21264 ) | ( ~n21263 & n21264 ) ;
  assign n21260 = x160 & ~n2539 ;
  assign n21261 = ~n9069 & n21260 ;
  assign n21259 = n13611 ^ n3240 ^ 1'b0 ;
  assign n21262 = n21261 ^ n21259 ^ n13867 ;
  assign n21266 = n21265 ^ n21262 ^ 1'b0 ;
  assign n21267 = n13657 ^ n6523 ^ 1'b0 ;
  assign n21268 = n16856 ^ n7196 ^ n2275 ;
  assign n21269 = ( n1097 & ~n9244 ) | ( n1097 & n10495 ) | ( ~n9244 & n10495 ) ;
  assign n21270 = ( n17118 & ~n21268 ) | ( n17118 & n21269 ) | ( ~n21268 & n21269 ) ;
  assign n21271 = n18642 ^ n12497 ^ n6435 ;
  assign n21272 = n13999 | n21271 ;
  assign n21273 = ~n10618 & n19793 ;
  assign n21274 = n19393 & n21273 ;
  assign n21275 = n21272 & ~n21274 ;
  assign n21276 = n21275 ^ n3948 ^ 1'b0 ;
  assign n21277 = n7100 ^ n2019 ^ 1'b0 ;
  assign n21278 = n21277 ^ n12813 ^ 1'b0 ;
  assign n21279 = n21278 ^ n11718 ^ n9613 ;
  assign n21280 = n17715 ^ n3895 ^ 1'b0 ;
  assign n21282 = ( n6310 & n6942 ) | ( n6310 & n18051 ) | ( n6942 & n18051 ) ;
  assign n21283 = ( n9988 & n21199 ) | ( n9988 & ~n21282 ) | ( n21199 & ~n21282 ) ;
  assign n21281 = ( n7686 & n9878 ) | ( n7686 & ~n11059 ) | ( n9878 & ~n11059 ) ;
  assign n21284 = n21283 ^ n21281 ^ 1'b0 ;
  assign n21285 = n14098 | n21284 ;
  assign n21286 = n18172 | n18697 ;
  assign n21287 = n21286 ^ n9187 ^ 1'b0 ;
  assign n21292 = n15259 ^ n8199 ^ n882 ;
  assign n21288 = n2722 & ~n13461 ;
  assign n21289 = n21288 ^ n1287 ^ 1'b0 ;
  assign n21290 = n21289 ^ n19248 ^ n10767 ;
  assign n21291 = n21290 ^ n16266 ^ n5893 ;
  assign n21293 = n21292 ^ n21291 ^ n8187 ;
  assign n21294 = n17864 ^ n16961 ^ n15517 ;
  assign n21295 = n18751 ^ n7373 ^ n1909 ;
  assign n21296 = ~n5944 & n8386 ;
  assign n21297 = n2265 & n21296 ;
  assign n21298 = n6617 ^ n1813 ^ n375 ;
  assign n21299 = n11127 ^ n2871 ^ 1'b0 ;
  assign n21300 = n21298 & n21299 ;
  assign n21301 = ~n11061 & n21300 ;
  assign n21302 = ~n16809 & n21301 ;
  assign n21303 = n13830 ^ n1449 ^ n397 ;
  assign n21304 = n21303 ^ n2477 ^ n530 ;
  assign n21305 = n21304 ^ n4124 ^ 1'b0 ;
  assign n21306 = n18044 ^ n14777 ^ n10523 ;
  assign n21307 = n2213 ^ n430 ^ 1'b0 ;
  assign n21308 = n21306 | n21307 ;
  assign n21309 = ( ~n9169 & n9677 ) | ( ~n9169 & n21308 ) | ( n9677 & n21308 ) ;
  assign n21310 = n21309 ^ n12249 ^ n8909 ;
  assign n21311 = n21310 ^ n14304 ^ n13408 ;
  assign n21312 = n275 & ~n10466 ;
  assign n21313 = n21312 ^ n3829 ^ 1'b0 ;
  assign n21314 = n21313 ^ n8790 ^ n7311 ;
  assign n21315 = n7311 ^ n7220 ^ 1'b0 ;
  assign n21316 = n1256 & ~n21315 ;
  assign n21317 = n21316 ^ n19452 ^ n1911 ;
  assign n21318 = ( n2971 & n3092 ) | ( n2971 & ~n3643 ) | ( n3092 & ~n3643 ) ;
  assign n21319 = n21318 ^ n18190 ^ n12503 ;
  assign n21320 = n15284 ^ n8551 ^ 1'b0 ;
  assign n21321 = n18322 ^ n7072 ^ n1903 ;
  assign n21322 = n21321 ^ n3997 ^ n1768 ;
  assign n21323 = ( x79 & n8691 ) | ( x79 & n21322 ) | ( n8691 & n21322 ) ;
  assign n21324 = n21323 ^ n6379 ^ 1'b0 ;
  assign n21325 = ~n21320 & n21324 ;
  assign n21326 = ~n21319 & n21325 ;
  assign n21327 = ( ~x125 & n723 ) | ( ~x125 & n2247 ) | ( n723 & n2247 ) ;
  assign n21328 = ( n10130 & ~n11780 ) | ( n10130 & n21327 ) | ( ~n11780 & n21327 ) ;
  assign n21329 = ( n15959 & ~n20399 ) | ( n15959 & n21328 ) | ( ~n20399 & n21328 ) ;
  assign n21330 = n21329 ^ n7890 ^ x109 ;
  assign n21331 = ( ~n932 & n6261 ) | ( ~n932 & n13421 ) | ( n6261 & n13421 ) ;
  assign n21332 = n18947 ^ n10897 ^ n9000 ;
  assign n21333 = n21332 ^ n11307 ^ n4950 ;
  assign n21334 = n19210 ^ n10506 ^ n1593 ;
  assign n21335 = ( n3952 & ~n21333 ) | ( n3952 & n21334 ) | ( ~n21333 & n21334 ) ;
  assign n21336 = n5832 & n8557 ;
  assign n21337 = n21336 ^ n12603 ^ 1'b0 ;
  assign n21338 = n1961 | n21337 ;
  assign n21339 = x231 & ~n21338 ;
  assign n21340 = ~x20 & n21339 ;
  assign n21341 = n4333 ^ n2273 ^ 1'b0 ;
  assign n21342 = ~n14932 & n21341 ;
  assign n21343 = n21342 ^ n12804 ^ n2280 ;
  assign n21344 = ~n10779 & n11055 ;
  assign n21345 = n21344 ^ n15298 ^ 1'b0 ;
  assign n21346 = n13890 ^ n9592 ^ n708 ;
  assign n21347 = ( ~n5786 & n21345 ) | ( ~n5786 & n21346 ) | ( n21345 & n21346 ) ;
  assign n21348 = ( ~x196 & n6521 ) | ( ~x196 & n7888 ) | ( n6521 & n7888 ) ;
  assign n21349 = n21348 ^ n12931 ^ 1'b0 ;
  assign n21350 = n12084 ^ n4371 ^ n2839 ;
  assign n21351 = n21350 ^ n12308 ^ n7375 ;
  assign n21352 = n21351 ^ n16820 ^ 1'b0 ;
  assign n21357 = n13955 ^ n9583 ^ n7766 ;
  assign n21355 = ( ~n5882 & n7886 ) | ( ~n5882 & n19271 ) | ( n7886 & n19271 ) ;
  assign n21356 = n21355 ^ n9150 ^ n2468 ;
  assign n21353 = n3962 | n5923 ;
  assign n21354 = n13394 & ~n21353 ;
  assign n21358 = n21357 ^ n21356 ^ n21354 ;
  assign n21359 = ( n5229 & n6531 ) | ( n5229 & ~n10148 ) | ( n6531 & ~n10148 ) ;
  assign n21360 = n21359 ^ n12900 ^ n12430 ;
  assign n21361 = n21360 ^ n13705 ^ 1'b0 ;
  assign n21362 = n3583 & ~n21361 ;
  assign n21363 = n7954 & n10312 ;
  assign n21364 = n21363 ^ n7489 ^ 1'b0 ;
  assign n21365 = n11334 ^ n2697 ^ x22 ;
  assign n21366 = n21365 ^ n17339 ^ 1'b0 ;
  assign n21367 = n6151 & ~n21366 ;
  assign n21368 = n12102 & n21031 ;
  assign n21369 = ( n2084 & n19969 ) | ( n2084 & ~n21368 ) | ( n19969 & ~n21368 ) ;
  assign n21370 = ( n7322 & ~n21367 ) | ( n7322 & n21369 ) | ( ~n21367 & n21369 ) ;
  assign n21371 = n19936 ^ n17479 ^ n4396 ;
  assign n21372 = ( n3606 & ~n7741 ) | ( n3606 & n12920 ) | ( ~n7741 & n12920 ) ;
  assign n21373 = n21372 ^ n17074 ^ n11905 ;
  assign n21374 = ( n12454 & n21371 ) | ( n12454 & ~n21373 ) | ( n21371 & ~n21373 ) ;
  assign n21375 = n9480 & ~n12192 ;
  assign n21376 = n15392 ^ n8494 ^ n5418 ;
  assign n21377 = n7452 ^ n3208 ^ 1'b0 ;
  assign n21378 = ( ~n2795 & n21376 ) | ( ~n2795 & n21377 ) | ( n21376 & n21377 ) ;
  assign n21379 = n14528 ^ n12000 ^ n11913 ;
  assign n21381 = n7971 & n9972 ;
  assign n21380 = n14549 ^ n9226 ^ n8839 ;
  assign n21382 = n21381 ^ n21380 ^ n5990 ;
  assign n21383 = ( n6992 & n17666 ) | ( n6992 & ~n21382 ) | ( n17666 & ~n21382 ) ;
  assign n21384 = ~n12117 & n21383 ;
  assign n21386 = n15983 ^ n7798 ^ n1500 ;
  assign n21385 = ~n8930 & n10603 ;
  assign n21387 = n21386 ^ n21385 ^ 1'b0 ;
  assign n21388 = n9600 ^ n8562 ^ n4555 ;
  assign n21389 = ( n1354 & n10128 ) | ( n1354 & ~n21388 ) | ( n10128 & ~n21388 ) ;
  assign n21390 = ( n5748 & ~n19989 ) | ( n5748 & n21389 ) | ( ~n19989 & n21389 ) ;
  assign n21391 = ( ~n2519 & n3548 ) | ( ~n2519 & n20773 ) | ( n3548 & n20773 ) ;
  assign n21392 = ( n9958 & n19800 ) | ( n9958 & ~n19882 ) | ( n19800 & ~n19882 ) ;
  assign n21394 = n1948 & ~n19599 ;
  assign n21395 = n21394 ^ n13285 ^ 1'b0 ;
  assign n21393 = ~n4299 & n5324 ;
  assign n21396 = n21395 ^ n21393 ^ 1'b0 ;
  assign n21397 = ~n12238 & n14736 ;
  assign n21398 = ~n15333 & n21397 ;
  assign n21399 = n10840 & ~n21398 ;
  assign n21400 = n15362 ^ n5920 ^ 1'b0 ;
  assign n21401 = ~n2594 & n2607 ;
  assign n21402 = n16801 & n21401 ;
  assign n21403 = n18795 | n21402 ;
  assign n21404 = n21403 ^ n4848 ^ 1'b0 ;
  assign n21405 = n7271 & n8992 ;
  assign n21406 = ( n1518 & n19949 ) | ( n1518 & n21405 ) | ( n19949 & n21405 ) ;
  assign n21407 = ( n2735 & ~n20041 ) | ( n2735 & n21406 ) | ( ~n20041 & n21406 ) ;
  assign n21408 = n21407 ^ n17487 ^ n8997 ;
  assign n21409 = n13615 & ~n15721 ;
  assign n21410 = ~x22 & n1614 ;
  assign n21411 = ( n956 & n4404 ) | ( n956 & ~n4608 ) | ( n4404 & ~n4608 ) ;
  assign n21412 = n21410 & ~n21411 ;
  assign n21413 = n14055 & ~n16138 ;
  assign n21414 = ( n2607 & n3784 ) | ( n2607 & n12569 ) | ( n3784 & n12569 ) ;
  assign n21415 = n21414 ^ n8716 ^ 1'b0 ;
  assign n21416 = n16321 ^ n15689 ^ 1'b0 ;
  assign n21417 = n13481 & n21416 ;
  assign n21420 = n13731 ^ n4428 ^ n1769 ;
  assign n21418 = n3575 & n3981 ;
  assign n21419 = ~n6327 & n21418 ;
  assign n21421 = n21420 ^ n21419 ^ 1'b0 ;
  assign n21422 = ~n17323 & n21421 ;
  assign n21423 = ( n606 & ~n1686 ) | ( n606 & n3950 ) | ( ~n1686 & n3950 ) ;
  assign n21424 = n4526 & n21423 ;
  assign n21425 = n21424 ^ n7910 ^ 1'b0 ;
  assign n21426 = ( n7667 & n14533 ) | ( n7667 & ~n21425 ) | ( n14533 & ~n21425 ) ;
  assign n21427 = n10676 | n21426 ;
  assign n21428 = n9030 ^ n7123 ^ n6495 ;
  assign n21429 = n19642 ^ n8674 ^ 1'b0 ;
  assign n21430 = n21429 ^ n19224 ^ 1'b0 ;
  assign n21431 = n21430 ^ n16408 ^ n5260 ;
  assign n21432 = x55 & n669 ;
  assign n21433 = n8223 & n21432 ;
  assign n21434 = ~n7148 & n15291 ;
  assign n21435 = ~n2454 & n21434 ;
  assign n21436 = n16227 & n21435 ;
  assign n21437 = n19590 ^ n11159 ^ n6990 ;
  assign n21439 = x55 & n3793 ;
  assign n21440 = ~n2248 & n21439 ;
  assign n21438 = n7004 & ~n8193 ;
  assign n21441 = n21440 ^ n21438 ^ 1'b0 ;
  assign n21442 = n11147 ^ n6068 ^ n561 ;
  assign n21443 = n19658 ^ n9822 ^ n4627 ;
  assign n21444 = n21442 & n21443 ;
  assign n21445 = n480 & ~n21444 ;
  assign n21446 = n14222 ^ n9746 ^ n1267 ;
  assign n21447 = n3626 ^ n938 ^ 1'b0 ;
  assign n21448 = n846 & n5037 ;
  assign n21449 = n21448 ^ n5324 ^ 1'b0 ;
  assign n21450 = ( ~n6642 & n14601 ) | ( ~n6642 & n21449 ) | ( n14601 & n21449 ) ;
  assign n21451 = n21450 ^ n2294 ^ 1'b0 ;
  assign n21452 = ( n4955 & n21447 ) | ( n4955 & n21451 ) | ( n21447 & n21451 ) ;
  assign n21453 = ( n2192 & n14502 ) | ( n2192 & ~n21452 ) | ( n14502 & ~n21452 ) ;
  assign n21454 = n21453 ^ n11306 ^ n8389 ;
  assign n21455 = n9949 ^ n5526 ^ 1'b0 ;
  assign n21456 = n10248 & ~n21455 ;
  assign n21457 = n15424 ^ n9186 ^ 1'b0 ;
  assign n21458 = n21457 ^ n12063 ^ n4503 ;
  assign n21459 = ( n14586 & n21456 ) | ( n14586 & ~n21458 ) | ( n21456 & ~n21458 ) ;
  assign n21460 = ~x146 & n15412 ;
  assign n21461 = n1491 & n21460 ;
  assign n21462 = n1271 & n21461 ;
  assign n21463 = ~n12118 & n21462 ;
  assign n21464 = n17420 ^ n10974 ^ n8182 ;
  assign n21465 = n18527 ^ n8139 ^ 1'b0 ;
  assign n21466 = n9239 ^ n8632 ^ n2206 ;
  assign n21467 = n21466 ^ n4995 ^ n1050 ;
  assign n21468 = ( x37 & ~n9919 ) | ( x37 & n21467 ) | ( ~n9919 & n21467 ) ;
  assign n21469 = n18973 ^ n12707 ^ n8434 ;
  assign n21470 = ( ~n8419 & n10246 ) | ( ~n8419 & n21469 ) | ( n10246 & n21469 ) ;
  assign n21471 = n11620 ^ n4181 ^ 1'b0 ;
  assign n21472 = ( ~n482 & n2342 ) | ( ~n482 & n21471 ) | ( n2342 & n21471 ) ;
  assign n21473 = n14630 ^ n8233 ^ 1'b0 ;
  assign n21474 = ( n6062 & ~n7721 ) | ( n6062 & n13494 ) | ( ~n7721 & n13494 ) ;
  assign n21475 = ( ~n10945 & n11160 ) | ( ~n10945 & n21474 ) | ( n11160 & n21474 ) ;
  assign n21476 = ( ~n2526 & n21473 ) | ( ~n2526 & n21475 ) | ( n21473 & n21475 ) ;
  assign n21477 = n5520 ^ n3390 ^ x120 ;
  assign n21478 = n13347 ^ n662 ^ 1'b0 ;
  assign n21479 = n7285 & ~n21478 ;
  assign n21480 = n9807 & n21479 ;
  assign n21481 = n21477 & n21480 ;
  assign n21482 = n16250 ^ n9903 ^ n4888 ;
  assign n21483 = ( n3210 & n8272 ) | ( n3210 & n19029 ) | ( n8272 & n19029 ) ;
  assign n21484 = n13498 ^ n10248 ^ 1'b0 ;
  assign n21485 = ~n21483 & n21484 ;
  assign n21486 = n20353 ^ n9971 ^ 1'b0 ;
  assign n21487 = ~n13556 & n21486 ;
  assign n21488 = ( n21482 & n21485 ) | ( n21482 & n21487 ) | ( n21485 & n21487 ) ;
  assign n21489 = ( n9049 & n20637 ) | ( n9049 & n21488 ) | ( n20637 & n21488 ) ;
  assign n21490 = n4748 & n21489 ;
  assign n21491 = n6992 ^ n2849 ^ n1714 ;
  assign n21492 = n21491 ^ n9951 ^ 1'b0 ;
  assign n21493 = ~n21490 & n21492 ;
  assign n21494 = n9032 ^ n7296 ^ n7029 ;
  assign n21495 = n21494 ^ n2677 ^ 1'b0 ;
  assign n21496 = n21495 ^ n19585 ^ n12625 ;
  assign n21497 = n11797 ^ n6079 ^ n4136 ;
  assign n21498 = ( n15856 & ~n16091 ) | ( n15856 & n21497 ) | ( ~n16091 & n21497 ) ;
  assign n21499 = n21498 ^ n3368 ^ 1'b0 ;
  assign n21500 = n9603 ^ n3561 ^ 1'b0 ;
  assign n21501 = ( n6531 & n11171 ) | ( n6531 & ~n21500 ) | ( n11171 & ~n21500 ) ;
  assign n21502 = n13598 ^ n3782 ^ 1'b0 ;
  assign n21503 = n5119 & n21502 ;
  assign n21504 = ( n6638 & ~n10986 ) | ( n6638 & n21503 ) | ( ~n10986 & n21503 ) ;
  assign n21505 = n1293 | n2222 ;
  assign n21506 = n21505 ^ n7299 ^ 1'b0 ;
  assign n21507 = n21506 ^ n20229 ^ n1574 ;
  assign n21508 = n17188 ^ n13821 ^ n326 ;
  assign n21509 = n21508 ^ n15207 ^ n13878 ;
  assign n21510 = ( ~n5981 & n9327 ) | ( ~n5981 & n14172 ) | ( n9327 & n14172 ) ;
  assign n21511 = ( ~n3102 & n10974 ) | ( ~n3102 & n21031 ) | ( n10974 & n21031 ) ;
  assign n21512 = ( n5662 & n5887 ) | ( n5662 & n21511 ) | ( n5887 & n21511 ) ;
  assign n21513 = n21510 & ~n21512 ;
  assign n21514 = n3247 | n14960 ;
  assign n21515 = ( n2953 & n3681 ) | ( n2953 & ~n13779 ) | ( n3681 & ~n13779 ) ;
  assign n21516 = n2742 & ~n4825 ;
  assign n21517 = n1405 & n21516 ;
  assign n21518 = n10164 ^ n1768 ^ x149 ;
  assign n21519 = n21518 ^ n19614 ^ n12114 ;
  assign n21520 = ~n3241 & n7375 ;
  assign n21521 = ( x170 & n1894 ) | ( x170 & n10314 ) | ( n1894 & n10314 ) ;
  assign n21522 = ~n15388 & n19937 ;
  assign n21523 = n12889 ^ n6702 ^ n1144 ;
  assign n21524 = n12230 ^ n6117 ^ 1'b0 ;
  assign n21525 = n13674 | n21524 ;
  assign n21526 = n21525 ^ n10112 ^ n3534 ;
  assign n21527 = ( ~n13422 & n21523 ) | ( ~n13422 & n21526 ) | ( n21523 & n21526 ) ;
  assign n21528 = n463 | n1886 ;
  assign n21529 = n13384 ^ n11468 ^ n5558 ;
  assign n21530 = n21529 ^ n10930 ^ n10661 ;
  assign n21531 = ( ~n1101 & n21328 ) | ( ~n1101 & n21530 ) | ( n21328 & n21530 ) ;
  assign n21539 = n9295 ^ n6942 ^ n3050 ;
  assign n21532 = n8895 ^ n5058 ^ n2239 ;
  assign n21533 = n5358 ^ n616 ^ x42 ;
  assign n21534 = n21533 ^ n19684 ^ 1'b0 ;
  assign n21535 = ( n6488 & n18001 ) | ( n6488 & n21534 ) | ( n18001 & n21534 ) ;
  assign n21536 = n21532 | n21535 ;
  assign n21537 = n21536 ^ n4888 ^ 1'b0 ;
  assign n21538 = ~n12024 & n21537 ;
  assign n21540 = n21539 ^ n21538 ^ n16604 ;
  assign n21541 = n12170 | n21540 ;
  assign n21542 = n21541 ^ n4277 ^ x140 ;
  assign n21543 = ( n1970 & ~n8799 ) | ( n1970 & n10733 ) | ( ~n8799 & n10733 ) ;
  assign n21544 = ( n12409 & ~n18020 ) | ( n12409 & n21543 ) | ( ~n18020 & n21543 ) ;
  assign n21545 = n4530 & ~n10065 ;
  assign n21546 = n14334 & ~n21545 ;
  assign n21547 = n21546 ^ n18053 ^ n16405 ;
  assign n21548 = n8124 ^ n7120 ^ n6935 ;
  assign n21549 = n9514 ^ n6700 ^ n859 ;
  assign n21550 = n21549 ^ x175 ^ 1'b0 ;
  assign n21551 = ( n9020 & n18689 ) | ( n9020 & n21550 ) | ( n18689 & n21550 ) ;
  assign n21552 = ( n10604 & n14139 ) | ( n10604 & ~n17476 ) | ( n14139 & ~n17476 ) ;
  assign n21553 = ( n6774 & ~n9487 ) | ( n6774 & n21552 ) | ( ~n9487 & n21552 ) ;
  assign n21554 = ( n13382 & n13511 ) | ( n13382 & ~n21553 ) | ( n13511 & ~n21553 ) ;
  assign n21555 = n8538 ^ n4422 ^ 1'b0 ;
  assign n21556 = ~n10740 & n21555 ;
  assign n21557 = n1355 | n5943 ;
  assign n21558 = n6184 | n21557 ;
  assign n21559 = ( n4025 & n4271 ) | ( n4025 & n21558 ) | ( n4271 & n21558 ) ;
  assign n21560 = n20598 ^ n3990 ^ 1'b0 ;
  assign n21561 = ~n21559 & n21560 ;
  assign n21562 = n16742 ^ n12237 ^ 1'b0 ;
  assign n21563 = ~n14755 & n21562 ;
  assign n21564 = n21563 ^ n9408 ^ 1'b0 ;
  assign n21565 = n317 | n2835 ;
  assign n21566 = n18097 & n21565 ;
  assign n21567 = ~n8422 & n21566 ;
  assign n21568 = n449 | n1486 ;
  assign n21569 = n1752 | n21568 ;
  assign n21570 = n21569 ^ n13217 ^ 1'b0 ;
  assign n21571 = ( ~n8455 & n12912 ) | ( ~n8455 & n15143 ) | ( n12912 & n15143 ) ;
  assign n21572 = ( ~n14958 & n21570 ) | ( ~n14958 & n21571 ) | ( n21570 & n21571 ) ;
  assign n21573 = ( n9057 & n12948 ) | ( n9057 & ~n13345 ) | ( n12948 & ~n13345 ) ;
  assign n21574 = n21573 ^ n505 ^ 1'b0 ;
  assign n21576 = n4926 | n6268 ;
  assign n21577 = n21576 ^ n4110 ^ 1'b0 ;
  assign n21575 = ~n18207 & n19190 ;
  assign n21578 = n21577 ^ n21575 ^ 1'b0 ;
  assign n21579 = n8599 ^ n2840 ^ n1283 ;
  assign n21580 = ( n2245 & n11341 ) | ( n2245 & n21579 ) | ( n11341 & n21579 ) ;
  assign n21581 = n5394 | n13291 ;
  assign n21582 = n21581 ^ n9484 ^ 1'b0 ;
  assign n21583 = n21582 ^ n17822 ^ n1670 ;
  assign n21584 = n3025 & n3042 ;
  assign n21585 = n21584 ^ n7875 ^ 1'b0 ;
  assign n21586 = ~n21583 & n21585 ;
  assign n21587 = ( n752 & n6998 ) | ( n752 & n17564 ) | ( n6998 & n17564 ) ;
  assign n21588 = n5664 & n7832 ;
  assign n21589 = n21588 ^ n17974 ^ 1'b0 ;
  assign n21590 = n21589 ^ n11008 ^ n2895 ;
  assign n21591 = ( n18054 & n21587 ) | ( n18054 & n21590 ) | ( n21587 & n21590 ) ;
  assign n21592 = n6875 ^ n5343 ^ n489 ;
  assign n21593 = n7010 | n21592 ;
  assign n21599 = n7600 | n16534 ;
  assign n21600 = n21599 ^ n8393 ^ 1'b0 ;
  assign n21601 = n21600 ^ n15096 ^ n2851 ;
  assign n21594 = n1507 | n2186 ;
  assign n21595 = n18402 | n21594 ;
  assign n21596 = ( n3550 & n9097 ) | ( n3550 & n21595 ) | ( n9097 & n21595 ) ;
  assign n21597 = n21596 ^ n18539 ^ n4235 ;
  assign n21598 = n390 & ~n21597 ;
  assign n21602 = n21601 ^ n21598 ^ 1'b0 ;
  assign n21604 = n4635 ^ n3151 ^ 1'b0 ;
  assign n21603 = ( ~n854 & n10497 ) | ( ~n854 & n15129 ) | ( n10497 & n15129 ) ;
  assign n21605 = n21604 ^ n21603 ^ n15632 ;
  assign n21606 = n20669 ^ n13632 ^ n7907 ;
  assign n21607 = n3048 & n7641 ;
  assign n21608 = n21607 ^ n8411 ^ 1'b0 ;
  assign n21609 = n21608 ^ n11591 ^ n8840 ;
  assign n21610 = n21609 ^ n19776 ^ n9104 ;
  assign n21611 = ( n17882 & ~n21606 ) | ( n17882 & n21610 ) | ( ~n21606 & n21610 ) ;
  assign n21612 = ( x56 & n2705 ) | ( x56 & ~n18281 ) | ( n2705 & ~n18281 ) ;
  assign n21613 = ( n6148 & n7325 ) | ( n6148 & n10676 ) | ( n7325 & n10676 ) ;
  assign n21614 = n21613 ^ n4142 ^ 1'b0 ;
  assign n21615 = n18351 ^ n12562 ^ x175 ;
  assign n21616 = n21615 ^ n1574 ^ 1'b0 ;
  assign n21617 = ( n2006 & n8285 ) | ( n2006 & n12658 ) | ( n8285 & n12658 ) ;
  assign n21618 = n11265 ^ n5856 ^ 1'b0 ;
  assign n21619 = ~n5506 & n21618 ;
  assign n21620 = n16447 | n21533 ;
  assign n21621 = n408 & ~n21620 ;
  assign n21622 = n3048 & n3330 ;
  assign n21623 = n13862 | n21622 ;
  assign n21624 = n21621 & ~n21623 ;
  assign n21625 = ( n21617 & n21619 ) | ( n21617 & n21624 ) | ( n21619 & n21624 ) ;
  assign n21626 = n20776 ^ n5119 ^ 1'b0 ;
  assign n21627 = n21626 ^ n15626 ^ n4052 ;
  assign n21628 = n8998 ^ n8323 ^ n615 ;
  assign n21629 = n21628 ^ n17434 ^ n15923 ;
  assign n21630 = ( n12507 & ~n21627 ) | ( n12507 & n21629 ) | ( ~n21627 & n21629 ) ;
  assign n21631 = ( n4307 & n20075 ) | ( n4307 & n21630 ) | ( n20075 & n21630 ) ;
  assign n21632 = n18428 ^ n6363 ^ x243 ;
  assign n21633 = n3918 & n21632 ;
  assign n21634 = ( n4743 & n12471 ) | ( n4743 & n17082 ) | ( n12471 & n17082 ) ;
  assign n21635 = n13162 | n21634 ;
  assign n21636 = ( n325 & n7922 ) | ( n325 & ~n15526 ) | ( n7922 & ~n15526 ) ;
  assign n21637 = n21636 ^ n21274 ^ n7682 ;
  assign n21640 = ( n2397 & ~n6821 ) | ( n2397 & n18417 ) | ( ~n6821 & n18417 ) ;
  assign n21638 = ( ~n1875 & n10201 ) | ( ~n1875 & n11459 ) | ( n10201 & n11459 ) ;
  assign n21639 = n21638 ^ n4745 ^ n505 ;
  assign n21641 = n21640 ^ n21639 ^ n15119 ;
  assign n21642 = n15287 ^ n3052 ^ n1274 ;
  assign n21643 = n21642 ^ n14584 ^ n7050 ;
  assign n21644 = n21643 ^ n7830 ^ 1'b0 ;
  assign n21645 = n21644 ^ n19262 ^ n12966 ;
  assign n21646 = n10457 | n15496 ;
  assign n21647 = n21646 ^ n16219 ^ 1'b0 ;
  assign n21648 = ( x218 & n1639 ) | ( x218 & n19455 ) | ( n1639 & n19455 ) ;
  assign n21649 = n21648 ^ n1162 ^ 1'b0 ;
  assign n21650 = ~n10211 & n15972 ;
  assign n21651 = n6127 ^ n4942 ^ 1'b0 ;
  assign n21652 = ~n9857 & n21651 ;
  assign n21653 = ( x224 & ~n21650 ) | ( x224 & n21652 ) | ( ~n21650 & n21652 ) ;
  assign n21654 = n4004 & n21653 ;
  assign n21655 = ( n6442 & n11066 ) | ( n6442 & n15032 ) | ( n11066 & n15032 ) ;
  assign n21656 = n10108 ^ n6069 ^ 1'b0 ;
  assign n21657 = n11357 & ~n21656 ;
  assign n21658 = ( x113 & n8479 ) | ( x113 & ~n21657 ) | ( n8479 & ~n21657 ) ;
  assign n21659 = n20738 & n21658 ;
  assign n21660 = ~n19807 & n21659 ;
  assign n21661 = n12274 ^ n10577 ^ n1463 ;
  assign n21662 = ( n3452 & ~n17630 ) | ( n3452 & n21661 ) | ( ~n17630 & n21661 ) ;
  assign n21663 = n21662 ^ n3841 ^ 1'b0 ;
  assign n21666 = ~n1161 & n4297 ;
  assign n21667 = n3888 & n21666 ;
  assign n21664 = ( n4697 & n10566 ) | ( n4697 & n17144 ) | ( n10566 & n17144 ) ;
  assign n21665 = n21664 ^ n20150 ^ n16914 ;
  assign n21668 = n21667 ^ n21665 ^ n15654 ;
  assign n21669 = n21668 ^ n4710 ^ 1'b0 ;
  assign n21670 = ( n8117 & ~n14567 ) | ( n8117 & n17861 ) | ( ~n14567 & n17861 ) ;
  assign n21671 = ( n5410 & ~n9241 ) | ( n5410 & n11917 ) | ( ~n9241 & n11917 ) ;
  assign n21672 = n18784 | n18836 ;
  assign n21673 = n21671 & ~n21672 ;
  assign n21675 = ( n425 & ~n5846 ) | ( n425 & n8454 ) | ( ~n5846 & n8454 ) ;
  assign n21674 = ( n10279 & ~n16219 ) | ( n10279 & n16433 ) | ( ~n16219 & n16433 ) ;
  assign n21676 = n21675 ^ n21674 ^ n4879 ;
  assign n21677 = ( ~n4721 & n7601 ) | ( ~n4721 & n20728 ) | ( n7601 & n20728 ) ;
  assign n21678 = ( ~n6651 & n16046 ) | ( ~n6651 & n21442 ) | ( n16046 & n21442 ) ;
  assign n21679 = n21678 ^ n3181 ^ 1'b0 ;
  assign n21680 = n6572 & n21679 ;
  assign n21681 = n1899 & n21680 ;
  assign n21682 = ( ~n6271 & n21677 ) | ( ~n6271 & n21681 ) | ( n21677 & n21681 ) ;
  assign n21683 = n18200 ^ n7419 ^ 1'b0 ;
  assign n21685 = n15104 ^ n3594 ^ n3460 ;
  assign n21684 = ~n2472 & n19512 ;
  assign n21686 = n21685 ^ n21684 ^ 1'b0 ;
  assign n21687 = n12792 ^ n8196 ^ n6442 ;
  assign n21688 = ~n3418 & n21687 ;
  assign n21689 = n21688 ^ n3030 ^ 1'b0 ;
  assign n21690 = ~n6073 & n10741 ;
  assign n21691 = ( ~n3497 & n8601 ) | ( ~n3497 & n13749 ) | ( n8601 & n13749 ) ;
  assign n21692 = n21691 ^ n10634 ^ 1'b0 ;
  assign n21693 = ( n1729 & n3820 ) | ( n1729 & ~n9571 ) | ( n3820 & ~n9571 ) ;
  assign n21694 = n5445 ^ n3117 ^ 1'b0 ;
  assign n21695 = n3190 & ~n21694 ;
  assign n21696 = n21693 & n21695 ;
  assign n21698 = ~n3342 & n4438 ;
  assign n21699 = ~n8138 & n21698 ;
  assign n21700 = n21699 ^ n12362 ^ n12200 ;
  assign n21697 = n12663 ^ n7392 ^ 1'b0 ;
  assign n21701 = n21700 ^ n21697 ^ n2916 ;
  assign n21702 = ( n1027 & n3743 ) | ( n1027 & n15158 ) | ( n3743 & n15158 ) ;
  assign n21703 = n21702 ^ n9558 ^ 1'b0 ;
  assign n21704 = n12834 & ~n21703 ;
  assign n21705 = ( n2904 & ~n7807 ) | ( n2904 & n8885 ) | ( ~n7807 & n8885 ) ;
  assign n21706 = n21705 ^ n21116 ^ n17812 ;
  assign n21707 = n15395 ^ n6260 ^ n5857 ;
  assign n21708 = n21707 ^ n9966 ^ 1'b0 ;
  assign n21709 = ~n2679 & n21708 ;
  assign n21713 = n11553 ^ n11155 ^ n4750 ;
  assign n21711 = ( n3577 & n13302 ) | ( n3577 & ~n15660 ) | ( n13302 & ~n15660 ) ;
  assign n21712 = n21711 ^ n11569 ^ x134 ;
  assign n21710 = n16158 ^ n12258 ^ n6359 ;
  assign n21714 = n21713 ^ n21712 ^ n21710 ;
  assign n21715 = n20182 ^ n13651 ^ n3266 ;
  assign n21716 = n16238 ^ n2154 ^ n1493 ;
  assign n21717 = n6801 & n14861 ;
  assign n21718 = n21717 ^ n12059 ^ 1'b0 ;
  assign n21719 = n5818 & n21718 ;
  assign n21720 = ~n15911 & n21719 ;
  assign n21721 = ~n21110 & n21720 ;
  assign n21722 = n8441 ^ n8088 ^ n1025 ;
  assign n21723 = n21722 ^ n5567 ^ 1'b0 ;
  assign n21724 = ( ~n6034 & n12486 ) | ( ~n6034 & n21723 ) | ( n12486 & n21723 ) ;
  assign n21725 = n15294 ^ n3956 ^ n668 ;
  assign n21726 = ( n987 & ~n1768 ) | ( n987 & n5033 ) | ( ~n1768 & n5033 ) ;
  assign n21727 = n21726 ^ n6995 ^ 1'b0 ;
  assign n21728 = ~n21725 & n21727 ;
  assign n21733 = ( n3932 & ~n9639 ) | ( n3932 & n9646 ) | ( ~n9639 & n9646 ) ;
  assign n21734 = n21733 ^ n15693 ^ n5412 ;
  assign n21730 = n12053 ^ n4047 ^ n939 ;
  assign n21731 = n21730 ^ n12416 ^ 1'b0 ;
  assign n21729 = x41 & ~n2393 ;
  assign n21732 = n21731 ^ n21729 ^ n12282 ;
  assign n21735 = n21734 ^ n21732 ^ n10241 ;
  assign n21742 = n7537 ^ n4177 ^ n2706 ;
  assign n21738 = ( n6017 & n8510 ) | ( n6017 & n8592 ) | ( n8510 & n8592 ) ;
  assign n21739 = ( n421 & ~n5350 ) | ( n421 & n7442 ) | ( ~n5350 & n7442 ) ;
  assign n21740 = n21739 ^ n3615 ^ 1'b0 ;
  assign n21741 = ~n21738 & n21740 ;
  assign n21736 = n11914 ^ n7801 ^ 1'b0 ;
  assign n21737 = n18016 & ~n21736 ;
  assign n21743 = n21742 ^ n21741 ^ n21737 ;
  assign n21744 = n6193 & n16172 ;
  assign n21745 = n7756 ^ n5955 ^ n5097 ;
  assign n21746 = ( n1809 & n12807 ) | ( n1809 & ~n21745 ) | ( n12807 & ~n21745 ) ;
  assign n21747 = n3822 & ~n5166 ;
  assign n21748 = ( n519 & ~n12559 ) | ( n519 & n21747 ) | ( ~n12559 & n21747 ) ;
  assign n21749 = n15168 ^ n9257 ^ 1'b0 ;
  assign n21750 = n21748 | n21749 ;
  assign n21754 = ( ~n1754 & n8676 ) | ( ~n1754 & n8772 ) | ( n8676 & n8772 ) ;
  assign n21751 = n9079 & ~n13823 ;
  assign n21752 = ( n6895 & ~n10794 ) | ( n6895 & n21751 ) | ( ~n10794 & n21751 ) ;
  assign n21753 = n2152 & ~n21752 ;
  assign n21755 = n21754 ^ n21753 ^ 1'b0 ;
  assign n21756 = ( n3353 & ~n4093 ) | ( n3353 & n8576 ) | ( ~n4093 & n8576 ) ;
  assign n21757 = ( n4669 & n5134 ) | ( n4669 & ~n16515 ) | ( n5134 & ~n16515 ) ;
  assign n21758 = ( n8061 & n21756 ) | ( n8061 & n21757 ) | ( n21756 & n21757 ) ;
  assign n21759 = n9753 & ~n16745 ;
  assign n21760 = n20470 & n21759 ;
  assign n21762 = n10312 ^ n6942 ^ 1'b0 ;
  assign n21761 = n1924 & ~n13662 ;
  assign n21763 = n21762 ^ n21761 ^ n4853 ;
  assign n21764 = ( n4807 & n21760 ) | ( n4807 & n21763 ) | ( n21760 & n21763 ) ;
  assign n21765 = ( n6591 & ~n9640 ) | ( n6591 & n11893 ) | ( ~n9640 & n11893 ) ;
  assign n21766 = ( n677 & n10776 ) | ( n677 & ~n21765 ) | ( n10776 & ~n21765 ) ;
  assign n21767 = n13042 ^ n5344 ^ n4136 ;
  assign n21768 = ( n3463 & n9529 ) | ( n3463 & n9579 ) | ( n9529 & n9579 ) ;
  assign n21769 = ( n418 & n2092 ) | ( n418 & n2529 ) | ( n2092 & n2529 ) ;
  assign n21770 = x23 & ~n21769 ;
  assign n21771 = n4109 & n21770 ;
  assign n21772 = ( n2667 & ~n10771 ) | ( n2667 & n21771 ) | ( ~n10771 & n21771 ) ;
  assign n21773 = n21768 | n21772 ;
  assign n21774 = n21773 ^ n6814 ^ 1'b0 ;
  assign n21775 = ( n6089 & n21767 ) | ( n6089 & n21774 ) | ( n21767 & n21774 ) ;
  assign n21776 = ( n10823 & n13496 ) | ( n10823 & ~n14037 ) | ( n13496 & ~n14037 ) ;
  assign n21777 = n21776 ^ n20567 ^ n11694 ;
  assign n21778 = n21777 ^ n16197 ^ n16071 ;
  assign n21779 = n12973 & ~n19718 ;
  assign n21780 = n5925 & n21779 ;
  assign n21782 = n4788 & ~n12328 ;
  assign n21781 = n10578 ^ n7573 ^ n6708 ;
  assign n21783 = n21782 ^ n21781 ^ 1'b0 ;
  assign n21784 = ~n21780 & n21783 ;
  assign n21785 = n17604 ^ n7054 ^ n4867 ;
  assign n21786 = ~n7722 & n21785 ;
  assign n21787 = n4417 & n21786 ;
  assign n21788 = ( n3599 & n4438 ) | ( n3599 & ~n21787 ) | ( n4438 & ~n21787 ) ;
  assign n21790 = n2745 & ~n6027 ;
  assign n21789 = n11631 ^ n5524 ^ n3638 ;
  assign n21791 = n21790 ^ n21789 ^ 1'b0 ;
  assign n21792 = ~n2631 & n16357 ;
  assign n21793 = n21792 ^ n10913 ^ 1'b0 ;
  assign n21794 = ( ~n1957 & n21791 ) | ( ~n1957 & n21793 ) | ( n21791 & n21793 ) ;
  assign n21795 = n20056 ^ n17639 ^ 1'b0 ;
  assign n21796 = ~n19651 & n21795 ;
  assign n21797 = n21139 ^ n15503 ^ n5210 ;
  assign n21801 = n4855 & ~n6963 ;
  assign n21802 = ~n9810 & n21801 ;
  assign n21798 = x19 | n7254 ;
  assign n21799 = ( n9962 & ~n10642 ) | ( n9962 & n11244 ) | ( ~n10642 & n11244 ) ;
  assign n21800 = n21798 & ~n21799 ;
  assign n21803 = n21802 ^ n21800 ^ 1'b0 ;
  assign n21804 = n18749 ^ n16928 ^ n16228 ;
  assign n21805 = n21804 ^ n1278 ^ 1'b0 ;
  assign n21807 = n10910 ^ n10074 ^ 1'b0 ;
  assign n21808 = n9011 ^ n7795 ^ n5171 ;
  assign n21809 = n21808 ^ n8218 ^ 1'b0 ;
  assign n21810 = ~n2823 & n21809 ;
  assign n21811 = n21810 ^ n10479 ^ 1'b0 ;
  assign n21812 = n21807 & n21811 ;
  assign n21806 = ( n17203 & ~n19843 ) | ( n17203 & n20584 ) | ( ~n19843 & n20584 ) ;
  assign n21813 = n21812 ^ n21806 ^ n15457 ;
  assign n21814 = ( n6135 & n14572 ) | ( n6135 & ~n16717 ) | ( n14572 & ~n16717 ) ;
  assign n21816 = n1356 ^ n971 ^ 1'b0 ;
  assign n21815 = n16706 & ~n19978 ;
  assign n21817 = n21816 ^ n21815 ^ 1'b0 ;
  assign n21818 = n9449 ^ n1015 ^ 1'b0 ;
  assign n21819 = n8676 & n21818 ;
  assign n21820 = n21819 ^ n3517 ^ n523 ;
  assign n21821 = n21820 ^ n20040 ^ 1'b0 ;
  assign n21822 = ( n877 & ~n11597 ) | ( n877 & n21821 ) | ( ~n11597 & n21821 ) ;
  assign n21823 = n21822 ^ n3963 ^ n3630 ;
  assign n21824 = ( n7160 & n16313 ) | ( n7160 & n21823 ) | ( n16313 & n21823 ) ;
  assign n21825 = n11802 ^ n6058 ^ n4605 ;
  assign n21826 = n13845 & ~n15110 ;
  assign n21827 = n21825 & ~n21826 ;
  assign n21828 = n13899 ^ n653 ^ 1'b0 ;
  assign n21829 = n6301 | n21828 ;
  assign n21830 = n7529 | n13294 ;
  assign n21831 = n21830 ^ n17824 ^ 1'b0 ;
  assign n21832 = n21829 | n21831 ;
  assign n21833 = n20829 & ~n21832 ;
  assign n21834 = ~n3362 & n21833 ;
  assign n21835 = ( n6507 & n7037 ) | ( n6507 & n7814 ) | ( n7037 & n7814 ) ;
  assign n21836 = n10213 ^ n2977 ^ n593 ;
  assign n21837 = ( n7286 & n8345 ) | ( n7286 & ~n21836 ) | ( n8345 & ~n21836 ) ;
  assign n21838 = ( n1902 & ~n21835 ) | ( n1902 & n21837 ) | ( ~n21835 & n21837 ) ;
  assign n21841 = ~n11062 & n13929 ;
  assign n21842 = ~n13584 & n21841 ;
  assign n21839 = ( n2059 & n4616 ) | ( n2059 & n20348 ) | ( n4616 & n20348 ) ;
  assign n21840 = ( n12031 & n14610 ) | ( n12031 & ~n21839 ) | ( n14610 & ~n21839 ) ;
  assign n21843 = n21842 ^ n21840 ^ 1'b0 ;
  assign n21844 = ( ~n17151 & n17706 ) | ( ~n17151 & n19492 ) | ( n17706 & n19492 ) ;
  assign n21845 = ( n5220 & ~n8071 ) | ( n5220 & n12361 ) | ( ~n8071 & n12361 ) ;
  assign n21847 = n15242 ^ n579 ^ n463 ;
  assign n21848 = n21847 ^ n19172 ^ n17765 ;
  assign n21846 = n1672 & ~n11373 ;
  assign n21849 = n21848 ^ n21846 ^ 1'b0 ;
  assign n21850 = ~n459 & n8827 ;
  assign n21851 = ~n7187 & n21850 ;
  assign n21852 = n21851 ^ n12883 ^ n11965 ;
  assign n21853 = n6557 & n7901 ;
  assign n21854 = n7615 & n21853 ;
  assign n21855 = ( ~n572 & n18810 ) | ( ~n572 & n21854 ) | ( n18810 & n21854 ) ;
  assign n21856 = ( n1009 & n21852 ) | ( n1009 & ~n21855 ) | ( n21852 & ~n21855 ) ;
  assign n21857 = n8008 ^ n6341 ^ n4292 ;
  assign n21858 = n21857 ^ n18854 ^ n4166 ;
  assign n21859 = ( n575 & n13773 ) | ( n575 & n21858 ) | ( n13773 & n21858 ) ;
  assign n21860 = ( n8846 & n11501 ) | ( n8846 & ~n15962 ) | ( n11501 & ~n15962 ) ;
  assign n21861 = n17352 ^ n17189 ^ 1'b0 ;
  assign n21862 = n18110 ^ n10672 ^ 1'b0 ;
  assign n21863 = ~n6398 & n21862 ;
  assign n21864 = n7758 & ~n16922 ;
  assign n21866 = ~n664 & n3397 ;
  assign n21867 = n21866 ^ n18489 ^ n4991 ;
  assign n21865 = ~n3383 & n14678 ;
  assign n21868 = n21867 ^ n21865 ^ 1'b0 ;
  assign n21869 = n7522 ^ n5776 ^ n1536 ;
  assign n21870 = n21869 ^ n13555 ^ n3721 ;
  assign n21871 = n8046 & n21870 ;
  assign n21872 = n21871 ^ n9546 ^ 1'b0 ;
  assign n21873 = ( n6021 & ~n10242 ) | ( n6021 & n21872 ) | ( ~n10242 & n21872 ) ;
  assign n21874 = ( n7110 & ~n7788 ) | ( n7110 & n9114 ) | ( ~n7788 & n9114 ) ;
  assign n21875 = ( n1664 & ~n3526 ) | ( n1664 & n21874 ) | ( ~n3526 & n21874 ) ;
  assign n21876 = n6868 & n21875 ;
  assign n21877 = n19729 ^ n12728 ^ 1'b0 ;
  assign n21878 = ( ~n456 & n1853 ) | ( ~n456 & n5761 ) | ( n1853 & n5761 ) ;
  assign n21879 = ( ~n11119 & n12919 ) | ( ~n11119 & n21878 ) | ( n12919 & n21878 ) ;
  assign n21880 = n6372 & n8649 ;
  assign n21881 = ( ~n1120 & n3319 ) | ( ~n1120 & n21880 ) | ( n3319 & n21880 ) ;
  assign n21888 = n5554 ^ n5069 ^ n3489 ;
  assign n21882 = n10243 ^ n3649 ^ 1'b0 ;
  assign n21883 = n18257 & ~n21882 ;
  assign n21884 = n1080 ^ n470 ^ 1'b0 ;
  assign n21885 = ~n12032 & n21884 ;
  assign n21886 = ~n9044 & n21885 ;
  assign n21887 = n21883 & ~n21886 ;
  assign n21889 = n21888 ^ n21887 ^ 1'b0 ;
  assign n21890 = n21889 ^ n5795 ^ n2317 ;
  assign n21891 = ( n3814 & n13982 ) | ( n3814 & ~n21890 ) | ( n13982 & ~n21890 ) ;
  assign n21892 = n14405 ^ n8052 ^ 1'b0 ;
  assign n21893 = n17188 & ~n21892 ;
  assign n21894 = n16892 ^ n4922 ^ 1'b0 ;
  assign n21895 = n1958 & n21894 ;
  assign n21896 = n21895 ^ n16686 ^ 1'b0 ;
  assign n21897 = ( n6843 & ~n9991 ) | ( n6843 & n14282 ) | ( ~n9991 & n14282 ) ;
  assign n21898 = n21897 ^ n20377 ^ 1'b0 ;
  assign n21899 = ( ~n10572 & n21444 ) | ( ~n10572 & n21898 ) | ( n21444 & n21898 ) ;
  assign n21900 = n15345 ^ n13358 ^ n3837 ;
  assign n21901 = ( n3541 & ~n13027 ) | ( n3541 & n21900 ) | ( ~n13027 & n21900 ) ;
  assign n21902 = n8401 ^ n3674 ^ n899 ;
  assign n21903 = ( ~n4703 & n17462 ) | ( ~n4703 & n21902 ) | ( n17462 & n21902 ) ;
  assign n21904 = ( n3754 & n14459 ) | ( n3754 & n21903 ) | ( n14459 & n21903 ) ;
  assign n21905 = n16881 & ~n21532 ;
  assign n21906 = ~n16181 & n21905 ;
  assign n21907 = ( ~n887 & n17821 ) | ( ~n887 & n21906 ) | ( n17821 & n21906 ) ;
  assign n21908 = ( ~n5133 & n5467 ) | ( ~n5133 & n18351 ) | ( n5467 & n18351 ) ;
  assign n21909 = n21908 ^ n11361 ^ 1'b0 ;
  assign n21910 = ~n9729 & n21909 ;
  assign n21911 = n21910 ^ n4782 ^ n2547 ;
  assign n21912 = n6143 & n21911 ;
  assign n21913 = n21912 ^ n5558 ^ 1'b0 ;
  assign n21914 = ~n707 & n18963 ;
  assign n21915 = n21914 ^ n14026 ^ 1'b0 ;
  assign n21916 = n759 & n18613 ;
  assign n21917 = n1290 & n21916 ;
  assign n21918 = n13234 ^ n9575 ^ n4807 ;
  assign n21919 = n20336 | n21918 ;
  assign n21920 = n21919 ^ x6 ^ 1'b0 ;
  assign n21921 = n21920 ^ n4075 ^ 1'b0 ;
  assign n21922 = n21917 | n21921 ;
  assign n21924 = ( n2162 & n14112 ) | ( n2162 & n19172 ) | ( n14112 & n19172 ) ;
  assign n21923 = n1785 & ~n19875 ;
  assign n21925 = n21924 ^ n21923 ^ 1'b0 ;
  assign n21926 = ( n913 & n7191 ) | ( n913 & ~n9740 ) | ( n7191 & ~n9740 ) ;
  assign n21927 = ~n2382 & n5415 ;
  assign n21928 = ( n13786 & ~n14004 ) | ( n13786 & n21927 ) | ( ~n14004 & n21927 ) ;
  assign n21930 = ( n7189 & n16518 ) | ( n7189 & n17012 ) | ( n16518 & n17012 ) ;
  assign n21931 = n21930 ^ n14446 ^ n12082 ;
  assign n21929 = n11713 ^ n728 ^ 1'b0 ;
  assign n21932 = n21931 ^ n21929 ^ n4198 ;
  assign n21933 = n19455 ^ n11730 ^ 1'b0 ;
  assign n21934 = n20958 ^ n16551 ^ n1516 ;
  assign n21935 = n2268 & n21869 ;
  assign n21936 = ~n20553 & n21935 ;
  assign n21937 = ( ~n1712 & n21934 ) | ( ~n1712 & n21936 ) | ( n21934 & n21936 ) ;
  assign n21938 = ( n7905 & ~n19402 ) | ( n7905 & n21937 ) | ( ~n19402 & n21937 ) ;
  assign n21939 = ( n1444 & ~n10319 ) | ( n1444 & n19013 ) | ( ~n10319 & n19013 ) ;
  assign n21940 = ( ~n13073 & n13080 ) | ( ~n13073 & n20207 ) | ( n13080 & n20207 ) ;
  assign n21941 = n5011 ^ n1594 ^ n563 ;
  assign n21942 = ( n15615 & ~n19216 ) | ( n15615 & n21941 ) | ( ~n19216 & n21941 ) ;
  assign n21943 = n14421 ^ n7967 ^ x3 ;
  assign n21944 = ( n4639 & ~n6918 ) | ( n4639 & n7116 ) | ( ~n6918 & n7116 ) ;
  assign n21945 = ( ~n8551 & n21943 ) | ( ~n8551 & n21944 ) | ( n21943 & n21944 ) ;
  assign n21946 = n21945 ^ n7082 ^ 1'b0 ;
  assign n21947 = n7452 | n21946 ;
  assign n21948 = ~n6493 & n15845 ;
  assign n21949 = ~n11218 & n21948 ;
  assign n21950 = n8342 ^ n7022 ^ n4072 ;
  assign n21951 = ( n3678 & n4376 ) | ( n3678 & n13921 ) | ( n4376 & n13921 ) ;
  assign n21952 = n21951 ^ n4930 ^ n4820 ;
  assign n21953 = ( ~n7297 & n21950 ) | ( ~n7297 & n21952 ) | ( n21950 & n21952 ) ;
  assign n21954 = n7307 ^ n6302 ^ 1'b0 ;
  assign n21955 = n21954 ^ n12886 ^ n12008 ;
  assign n21956 = n5608 & n7667 ;
  assign n21957 = n16742 & n21956 ;
  assign n21958 = ( ~n5343 & n12023 ) | ( ~n5343 & n21957 ) | ( n12023 & n21957 ) ;
  assign n21959 = ( x173 & n17107 ) | ( x173 & n21958 ) | ( n17107 & n21958 ) ;
  assign n21960 = ~n12016 & n18233 ;
  assign n21961 = n21960 ^ n16914 ^ 1'b0 ;
  assign n21962 = n1600 & ~n5870 ;
  assign n21963 = n15283 & n21962 ;
  assign n21964 = n5688 & n17681 ;
  assign n21965 = ( ~n2050 & n10573 ) | ( ~n2050 & n15063 ) | ( n10573 & n15063 ) ;
  assign n21966 = ( n2878 & ~n9944 ) | ( n2878 & n10449 ) | ( ~n9944 & n10449 ) ;
  assign n21967 = n3245 ^ n987 ^ 1'b0 ;
  assign n21968 = n21966 & n21967 ;
  assign n21971 = n5975 & n21950 ;
  assign n21972 = n3854 & n21971 ;
  assign n21969 = ( n7361 & ~n14379 ) | ( n7361 & n19086 ) | ( ~n14379 & n19086 ) ;
  assign n21970 = ( n3231 & ~n13773 ) | ( n3231 & n21969 ) | ( ~n13773 & n21969 ) ;
  assign n21973 = n21972 ^ n21970 ^ 1'b0 ;
  assign n21974 = ~n7022 & n21973 ;
  assign n21975 = n9531 ^ n7112 ^ n5620 ;
  assign n21976 = n21975 ^ n20546 ^ n16807 ;
  assign n21977 = ( n17595 & n21974 ) | ( n17595 & n21976 ) | ( n21974 & n21976 ) ;
  assign n21978 = n14270 & ~n17998 ;
  assign n21979 = n17722 ^ n11007 ^ n9077 ;
  assign n21980 = n21979 ^ n20875 ^ n9420 ;
  assign n21981 = n21980 ^ n21368 ^ n8916 ;
  assign n21982 = n5503 ^ n1125 ^ x48 ;
  assign n21983 = n21982 ^ n8582 ^ 1'b0 ;
  assign n21984 = ( ~n14046 & n21981 ) | ( ~n14046 & n21983 ) | ( n21981 & n21983 ) ;
  assign n21989 = n10651 ^ n9602 ^ n3453 ;
  assign n21985 = ( n1431 & n6414 ) | ( n1431 & ~n9673 ) | ( n6414 & ~n9673 ) ;
  assign n21986 = n21985 ^ n21238 ^ n15252 ;
  assign n21987 = n4062 | n21986 ;
  assign n21988 = n1843 | n21987 ;
  assign n21990 = n21989 ^ n21988 ^ n8976 ;
  assign n21998 = ( n2077 & n8585 ) | ( n2077 & ~n12886 ) | ( n8585 & ~n12886 ) ;
  assign n21991 = n3439 & n5863 ;
  assign n21992 = n9896 | n21991 ;
  assign n21993 = n21992 ^ n14209 ^ 1'b0 ;
  assign n21994 = n1299 ^ n882 ^ n379 ;
  assign n21995 = ( n14513 & n18629 ) | ( n14513 & n21994 ) | ( n18629 & n21994 ) ;
  assign n21996 = n21995 ^ n16883 ^ n4570 ;
  assign n21997 = ( ~n21869 & n21993 ) | ( ~n21869 & n21996 ) | ( n21993 & n21996 ) ;
  assign n21999 = n21998 ^ n21997 ^ n16657 ;
  assign n22000 = n19046 ^ n5142 ^ 1'b0 ;
  assign n22001 = n9255 & n22000 ;
  assign n22002 = n1753 & n2366 ;
  assign n22003 = n22002 ^ n9980 ^ n5556 ;
  assign n22004 = n8554 | n22003 ;
  assign n22005 = n22004 ^ n6236 ^ 1'b0 ;
  assign n22006 = n12476 ^ n9790 ^ n9145 ;
  assign n22007 = n2650 & ~n10787 ;
  assign n22008 = n22007 ^ n17519 ^ 1'b0 ;
  assign n22009 = ( n550 & n3157 ) | ( n550 & n5926 ) | ( n3157 & n5926 ) ;
  assign n22010 = ( n5163 & n13011 ) | ( n5163 & n22009 ) | ( n13011 & n22009 ) ;
  assign n22011 = n22010 ^ n8679 ^ n4633 ;
  assign n22012 = x151 | n6467 ;
  assign n22013 = n22012 ^ n14244 ^ n9866 ;
  assign n22014 = ( n5614 & n11594 ) | ( n5614 & n21948 ) | ( n11594 & n21948 ) ;
  assign n22015 = ( n4115 & ~n22013 ) | ( n4115 & n22014 ) | ( ~n22013 & n22014 ) ;
  assign n22016 = ( n13715 & n15993 ) | ( n13715 & n22015 ) | ( n15993 & n22015 ) ;
  assign n22017 = ( n12823 & ~n16029 ) | ( n12823 & n16420 ) | ( ~n16029 & n16420 ) ;
  assign n22018 = n22017 ^ n9292 ^ 1'b0 ;
  assign n22019 = n6185 ^ n1050 ^ 1'b0 ;
  assign n22020 = n6976 | n22019 ;
  assign n22021 = n22020 ^ n14292 ^ n12388 ;
  assign n22022 = n1068 & n16569 ;
  assign n22023 = n22022 ^ n12236 ^ 1'b0 ;
  assign n22024 = n22023 ^ n279 ^ 1'b0 ;
  assign n22025 = n7568 & n22024 ;
  assign n22026 = n6622 & n8339 ;
  assign n22027 = ~n582 & n22026 ;
  assign n22028 = ( x3 & n14883 ) | ( x3 & ~n19693 ) | ( n14883 & ~n19693 ) ;
  assign n22029 = ( n1115 & n8994 ) | ( n1115 & ~n22028 ) | ( n8994 & ~n22028 ) ;
  assign n22030 = n22029 ^ n9522 ^ n5838 ;
  assign n22031 = ~n22027 & n22030 ;
  assign n22032 = ~n22025 & n22031 ;
  assign n22033 = ( n16835 & ~n20627 ) | ( n16835 & n21675 ) | ( ~n20627 & n21675 ) ;
  assign n22034 = n8313 ^ n908 ^ 1'b0 ;
  assign n22035 = n10955 ^ n6717 ^ 1'b0 ;
  assign n22036 = ( ~n4890 & n22034 ) | ( ~n4890 & n22035 ) | ( n22034 & n22035 ) ;
  assign n22037 = ( n5465 & ~n22033 ) | ( n5465 & n22036 ) | ( ~n22033 & n22036 ) ;
  assign n22038 = n7120 ^ n3266 ^ 1'b0 ;
  assign n22039 = ( ~n13577 & n21920 ) | ( ~n13577 & n22038 ) | ( n21920 & n22038 ) ;
  assign n22040 = ( n1359 & n17783 ) | ( n1359 & n22039 ) | ( n17783 & n22039 ) ;
  assign n22041 = n20423 ^ n11336 ^ n4045 ;
  assign n22042 = n4520 | n7021 ;
  assign n22043 = n22042 ^ n11577 ^ 1'b0 ;
  assign n22044 = ( n3877 & n22041 ) | ( n3877 & n22043 ) | ( n22041 & n22043 ) ;
  assign n22045 = ( ~x194 & n13974 ) | ( ~x194 & n22044 ) | ( n13974 & n22044 ) ;
  assign n22046 = n21158 ^ n17564 ^ n5540 ;
  assign n22047 = n3916 | n12391 ;
  assign n22048 = ( n9792 & n22046 ) | ( n9792 & ~n22047 ) | ( n22046 & ~n22047 ) ;
  assign n22049 = n19737 ^ n18672 ^ n18365 ;
  assign n22050 = n7886 | n22049 ;
  assign n22051 = n17174 & ~n22050 ;
  assign n22052 = n6120 ^ n2463 ^ 1'b0 ;
  assign n22053 = n22052 ^ n19271 ^ n8834 ;
  assign n22054 = n12296 ^ n6545 ^ n1158 ;
  assign n22055 = n19853 ^ n9901 ^ n4717 ;
  assign n22056 = n22055 ^ n17743 ^ n7900 ;
  assign n22057 = ~n2389 & n3901 ;
  assign n22058 = n6833 & n22057 ;
  assign n22059 = ( ~n4849 & n13755 ) | ( ~n4849 & n22058 ) | ( n13755 & n22058 ) ;
  assign n22060 = n15788 ^ n14158 ^ n7120 ;
  assign n22061 = n4434 ^ n967 ^ 1'b0 ;
  assign n22062 = n11376 | n22061 ;
  assign n22063 = n18679 ^ n18221 ^ n9765 ;
  assign n22064 = n22063 ^ n861 ^ 1'b0 ;
  assign n22065 = ( n9123 & n22062 ) | ( n9123 & ~n22064 ) | ( n22062 & ~n22064 ) ;
  assign n22066 = n1121 & n8315 ;
  assign n22067 = ~n6097 & n8288 ;
  assign n22068 = n22067 ^ n13354 ^ n3193 ;
  assign n22069 = ( ~n384 & n20467 ) | ( ~n384 & n22068 ) | ( n20467 & n22068 ) ;
  assign n22070 = n22069 ^ n6235 ^ n4350 ;
  assign n22071 = ~n22066 & n22070 ;
  assign n22072 = n13497 ^ n1119 ^ 1'b0 ;
  assign n22073 = ~n10178 & n22072 ;
  assign n22074 = n22073 ^ n9117 ^ n722 ;
  assign n22075 = n10248 ^ n8239 ^ n1299 ;
  assign n22076 = n8742 | n12750 ;
  assign n22077 = n22075 & ~n22076 ;
  assign n22078 = ( n10914 & ~n14549 ) | ( n10914 & n22077 ) | ( ~n14549 & n22077 ) ;
  assign n22079 = ( ~n4422 & n7988 ) | ( ~n4422 & n22078 ) | ( n7988 & n22078 ) ;
  assign n22080 = ( x32 & n836 ) | ( x32 & n5878 ) | ( n836 & n5878 ) ;
  assign n22081 = n22080 ^ n20116 ^ 1'b0 ;
  assign n22082 = ( ~n11601 & n16964 ) | ( ~n11601 & n22081 ) | ( n16964 & n22081 ) ;
  assign n22083 = n19494 ^ n12912 ^ n12564 ;
  assign n22084 = n22083 ^ n16548 ^ n3269 ;
  assign n22085 = n7628 & ~n10280 ;
  assign n22086 = ~n19679 & n22085 ;
  assign n22088 = n6083 & n7818 ;
  assign n22089 = n22088 ^ n21829 ^ 1'b0 ;
  assign n22087 = n14844 ^ n12595 ^ n7592 ;
  assign n22090 = n22089 ^ n22087 ^ 1'b0 ;
  assign n22091 = ( ~x158 & n563 ) | ( ~x158 & n4256 ) | ( n563 & n4256 ) ;
  assign n22092 = ( n5346 & n13125 ) | ( n5346 & n21447 ) | ( n13125 & n21447 ) ;
  assign n22094 = ( n1233 & n5910 ) | ( n1233 & ~n7830 ) | ( n5910 & ~n7830 ) ;
  assign n22095 = n22094 ^ n4625 ^ n2417 ;
  assign n22093 = ~n673 & n6182 ;
  assign n22096 = n22095 ^ n22093 ^ 1'b0 ;
  assign n22097 = ( n12335 & n17748 ) | ( n12335 & n22096 ) | ( n17748 & n22096 ) ;
  assign n22098 = ( n22091 & n22092 ) | ( n22091 & ~n22097 ) | ( n22092 & ~n22097 ) ;
  assign n22099 = n5613 ^ n418 ^ 1'b0 ;
  assign n22100 = ~n8173 & n22099 ;
  assign n22101 = n22100 ^ n7873 ^ n5100 ;
  assign n22102 = n22101 ^ n14266 ^ 1'b0 ;
  assign n22103 = n12182 & n22102 ;
  assign n22104 = ( n9412 & n10453 ) | ( n9412 & ~n22103 ) | ( n10453 & ~n22103 ) ;
  assign n22105 = n2184 | n12826 ;
  assign n22106 = n22105 ^ n9422 ^ 1'b0 ;
  assign n22107 = n2533 & n16268 ;
  assign n22108 = n22107 ^ n14893 ^ 1'b0 ;
  assign n22109 = ( ~n6985 & n15108 ) | ( ~n6985 & n22108 ) | ( n15108 & n22108 ) ;
  assign n22110 = n22109 ^ n9160 ^ n3340 ;
  assign n22111 = n14505 ^ n4855 ^ 1'b0 ;
  assign n22112 = n4805 & ~n22111 ;
  assign n22113 = n11663 & n22112 ;
  assign n22114 = n22113 ^ n20524 ^ n19526 ;
  assign n22118 = n7044 ^ n3481 ^ n719 ;
  assign n22116 = n11126 ^ n11023 ^ 1'b0 ;
  assign n22117 = n6040 | n22116 ;
  assign n22115 = ~n6945 & n12688 ;
  assign n22119 = n22118 ^ n22117 ^ n22115 ;
  assign n22120 = ( n11133 & n22114 ) | ( n11133 & n22119 ) | ( n22114 & n22119 ) ;
  assign n22122 = ( n10702 & n11603 ) | ( n10702 & ~n11970 ) | ( n11603 & ~n11970 ) ;
  assign n22123 = ( n10391 & ~n19579 ) | ( n10391 & n22122 ) | ( ~n19579 & n22122 ) ;
  assign n22121 = ( n568 & ~n3050 ) | ( n568 & n8544 ) | ( ~n3050 & n8544 ) ;
  assign n22124 = n22123 ^ n22121 ^ n21596 ;
  assign n22125 = n10506 ^ n9471 ^ 1'b0 ;
  assign n22126 = n14572 & n22125 ;
  assign n22127 = n5597 & n9606 ;
  assign n22128 = n22127 ^ n15315 ^ 1'b0 ;
  assign n22129 = ( n2217 & n8813 ) | ( n2217 & ~n22128 ) | ( n8813 & ~n22128 ) ;
  assign n22130 = ( ~n6110 & n8750 ) | ( ~n6110 & n12890 ) | ( n8750 & n12890 ) ;
  assign n22132 = n1076 | n2559 ;
  assign n22131 = n10731 ^ n9740 ^ 1'b0 ;
  assign n22133 = n22132 ^ n22131 ^ n7187 ;
  assign n22134 = ~n22130 & n22133 ;
  assign n22135 = n7245 & ~n10749 ;
  assign n22136 = n7972 & n22135 ;
  assign n22137 = n12260 ^ n3808 ^ n2581 ;
  assign n22138 = ( x70 & n4323 ) | ( x70 & n22137 ) | ( n4323 & n22137 ) ;
  assign n22140 = n15949 ^ n6338 ^ n1583 ;
  assign n22139 = ( n8585 & ~n9999 ) | ( n8585 & n14402 ) | ( ~n9999 & n14402 ) ;
  assign n22141 = n22140 ^ n22139 ^ n10708 ;
  assign n22142 = ( n22136 & n22138 ) | ( n22136 & n22141 ) | ( n22138 & n22141 ) ;
  assign n22143 = n22142 ^ n6547 ^ 1'b0 ;
  assign n22144 = n15959 ^ n1954 ^ 1'b0 ;
  assign n22145 = n6216 | n22144 ;
  assign n22146 = n22145 ^ n18810 ^ n6871 ;
  assign n22147 = n20022 ^ n18096 ^ n13535 ;
  assign n22149 = n2762 | n13693 ;
  assign n22148 = n12268 ^ n5108 ^ 1'b0 ;
  assign n22150 = n22149 ^ n22148 ^ n2956 ;
  assign n22151 = n22150 ^ n15215 ^ n9112 ;
  assign n22152 = n21032 ^ n20553 ^ n17695 ;
  assign n22153 = n22152 ^ n10794 ^ n7476 ;
  assign n22154 = ( x29 & n4673 ) | ( x29 & n22132 ) | ( n4673 & n22132 ) ;
  assign n22155 = n12092 & ~n22154 ;
  assign n22156 = n22155 ^ n19422 ^ 1'b0 ;
  assign n22157 = n22156 ^ n2379 ^ 1'b0 ;
  assign n22158 = n22157 ^ n5658 ^ 1'b0 ;
  assign n22159 = n21549 | n22158 ;
  assign n22160 = n11251 ^ n4639 ^ 1'b0 ;
  assign n22161 = ~n22159 & n22160 ;
  assign n22162 = ( n5335 & n6237 ) | ( n5335 & n9638 ) | ( n6237 & n9638 ) ;
  assign n22163 = n10434 ^ n5213 ^ n5169 ;
  assign n22164 = n22163 ^ n10982 ^ n7924 ;
  assign n22165 = n10422 | n22164 ;
  assign n22166 = n6182 | n22165 ;
  assign n22181 = n21435 ^ n14296 ^ n4190 ;
  assign n22182 = n22181 ^ n3435 ^ 1'b0 ;
  assign n22167 = n9712 ^ n9291 ^ n1752 ;
  assign n22168 = ( n4217 & n6855 ) | ( n4217 & ~n22167 ) | ( n6855 & ~n22167 ) ;
  assign n22169 = n10573 ^ n9918 ^ 1'b0 ;
  assign n22170 = n22169 ^ n8644 ^ n7302 ;
  assign n22171 = n22170 ^ n17838 ^ n17180 ;
  assign n22172 = n455 | n19130 ;
  assign n22173 = ( ~n17704 & n22171 ) | ( ~n17704 & n22172 ) | ( n22171 & n22172 ) ;
  assign n22176 = ( n4014 & n11556 ) | ( n4014 & n15368 ) | ( n11556 & n15368 ) ;
  assign n22174 = n12998 ^ n8793 ^ 1'b0 ;
  assign n22175 = n4462 & n22174 ;
  assign n22177 = n22176 ^ n22175 ^ 1'b0 ;
  assign n22178 = ~n22173 & n22177 ;
  assign n22179 = ( ~x203 & n752 ) | ( ~x203 & n22178 ) | ( n752 & n22178 ) ;
  assign n22180 = ( ~n15281 & n22168 ) | ( ~n15281 & n22179 ) | ( n22168 & n22179 ) ;
  assign n22183 = n22182 ^ n22180 ^ n3235 ;
  assign n22184 = ( n2101 & n2271 ) | ( n2101 & ~n8669 ) | ( n2271 & ~n8669 ) ;
  assign n22185 = n14675 ^ n1222 ^ 1'b0 ;
  assign n22186 = n19070 | n22185 ;
  assign n22187 = n22186 ^ n20260 ^ 1'b0 ;
  assign n22188 = ~n22184 & n22187 ;
  assign n22189 = ( ~n5745 & n8819 ) | ( ~n5745 & n22188 ) | ( n8819 & n22188 ) ;
  assign n22190 = n13701 | n19047 ;
  assign n22191 = n14518 ^ n4200 ^ 1'b0 ;
  assign n22192 = ~n22190 & n22191 ;
  assign n22193 = n13514 ^ n6695 ^ n4605 ;
  assign n22194 = ( n18148 & ~n22192 ) | ( n18148 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n22195 = ( ~n3303 & n9270 ) | ( ~n3303 & n16081 ) | ( n9270 & n16081 ) ;
  assign n22196 = ( n9816 & n15073 ) | ( n9816 & ~n22195 ) | ( n15073 & ~n22195 ) ;
  assign n22202 = ( ~n4955 & n12232 ) | ( ~n4955 & n14471 ) | ( n12232 & n14471 ) ;
  assign n22203 = n22202 ^ n11919 ^ n9505 ;
  assign n22197 = ( n5769 & ~n9361 ) | ( n5769 & n11773 ) | ( ~n9361 & n11773 ) ;
  assign n22198 = ( n4736 & ~n9383 ) | ( n4736 & n22197 ) | ( ~n9383 & n22197 ) ;
  assign n22199 = n14282 & ~n22198 ;
  assign n22200 = ~n19030 & n22199 ;
  assign n22201 = n4156 | n22200 ;
  assign n22204 = n22203 ^ n22201 ^ 1'b0 ;
  assign n22205 = n4092 & ~n22204 ;
  assign n22206 = n22196 & n22205 ;
  assign n22207 = ~n13768 & n21477 ;
  assign n22209 = n15534 ^ n5445 ^ n2270 ;
  assign n22208 = n4790 | n11483 ;
  assign n22210 = n22209 ^ n22208 ^ 1'b0 ;
  assign n22211 = n15224 ^ n9687 ^ 1'b0 ;
  assign n22212 = n22211 ^ n20596 ^ n3106 ;
  assign n22215 = ( n6317 & n8626 ) | ( n6317 & n9515 ) | ( n8626 & n9515 ) ;
  assign n22213 = n7080 ^ n4288 ^ n3713 ;
  assign n22214 = n22213 ^ n7560 ^ n5435 ;
  assign n22216 = n22215 ^ n22214 ^ n5115 ;
  assign n22218 = n7668 ^ n3504 ^ x68 ;
  assign n22219 = ( n5884 & n8403 ) | ( n5884 & ~n22218 ) | ( n8403 & ~n22218 ) ;
  assign n22217 = n16810 ^ n1284 ^ n889 ;
  assign n22220 = n22219 ^ n22217 ^ n9751 ;
  assign n22222 = ( ~n1499 & n9065 ) | ( ~n1499 & n9571 ) | ( n9065 & n9571 ) ;
  assign n22223 = ~n17174 & n22222 ;
  assign n22224 = n22223 ^ n21685 ^ 1'b0 ;
  assign n22221 = ( n4594 & ~n6614 ) | ( n4594 & n6659 ) | ( ~n6614 & n6659 ) ;
  assign n22225 = n22224 ^ n22221 ^ n11400 ;
  assign n22226 = n15298 ^ n7105 ^ 1'b0 ;
  assign n22227 = ~n742 & n22226 ;
  assign n22228 = ( n7689 & n9261 ) | ( n7689 & n22227 ) | ( n9261 & n22227 ) ;
  assign n22229 = x149 & n22228 ;
  assign n22230 = ~n3022 & n3303 ;
  assign n22231 = ( n5763 & ~n16043 ) | ( n5763 & n22230 ) | ( ~n16043 & n22230 ) ;
  assign n22232 = n20103 ^ n19628 ^ n19293 ;
  assign n22233 = n2865 ^ n1293 ^ n1242 ;
  assign n22234 = n22233 ^ n9398 ^ n7479 ;
  assign n22235 = n22234 ^ n8267 ^ n2231 ;
  assign n22236 = n22235 ^ n4842 ^ n2068 ;
  assign n22237 = n22236 ^ n8848 ^ 1'b0 ;
  assign n22238 = n17560 & ~n22237 ;
  assign n22245 = ( n2348 & n4811 ) | ( n2348 & n20997 ) | ( n4811 & n20997 ) ;
  assign n22239 = ~n5098 & n11768 ;
  assign n22240 = n22239 ^ n3343 ^ 1'b0 ;
  assign n22241 = n1448 | n22240 ;
  assign n22242 = n22241 ^ n11461 ^ 1'b0 ;
  assign n22243 = ( n6783 & n8462 ) | ( n6783 & ~n22242 ) | ( n8462 & ~n22242 ) ;
  assign n22244 = n22243 ^ n10287 ^ n5930 ;
  assign n22246 = n22245 ^ n22244 ^ n2217 ;
  assign n22247 = ( n4328 & ~n6049 ) | ( n4328 & n7345 ) | ( ~n6049 & n7345 ) ;
  assign n22248 = n22247 ^ n20432 ^ n19349 ;
  assign n22252 = n10570 ^ n3636 ^ 1'b0 ;
  assign n22253 = ~n6123 & n22252 ;
  assign n22249 = ( n942 & n4205 ) | ( n942 & ~n4245 ) | ( n4205 & ~n4245 ) ;
  assign n22250 = n22249 ^ n10016 ^ x86 ;
  assign n22251 = n22250 ^ n8777 ^ n7808 ;
  assign n22254 = n22253 ^ n22251 ^ 1'b0 ;
  assign n22255 = n22248 & ~n22254 ;
  assign n22256 = ( n3010 & ~n3248 ) | ( n3010 & n19764 ) | ( ~n3248 & n19764 ) ;
  assign n22257 = ( n4826 & ~n18162 ) | ( n4826 & n22256 ) | ( ~n18162 & n22256 ) ;
  assign n22258 = n22257 ^ n22030 ^ 1'b0 ;
  assign n22259 = n14549 ^ n8137 ^ n6093 ;
  assign n22260 = n2754 & n22259 ;
  assign n22261 = n9085 & n22260 ;
  assign n22262 = n22261 ^ n14828 ^ 1'b0 ;
  assign n22263 = n2089 & ~n22262 ;
  assign n22264 = n16312 & n22263 ;
  assign n22265 = ~n7277 & n7821 ;
  assign n22266 = n12598 & n22265 ;
  assign n22267 = n22266 ^ n874 ^ 1'b0 ;
  assign n22268 = x6 & n6998 ;
  assign n22269 = n22268 ^ n5939 ^ 1'b0 ;
  assign n22270 = ( n6403 & n21050 ) | ( n6403 & ~n22269 ) | ( n21050 & ~n22269 ) ;
  assign n22271 = ( ~n9659 & n11695 ) | ( ~n9659 & n19219 ) | ( n11695 & n19219 ) ;
  assign n22272 = ( n6023 & n11217 ) | ( n6023 & ~n22271 ) | ( n11217 & ~n22271 ) ;
  assign n22273 = n12553 & ~n22272 ;
  assign n22274 = ( n7462 & ~n22270 ) | ( n7462 & n22273 ) | ( ~n22270 & n22273 ) ;
  assign n22275 = ( n4422 & n5843 ) | ( n4422 & n10739 ) | ( n5843 & n10739 ) ;
  assign n22276 = ~n15405 & n16180 ;
  assign n22277 = n22275 & ~n22276 ;
  assign n22278 = n19114 ^ n17056 ^ n13858 ;
  assign n22279 = ( n1120 & ~n10317 ) | ( n1120 & n10737 ) | ( ~n10317 & n10737 ) ;
  assign n22280 = n22279 ^ n14837 ^ 1'b0 ;
  assign n22281 = ( n21798 & ~n22278 ) | ( n21798 & n22280 ) | ( ~n22278 & n22280 ) ;
  assign n22282 = n16266 ^ n5945 ^ x45 ;
  assign n22283 = ( ~n12069 & n14569 ) | ( ~n12069 & n22282 ) | ( n14569 & n22282 ) ;
  assign n22284 = n15501 ^ n11276 ^ n1217 ;
  assign n22285 = n12588 ^ n11875 ^ 1'b0 ;
  assign n22286 = n8436 & ~n22285 ;
  assign n22287 = ( ~n7768 & n10652 ) | ( ~n7768 & n22286 ) | ( n10652 & n22286 ) ;
  assign n22288 = ( ~n2688 & n11803 ) | ( ~n2688 & n22287 ) | ( n11803 & n22287 ) ;
  assign n22289 = n22288 ^ n21208 ^ n12009 ;
  assign n22290 = n5806 ^ n1924 ^ n1321 ;
  assign n22291 = ( n1479 & n11725 ) | ( n1479 & n22290 ) | ( n11725 & n22290 ) ;
  assign n22292 = ( ~n16391 & n17234 ) | ( ~n16391 & n18467 ) | ( n17234 & n18467 ) ;
  assign n22293 = ( n763 & n7967 ) | ( n763 & ~n10398 ) | ( n7967 & ~n10398 ) ;
  assign n22294 = n1729 & ~n22293 ;
  assign n22295 = n4787 & n22294 ;
  assign n22296 = n14630 ^ n13531 ^ n10495 ;
  assign n22297 = n325 | n22296 ;
  assign n22298 = ( x239 & n17140 ) | ( x239 & ~n22297 ) | ( n17140 & ~n22297 ) ;
  assign n22299 = ~n1416 & n14654 ;
  assign n22300 = n18691 & n22299 ;
  assign n22301 = n22300 ^ n6877 ^ 1'b0 ;
  assign n22302 = n11298 ^ n7338 ^ 1'b0 ;
  assign n22303 = n7807 & ~n22302 ;
  assign n22304 = ( ~n7423 & n14713 ) | ( ~n7423 & n16487 ) | ( n14713 & n16487 ) ;
  assign n22305 = n10150 & n13937 ;
  assign n22306 = ~n22304 & n22305 ;
  assign n22307 = ( n2749 & ~n6491 ) | ( n2749 & n13304 ) | ( ~n6491 & n13304 ) ;
  assign n22308 = ( n4304 & n14648 ) | ( n4304 & ~n22307 ) | ( n14648 & ~n22307 ) ;
  assign n22309 = ( ~n2377 & n14438 ) | ( ~n2377 & n22308 ) | ( n14438 & n22308 ) ;
  assign n22310 = ( x166 & n6368 ) | ( x166 & n8136 ) | ( n6368 & n8136 ) ;
  assign n22311 = ( n1977 & n3038 ) | ( n1977 & ~n6633 ) | ( n3038 & ~n6633 ) ;
  assign n22312 = ( n4186 & n16373 ) | ( n4186 & n22311 ) | ( n16373 & n22311 ) ;
  assign n22313 = n7736 ^ n5338 ^ n1125 ;
  assign n22314 = ( n22310 & n22312 ) | ( n22310 & ~n22313 ) | ( n22312 & ~n22313 ) ;
  assign n22315 = n22314 ^ n21308 ^ 1'b0 ;
  assign n22316 = n9591 ^ n8757 ^ 1'b0 ;
  assign n22317 = ( n3356 & ~n5609 ) | ( n3356 & n22316 ) | ( ~n5609 & n22316 ) ;
  assign n22318 = n22317 ^ n846 ^ 1'b0 ;
  assign n22319 = n16480 | n22318 ;
  assign n22320 = n17414 & ~n20427 ;
  assign n22321 = n22319 & n22320 ;
  assign n22327 = n4507 & ~n5613 ;
  assign n22328 = n22327 ^ n3686 ^ 1'b0 ;
  assign n22329 = ~n18417 & n22328 ;
  assign n22330 = n16004 & n22329 ;
  assign n22322 = n9306 ^ n7746 ^ 1'b0 ;
  assign n22323 = n14495 & ~n22322 ;
  assign n22324 = ~n9692 & n17141 ;
  assign n22325 = ~n22323 & n22324 ;
  assign n22326 = n22325 ^ n17198 ^ n12075 ;
  assign n22331 = n22330 ^ n22326 ^ n1140 ;
  assign n22332 = ( n6087 & ~n11252 ) | ( n6087 & n13232 ) | ( ~n11252 & n13232 ) ;
  assign n22333 = n3448 | n7018 ;
  assign n22334 = n22333 ^ n3306 ^ 1'b0 ;
  assign n22335 = n21767 ^ n3781 ^ n3399 ;
  assign n22336 = n22335 ^ n15034 ^ 1'b0 ;
  assign n22337 = ( n9380 & n22334 ) | ( n9380 & n22336 ) | ( n22334 & n22336 ) ;
  assign n22338 = n19293 & n22337 ;
  assign n22339 = n22338 ^ n12250 ^ n1999 ;
  assign n22340 = ( n7515 & n22332 ) | ( n7515 & n22339 ) | ( n22332 & n22339 ) ;
  assign n22341 = n16589 | n21304 ;
  assign n22342 = n19818 ^ n10945 ^ n10796 ;
  assign n22343 = n9812 ^ n5797 ^ 1'b0 ;
  assign n22344 = n22343 ^ n10896 ^ n5863 ;
  assign n22345 = n22344 ^ n11277 ^ x121 ;
  assign n22346 = n846 & n1537 ;
  assign n22347 = n22346 ^ n961 ^ 1'b0 ;
  assign n22348 = n3731 | n22240 ;
  assign n22349 = n22348 ^ n4865 ^ x110 ;
  assign n22350 = n21053 ^ n7758 ^ n3285 ;
  assign n22351 = n604 | n778 ;
  assign n22352 = n1583 & ~n22351 ;
  assign n22353 = n22352 ^ n1622 ^ 1'b0 ;
  assign n22354 = n1429 & ~n13512 ;
  assign n22355 = n2245 & n22354 ;
  assign n22356 = n5208 & n22355 ;
  assign n22357 = n22356 ^ n1631 ^ 1'b0 ;
  assign n22358 = n9303 & n22357 ;
  assign n22359 = n22358 ^ n2668 ^ 1'b0 ;
  assign n22360 = n7674 & ~n8464 ;
  assign n22361 = ~n15902 & n22360 ;
  assign n22362 = n2708 | n7965 ;
  assign n22363 = ( n1040 & ~n11079 ) | ( n1040 & n22362 ) | ( ~n11079 & n22362 ) ;
  assign n22364 = n11863 ^ n3245 ^ 1'b0 ;
  assign n22365 = ~n22363 & n22364 ;
  assign n22366 = n8076 ^ n3904 ^ 1'b0 ;
  assign n22367 = n7834 & n22366 ;
  assign n22368 = n22367 ^ n6660 ^ 1'b0 ;
  assign n22369 = ( n1558 & ~n2294 ) | ( n1558 & n15696 ) | ( ~n2294 & n15696 ) ;
  assign n22370 = ( n4916 & n19512 ) | ( n4916 & n22369 ) | ( n19512 & n22369 ) ;
  assign n22372 = n8175 ^ n6919 ^ n1358 ;
  assign n22371 = n9694 ^ n7329 ^ x127 ;
  assign n22373 = n22372 ^ n22371 ^ n20515 ;
  assign n22374 = ( ~n8714 & n14266 ) | ( ~n8714 & n22373 ) | ( n14266 & n22373 ) ;
  assign n22375 = n3599 ^ n374 ^ x97 ;
  assign n22376 = ( n3684 & n6048 ) | ( n3684 & ~n18699 ) | ( n6048 & ~n18699 ) ;
  assign n22377 = n287 & ~n22376 ;
  assign n22378 = n14282 ^ n1771 ^ 1'b0 ;
  assign n22379 = ~n2848 & n22378 ;
  assign n22380 = ~n18896 & n22379 ;
  assign n22381 = n22380 ^ n18994 ^ 1'b0 ;
  assign n22382 = ~n752 & n9443 ;
  assign n22383 = n4475 | n22382 ;
  assign n22385 = ( ~n8833 & n10573 ) | ( ~n8833 & n14516 ) | ( n10573 & n14516 ) ;
  assign n22384 = n9066 ^ n347 ^ 1'b0 ;
  assign n22386 = n22385 ^ n22384 ^ n3538 ;
  assign n22387 = n10923 ^ n1612 ^ 1'b0 ;
  assign n22388 = n22386 & ~n22387 ;
  assign n22389 = n18612 & ~n22388 ;
  assign n22390 = n7508 ^ n3219 ^ 1'b0 ;
  assign n22391 = n9557 & n22390 ;
  assign n22392 = n22391 ^ n10439 ^ n2765 ;
  assign n22393 = n20423 ^ n19624 ^ 1'b0 ;
  assign n22394 = n22393 ^ n18554 ^ 1'b0 ;
  assign n22395 = n22392 & ~n22394 ;
  assign n22396 = n21969 ^ n15777 ^ n9965 ;
  assign n22397 = ( ~n4093 & n10649 ) | ( ~n4093 & n20969 ) | ( n10649 & n20969 ) ;
  assign n22398 = n22397 ^ n12635 ^ n7553 ;
  assign n22399 = ( ~x84 & n22396 ) | ( ~x84 & n22398 ) | ( n22396 & n22398 ) ;
  assign n22404 = n7741 ^ n3961 ^ n1297 ;
  assign n22400 = n7574 ^ n909 ^ 1'b0 ;
  assign n22401 = ~n1791 & n22400 ;
  assign n22402 = n22401 ^ n15274 ^ n5523 ;
  assign n22403 = n22402 ^ n20234 ^ n1672 ;
  assign n22405 = n22404 ^ n22403 ^ n16518 ;
  assign n22406 = n7277 | n14945 ;
  assign n22407 = n13961 ^ n3209 ^ n681 ;
  assign n22408 = n20829 ^ n11164 ^ n10296 ;
  assign n22409 = n19115 ^ n4288 ^ 1'b0 ;
  assign n22410 = n8226 & n22409 ;
  assign n22411 = ( x219 & n3749 ) | ( x219 & n22410 ) | ( n3749 & n22410 ) ;
  assign n22414 = n8400 & n17955 ;
  assign n22415 = ~n4507 & n22414 ;
  assign n22412 = ( n1149 & ~n1523 ) | ( n1149 & n5300 ) | ( ~n1523 & n5300 ) ;
  assign n22413 = n22412 ^ n9361 ^ 1'b0 ;
  assign n22416 = n22415 ^ n22413 ^ n14296 ;
  assign n22417 = ( n3889 & n22411 ) | ( n3889 & n22416 ) | ( n22411 & n22416 ) ;
  assign n22418 = n22417 ^ n22140 ^ n8851 ;
  assign n22419 = ( n22407 & ~n22408 ) | ( n22407 & n22418 ) | ( ~n22408 & n22418 ) ;
  assign n22420 = ( n1326 & n11787 ) | ( n1326 & ~n22066 ) | ( n11787 & ~n22066 ) ;
  assign n22421 = ~n6593 & n7775 ;
  assign n22422 = ~n2454 & n22421 ;
  assign n22423 = n22422 ^ n13762 ^ n830 ;
  assign n22424 = n17183 ^ n6666 ^ 1'b0 ;
  assign n22425 = ( n2113 & ~n14594 ) | ( n2113 & n22424 ) | ( ~n14594 & n22424 ) ;
  assign n22426 = ( n3816 & ~n12272 ) | ( n3816 & n22425 ) | ( ~n12272 & n22425 ) ;
  assign n22427 = n22426 ^ n13386 ^ 1'b0 ;
  assign n22428 = n14419 & ~n16885 ;
  assign n22429 = n22428 ^ n3524 ^ 1'b0 ;
  assign n22430 = ( n2152 & ~n22427 ) | ( n2152 & n22429 ) | ( ~n22427 & n22429 ) ;
  assign n22431 = ~n8375 & n21348 ;
  assign n22432 = n16667 & n22431 ;
  assign n22433 = n22432 ^ n2075 ^ n1697 ;
  assign n22434 = n21657 ^ n20380 ^ n1194 ;
  assign n22435 = n22434 ^ n7378 ^ 1'b0 ;
  assign n22436 = n22433 & n22435 ;
  assign n22437 = n22436 ^ n15932 ^ 1'b0 ;
  assign n22438 = n1632 | n3629 ;
  assign n22439 = n12564 & ~n22438 ;
  assign n22440 = ( n10929 & n13244 ) | ( n10929 & ~n17574 ) | ( n13244 & ~n17574 ) ;
  assign n22441 = n22440 ^ n3385 ^ 1'b0 ;
  assign n22442 = ~n20107 & n22441 ;
  assign n22443 = n22442 ^ n13774 ^ n10929 ;
  assign n22444 = n16532 ^ n14278 ^ n13002 ;
  assign n22445 = n13361 ^ n5024 ^ n2756 ;
  assign n22446 = n11365 ^ n778 ^ 1'b0 ;
  assign n22447 = ( n2441 & ~n12230 ) | ( n2441 & n22446 ) | ( ~n12230 & n22446 ) ;
  assign n22448 = ( n1758 & ~n4916 ) | ( n1758 & n6917 ) | ( ~n4916 & n6917 ) ;
  assign n22449 = ( n7506 & n8226 ) | ( n7506 & n22448 ) | ( n8226 & n22448 ) ;
  assign n22450 = ( n3716 & n10062 ) | ( n3716 & ~n22449 ) | ( n10062 & ~n22449 ) ;
  assign n22451 = n22450 ^ n13009 ^ n301 ;
  assign n22452 = n981 & ~n4586 ;
  assign n22453 = ~n4674 & n22452 ;
  assign n22454 = n22453 ^ n5255 ^ 1'b0 ;
  assign n22455 = n12965 | n22454 ;
  assign n22456 = ~n1400 & n11934 ;
  assign n22457 = n19897 ^ n9861 ^ 1'b0 ;
  assign n22458 = ~n22456 & n22457 ;
  assign n22459 = n22458 ^ n17434 ^ n5017 ;
  assign n22460 = n13530 | n17265 ;
  assign n22469 = n21460 ^ n7720 ^ 1'b0 ;
  assign n22470 = n2670 & n22469 ;
  assign n22462 = x57 & n1125 ;
  assign n22463 = n13589 & ~n22462 ;
  assign n22464 = ~n5824 & n22463 ;
  assign n22465 = n16254 ^ n8367 ^ n1379 ;
  assign n22466 = ( n14202 & n22464 ) | ( n14202 & ~n22465 ) | ( n22464 & ~n22465 ) ;
  assign n22461 = ( ~n599 & n5083 ) | ( ~n599 & n20941 ) | ( n5083 & n20941 ) ;
  assign n22467 = n22466 ^ n22461 ^ n19617 ;
  assign n22468 = n22467 ^ n5909 ^ 1'b0 ;
  assign n22471 = n22470 ^ n22468 ^ n511 ;
  assign n22472 = n3050 & n3753 ;
  assign n22473 = n9214 & n22472 ;
  assign n22474 = n22473 ^ n7045 ^ 1'b0 ;
  assign n22475 = ( n14047 & n18576 ) | ( n14047 & ~n22474 ) | ( n18576 & ~n22474 ) ;
  assign n22476 = n1712 | n17502 ;
  assign n22477 = n7407 & ~n22476 ;
  assign n22478 = n14016 ^ n12804 ^ n8906 ;
  assign n22479 = ~n3420 & n22478 ;
  assign n22480 = ( ~n5932 & n7689 ) | ( ~n5932 & n19198 ) | ( n7689 & n19198 ) ;
  assign n22481 = n9385 & n22062 ;
  assign n22482 = n18207 ^ n14813 ^ 1'b0 ;
  assign n22483 = n18036 & ~n22482 ;
  assign n22484 = n2538 ^ n501 ^ 1'b0 ;
  assign n22485 = ( n2200 & ~n14629 ) | ( n2200 & n16111 ) | ( ~n14629 & n16111 ) ;
  assign n22486 = n10766 ^ n8571 ^ n1860 ;
  assign n22487 = n22486 ^ n19888 ^ n4283 ;
  assign n22488 = ( n7903 & n22485 ) | ( n7903 & ~n22487 ) | ( n22485 & ~n22487 ) ;
  assign n22489 = n22484 & n22488 ;
  assign n22490 = n14140 ^ n1352 ^ 1'b0 ;
  assign n22491 = n1599 | n22490 ;
  assign n22492 = ( n3977 & n22489 ) | ( n3977 & n22491 ) | ( n22489 & n22491 ) ;
  assign n22493 = n5521 & ~n8175 ;
  assign n22494 = n5271 & n22493 ;
  assign n22495 = n22494 ^ n9899 ^ n2696 ;
  assign n22496 = n2854 & n4301 ;
  assign n22497 = n22496 ^ n12592 ^ 1'b0 ;
  assign n22498 = n22497 ^ n9130 ^ n8829 ;
  assign n22499 = n1007 & n7876 ;
  assign n22500 = ~n4888 & n22499 ;
  assign n22501 = ( n10907 & n19092 ) | ( n10907 & ~n22500 ) | ( n19092 & ~n22500 ) ;
  assign n22502 = ( n13640 & ~n17211 ) | ( n13640 & n22501 ) | ( ~n17211 & n22501 ) ;
  assign n22503 = ( ~n1835 & n22498 ) | ( ~n1835 & n22502 ) | ( n22498 & n22502 ) ;
  assign n22504 = n6911 ^ n2271 ^ 1'b0 ;
  assign n22505 = n538 | n22504 ;
  assign n22506 = n13992 ^ n6021 ^ n3595 ;
  assign n22507 = ( n5106 & ~n11946 ) | ( n5106 & n22506 ) | ( ~n11946 & n22506 ) ;
  assign n22508 = n22507 ^ n12151 ^ n3244 ;
  assign n22509 = ( n3125 & ~n11526 ) | ( n3125 & n18360 ) | ( ~n11526 & n18360 ) ;
  assign n22510 = n19309 & ~n22509 ;
  assign n22511 = ( n22505 & n22508 ) | ( n22505 & ~n22510 ) | ( n22508 & ~n22510 ) ;
  assign n22512 = ( n5475 & n8712 ) | ( n5475 & n16855 ) | ( n8712 & n16855 ) ;
  assign n22513 = ( n15116 & n20101 ) | ( n15116 & n22512 ) | ( n20101 & n22512 ) ;
  assign n22514 = n271 | n10370 ;
  assign n22519 = ( ~x202 & n2075 ) | ( ~x202 & n3298 ) | ( n2075 & n3298 ) ;
  assign n22516 = n18114 ^ x134 ^ 1'b0 ;
  assign n22517 = n13609 & n22516 ;
  assign n22515 = ( n306 & n7197 ) | ( n306 & n8543 ) | ( n7197 & n8543 ) ;
  assign n22518 = n22517 ^ n22515 ^ n8167 ;
  assign n22520 = n22519 ^ n22518 ^ 1'b0 ;
  assign n22521 = ~n12379 & n22520 ;
  assign n22523 = ~n8037 & n9368 ;
  assign n22524 = ( n4175 & n8830 ) | ( n4175 & ~n19156 ) | ( n8830 & ~n19156 ) ;
  assign n22525 = n22524 ^ n10549 ^ 1'b0 ;
  assign n22526 = n6284 & n22525 ;
  assign n22527 = n14580 | n22526 ;
  assign n22528 = ( n1345 & n6645 ) | ( n1345 & ~n22527 ) | ( n6645 & ~n22527 ) ;
  assign n22529 = ( n12852 & n22523 ) | ( n12852 & ~n22528 ) | ( n22523 & ~n22528 ) ;
  assign n22522 = n7948 ^ n612 ^ 1'b0 ;
  assign n22530 = n22529 ^ n22522 ^ n4702 ;
  assign n22531 = ( n20446 & ~n22521 ) | ( n20446 & n22530 ) | ( ~n22521 & n22530 ) ;
  assign n22537 = ~n1017 & n10265 ;
  assign n22532 = n11336 & n12924 ;
  assign n22533 = n1995 & ~n22532 ;
  assign n22534 = n22533 ^ n9735 ^ 1'b0 ;
  assign n22535 = n22534 ^ n4159 ^ 1'b0 ;
  assign n22536 = n22535 ^ n4703 ^ 1'b0 ;
  assign n22538 = n22537 ^ n22536 ^ n12200 ;
  assign n22539 = n8085 & n12707 ;
  assign n22540 = ( n9339 & n10161 ) | ( n9339 & n11072 ) | ( n10161 & n11072 ) ;
  assign n22541 = ~n8585 & n22540 ;
  assign n22542 = n22539 & ~n22541 ;
  assign n22543 = ~n18194 & n18539 ;
  assign n22544 = n22543 ^ n5205 ^ 1'b0 ;
  assign n22545 = ( n4883 & n15167 ) | ( n4883 & n22544 ) | ( n15167 & n22544 ) ;
  assign n22546 = n8980 | n22545 ;
  assign n22547 = n2518 ^ n1530 ^ 1'b0 ;
  assign n22548 = n9516 & n22547 ;
  assign n22549 = n4106 & n21819 ;
  assign n22550 = n8246 & n22549 ;
  assign n22551 = ( n5830 & ~n8902 ) | ( n5830 & n13460 ) | ( ~n8902 & n13460 ) ;
  assign n22553 = n4460 ^ n4221 ^ 1'b0 ;
  assign n22552 = n7829 & ~n12052 ;
  assign n22554 = n22553 ^ n22552 ^ 1'b0 ;
  assign n22555 = n22554 ^ n17482 ^ n11365 ;
  assign n22556 = ( n2520 & n22551 ) | ( n2520 & n22555 ) | ( n22551 & n22555 ) ;
  assign n22557 = n9000 ^ n8697 ^ n3605 ;
  assign n22558 = n15808 & ~n22557 ;
  assign n22559 = n22556 & n22558 ;
  assign n22560 = n4796 ^ n274 ^ 1'b0 ;
  assign n22561 = n4396 | n22560 ;
  assign n22562 = ( ~n2590 & n4757 ) | ( ~n2590 & n17964 ) | ( n4757 & n17964 ) ;
  assign n22563 = ~n22561 & n22562 ;
  assign n22564 = n20308 ^ n6996 ^ 1'b0 ;
  assign n22565 = n22563 & ~n22564 ;
  assign n22569 = ( ~n4032 & n14127 ) | ( ~n4032 & n15416 ) | ( n14127 & n15416 ) ;
  assign n22566 = n1813 & ~n13361 ;
  assign n22567 = n22566 ^ n12909 ^ n9255 ;
  assign n22568 = ( ~n13597 & n15243 ) | ( ~n13597 & n22567 ) | ( n15243 & n22567 ) ;
  assign n22570 = n22569 ^ n22568 ^ n7227 ;
  assign n22571 = ( n2849 & n3553 ) | ( n2849 & n3894 ) | ( n3553 & n3894 ) ;
  assign n22572 = n5931 & n10334 ;
  assign n22573 = n22572 ^ n5445 ^ 1'b0 ;
  assign n22574 = ( n12952 & n22571 ) | ( n12952 & n22573 ) | ( n22571 & n22573 ) ;
  assign n22576 = n13775 ^ n12827 ^ 1'b0 ;
  assign n22575 = n10548 & n16385 ;
  assign n22577 = n22576 ^ n22575 ^ 1'b0 ;
  assign n22578 = ( n2052 & ~n9086 ) | ( n2052 & n15980 ) | ( ~n9086 & n15980 ) ;
  assign n22579 = ( ~n3510 & n20958 ) | ( ~n3510 & n22578 ) | ( n20958 & n22578 ) ;
  assign n22580 = ( ~n345 & n9171 ) | ( ~n345 & n22579 ) | ( n9171 & n22579 ) ;
  assign n22581 = n11107 ^ n8947 ^ 1'b0 ;
  assign n22582 = n15452 ^ n8001 ^ n3879 ;
  assign n22583 = ( n318 & n2286 ) | ( n318 & n22582 ) | ( n2286 & n22582 ) ;
  assign n22584 = n511 & n16203 ;
  assign n22585 = n5335 & n22584 ;
  assign n22586 = ~n15395 & n22585 ;
  assign n22587 = n4357 & ~n19978 ;
  assign n22588 = n11658 ^ n6833 ^ n1271 ;
  assign n22594 = n10947 ^ n2116 ^ 1'b0 ;
  assign n22595 = ( ~n2871 & n7938 ) | ( ~n2871 & n22594 ) | ( n7938 & n22594 ) ;
  assign n22589 = n10157 ^ n10152 ^ n7640 ;
  assign n22590 = n22186 ^ n10331 ^ 1'b0 ;
  assign n22591 = n1727 & n22590 ;
  assign n22592 = n22589 & n22591 ;
  assign n22593 = ~n3323 & n22592 ;
  assign n22596 = n22595 ^ n22593 ^ n16631 ;
  assign n22605 = n5452 ^ n846 ^ 1'b0 ;
  assign n22606 = n4910 & ~n22605 ;
  assign n22603 = n8171 ^ n5780 ^ x220 ;
  assign n22600 = ( ~n3551 & n3910 ) | ( ~n3551 & n9169 ) | ( n3910 & n9169 ) ;
  assign n22597 = n7384 ^ n6253 ^ 1'b0 ;
  assign n22598 = n1997 & ~n22597 ;
  assign n22599 = n22598 ^ n6680 ^ 1'b0 ;
  assign n22601 = n22600 ^ n22599 ^ 1'b0 ;
  assign n22602 = n2871 & n22601 ;
  assign n22604 = n22603 ^ n22602 ^ 1'b0 ;
  assign n22607 = n22606 ^ n22604 ^ n3592 ;
  assign n22608 = n17844 ^ n16152 ^ n1027 ;
  assign n22617 = n4969 ^ n3977 ^ n3819 ;
  assign n22618 = ~n16531 & n22617 ;
  assign n22619 = n22618 ^ n7562 ^ 1'b0 ;
  assign n22609 = n18653 ^ n4862 ^ 1'b0 ;
  assign n22610 = n13660 | n22609 ;
  assign n22611 = ( n1884 & n19946 ) | ( n1884 & ~n22610 ) | ( n19946 & ~n22610 ) ;
  assign n22613 = ( n4465 & n5445 ) | ( n4465 & ~n10114 ) | ( n5445 & ~n10114 ) ;
  assign n22614 = ( n838 & ~n2798 ) | ( n838 & n22613 ) | ( ~n2798 & n22613 ) ;
  assign n22612 = ~n6249 & n20476 ;
  assign n22615 = n22614 ^ n22612 ^ 1'b0 ;
  assign n22616 = n22611 & n22615 ;
  assign n22620 = n22619 ^ n22616 ^ 1'b0 ;
  assign n22631 = n20985 ^ n15175 ^ n5706 ;
  assign n22621 = ( n3331 & ~n4870 ) | ( n3331 & n13921 ) | ( ~n4870 & n13921 ) ;
  assign n22622 = ( n6124 & ~n6834 ) | ( n6124 & n22621 ) | ( ~n6834 & n22621 ) ;
  assign n22623 = n22622 ^ n13642 ^ n3838 ;
  assign n22624 = ( n7031 & ~n10823 ) | ( n7031 & n22623 ) | ( ~n10823 & n22623 ) ;
  assign n22625 = n8895 ^ n5241 ^ 1'b0 ;
  assign n22626 = ( n677 & n17081 ) | ( n677 & n22625 ) | ( n17081 & n22625 ) ;
  assign n22627 = n22626 ^ n8058 ^ 1'b0 ;
  assign n22628 = n4444 & ~n22627 ;
  assign n22629 = ( n5980 & ~n6919 ) | ( n5980 & n22628 ) | ( ~n6919 & n22628 ) ;
  assign n22630 = ( n8451 & n22624 ) | ( n8451 & ~n22629 ) | ( n22624 & ~n22629 ) ;
  assign n22632 = n22631 ^ n22630 ^ 1'b0 ;
  assign n22633 = n2779 | n22632 ;
  assign n22634 = n19831 ^ n14233 ^ n13466 ;
  assign n22635 = n13066 ^ n3178 ^ n2044 ;
  assign n22636 = n3853 & ~n22635 ;
  assign n22637 = ( ~n1204 & n11507 ) | ( ~n1204 & n16212 ) | ( n11507 & n16212 ) ;
  assign n22638 = ~n21886 & n22637 ;
  assign n22639 = ~n22636 & n22638 ;
  assign n22640 = ( n10474 & n10538 ) | ( n10474 & n15926 ) | ( n10538 & n15926 ) ;
  assign n22641 = x66 & n22640 ;
  assign n22642 = n18101 ^ n17304 ^ n1616 ;
  assign n22643 = n22642 ^ n20534 ^ 1'b0 ;
  assign n22644 = ~n15293 & n22643 ;
  assign n22645 = n22644 ^ n12272 ^ n860 ;
  assign n22646 = ( n7252 & ~n11338 ) | ( n7252 & n11745 ) | ( ~n11338 & n11745 ) ;
  assign n22647 = n11114 & n20313 ;
  assign n22648 = n22647 ^ n9691 ^ 1'b0 ;
  assign n22649 = ( ~n6298 & n22646 ) | ( ~n6298 & n22648 ) | ( n22646 & n22648 ) ;
  assign n22650 = n4366 ^ n3292 ^ n1009 ;
  assign n22651 = n22650 ^ n5672 ^ 1'b0 ;
  assign n22652 = ~n2521 & n22651 ;
  assign n22653 = n12773 ^ n9590 ^ n4337 ;
  assign n22654 = n7419 ^ n2525 ^ 1'b0 ;
  assign n22655 = ( n5618 & n21518 ) | ( n5618 & n22654 ) | ( n21518 & n22654 ) ;
  assign n22656 = ( ~n13131 & n22653 ) | ( ~n13131 & n22655 ) | ( n22653 & n22655 ) ;
  assign n22657 = n21023 ^ n19071 ^ 1'b0 ;
  assign n22658 = ~n13234 & n22163 ;
  assign n22659 = n22658 ^ n16581 ^ 1'b0 ;
  assign n22660 = n19850 ^ n9004 ^ 1'b0 ;
  assign n22661 = ~n7605 & n21352 ;
  assign n22662 = n21725 ^ n20672 ^ n15405 ;
  assign n22663 = n14950 ^ n10353 ^ 1'b0 ;
  assign n22664 = ~n3185 & n7449 ;
  assign n22665 = n22664 ^ x179 ^ 1'b0 ;
  assign n22666 = ( n9170 & n9358 ) | ( n9170 & n22665 ) | ( n9358 & n22665 ) ;
  assign n22667 = ( ~n6338 & n20062 ) | ( ~n6338 & n22666 ) | ( n20062 & n22666 ) ;
  assign n22668 = n22667 ^ n17241 ^ n7972 ;
  assign n22669 = n17748 ^ n14998 ^ n7888 ;
  assign n22670 = n9292 ^ n3849 ^ 1'b0 ;
  assign n22671 = ( n1599 & n3566 ) | ( n1599 & ~n22670 ) | ( n3566 & ~n22670 ) ;
  assign n22672 = n13733 ^ n8510 ^ n4472 ;
  assign n22673 = ~n22671 & n22672 ;
  assign n22674 = ( n6252 & n19358 ) | ( n6252 & ~n22673 ) | ( n19358 & ~n22673 ) ;
  assign n22675 = ( n1917 & n2376 ) | ( n1917 & ~n7987 ) | ( n2376 & ~n7987 ) ;
  assign n22676 = n10335 & ~n18786 ;
  assign n22677 = n22676 ^ n1845 ^ n1350 ;
  assign n22678 = ( n22613 & n22675 ) | ( n22613 & ~n22677 ) | ( n22675 & ~n22677 ) ;
  assign n22679 = n7039 | n8106 ;
  assign n22680 = n17155 | n22679 ;
  assign n22681 = ~n5858 & n15318 ;
  assign n22682 = n22681 ^ n4365 ^ 1'b0 ;
  assign n22683 = ~n15407 & n17370 ;
  assign n22684 = ~n22682 & n22683 ;
  assign n22685 = n15016 ^ n6245 ^ 1'b0 ;
  assign n22686 = ( n3628 & ~n9039 ) | ( n3628 & n11462 ) | ( ~n9039 & n11462 ) ;
  assign n22687 = n22686 ^ n7112 ^ 1'b0 ;
  assign n22688 = ~n14394 & n22687 ;
  assign n22689 = n22685 & n22688 ;
  assign n22690 = ( n5553 & ~n6088 ) | ( n5553 & n7066 ) | ( ~n6088 & n7066 ) ;
  assign n22691 = n22690 ^ n18638 ^ n17231 ;
  assign n22692 = n8663 | n18946 ;
  assign n22693 = n14523 & ~n22692 ;
  assign n22694 = n3169 & ~n11734 ;
  assign n22695 = n22694 ^ n7473 ^ 1'b0 ;
  assign n22696 = n8526 | n19548 ;
  assign n22697 = ( n4464 & n4691 ) | ( n4464 & ~n6994 ) | ( n4691 & ~n6994 ) ;
  assign n22698 = n22697 ^ n20567 ^ n8307 ;
  assign n22699 = n18171 ^ n15498 ^ n12376 ;
  assign n22701 = n20552 ^ n4926 ^ 1'b0 ;
  assign n22700 = ( ~n1594 & n9740 ) | ( ~n1594 & n13073 ) | ( n9740 & n13073 ) ;
  assign n22702 = n22701 ^ n22700 ^ n9331 ;
  assign n22703 = ( n1578 & ~n11716 ) | ( n1578 & n22702 ) | ( ~n11716 & n22702 ) ;
  assign n22704 = n772 | n18768 ;
  assign n22705 = n22704 ^ n9697 ^ 1'b0 ;
  assign n22706 = n20885 ^ n11485 ^ 1'b0 ;
  assign n22707 = ~n22705 & n22706 ;
  assign n22708 = n21525 ^ n8774 ^ n6535 ;
  assign n22709 = n22708 ^ n11178 ^ x173 ;
  assign n22710 = ( n1227 & n21420 ) | ( n1227 & n21664 ) | ( n21420 & n21664 ) ;
  assign n22711 = ( ~n3878 & n17278 ) | ( ~n3878 & n22710 ) | ( n17278 & n22710 ) ;
  assign n22712 = n5776 & ~n7968 ;
  assign n22713 = n1647 & n22712 ;
  assign n22718 = ( n4468 & n6980 ) | ( n4468 & n8537 ) | ( n6980 & n8537 ) ;
  assign n22714 = n9383 ^ n8505 ^ n4090 ;
  assign n22715 = n19078 ^ n5174 ^ 1'b0 ;
  assign n22716 = n7449 & ~n22715 ;
  assign n22717 = n22714 & n22716 ;
  assign n22719 = n22718 ^ n22717 ^ 1'b0 ;
  assign n22720 = ( n16757 & n22713 ) | ( n16757 & ~n22719 ) | ( n22713 & ~n22719 ) ;
  assign n22721 = n14508 | n22720 ;
  assign n22722 = n22721 ^ n993 ^ 1'b0 ;
  assign n22723 = ( n1947 & n12560 ) | ( n1947 & n22434 ) | ( n12560 & n22434 ) ;
  assign n22725 = n2979 & n19941 ;
  assign n22726 = n22725 ^ n14731 ^ n1729 ;
  assign n22727 = n22726 ^ n606 ^ 1'b0 ;
  assign n22724 = ( ~n2614 & n9385 ) | ( ~n2614 & n12427 ) | ( n9385 & n12427 ) ;
  assign n22728 = n22727 ^ n22724 ^ 1'b0 ;
  assign n22729 = n22728 ^ n14988 ^ 1'b0 ;
  assign n22730 = ~x10 & n16216 ;
  assign n22731 = ( n7188 & n13709 ) | ( n7188 & n22730 ) | ( n13709 & n22730 ) ;
  assign n22732 = n15475 ^ n3769 ^ 1'b0 ;
  assign n22733 = ~n7527 & n22732 ;
  assign n22734 = n3034 | n13698 ;
  assign n22735 = n22733 | n22734 ;
  assign n22736 = n5326 & ~n22735 ;
  assign n22737 = ( n3171 & ~n7154 ) | ( n3171 & n8953 ) | ( ~n7154 & n8953 ) ;
  assign n22738 = ( n1893 & n7207 ) | ( n1893 & n22737 ) | ( n7207 & n22737 ) ;
  assign n22739 = x76 & ~n7279 ;
  assign n22740 = n17336 ^ n958 ^ n482 ;
  assign n22741 = ( n7905 & n22739 ) | ( n7905 & n22740 ) | ( n22739 & n22740 ) ;
  assign n22742 = ( ~n1264 & n2995 ) | ( ~n1264 & n3922 ) | ( n2995 & n3922 ) ;
  assign n22743 = n22742 ^ n20765 ^ n821 ;
  assign n22744 = n1477 & ~n22743 ;
  assign n22745 = n22744 ^ n17458 ^ 1'b0 ;
  assign n22746 = n22745 ^ n17210 ^ n8087 ;
  assign n22747 = n1898 & n21448 ;
  assign n22748 = n5918 | n22747 ;
  assign n22749 = n22748 ^ n20376 ^ 1'b0 ;
  assign n22750 = n10381 | n16432 ;
  assign n22751 = n2586 & n22750 ;
  assign n22752 = ~n11558 & n22751 ;
  assign n22753 = ( n9403 & n17496 ) | ( n9403 & n22752 ) | ( n17496 & n22752 ) ;
  assign n22754 = ( ~n1924 & n5297 ) | ( ~n1924 & n14793 ) | ( n5297 & n14793 ) ;
  assign n22755 = n22754 ^ n650 ^ 1'b0 ;
  assign n22756 = n8606 & n22755 ;
  assign n22757 = n22756 ^ n19385 ^ n18905 ;
  assign n22758 = n15591 ^ n12443 ^ n4866 ;
  assign n22759 = n15002 ^ n8956 ^ 1'b0 ;
  assign n22760 = n6886 | n22759 ;
  assign n22761 = n7365 | n22760 ;
  assign n22762 = n10814 | n22761 ;
  assign n22763 = ( ~n1189 & n11695 ) | ( ~n1189 & n22762 ) | ( n11695 & n22762 ) ;
  assign n22764 = n22763 ^ n19739 ^ n3729 ;
  assign n22765 = ~n673 & n1168 ;
  assign n22766 = n22765 ^ n14934 ^ 1'b0 ;
  assign n22767 = n12484 | n22766 ;
  assign n22768 = n22767 ^ n897 ^ 1'b0 ;
  assign n22769 = n6908 & ~n22768 ;
  assign n22770 = ( n5833 & n21060 ) | ( n5833 & ~n22769 ) | ( n21060 & ~n22769 ) ;
  assign n22771 = n22770 ^ n14773 ^ n13639 ;
  assign n22772 = n5744 | n10065 ;
  assign n22773 = n22772 ^ x137 ^ 1'b0 ;
  assign n22774 = n15113 & ~n15756 ;
  assign n22775 = n22774 ^ n7885 ^ 1'b0 ;
  assign n22776 = n15543 ^ n2931 ^ 1'b0 ;
  assign n22777 = n8676 ^ n3221 ^ 1'b0 ;
  assign n22778 = ( n2192 & n7267 ) | ( n2192 & ~n11507 ) | ( n7267 & ~n11507 ) ;
  assign n22779 = n1632 | n17561 ;
  assign n22780 = ( ~n22777 & n22778 ) | ( ~n22777 & n22779 ) | ( n22778 & n22779 ) ;
  assign n22781 = ~n17864 & n22780 ;
  assign n22782 = ( n11916 & n22776 ) | ( n11916 & ~n22781 ) | ( n22776 & ~n22781 ) ;
  assign n22786 = n14669 ^ n11751 ^ 1'b0 ;
  assign n22787 = n13641 & n22786 ;
  assign n22788 = ( n10384 & ~n18120 ) | ( n10384 & n22787 ) | ( ~n18120 & n22787 ) ;
  assign n22783 = n8087 ^ n1436 ^ 1'b0 ;
  assign n22784 = n14382 ^ n5774 ^ 1'b0 ;
  assign n22785 = n22783 | n22784 ;
  assign n22789 = n22788 ^ n22785 ^ n1824 ;
  assign n22790 = n11397 ^ n10549 ^ n1007 ;
  assign n22791 = n22790 ^ n16356 ^ n11599 ;
  assign n22792 = n17227 ^ n12914 ^ 1'b0 ;
  assign n22793 = n2856 & n22792 ;
  assign n22794 = n9396 ^ n3690 ^ n1809 ;
  assign n22795 = n21162 ^ n13991 ^ n11956 ;
  assign n22796 = n537 & n16936 ;
  assign n22797 = n22796 ^ n11942 ^ 1'b0 ;
  assign n22798 = ( n11764 & n22795 ) | ( n11764 & n22797 ) | ( n22795 & n22797 ) ;
  assign n22799 = x57 & ~n10402 ;
  assign n22802 = n12064 ^ n1257 ^ 1'b0 ;
  assign n22803 = n16439 ^ n9956 ^ 1'b0 ;
  assign n22804 = n22802 & n22803 ;
  assign n22800 = n1400 & n18261 ;
  assign n22801 = n22800 ^ n9521 ^ 1'b0 ;
  assign n22805 = n22804 ^ n22801 ^ n2594 ;
  assign n22806 = n19217 ^ n6171 ^ 1'b0 ;
  assign n22807 = ~n6437 & n22806 ;
  assign n22808 = ( n11730 & n13092 ) | ( n11730 & n22807 ) | ( n13092 & n22807 ) ;
  assign n22809 = ~n3857 & n6299 ;
  assign n22810 = ( ~n7547 & n22506 ) | ( ~n7547 & n22809 ) | ( n22506 & n22809 ) ;
  assign n22811 = n16272 ^ n513 ^ 1'b0 ;
  assign n22812 = n22811 ^ n6834 ^ n5829 ;
  assign n22813 = n20728 & n22812 ;
  assign n22814 = ~n10464 & n22813 ;
  assign n22815 = n10404 | n13413 ;
  assign n22816 = n15032 ^ n6038 ^ 1'b0 ;
  assign n22818 = n16612 ^ n3386 ^ 1'b0 ;
  assign n22819 = ~n7798 & n22818 ;
  assign n22817 = x111 & ~n17801 ;
  assign n22820 = n22819 ^ n22817 ^ 1'b0 ;
  assign n22821 = ~n22816 & n22820 ;
  assign n22823 = ~n1106 & n18159 ;
  assign n22824 = n22823 ^ n13037 ^ 1'b0 ;
  assign n22822 = n13012 ^ n7955 ^ n4924 ;
  assign n22825 = n22824 ^ n22822 ^ n14413 ;
  assign n22826 = n22825 ^ n19934 ^ 1'b0 ;
  assign n22827 = n12675 & n22826 ;
  assign n22828 = ( n5227 & n6521 ) | ( n5227 & ~n15331 ) | ( n6521 & ~n15331 ) ;
  assign n22829 = ( n2268 & ~n14364 ) | ( n2268 & n16838 ) | ( ~n14364 & n16838 ) ;
  assign n22833 = x75 & ~n10711 ;
  assign n22834 = n3581 & n22833 ;
  assign n22835 = n22834 ^ n10516 ^ 1'b0 ;
  assign n22832 = n11573 ^ n7530 ^ n2797 ;
  assign n22830 = n21248 ^ n10513 ^ 1'b0 ;
  assign n22831 = n22830 ^ n3158 ^ n367 ;
  assign n22836 = n22835 ^ n22832 ^ n22831 ;
  assign n22837 = ~n14706 & n22836 ;
  assign n22838 = ~n2745 & n22837 ;
  assign n22839 = ( n4179 & n5142 ) | ( n4179 & n11908 ) | ( n5142 & n11908 ) ;
  assign n22841 = n6470 ^ n3673 ^ n3238 ;
  assign n22842 = ( n2113 & ~n7388 ) | ( n2113 & n22841 ) | ( ~n7388 & n22841 ) ;
  assign n22843 = ( n15507 & n21236 ) | ( n15507 & n22842 ) | ( n21236 & n22842 ) ;
  assign n22840 = ~n1657 & n13883 ;
  assign n22844 = n22843 ^ n22840 ^ 1'b0 ;
  assign n22845 = ~n13639 & n22844 ;
  assign n22846 = n17523 ^ n16246 ^ 1'b0 ;
  assign n22847 = ~n16826 & n22846 ;
  assign n22848 = n8854 ^ n7169 ^ n6603 ;
  assign n22849 = ~n12388 & n22848 ;
  assign n22850 = n21980 ^ n11265 ^ n5344 ;
  assign n22851 = ( n13111 & n22523 ) | ( n13111 & n22850 ) | ( n22523 & n22850 ) ;
  assign n22861 = ~x71 & n13625 ;
  assign n22862 = n22861 ^ n11313 ^ 1'b0 ;
  assign n22860 = n1514 ^ x29 ^ 1'b0 ;
  assign n22857 = n14047 ^ n6687 ^ 1'b0 ;
  assign n22858 = n7027 & ~n22857 ;
  assign n22855 = n13696 ^ n9481 ^ 1'b0 ;
  assign n22856 = n3632 & n22855 ;
  assign n22859 = n22858 ^ n22856 ^ 1'b0 ;
  assign n22863 = n22862 ^ n22860 ^ n22859 ;
  assign n22852 = n21298 ^ n6122 ^ 1'b0 ;
  assign n22853 = n10227 & n22852 ;
  assign n22854 = ( n5265 & n15175 ) | ( n5265 & n22853 ) | ( n15175 & n22853 ) ;
  assign n22864 = n22863 ^ n22854 ^ n14359 ;
  assign n22865 = n13371 ^ n10060 ^ n2224 ;
  assign n22866 = n22865 ^ n16767 ^ 1'b0 ;
  assign n22870 = n2076 ^ n1503 ^ 1'b0 ;
  assign n22869 = n14665 ^ n8458 ^ n2540 ;
  assign n22867 = n2176 & ~n5563 ;
  assign n22868 = n22867 ^ n14528 ^ 1'b0 ;
  assign n22871 = n22870 ^ n22869 ^ n22868 ;
  assign n22872 = n15716 ^ n7691 ^ 1'b0 ;
  assign n22873 = ( ~n9558 & n20230 ) | ( ~n9558 & n22872 ) | ( n20230 & n22872 ) ;
  assign n22874 = ( n11192 & ~n12404 ) | ( n11192 & n17822 ) | ( ~n12404 & n17822 ) ;
  assign n22875 = ~n3458 & n22874 ;
  assign n22876 = ~n6284 & n22875 ;
  assign n22877 = ( n2732 & n4064 ) | ( n2732 & ~n6230 ) | ( n4064 & ~n6230 ) ;
  assign n22878 = n22877 ^ n21426 ^ n13417 ;
  assign n22879 = ( ~n2676 & n5132 ) | ( ~n2676 & n7328 ) | ( n5132 & n7328 ) ;
  assign n22880 = n15592 & ~n22879 ;
  assign n22881 = n13212 ^ n3253 ^ 1'b0 ;
  assign n22882 = n4398 ^ n2353 ^ n1464 ;
  assign n22883 = n18688 ^ n3906 ^ 1'b0 ;
  assign n22884 = n22882 | n22883 ;
  assign n22885 = n22881 & ~n22884 ;
  assign n22886 = ( ~n14195 & n17739 ) | ( ~n14195 & n22885 ) | ( n17739 & n22885 ) ;
  assign n22887 = n10033 & n20943 ;
  assign n22888 = ( n12419 & n19271 ) | ( n12419 & n22887 ) | ( n19271 & n22887 ) ;
  assign n22889 = ( ~n10222 & n15199 ) | ( ~n10222 & n22888 ) | ( n15199 & n22888 ) ;
  assign n22891 = n18079 ^ n8189 ^ 1'b0 ;
  assign n22890 = n16836 ^ n10223 ^ n8941 ;
  assign n22892 = n22891 ^ n22890 ^ 1'b0 ;
  assign n22893 = n13815 & ~n15431 ;
  assign n22894 = n15133 & ~n19588 ;
  assign n22895 = ( n3408 & n14859 ) | ( n3408 & ~n22894 ) | ( n14859 & ~n22894 ) ;
  assign n22896 = ( n8128 & ~n10477 ) | ( n8128 & n15949 ) | ( ~n10477 & n15949 ) ;
  assign n22899 = n1156 & ~n1500 ;
  assign n22897 = n7098 & ~n7415 ;
  assign n22898 = ~n7273 & n22897 ;
  assign n22900 = n22899 ^ n22898 ^ n3366 ;
  assign n22901 = n22900 ^ n14252 ^ 1'b0 ;
  assign n22902 = ( n1236 & n5910 ) | ( n1236 & n22901 ) | ( n5910 & n22901 ) ;
  assign n22903 = n9067 ^ n4684 ^ 1'b0 ;
  assign n22904 = n6685 & ~n22903 ;
  assign n22905 = n22904 ^ n15827 ^ n12206 ;
  assign n22906 = ( n2428 & ~n15361 ) | ( n2428 & n22905 ) | ( ~n15361 & n22905 ) ;
  assign n22907 = n17387 ^ n14459 ^ n2939 ;
  assign n22908 = n22907 ^ n13017 ^ n3733 ;
  assign n22909 = n22332 ^ n22025 ^ n3267 ;
  assign n22910 = n785 | n13866 ;
  assign n22911 = n22909 | n22910 ;
  assign n22912 = n5955 ^ x114 ^ 1'b0 ;
  assign n22913 = n3245 ^ n2539 ^ 1'b0 ;
  assign n22914 = ( n5519 & n21262 ) | ( n5519 & ~n22913 ) | ( n21262 & ~n22913 ) ;
  assign n22915 = ( n8267 & ~n14628 ) | ( n8267 & n18569 ) | ( ~n14628 & n18569 ) ;
  assign n22916 = n22915 ^ n8814 ^ n488 ;
  assign n22917 = n4418 | n22916 ;
  assign n22918 = n22917 ^ n5467 ^ 1'b0 ;
  assign n22928 = n15192 ^ n8803 ^ n4557 ;
  assign n22919 = ( n1376 & n5102 ) | ( n1376 & n6242 ) | ( n5102 & n6242 ) ;
  assign n22922 = ( n1619 & ~n3319 ) | ( n1619 & n10856 ) | ( ~n3319 & n10856 ) ;
  assign n22920 = n3316 & ~n7757 ;
  assign n22921 = n22920 ^ n15383 ^ x102 ;
  assign n22923 = n22922 ^ n22921 ^ 1'b0 ;
  assign n22924 = n22923 ^ n13665 ^ 1'b0 ;
  assign n22925 = n14340 | n22924 ;
  assign n22926 = n22919 & ~n22925 ;
  assign n22927 = ~n6200 & n22926 ;
  assign n22929 = n22928 ^ n22927 ^ 1'b0 ;
  assign n22931 = n9614 ^ x146 ^ 1'b0 ;
  assign n22930 = ( n327 & n1663 ) | ( n327 & ~n1748 ) | ( n1663 & ~n1748 ) ;
  assign n22932 = n22931 ^ n22930 ^ n5084 ;
  assign n22933 = n17877 ^ n15883 ^ 1'b0 ;
  assign n22934 = n22932 | n22933 ;
  assign n22935 = n22934 ^ n5705 ^ 1'b0 ;
  assign n22936 = n22935 ^ n19179 ^ n14857 ;
  assign n22937 = n20086 ^ n1958 ^ n1753 ;
  assign n22938 = n15218 & ~n22937 ;
  assign n22939 = n22938 ^ n5614 ^ 1'b0 ;
  assign n22943 = n7764 & ~n13369 ;
  assign n22940 = ( n4967 & n7909 ) | ( n4967 & n16567 ) | ( n7909 & n16567 ) ;
  assign n22941 = n11579 | n22940 ;
  assign n22942 = ( ~n6813 & n14296 ) | ( ~n6813 & n22941 ) | ( n14296 & n22941 ) ;
  assign n22944 = n22943 ^ n22942 ^ 1'b0 ;
  assign n22945 = n5911 & n11860 ;
  assign n22947 = n7738 ^ n7065 ^ n6316 ;
  assign n22946 = n13562 | n16567 ;
  assign n22948 = n22947 ^ n22946 ^ 1'b0 ;
  assign n22949 = ( ~n3572 & n18010 ) | ( ~n3572 & n22948 ) | ( n18010 & n22948 ) ;
  assign n22950 = n22949 ^ n18962 ^ 1'b0 ;
  assign n22951 = n9586 ^ n3757 ^ 1'b0 ;
  assign n22952 = x250 & ~n22951 ;
  assign n22953 = ( n6199 & n13482 ) | ( n6199 & ~n22952 ) | ( n13482 & ~n22952 ) ;
  assign n22954 = n22953 ^ n6571 ^ n6231 ;
  assign n22955 = n5613 ^ n264 ^ 1'b0 ;
  assign n22956 = ( n8916 & n11021 ) | ( n8916 & n22955 ) | ( n11021 & n22955 ) ;
  assign n22957 = n18835 ^ n17387 ^ n1616 ;
  assign n22958 = n22957 ^ n6503 ^ n5933 ;
  assign n22959 = n13058 ^ n10859 ^ 1'b0 ;
  assign n22960 = n22900 ^ n15004 ^ n7475 ;
  assign n22961 = n22959 | n22960 ;
  assign n22962 = n22877 & ~n22961 ;
  assign n22963 = n22962 ^ n19962 ^ n4445 ;
  assign n22964 = ( n3126 & ~n3492 ) | ( n3126 & n6259 ) | ( ~n3492 & n6259 ) ;
  assign n22965 = n22964 ^ n3800 ^ 1'b0 ;
  assign n22966 = n8981 & n22965 ;
  assign n22967 = n8981 ^ n783 ^ 1'b0 ;
  assign n22968 = ~n20135 & n22967 ;
  assign n22969 = ( ~n817 & n3404 ) | ( ~n817 & n6148 ) | ( n3404 & n6148 ) ;
  assign n22970 = n2996 | n22969 ;
  assign n22971 = n16586 ^ n10096 ^ 1'b0 ;
  assign n22972 = n22971 ^ n17900 ^ n15269 ;
  assign n22973 = n530 | n22972 ;
  assign n22974 = n22973 ^ n11802 ^ 1'b0 ;
  assign n22975 = n8448 ^ n2353 ^ 1'b0 ;
  assign n22976 = n7934 ^ n6391 ^ 1'b0 ;
  assign n22977 = n22975 | n22976 ;
  assign n22978 = n13387 ^ n7959 ^ 1'b0 ;
  assign n22979 = n7862 & ~n22978 ;
  assign n22980 = ( n3735 & ~n9718 ) | ( n3735 & n22979 ) | ( ~n9718 & n22979 ) ;
  assign n22981 = ( n8908 & ~n9361 ) | ( n8908 & n17323 ) | ( ~n9361 & n17323 ) ;
  assign n22982 = ( n4147 & n8882 ) | ( n4147 & ~n22981 ) | ( n8882 & ~n22981 ) ;
  assign n22983 = n6654 ^ n3966 ^ 1'b0 ;
  assign n22984 = ( n7727 & n22982 ) | ( n7727 & n22983 ) | ( n22982 & n22983 ) ;
  assign n22986 = n11236 | n16823 ;
  assign n22987 = n12142 & ~n22986 ;
  assign n22985 = ( n1017 & ~n13800 ) | ( n1017 & n22391 ) | ( ~n13800 & n22391 ) ;
  assign n22988 = n22987 ^ n22985 ^ n11167 ;
  assign n22989 = n9530 ^ n4223 ^ n342 ;
  assign n22990 = ( n10309 & n12337 ) | ( n10309 & n22989 ) | ( n12337 & n22989 ) ;
  assign n22991 = n21483 ^ n17873 ^ 1'b0 ;
  assign n22992 = ( ~n592 & n5092 ) | ( ~n592 & n14122 ) | ( n5092 & n14122 ) ;
  assign n22993 = n22991 | n22992 ;
  assign n22994 = n20870 & ~n22993 ;
  assign n22995 = n20389 ^ x5 ^ 1'b0 ;
  assign n22996 = x82 & ~n22995 ;
  assign n22997 = ~n8977 & n22996 ;
  assign n22998 = ( n8790 & ~n12136 ) | ( n8790 & n22997 ) | ( ~n12136 & n22997 ) ;
  assign n22999 = n3715 & n11426 ;
  assign n23004 = n15010 ^ n974 ^ 1'b0 ;
  assign n23000 = ( n8466 & n13319 ) | ( n8466 & n21854 ) | ( n13319 & n21854 ) ;
  assign n23001 = n12630 ^ n3008 ^ 1'b0 ;
  assign n23002 = n19309 & ~n23001 ;
  assign n23003 = n23000 & n23002 ;
  assign n23005 = n23004 ^ n23003 ^ n3580 ;
  assign n23006 = n2955 | n12744 ;
  assign n23007 = n12695 ^ n12010 ^ 1'b0 ;
  assign n23008 = n9879 & n23007 ;
  assign n23009 = ( n2925 & ~n12034 ) | ( n2925 & n12991 ) | ( ~n12034 & n12991 ) ;
  assign n23010 = ( n9677 & ~n17513 ) | ( n9677 & n20985 ) | ( ~n17513 & n20985 ) ;
  assign n23011 = ( n9146 & n12936 ) | ( n9146 & n23010 ) | ( n12936 & n23010 ) ;
  assign n23012 = n6436 ^ n2955 ^ 1'b0 ;
  assign n23013 = ~n23011 & n23012 ;
  assign n23014 = ( n13747 & n18886 ) | ( n13747 & n23013 ) | ( n18886 & n23013 ) ;
  assign n23015 = n12995 ^ n8474 ^ 1'b0 ;
  assign n23016 = n15478 ^ n13878 ^ n5192 ;
  assign n23017 = n23016 ^ n16574 ^ n13983 ;
  assign n23018 = n11442 ^ n2210 ^ n1340 ;
  assign n23019 = n5249 ^ n706 ^ 1'b0 ;
  assign n23020 = ~n23018 & n23019 ;
  assign n23021 = n23017 & n23020 ;
  assign n23022 = n16379 & ~n18325 ;
  assign n23023 = n23022 ^ n14800 ^ 1'b0 ;
  assign n23024 = n5340 & ~n23023 ;
  assign n23025 = ~n23021 & n23024 ;
  assign n23026 = n22964 ^ n20182 ^ n11450 ;
  assign n23027 = n23026 ^ n15316 ^ n11529 ;
  assign n23028 = ~n9691 & n18029 ;
  assign n23029 = n23028 ^ n14399 ^ 1'b0 ;
  assign n23031 = x97 & n17088 ;
  assign n23032 = n23031 ^ n6019 ^ 1'b0 ;
  assign n23030 = n14444 ^ n13387 ^ n6960 ;
  assign n23033 = n23032 ^ n23030 ^ n14374 ;
  assign n23034 = n17262 ^ n14537 ^ 1'b0 ;
  assign n23035 = n23033 | n23034 ;
  assign n23036 = n6861 & n20112 ;
  assign n23037 = n23036 ^ n11030 ^ n4089 ;
  assign n23038 = n18659 & ~n23037 ;
  assign n23039 = n12236 & n23038 ;
  assign n23040 = ( n12260 & n12577 ) | ( n12260 & ~n13582 ) | ( n12577 & ~n13582 ) ;
  assign n23041 = n14742 ^ n1101 ^ 1'b0 ;
  assign n23042 = ( n1905 & ~n23040 ) | ( n1905 & n23041 ) | ( ~n23040 & n23041 ) ;
  assign n23043 = n17521 ^ n9044 ^ 1'b0 ;
  assign n23044 = n948 | n23043 ;
  assign n23045 = n4126 ^ n3523 ^ 1'b0 ;
  assign n23046 = ~n1807 & n4579 ;
  assign n23047 = n23046 ^ n10235 ^ 1'b0 ;
  assign n23048 = ( n2240 & n3048 ) | ( n2240 & ~n23047 ) | ( n3048 & ~n23047 ) ;
  assign n23049 = ( ~n5951 & n6398 ) | ( ~n5951 & n7858 ) | ( n6398 & n7858 ) ;
  assign n23050 = ~n352 & n11976 ;
  assign n23051 = ~n21804 & n23050 ;
  assign n23052 = ( n20558 & ~n23049 ) | ( n20558 & n23051 ) | ( ~n23049 & n23051 ) ;
  assign n23053 = n23052 ^ n21685 ^ n18058 ;
  assign n23054 = ( n10356 & n23048 ) | ( n10356 & n23053 ) | ( n23048 & n23053 ) ;
  assign n23057 = n14917 ^ n10432 ^ n574 ;
  assign n23058 = n1099 | n23057 ;
  assign n23055 = n13342 ^ n1418 ^ 1'b0 ;
  assign n23056 = n11769 | n23055 ;
  assign n23059 = n23058 ^ n23056 ^ n21509 ;
  assign n23060 = ( ~n3270 & n17217 ) | ( ~n3270 & n17810 ) | ( n17217 & n17810 ) ;
  assign n23061 = n4554 ^ n3363 ^ n1666 ;
  assign n23062 = n21405 & ~n23061 ;
  assign n23063 = n23062 ^ n12726 ^ 1'b0 ;
  assign n23064 = n21859 ^ n17513 ^ n1140 ;
  assign n23067 = n7442 ^ n4774 ^ n379 ;
  assign n23068 = ( n1680 & n3542 ) | ( n1680 & n23067 ) | ( n3542 & n23067 ) ;
  assign n23066 = n15317 ^ n13888 ^ n1850 ;
  assign n23069 = n23068 ^ n23066 ^ 1'b0 ;
  assign n23065 = n19614 ^ n9412 ^ n7867 ;
  assign n23070 = n23069 ^ n23065 ^ n13200 ;
  assign n23071 = n23070 ^ n16166 ^ n9428 ;
  assign n23072 = n4837 | n18149 ;
  assign n23073 = n16726 | n23072 ;
  assign n23074 = n4234 ^ n2113 ^ 1'b0 ;
  assign n23075 = n20307 ^ n20100 ^ 1'b0 ;
  assign n23076 = n23074 & ~n23075 ;
  assign n23077 = n18592 ^ n6088 ^ 1'b0 ;
  assign n23078 = n23076 & n23077 ;
  assign n23085 = n7362 & ~n13500 ;
  assign n23081 = n6364 ^ n6052 ^ n2036 ;
  assign n23082 = ( n3927 & n19106 ) | ( n3927 & n23081 ) | ( n19106 & n23081 ) ;
  assign n23083 = n15905 & n23082 ;
  assign n23084 = n19640 & n23083 ;
  assign n23079 = n9144 ^ n2189 ^ 1'b0 ;
  assign n23080 = n23079 ^ n21083 ^ n1561 ;
  assign n23086 = n23085 ^ n23084 ^ n23080 ;
  assign n23092 = n14410 & ~n15825 ;
  assign n23093 = ~n8239 & n23092 ;
  assign n23091 = n21604 ^ n8411 ^ n1126 ;
  assign n23087 = n9530 ^ n5878 ^ 1'b0 ;
  assign n23088 = ( n5533 & ~n16996 ) | ( n5533 & n23087 ) | ( ~n16996 & n23087 ) ;
  assign n23089 = n23088 ^ n12988 ^ n10374 ;
  assign n23090 = ( n6242 & n13983 ) | ( n6242 & ~n23089 ) | ( n13983 & ~n23089 ) ;
  assign n23094 = n23093 ^ n23091 ^ n23090 ;
  assign n23095 = ~n843 & n9102 ;
  assign n23096 = n11927 | n23095 ;
  assign n23097 = n11160 | n23096 ;
  assign n23098 = ( n1707 & n12499 ) | ( n1707 & n20271 ) | ( n12499 & n20271 ) ;
  assign n23099 = n21458 & ~n23098 ;
  assign n23100 = ( ~n3173 & n3719 ) | ( ~n3173 & n23099 ) | ( n3719 & n23099 ) ;
  assign n23101 = n12826 ^ n8574 ^ n750 ;
  assign n23102 = n8519 & n16892 ;
  assign n23103 = n2548 & ~n23102 ;
  assign n23104 = n23103 ^ n5074 ^ n2550 ;
  assign n23105 = n5192 | n13194 ;
  assign n23106 = ( n505 & n3347 ) | ( n505 & ~n3449 ) | ( n3347 & ~n3449 ) ;
  assign n23107 = n23106 ^ n3794 ^ 1'b0 ;
  assign n23108 = n10419 & ~n23107 ;
  assign n23109 = n2124 & n17879 ;
  assign n23110 = ~n17425 & n23109 ;
  assign n23111 = ~n5663 & n7488 ;
  assign n23112 = n23111 ^ n18538 ^ 1'b0 ;
  assign n23113 = ~n11513 & n22881 ;
  assign n23114 = n23113 ^ n19110 ^ 1'b0 ;
  assign n23115 = n18431 & n23114 ;
  assign n23116 = n17392 & ~n23115 ;
  assign n23117 = n23116 ^ n20268 ^ 1'b0 ;
  assign n23123 = x51 & n12170 ;
  assign n23124 = n23123 ^ n14355 ^ n3879 ;
  assign n23122 = n1383 & n20477 ;
  assign n23125 = n23124 ^ n23122 ^ 1'b0 ;
  assign n23126 = n2833 & n14080 ;
  assign n23127 = n23125 & n23126 ;
  assign n23118 = n2691 | n6938 ;
  assign n23119 = n2365 | n23118 ;
  assign n23120 = n23119 ^ n8455 ^ n8158 ;
  assign n23121 = n23120 ^ n15560 ^ 1'b0 ;
  assign n23128 = n23127 ^ n23121 ^ n13813 ;
  assign n23130 = n15533 ^ n14304 ^ 1'b0 ;
  assign n23129 = n12440 ^ n10277 ^ n5527 ;
  assign n23131 = n23130 ^ n23129 ^ n10881 ;
  assign n23134 = n12901 ^ n7809 ^ n6875 ;
  assign n23135 = n23134 ^ n10701 ^ n2516 ;
  assign n23132 = n15616 ^ x7 ^ 1'b0 ;
  assign n23133 = n4009 & n23132 ;
  assign n23136 = n23135 ^ n23133 ^ n7810 ;
  assign n23137 = ( n1215 & n18631 ) | ( n1215 & n23136 ) | ( n18631 & n23136 ) ;
  assign n23138 = ~n4959 & n19274 ;
  assign n23139 = ( n8601 & n11904 ) | ( n8601 & ~n23138 ) | ( n11904 & ~n23138 ) ;
  assign n23140 = ( n6389 & n8252 ) | ( n6389 & ~n19203 ) | ( n8252 & ~n19203 ) ;
  assign n23141 = n8617 ^ n1511 ^ 1'b0 ;
  assign n23142 = n4145 & ~n8053 ;
  assign n23143 = n1200 & n23142 ;
  assign n23144 = ( ~x97 & n546 ) | ( ~x97 & n2455 ) | ( n546 & n2455 ) ;
  assign n23145 = ( n23141 & n23143 ) | ( n23141 & n23144 ) | ( n23143 & n23144 ) ;
  assign n23146 = n4336 & n22996 ;
  assign n23147 = x242 & n3126 ;
  assign n23148 = ( n20462 & n21083 ) | ( n20462 & n23147 ) | ( n21083 & n23147 ) ;
  assign n23152 = ( n6523 & ~n13747 ) | ( n6523 & n18388 ) | ( ~n13747 & n18388 ) ;
  assign n23150 = ( n3162 & ~n9901 ) | ( n3162 & n18341 ) | ( ~n9901 & n18341 ) ;
  assign n23149 = ( ~n6124 & n6475 ) | ( ~n6124 & n8374 ) | ( n6475 & n8374 ) ;
  assign n23151 = n23150 ^ n23149 ^ 1'b0 ;
  assign n23153 = n23152 ^ n23151 ^ 1'b0 ;
  assign n23154 = n23148 & ~n23153 ;
  assign n23155 = n10032 ^ n9594 ^ n5304 ;
  assign n23156 = ( n2290 & n12049 ) | ( n2290 & ~n14736 ) | ( n12049 & ~n14736 ) ;
  assign n23157 = n23156 ^ n11493 ^ n7404 ;
  assign n23158 = ~n2823 & n23157 ;
  assign n23159 = n19044 ^ n2804 ^ n1914 ;
  assign n23160 = ( n12728 & n15252 ) | ( n12728 & n23159 ) | ( n15252 & n23159 ) ;
  assign n23161 = n10685 & ~n12188 ;
  assign n23162 = ( n1579 & n3021 ) | ( n1579 & n23161 ) | ( n3021 & n23161 ) ;
  assign n23163 = n23162 ^ n4306 ^ n2137 ;
  assign n23164 = n23163 ^ n15825 ^ x5 ;
  assign n23171 = ~n2965 & n3626 ;
  assign n23172 = n1299 & n23171 ;
  assign n23170 = ( n799 & n13310 ) | ( n799 & ~n15510 ) | ( n13310 & ~n15510 ) ;
  assign n23173 = n23172 ^ n23170 ^ 1'b0 ;
  assign n23174 = n3628 & ~n23173 ;
  assign n23175 = n11976 & n23174 ;
  assign n23169 = n7736 ^ n4791 ^ n3605 ;
  assign n23165 = n12510 ^ n6736 ^ 1'b0 ;
  assign n23166 = n7445 & ~n23165 ;
  assign n23167 = n7870 ^ n1378 ^ 1'b0 ;
  assign n23168 = n23166 & ~n23167 ;
  assign n23176 = n23175 ^ n23169 ^ n23168 ;
  assign n23177 = n4697 ^ n2644 ^ 1'b0 ;
  assign n23178 = n3763 & n23177 ;
  assign n23179 = n9519 & n23178 ;
  assign n23180 = n23179 ^ n22745 ^ 1'b0 ;
  assign n23181 = n9574 ^ n1799 ^ 1'b0 ;
  assign n23182 = n2096 | n23181 ;
  assign n23183 = ( n10189 & n17397 ) | ( n10189 & ~n23182 ) | ( n17397 & ~n23182 ) ;
  assign n23184 = n7594 ^ n5358 ^ n621 ;
  assign n23185 = n1924 & n10250 ;
  assign n23186 = n23184 & n23185 ;
  assign n23187 = ( ~n7182 & n20838 ) | ( ~n7182 & n23186 ) | ( n20838 & n23186 ) ;
  assign n23188 = n14473 ^ n7442 ^ n6380 ;
  assign n23189 = n23188 ^ n4524 ^ 1'b0 ;
  assign n23190 = ~n20466 & n23189 ;
  assign n23191 = n8064 & n23190 ;
  assign n23192 = n22130 & n23191 ;
  assign n23193 = n23192 ^ n19499 ^ n9605 ;
  assign n23194 = ~n23187 & n23193 ;
  assign n23195 = ~n23183 & n23194 ;
  assign n23196 = n15882 ^ n10804 ^ 1'b0 ;
  assign n23197 = ~n8014 & n23196 ;
  assign n23198 = n23197 ^ n17569 ^ n15765 ;
  assign n23199 = ( n3555 & n7840 ) | ( n3555 & ~n8794 ) | ( n7840 & ~n8794 ) ;
  assign n23200 = ( n14063 & ~n22107 ) | ( n14063 & n23199 ) | ( ~n22107 & n23199 ) ;
  assign n23201 = n3306 ^ n2318 ^ x173 ;
  assign n23202 = ( n14057 & n23200 ) | ( n14057 & ~n23201 ) | ( n23200 & ~n23201 ) ;
  assign n23203 = n21847 ^ n17848 ^ 1'b0 ;
  assign n23204 = n7713 | n8554 ;
  assign n23205 = ( ~n7031 & n20533 ) | ( ~n7031 & n23204 ) | ( n20533 & n23204 ) ;
  assign n23206 = ( ~n3399 & n9012 ) | ( ~n3399 & n23205 ) | ( n9012 & n23205 ) ;
  assign n23207 = n19795 ^ n16543 ^ 1'b0 ;
  assign n23208 = n16538 ^ n4823 ^ n1967 ;
  assign n23209 = n1809 & ~n9403 ;
  assign n23212 = ~n6428 & n8881 ;
  assign n23213 = n23212 ^ n3374 ^ 1'b0 ;
  assign n23214 = n15284 ^ n1947 ^ 1'b0 ;
  assign n23215 = ~n23213 & n23214 ;
  assign n23210 = ~n325 & n13416 ;
  assign n23211 = n23210 ^ n19107 ^ 1'b0 ;
  assign n23216 = n23215 ^ n23211 ^ n3706 ;
  assign n23217 = ( ~n15563 & n23209 ) | ( ~n15563 & n23216 ) | ( n23209 & n23216 ) ;
  assign n23218 = ( n7494 & n23208 ) | ( n7494 & n23217 ) | ( n23208 & n23217 ) ;
  assign n23219 = n20083 ^ n7531 ^ n1231 ;
  assign n23220 = ~n6227 & n8648 ;
  assign n23221 = n8610 & n23220 ;
  assign n23222 = ( n10942 & n18729 ) | ( n10942 & ~n23221 ) | ( n18729 & ~n23221 ) ;
  assign n23223 = ( n11007 & ~n17548 ) | ( n11007 & n23222 ) | ( ~n17548 & n23222 ) ;
  assign n23224 = ( n2935 & n23219 ) | ( n2935 & ~n23223 ) | ( n23219 & ~n23223 ) ;
  assign n23226 = n1987 & ~n13403 ;
  assign n23225 = ( n1459 & n2447 ) | ( n1459 & n3945 ) | ( n2447 & n3945 ) ;
  assign n23227 = n23226 ^ n23225 ^ n9885 ;
  assign n23228 = ( n312 & n1455 ) | ( n312 & ~n19888 ) | ( n1455 & ~n19888 ) ;
  assign n23229 = n21101 ^ n10749 ^ n2399 ;
  assign n23230 = n17451 & ~n23229 ;
  assign n23231 = n943 | n9610 ;
  assign n23232 = n10228 ^ n8551 ^ 1'b0 ;
  assign n23233 = n4540 | n23232 ;
  assign n23234 = n14487 ^ n9394 ^ n933 ;
  assign n23235 = n23234 ^ n7651 ^ n4384 ;
  assign n23236 = ( ~n23231 & n23233 ) | ( ~n23231 & n23235 ) | ( n23233 & n23235 ) ;
  assign n23237 = ~n1633 & n6341 ;
  assign n23238 = n23237 ^ n17864 ^ n15686 ;
  assign n23239 = n10378 | n15638 ;
  assign n23240 = n931 & n1536 ;
  assign n23241 = ~n20475 & n23240 ;
  assign n23242 = n5312 & n16303 ;
  assign n23243 = n23241 & n23242 ;
  assign n23256 = n827 | n2897 ;
  assign n23244 = ~n1313 & n7273 ;
  assign n23245 = n17868 & n23244 ;
  assign n23253 = ~n9061 & n13597 ;
  assign n23246 = n13474 ^ n8145 ^ n7066 ;
  assign n23247 = n23246 ^ n7331 ^ n3145 ;
  assign n23248 = ( x147 & ~n11444 ) | ( x147 & n23010 ) | ( ~n11444 & n23010 ) ;
  assign n23249 = n23248 ^ n2824 ^ 1'b0 ;
  assign n23250 = ~n10672 & n23249 ;
  assign n23251 = n12021 & n23250 ;
  assign n23252 = ~n23247 & n23251 ;
  assign n23254 = n23253 ^ n23252 ^ n10528 ;
  assign n23255 = n23245 | n23254 ;
  assign n23257 = n23256 ^ n23255 ^ 1'b0 ;
  assign n23258 = n13295 ^ n2342 ^ n1635 ;
  assign n23259 = n2315 & ~n3584 ;
  assign n23260 = n6359 & ~n18768 ;
  assign n23261 = ( n19630 & n23259 ) | ( n19630 & n23260 ) | ( n23259 & n23260 ) ;
  assign n23262 = n17408 ^ n6979 ^ 1'b0 ;
  assign n23263 = n6264 | n23262 ;
  assign n23264 = n19467 ^ n9725 ^ 1'b0 ;
  assign n23265 = n13605 ^ n11060 ^ 1'b0 ;
  assign n23266 = ( n8123 & ~n15491 ) | ( n8123 & n23265 ) | ( ~n15491 & n23265 ) ;
  assign n23267 = ( n17369 & n23264 ) | ( n17369 & ~n23266 ) | ( n23264 & ~n23266 ) ;
  assign n23268 = n22041 ^ n8662 ^ n4668 ;
  assign n23269 = ( n8722 & ~n22573 ) | ( n8722 & n23268 ) | ( ~n22573 & n23268 ) ;
  assign n23272 = ( n2486 & ~n11205 ) | ( n2486 & n12678 ) | ( ~n11205 & n12678 ) ;
  assign n23270 = ( n912 & ~n8948 ) | ( n912 & n10723 ) | ( ~n8948 & n10723 ) ;
  assign n23271 = ( n7620 & ~n12135 ) | ( n7620 & n23270 ) | ( ~n12135 & n23270 ) ;
  assign n23273 = n23272 ^ n23271 ^ n9910 ;
  assign n23274 = ( n2209 & n7088 ) | ( n2209 & ~n9003 ) | ( n7088 & ~n9003 ) ;
  assign n23275 = ~n6076 & n23274 ;
  assign n23276 = n10473 ^ n10169 ^ n4482 ;
  assign n23277 = n23276 ^ n16048 ^ 1'b0 ;
  assign n23278 = n12828 & ~n23277 ;
  assign n23279 = ~n23275 & n23278 ;
  assign n23282 = ( n1780 & n2033 ) | ( n1780 & n6653 ) | ( n2033 & n6653 ) ;
  assign n23280 = n4024 & ~n11316 ;
  assign n23281 = n14085 & n23280 ;
  assign n23283 = n23282 ^ n23281 ^ n8745 ;
  assign n23284 = n13750 & ~n23027 ;
  assign n23285 = n9563 ^ x183 ^ 1'b0 ;
  assign n23286 = n12782 ^ n9474 ^ 1'b0 ;
  assign n23287 = n9105 & ~n10568 ;
  assign n23288 = n18949 | n22313 ;
  assign n23289 = n23288 ^ n15333 ^ 1'b0 ;
  assign n23290 = ( n4165 & n16415 ) | ( n4165 & ~n22713 ) | ( n16415 & ~n22713 ) ;
  assign n23291 = ( n1048 & n4307 ) | ( n1048 & ~n9514 ) | ( n4307 & ~n9514 ) ;
  assign n23292 = n23291 ^ n10852 ^ 1'b0 ;
  assign n23293 = ( n3061 & n10843 ) | ( n3061 & ~n23292 ) | ( n10843 & ~n23292 ) ;
  assign n23294 = n23290 & ~n23293 ;
  assign n23295 = n23294 ^ n585 ^ 1'b0 ;
  assign n23296 = n23289 & n23295 ;
  assign n23297 = n23287 & n23296 ;
  assign n23298 = n23297 ^ n4279 ^ 1'b0 ;
  assign n23299 = ~n23286 & n23298 ;
  assign n23300 = ( n6770 & n13908 ) | ( n6770 & ~n18962 ) | ( n13908 & ~n18962 ) ;
  assign n23301 = n21821 ^ n2815 ^ n1218 ;
  assign n23302 = n2882 & n23301 ;
  assign n23303 = ~n23300 & n23302 ;
  assign n23304 = ( n5418 & ~n6701 ) | ( n5418 & n12485 ) | ( ~n6701 & n12485 ) ;
  assign n23305 = ( n6919 & n14507 ) | ( n6919 & ~n23304 ) | ( n14507 & ~n23304 ) ;
  assign n23306 = ( n421 & ~n7540 ) | ( n421 & n21395 ) | ( ~n7540 & n21395 ) ;
  assign n23308 = n14420 ^ n12753 ^ n10695 ;
  assign n23309 = n2430 & n23308 ;
  assign n23307 = n7376 & n9020 ;
  assign n23310 = n23309 ^ n23307 ^ 1'b0 ;
  assign n23311 = n23310 ^ n3922 ^ 1'b0 ;
  assign n23312 = n5006 | n20008 ;
  assign n23313 = n23312 ^ n8387 ^ 1'b0 ;
  assign n23314 = n22500 ^ n5074 ^ 1'b0 ;
  assign n23315 = ~n539 & n23314 ;
  assign n23316 = n23315 ^ n8494 ^ n6992 ;
  assign n23317 = n9332 ^ n5729 ^ 1'b0 ;
  assign n23318 = n21282 & ~n23317 ;
  assign n23319 = n3130 ^ n2296 ^ 1'b0 ;
  assign n23320 = ( n1164 & ~n23318 ) | ( n1164 & n23319 ) | ( ~n23318 & n23319 ) ;
  assign n23321 = n17452 ^ n8813 ^ 1'b0 ;
  assign n23322 = n7492 | n23321 ;
  assign n23323 = n15565 & ~n23322 ;
  assign n23324 = n21562 ^ n17845 ^ n3006 ;
  assign n23325 = n5208 ^ n3212 ^ n1392 ;
  assign n23326 = n23325 ^ n3944 ^ x154 ;
  assign n23327 = n12476 & ~n20016 ;
  assign n23328 = n23327 ^ n18613 ^ 1'b0 ;
  assign n23329 = n23328 ^ n15761 ^ n10310 ;
  assign n23330 = n5316 ^ n2272 ^ 1'b0 ;
  assign n23331 = ~n8061 & n23330 ;
  assign n23332 = n6125 & ~n18156 ;
  assign n23333 = ~n10625 & n23332 ;
  assign n23334 = ( ~n18554 & n23331 ) | ( ~n18554 & n23333 ) | ( n23331 & n23333 ) ;
  assign n23335 = n11727 & n20438 ;
  assign n23336 = n23335 ^ n1267 ^ 1'b0 ;
  assign n23337 = n1238 & ~n23336 ;
  assign n23338 = n16480 ^ n7678 ^ 1'b0 ;
  assign n23339 = ( n3672 & ~n18506 ) | ( n3672 & n23338 ) | ( ~n18506 & n23338 ) ;
  assign n23343 = ~n2360 & n6298 ;
  assign n23340 = n20782 ^ n16417 ^ n8072 ;
  assign n23341 = n6190 & ~n14074 ;
  assign n23342 = ( x3 & n23340 ) | ( x3 & n23341 ) | ( n23340 & n23341 ) ;
  assign n23344 = n23343 ^ n23342 ^ n11664 ;
  assign n23345 = n2003 | n6339 ;
  assign n23346 = n23345 ^ n21278 ^ 1'b0 ;
  assign n23347 = n6628 & ~n7982 ;
  assign n23348 = n5517 ^ n5493 ^ 1'b0 ;
  assign n23349 = n1503 & n23348 ;
  assign n23350 = n16094 | n23349 ;
  assign n23357 = n17972 ^ n15058 ^ n327 ;
  assign n23351 = n6678 ^ n4579 ^ n1109 ;
  assign n23352 = n10013 & ~n11847 ;
  assign n23353 = n23352 ^ x150 ^ 1'b0 ;
  assign n23354 = ( n7671 & n23351 ) | ( n7671 & n23353 ) | ( n23351 & n23353 ) ;
  assign n23355 = n259 | n23354 ;
  assign n23356 = n23355 ^ n10257 ^ 1'b0 ;
  assign n23358 = n23357 ^ n23356 ^ n3260 ;
  assign n23359 = n1752 ^ n1326 ^ 1'b0 ;
  assign n23360 = n11027 & n23359 ;
  assign n23361 = ~n620 & n23360 ;
  assign n23362 = n23361 ^ n22697 ^ 1'b0 ;
  assign n23363 = n13003 ^ n6697 ^ n1635 ;
  assign n23364 = n13162 ^ n9118 ^ n2406 ;
  assign n23365 = ( n3203 & n7664 ) | ( n3203 & n23364 ) | ( n7664 & n23364 ) ;
  assign n23366 = n14282 & ~n23365 ;
  assign n23367 = n23363 & n23366 ;
  assign n23368 = n13061 ^ n6919 ^ n5022 ;
  assign n23369 = n12007 ^ n7937 ^ n1222 ;
  assign n23370 = ( n1186 & n9582 ) | ( n1186 & n23369 ) | ( n9582 & n23369 ) ;
  assign n23371 = ( n4137 & n11410 ) | ( n4137 & ~n23370 ) | ( n11410 & ~n23370 ) ;
  assign n23372 = n23368 | n23371 ;
  assign n23373 = n23372 ^ n5613 ^ n5135 ;
  assign n23374 = n8802 ^ n8160 ^ n7645 ;
  assign n23375 = n23374 ^ n6230 ^ n2302 ;
  assign n23376 = ~n16410 & n23375 ;
  assign n23377 = n17733 & ~n23376 ;
  assign n23378 = n10436 & n12696 ;
  assign n23379 = ~n3726 & n23378 ;
  assign n23380 = ~n12353 & n13596 ;
  assign n23381 = n2502 | n23380 ;
  assign n23382 = n22443 | n23381 ;
  assign n23383 = n9869 ^ n3621 ^ n2306 ;
  assign n23384 = n23383 ^ n15690 ^ n11896 ;
  assign n23385 = n12783 & n20237 ;
  assign n23386 = n1406 & n4931 ;
  assign n23387 = ~n14468 & n23386 ;
  assign n23388 = n12238 & ~n23387 ;
  assign n23389 = ~n19922 & n23388 ;
  assign n23390 = n9195 ^ n2376 ^ n2362 ;
  assign n23391 = n23390 ^ n7917 ^ 1'b0 ;
  assign n23392 = ~n3106 & n23391 ;
  assign n23393 = n8886 ^ n838 ^ 1'b0 ;
  assign n23394 = ~n325 & n23393 ;
  assign n23395 = n23394 ^ n9822 ^ 1'b0 ;
  assign n23396 = n13077 ^ n4575 ^ 1'b0 ;
  assign n23397 = n17121 & ~n23396 ;
  assign n23398 = n4353 ^ n2895 ^ n1140 ;
  assign n23399 = n23398 ^ n7592 ^ n3202 ;
  assign n23400 = ( n23395 & ~n23397 ) | ( n23395 & n23399 ) | ( ~n23397 & n23399 ) ;
  assign n23401 = n23164 ^ n15453 ^ n11361 ;
  assign n23402 = n14887 ^ n3298 ^ n905 ;
  assign n23403 = n1428 & ~n17174 ;
  assign n23404 = n23402 & n23403 ;
  assign n23405 = ( n5166 & ~n10030 ) | ( n5166 & n20408 ) | ( ~n10030 & n20408 ) ;
  assign n23406 = n11301 ^ n8397 ^ n598 ;
  assign n23407 = n7050 ^ n5457 ^ 1'b0 ;
  assign n23408 = n531 & n23407 ;
  assign n23409 = n8308 ^ n4884 ^ n4850 ;
  assign n23410 = n23409 ^ n16080 ^ 1'b0 ;
  assign n23411 = n13042 ^ n4777 ^ x92 ;
  assign n23412 = n23411 ^ n6041 ^ 1'b0 ;
  assign n23413 = ~n3390 & n23412 ;
  assign n23414 = n2285 & n23413 ;
  assign n23415 = ~n23410 & n23414 ;
  assign n23416 = n23415 ^ n21820 ^ n4681 ;
  assign n23417 = n23416 ^ n6222 ^ 1'b0 ;
  assign n23418 = n6467 ^ n5863 ^ 1'b0 ;
  assign n23419 = n6311 | n23418 ;
  assign n23420 = n23419 ^ n4567 ^ n4092 ;
  assign n23421 = ( n13582 & n14837 ) | ( n13582 & n23420 ) | ( n14837 & n23420 ) ;
  assign n23422 = n23421 ^ n13912 ^ n7682 ;
  assign n23423 = n2942 ^ x86 ^ 1'b0 ;
  assign n23424 = ~n18078 & n23423 ;
  assign n23425 = n15513 ^ n11213 ^ 1'b0 ;
  assign n23426 = n23425 ^ n6961 ^ 1'b0 ;
  assign n23427 = n3701 & ~n23426 ;
  assign n23428 = ( n5919 & ~n10352 ) | ( n5919 & n14986 ) | ( ~n10352 & n14986 ) ;
  assign n23429 = n23428 ^ n7135 ^ 1'b0 ;
  assign n23430 = n6431 | n14553 ;
  assign n23431 = n13081 & ~n23430 ;
  assign n23432 = ( ~n17215 & n23429 ) | ( ~n17215 & n23431 ) | ( n23429 & n23431 ) ;
  assign n23433 = n1690 | n12447 ;
  assign n23434 = n23433 ^ n7366 ^ 1'b0 ;
  assign n23435 = ( n4357 & n5434 ) | ( n4357 & n7144 ) | ( n5434 & n7144 ) ;
  assign n23436 = n10948 | n23435 ;
  assign n23437 = n23436 ^ n17937 ^ 1'b0 ;
  assign n23442 = n15657 ^ n11721 ^ n5478 ;
  assign n23438 = n3326 ^ n1889 ^ 1'b0 ;
  assign n23439 = n7588 & ~n23438 ;
  assign n23440 = n23439 ^ n4644 ^ n922 ;
  assign n23441 = n23440 ^ n21252 ^ n15831 ;
  assign n23443 = n23442 ^ n23441 ^ n14195 ;
  assign n23444 = n7666 ^ n7099 ^ 1'b0 ;
  assign n23445 = n23444 ^ n17588 ^ n1236 ;
  assign n23455 = n21747 ^ n9312 ^ n717 ;
  assign n23456 = ( ~n4277 & n11287 ) | ( ~n4277 & n23455 ) | ( n11287 & n23455 ) ;
  assign n23457 = n23456 ^ n16057 ^ n14765 ;
  assign n23446 = x246 & n4471 ;
  assign n23447 = n23446 ^ n16638 ^ n2894 ;
  assign n23448 = n9583 ^ n6771 ^ 1'b0 ;
  assign n23449 = n12437 & n23448 ;
  assign n23450 = n3858 ^ n585 ^ 1'b0 ;
  assign n23451 = n811 | n23450 ;
  assign n23452 = ( n11660 & n23449 ) | ( n11660 & n23451 ) | ( n23449 & n23451 ) ;
  assign n23453 = ( n12325 & n13426 ) | ( n12325 & ~n23452 ) | ( n13426 & ~n23452 ) ;
  assign n23454 = ( n21572 & ~n23447 ) | ( n21572 & n23453 ) | ( ~n23447 & n23453 ) ;
  assign n23458 = n23457 ^ n23454 ^ n872 ;
  assign n23459 = n6445 & ~n16058 ;
  assign n23460 = n23459 ^ n9888 ^ 1'b0 ;
  assign n23461 = n23460 ^ n18217 ^ n14767 ;
  assign n23462 = ( n20623 & n22693 ) | ( n20623 & ~n23461 ) | ( n22693 & ~n23461 ) ;
  assign n23463 = n7900 & n8779 ;
  assign n23464 = n23463 ^ n6863 ^ 1'b0 ;
  assign n23465 = n17946 ^ n16010 ^ n1366 ;
  assign n23466 = ~n1754 & n23465 ;
  assign n23467 = n23466 ^ n21920 ^ 1'b0 ;
  assign n23468 = ( n4323 & n23464 ) | ( n4323 & n23467 ) | ( n23464 & n23467 ) ;
  assign n23469 = n5236 & n21086 ;
  assign n23470 = ( n4908 & n8982 ) | ( n4908 & n23469 ) | ( n8982 & n23469 ) ;
  assign n23473 = n10098 ^ n468 ^ 1'b0 ;
  assign n23471 = n14223 ^ n3883 ^ n2002 ;
  assign n23472 = n23471 ^ n7057 ^ 1'b0 ;
  assign n23474 = n23473 ^ n23472 ^ n22822 ;
  assign n23475 = n1241 | n2329 ;
  assign n23476 = n22770 | n23475 ;
  assign n23478 = ( n1215 & n3124 ) | ( n1215 & n5701 ) | ( n3124 & n5701 ) ;
  assign n23477 = n13144 & n22286 ;
  assign n23479 = n23478 ^ n23477 ^ 1'b0 ;
  assign n23480 = ( n1676 & ~n4795 ) | ( n1676 & n5188 ) | ( ~n4795 & n5188 ) ;
  assign n23481 = ~n10474 & n23480 ;
  assign n23482 = n23479 & n23481 ;
  assign n23483 = ( n771 & ~n13350 ) | ( n771 & n13474 ) | ( ~n13350 & n13474 ) ;
  assign n23484 = n13941 & n23483 ;
  assign n23485 = n16534 ^ n12381 ^ n7223 ;
  assign n23486 = ( n773 & n6326 ) | ( n773 & n13821 ) | ( n6326 & n13821 ) ;
  assign n23487 = n23486 ^ n6854 ^ 1'b0 ;
  assign n23488 = n12134 & n23487 ;
  assign n23489 = n23488 ^ n17162 ^ n7537 ;
  assign n23490 = n7412 ^ n5414 ^ 1'b0 ;
  assign n23491 = n23490 ^ n10590 ^ 1'b0 ;
  assign n23498 = n7206 ^ n3134 ^ n2041 ;
  assign n23492 = n896 & n6853 ;
  assign n23493 = ~n7218 & n23492 ;
  assign n23494 = n23493 ^ n8637 ^ 1'b0 ;
  assign n23495 = n3146 & ~n23494 ;
  assign n23496 = n1047 & n14667 ;
  assign n23497 = ~n23495 & n23496 ;
  assign n23499 = n23498 ^ n23497 ^ 1'b0 ;
  assign n23500 = n9228 ^ n6470 ^ n6317 ;
  assign n23501 = n23500 ^ n16480 ^ n8053 ;
  assign n23502 = ( n1380 & ~n8316 ) | ( n1380 & n23501 ) | ( ~n8316 & n23501 ) ;
  assign n23503 = n9744 ^ n9265 ^ 1'b0 ;
  assign n23504 = ~n10225 & n23503 ;
  assign n23505 = ~n19061 & n23504 ;
  assign n23506 = ( n13515 & n23502 ) | ( n13515 & n23505 ) | ( n23502 & n23505 ) ;
  assign n23507 = ( n4736 & ~n21359 ) | ( n4736 & n23506 ) | ( ~n21359 & n23506 ) ;
  assign n23508 = ( n5247 & n16544 ) | ( n5247 & n23507 ) | ( n16544 & n23507 ) ;
  assign n23509 = n9926 | n23471 ;
  assign n23510 = n11842 | n23509 ;
  assign n23511 = n6871 ^ n1712 ^ n1592 ;
  assign n23512 = ( n8916 & n23510 ) | ( n8916 & ~n23511 ) | ( n23510 & ~n23511 ) ;
  assign n23513 = ( ~n10048 & n13652 ) | ( ~n10048 & n23512 ) | ( n13652 & n23512 ) ;
  assign n23514 = n3122 | n22484 ;
  assign n23515 = ( n5985 & n9750 ) | ( n5985 & ~n15475 ) | ( n9750 & ~n15475 ) ;
  assign n23516 = n14726 ^ n5166 ^ n4856 ;
  assign n23517 = n23516 ^ n6776 ^ x4 ;
  assign n23518 = n23517 ^ n8184 ^ n1088 ;
  assign n23519 = n23518 ^ n7562 ^ 1'b0 ;
  assign n23520 = n20519 & n23334 ;
  assign n23521 = n20726 ^ n20587 ^ n3500 ;
  assign n23522 = n10106 | n16573 ;
  assign n23523 = n23522 ^ n6106 ^ 1'b0 ;
  assign n23524 = n4638 | n23523 ;
  assign n23525 = ( ~n21151 & n23521 ) | ( ~n21151 & n23524 ) | ( n23521 & n23524 ) ;
  assign n23526 = ( n2786 & n6222 ) | ( n2786 & n10845 ) | ( n6222 & n10845 ) ;
  assign n23527 = n23526 ^ n23199 ^ 1'b0 ;
  assign n23528 = x112 & ~n16540 ;
  assign n23529 = ~n22047 & n23528 ;
  assign n23530 = ( n2016 & n5591 ) | ( n2016 & ~n18436 ) | ( n5591 & ~n18436 ) ;
  assign n23532 = n15880 ^ n846 ^ 1'b0 ;
  assign n23531 = n4257 | n13978 ;
  assign n23533 = n23532 ^ n23531 ^ 1'b0 ;
  assign n23534 = ( ~n8925 & n23530 ) | ( ~n8925 & n23533 ) | ( n23530 & n23533 ) ;
  assign n23535 = n23188 ^ n17245 ^ n11071 ;
  assign n23536 = n21538 & n23535 ;
  assign n23537 = ( n3042 & n4474 ) | ( n3042 & ~n18479 ) | ( n4474 & ~n18479 ) ;
  assign n23538 = ~n5921 & n17950 ;
  assign n23539 = ~n3591 & n19624 ;
  assign n23540 = ( ~n20973 & n23538 ) | ( ~n20973 & n23539 ) | ( n23538 & n23539 ) ;
  assign n23541 = ( ~n257 & n6607 ) | ( ~n257 & n23540 ) | ( n6607 & n23540 ) ;
  assign n23542 = ( n15542 & n23537 ) | ( n15542 & ~n23541 ) | ( n23537 & ~n23541 ) ;
  assign n23543 = n20377 & n23542 ;
  assign n23544 = n587 & n23543 ;
  assign n23545 = n23544 ^ n13652 ^ 1'b0 ;
  assign n23546 = n15883 ^ n12012 ^ n11703 ;
  assign n23547 = n23546 ^ n18148 ^ n9855 ;
  assign n23548 = ( n10169 & ~n19729 ) | ( n10169 & n23547 ) | ( ~n19729 & n23547 ) ;
  assign n23549 = n12497 ^ n7259 ^ 1'b0 ;
  assign n23550 = n23549 ^ n11119 ^ n7066 ;
  assign n23551 = n10564 | n18860 ;
  assign n23553 = n7478 ^ n6648 ^ 1'b0 ;
  assign n23552 = n7300 | n9757 ;
  assign n23554 = n23553 ^ n23552 ^ 1'b0 ;
  assign n23555 = n22092 ^ n7049 ^ 1'b0 ;
  assign n23556 = n23555 ^ n15699 ^ 1'b0 ;
  assign n23558 = ( n841 & n11961 ) | ( n841 & ~n19205 ) | ( n11961 & ~n19205 ) ;
  assign n23557 = n3043 & ~n19493 ;
  assign n23559 = n23558 ^ n23557 ^ 1'b0 ;
  assign n23561 = n23106 ^ n2234 ^ n1856 ;
  assign n23562 = n23561 ^ n13577 ^ n5643 ;
  assign n23560 = n6012 & n16015 ;
  assign n23563 = n23562 ^ n23560 ^ 1'b0 ;
  assign n23570 = n3620 | n12117 ;
  assign n23571 = n10242 | n23570 ;
  assign n23566 = n3508 & n4472 ;
  assign n23567 = n23566 ^ n1518 ^ 1'b0 ;
  assign n23568 = n23567 ^ n10200 ^ n6230 ;
  assign n23564 = ( n4009 & n4858 ) | ( n4009 & ~n8092 ) | ( n4858 & ~n8092 ) ;
  assign n23565 = n23564 ^ n5449 ^ 1'b0 ;
  assign n23569 = n23568 ^ n23565 ^ n11384 ;
  assign n23572 = n23571 ^ n23569 ^ n10308 ;
  assign n23573 = n1973 ^ n561 ^ x212 ;
  assign n23574 = n23573 ^ n19625 ^ n8275 ;
  assign n23575 = n23574 ^ n23091 ^ n13510 ;
  assign n23577 = n5540 & ~n10109 ;
  assign n23578 = n23577 ^ n5808 ^ 1'b0 ;
  assign n23576 = ( n3828 & ~n13149 ) | ( n3828 & n23123 ) | ( ~n13149 & n23123 ) ;
  assign n23579 = n23578 ^ n23576 ^ n20040 ;
  assign n23580 = n23579 ^ n7045 ^ n3616 ;
  assign n23581 = n12601 ^ n3740 ^ n1104 ;
  assign n23582 = n12337 | n15967 ;
  assign n23583 = n23582 ^ n18994 ^ 1'b0 ;
  assign n23584 = n23318 ^ n8892 ^ x33 ;
  assign n23585 = n23584 ^ n13249 ^ n12151 ;
  assign n23586 = ( n2308 & n5596 ) | ( n2308 & ~n15724 ) | ( n5596 & ~n15724 ) ;
  assign n23587 = n16250 ^ n8519 ^ n5918 ;
  assign n23588 = ( n17212 & ~n19776 ) | ( n17212 & n23587 ) | ( ~n19776 & n23587 ) ;
  assign n23589 = n13941 ^ n11440 ^ n2372 ;
  assign n23590 = n23589 ^ n7523 ^ 1'b0 ;
  assign n23591 = ( n6591 & n8562 ) | ( n6591 & n8569 ) | ( n8562 & n8569 ) ;
  assign n23592 = n23591 ^ n18804 ^ n9320 ;
  assign n23593 = n23592 ^ n11232 ^ n2715 ;
  assign n23594 = n23593 ^ n16547 ^ 1'b0 ;
  assign n23595 = ( ~n8727 & n19583 ) | ( ~n8727 & n23594 ) | ( n19583 & n23594 ) ;
  assign n23596 = n12007 | n17048 ;
  assign n23597 = n23596 ^ n5259 ^ n2081 ;
  assign n23598 = ( n2110 & n5823 ) | ( n2110 & n15852 ) | ( n5823 & n15852 ) ;
  assign n23599 = n23598 ^ n13737 ^ n5996 ;
  assign n23600 = ( n14476 & ~n23597 ) | ( n14476 & n23599 ) | ( ~n23597 & n23599 ) ;
  assign n23601 = ~x87 & n12998 ;
  assign n23602 = n23601 ^ n17539 ^ 1'b0 ;
  assign n23603 = n10574 ^ n2296 ^ 1'b0 ;
  assign n23604 = ~n10808 & n23603 ;
  assign n23605 = n23604 ^ n16480 ^ n7178 ;
  assign n23606 = n23605 ^ n13385 ^ n3514 ;
  assign n23607 = n22140 ^ n16507 ^ 1'b0 ;
  assign n23608 = ~n12853 & n21049 ;
  assign n23609 = ~n23607 & n23608 ;
  assign n23610 = n1828 & n7100 ;
  assign n23611 = n23610 ^ n5974 ^ 1'b0 ;
  assign n23612 = ( n2426 & ~n3361 ) | ( n2426 & n11048 ) | ( ~n3361 & n11048 ) ;
  assign n23613 = n23612 ^ n5799 ^ 1'b0 ;
  assign n23614 = ( n1310 & n6959 ) | ( n1310 & ~n23613 ) | ( n6959 & ~n23613 ) ;
  assign n23615 = n23614 ^ n23495 ^ 1'b0 ;
  assign n23616 = ~n23611 & n23615 ;
  assign n23617 = n12992 ^ n1170 ^ 1'b0 ;
  assign n23618 = n16019 ^ n14633 ^ n10726 ;
  assign n23619 = n10047 | n15728 ;
  assign n23620 = ( n3412 & n8241 ) | ( n3412 & n15162 ) | ( n8241 & n15162 ) ;
  assign n23621 = ~n4998 & n8818 ;
  assign n23622 = n23621 ^ n14999 ^ 1'b0 ;
  assign n23623 = ~n23620 & n23622 ;
  assign n23624 = ~n23619 & n23623 ;
  assign n23625 = ( n12294 & ~n14186 ) | ( n12294 & n23624 ) | ( ~n14186 & n23624 ) ;
  assign n23628 = n12101 ^ n10216 ^ n8322 ;
  assign n23626 = n12792 ^ n8401 ^ n5358 ;
  assign n23627 = n22667 & n23626 ;
  assign n23629 = n23628 ^ n23627 ^ n5975 ;
  assign n23637 = ( ~n2851 & n7089 ) | ( ~n2851 & n11410 ) | ( n7089 & n11410 ) ;
  assign n23631 = ( ~n5611 & n7183 ) | ( ~n5611 & n16118 ) | ( n7183 & n16118 ) ;
  assign n23632 = n2231 & n23631 ;
  assign n23633 = ~n1206 & n23632 ;
  assign n23634 = ( n1587 & n12303 ) | ( n1587 & ~n23633 ) | ( n12303 & ~n23633 ) ;
  assign n23635 = n23634 ^ n12590 ^ n8701 ;
  assign n23630 = n16621 ^ n9002 ^ 1'b0 ;
  assign n23636 = n23635 ^ n23630 ^ n2701 ;
  assign n23638 = n23637 ^ n23636 ^ 1'b0 ;
  assign n23639 = n15034 ^ n2092 ^ 1'b0 ;
  assign n23640 = n23247 & ~n23639 ;
  assign n23641 = n23640 ^ n5077 ^ n1756 ;
  assign n23642 = n16936 & ~n23641 ;
  assign n23643 = n6429 & n23642 ;
  assign n23644 = ( n5020 & n7645 ) | ( n5020 & n18595 ) | ( n7645 & n18595 ) ;
  assign n23645 = n21986 ^ n2774 ^ 1'b0 ;
  assign n23646 = ~n23644 & n23645 ;
  assign n23647 = ~n8754 & n10209 ;
  assign n23648 = n9093 ^ n8819 ^ n5697 ;
  assign n23649 = n12249 ^ n7703 ^ 1'b0 ;
  assign n23650 = n23648 | n23649 ;
  assign n23652 = n1480 & n5197 ;
  assign n23653 = n1294 & n23652 ;
  assign n23651 = n12059 ^ n11378 ^ n5084 ;
  assign n23654 = n23653 ^ n23651 ^ 1'b0 ;
  assign n23655 = n23650 | n23654 ;
  assign n23656 = n7228 & n17034 ;
  assign n23657 = ( n2401 & n4433 ) | ( n2401 & ~n13515 ) | ( n4433 & ~n13515 ) ;
  assign n23658 = n23657 ^ n763 ^ 1'b0 ;
  assign n23659 = n5370 & ~n7461 ;
  assign n23660 = ~n5080 & n23659 ;
  assign n23661 = n5661 ^ n2313 ^ 1'b0 ;
  assign n23662 = n280 & n23661 ;
  assign n23663 = n23662 ^ n3493 ^ 1'b0 ;
  assign n23664 = n9023 & ~n11990 ;
  assign n23665 = n6404 | n8319 ;
  assign n23666 = ( n23663 & ~n23664 ) | ( n23663 & n23665 ) | ( ~n23664 & n23665 ) ;
  assign n23667 = ( ~n6394 & n23660 ) | ( ~n6394 & n23666 ) | ( n23660 & n23666 ) ;
  assign n23668 = n23667 ^ n18058 ^ n1299 ;
  assign n23669 = n23253 ^ n3824 ^ 1'b0 ;
  assign n23670 = n23669 ^ n3723 ^ 1'b0 ;
  assign n23671 = n20398 ^ n6505 ^ n6400 ;
  assign n23672 = n8432 & ~n23671 ;
  assign n23673 = n23672 ^ n8955 ^ 1'b0 ;
  assign n23674 = n8133 & ~n23673 ;
  assign n23675 = n23674 ^ n11149 ^ 1'b0 ;
  assign n23676 = n14357 ^ n7000 ^ 1'b0 ;
  assign n23677 = ( n14000 & ~n15478 ) | ( n14000 & n23676 ) | ( ~n15478 & n23676 ) ;
  assign n23678 = n16519 ^ n864 ^ 1'b0 ;
  assign n23679 = ~n13654 & n23678 ;
  assign n23680 = n12001 ^ n5290 ^ n765 ;
  assign n23681 = ~n1807 & n23680 ;
  assign n23682 = n12122 | n23681 ;
  assign n23683 = n23679 | n23682 ;
  assign n23686 = n4576 & n18778 ;
  assign n23684 = ~n4142 & n4952 ;
  assign n23685 = n8027 & n23684 ;
  assign n23687 = n23686 ^ n23685 ^ n10933 ;
  assign n23688 = n11545 & ~n23687 ;
  assign n23689 = n23688 ^ n6616 ^ 1'b0 ;
  assign n23690 = ( n11953 & n12801 ) | ( n11953 & n22249 ) | ( n12801 & n22249 ) ;
  assign n23691 = ( ~n7840 & n13803 ) | ( ~n7840 & n23690 ) | ( n13803 & n23690 ) ;
  assign n23692 = n6139 | n23691 ;
  assign n23693 = n23205 ^ n21975 ^ n7149 ;
  assign n23695 = n10439 ^ n5469 ^ n1730 ;
  assign n23694 = n16137 ^ n3154 ^ 1'b0 ;
  assign n23696 = n23695 ^ n23694 ^ 1'b0 ;
  assign n23697 = ( ~n974 & n7720 ) | ( ~n974 & n21456 ) | ( n7720 & n21456 ) ;
  assign n23699 = n8402 ^ n825 ^ 1'b0 ;
  assign n23700 = n6865 & ~n23699 ;
  assign n23698 = n17424 | n20535 ;
  assign n23701 = n23700 ^ n23698 ^ 1'b0 ;
  assign n23702 = n23697 & n23701 ;
  assign n23703 = n23702 ^ n19152 ^ 1'b0 ;
  assign n23704 = n10036 ^ n9976 ^ 1'b0 ;
  assign n23707 = n23226 ^ n17151 ^ n8016 ;
  assign n23705 = n2069 ^ n1903 ^ 1'b0 ;
  assign n23706 = n23705 ^ n13528 ^ n5613 ;
  assign n23708 = n23707 ^ n23706 ^ 1'b0 ;
  assign n23709 = ( n9412 & n13226 ) | ( n9412 & ~n23708 ) | ( n13226 & ~n23708 ) ;
  assign n23710 = n23709 ^ n14687 ^ 1'b0 ;
  assign n23711 = n23704 & n23710 ;
  assign n23712 = n15158 ^ n14195 ^ n4400 ;
  assign n23713 = n12779 & n23712 ;
  assign n23714 = ~n9057 & n23713 ;
  assign n23716 = n1509 ^ n1215 ^ 1'b0 ;
  assign n23717 = n3029 | n23716 ;
  assign n23715 = n10521 ^ n6767 ^ n3926 ;
  assign n23718 = n23717 ^ n23715 ^ n667 ;
  assign n23719 = n23718 ^ n11808 ^ n9651 ;
  assign n23720 = n13746 ^ n5952 ^ n5506 ;
  assign n23721 = n14394 ^ n10825 ^ n2115 ;
  assign n23722 = ( n2564 & ~n3871 ) | ( n2564 & n23721 ) | ( ~n3871 & n23721 ) ;
  assign n23723 = n18818 | n23722 ;
  assign n23724 = ( n3041 & n13015 ) | ( n3041 & ~n14226 ) | ( n13015 & ~n14226 ) ;
  assign n23725 = n23724 ^ n6915 ^ n6388 ;
  assign n23726 = n12013 ^ n5416 ^ 1'b0 ;
  assign n23727 = n23726 ^ n12812 ^ n615 ;
  assign n23728 = n23727 ^ n18200 ^ n10232 ;
  assign n23729 = n20566 ^ n17484 ^ n1853 ;
  assign n23730 = n8638 ^ n8411 ^ 1'b0 ;
  assign n23731 = n23730 ^ n23601 ^ n7630 ;
  assign n23732 = n23731 ^ n13661 ^ n6541 ;
  assign n23733 = ( n2677 & ~n8856 ) | ( n2677 & n13851 ) | ( ~n8856 & n13851 ) ;
  assign n23734 = n23495 ^ n23051 ^ 1'b0 ;
  assign n23736 = ~n10319 & n16063 ;
  assign n23737 = n18972 & n23736 ;
  assign n23735 = n20972 ^ n11573 ^ n5124 ;
  assign n23738 = n23737 ^ n23735 ^ n4884 ;
  assign n23739 = ( ~n3147 & n5141 ) | ( ~n3147 & n23738 ) | ( n5141 & n23738 ) ;
  assign n23740 = n859 & n23739 ;
  assign n23741 = n23734 & n23740 ;
  assign n23742 = n16907 & ~n23741 ;
  assign n23743 = n23742 ^ n18836 ^ 1'b0 ;
  assign n23744 = n18821 | n21539 ;
  assign n23745 = ( ~n4992 & n10739 ) | ( ~n4992 & n23744 ) | ( n10739 & n23744 ) ;
  assign n23746 = n10319 ^ n1747 ^ 1'b0 ;
  assign n23747 = n6524 | n22075 ;
  assign n23748 = n5534 | n23747 ;
  assign n23749 = n17425 & ~n23748 ;
  assign n23750 = n23746 & n23749 ;
  assign n23751 = ( ~n5652 & n12049 ) | ( ~n5652 & n23506 ) | ( n12049 & n23506 ) ;
  assign n23752 = n7668 ^ n3971 ^ n2654 ;
  assign n23753 = n23752 ^ n10903 ^ n6761 ;
  assign n23754 = n23753 ^ n17323 ^ n7316 ;
  assign n23755 = n10875 ^ n7568 ^ 1'b0 ;
  assign n23756 = n7687 & n16524 ;
  assign n23757 = n23755 & n23756 ;
  assign n23758 = n23124 ^ n10713 ^ 1'b0 ;
  assign n23759 = n23757 | n23758 ;
  assign n23761 = ( n7632 & n14613 ) | ( n7632 & ~n17321 ) | ( n14613 & ~n17321 ) ;
  assign n23762 = n23761 ^ n9927 ^ n5637 ;
  assign n23760 = n13633 | n19471 ;
  assign n23763 = n23762 ^ n23760 ^ 1'b0 ;
  assign n23764 = ( ~n23754 & n23759 ) | ( ~n23754 & n23763 ) | ( n23759 & n23763 ) ;
  assign n23765 = n11820 ^ n10796 ^ 1'b0 ;
  assign n23766 = n9170 & n23765 ;
  assign n23767 = ( n1319 & n23365 ) | ( n1319 & n23766 ) | ( n23365 & n23766 ) ;
  assign n23768 = n5550 ^ n2187 ^ n1218 ;
  assign n23769 = ( n3697 & n9533 ) | ( n3697 & ~n23768 ) | ( n9533 & ~n23768 ) ;
  assign n23770 = ( ~n5555 & n6052 ) | ( ~n5555 & n22456 ) | ( n6052 & n22456 ) ;
  assign n23771 = n12939 ^ n5564 ^ 1'b0 ;
  assign n23772 = n17626 & n23771 ;
  assign n23773 = n23772 ^ n22249 ^ 1'b0 ;
  assign n23774 = ( n15025 & ~n23241 ) | ( n15025 & n23773 ) | ( ~n23241 & n23773 ) ;
  assign n23775 = n23774 ^ n23763 ^ n1413 ;
  assign n23776 = n3045 | n5010 ;
  assign n23777 = ~n21554 & n23776 ;
  assign n23778 = n23777 ^ n14571 ^ 1'b0 ;
  assign n23779 = ( ~n1110 & n17817 ) | ( ~n1110 & n20630 ) | ( n17817 & n20630 ) ;
  assign n23782 = n2085 | n8126 ;
  assign n23783 = n23782 ^ n441 ^ 1'b0 ;
  assign n23784 = n23783 ^ n17979 ^ 1'b0 ;
  assign n23785 = n3125 | n23784 ;
  assign n23781 = n21367 & n21974 ;
  assign n23786 = n23785 ^ n23781 ^ 1'b0 ;
  assign n23780 = n12606 ^ n8303 ^ n597 ;
  assign n23787 = n23786 ^ n23780 ^ n5600 ;
  assign n23788 = n23787 ^ n7344 ^ 1'b0 ;
  assign n23789 = n6592 & n21622 ;
  assign n23790 = ( n7454 & n8477 ) | ( n7454 & n12600 ) | ( n8477 & n12600 ) ;
  assign n23791 = n14329 ^ n1751 ^ 1'b0 ;
  assign n23792 = n23790 & n23791 ;
  assign n23793 = n11228 & n18166 ;
  assign n23794 = ~n5391 & n23793 ;
  assign n23795 = ~n4523 & n18093 ;
  assign n23796 = n23795 ^ n9278 ^ 1'b0 ;
  assign n23797 = n736 | n14526 ;
  assign n23798 = n1957 & ~n23797 ;
  assign n23799 = n23798 ^ n6872 ^ 1'b0 ;
  assign n23800 = n23799 ^ n15460 ^ n2526 ;
  assign n23804 = ( n5500 & n13862 ) | ( n5500 & n16991 ) | ( n13862 & n16991 ) ;
  assign n23803 = n11548 ^ n4676 ^ n2145 ;
  assign n23805 = n23804 ^ n23803 ^ 1'b0 ;
  assign n23806 = ~n19063 & n23805 ;
  assign n23801 = n4090 ^ n3406 ^ n494 ;
  assign n23802 = ( n3911 & n12098 ) | ( n3911 & ~n23801 ) | ( n12098 & ~n23801 ) ;
  assign n23807 = n23806 ^ n23802 ^ 1'b0 ;
  assign n23808 = ( n1067 & n14026 ) | ( n1067 & ~n21158 ) | ( n14026 & ~n21158 ) ;
  assign n23809 = n14846 ^ n6733 ^ n490 ;
  assign n23810 = n23809 ^ n16352 ^ n4533 ;
  assign n23811 = n18938 & ~n23810 ;
  assign n23812 = n10276 ^ n4520 ^ 1'b0 ;
  assign n23814 = n22670 ^ n17339 ^ 1'b0 ;
  assign n23815 = n8454 | n23814 ;
  assign n23813 = ~n4152 & n13523 ;
  assign n23816 = n23815 ^ n23813 ^ 1'b0 ;
  assign n23817 = n13739 & ~n23816 ;
  assign n23818 = n6041 | n18120 ;
  assign n23819 = n23818 ^ n14133 ^ n4139 ;
  assign n23820 = n23068 ^ n652 ^ 1'b0 ;
  assign n23821 = n15724 ^ n14084 ^ n7084 ;
  assign n23822 = ( n8784 & ~n9081 ) | ( n8784 & n14602 ) | ( ~n9081 & n14602 ) ;
  assign n23823 = n23822 ^ n22097 ^ 1'b0 ;
  assign n23824 = ~n23821 & n23823 ;
  assign n23825 = n23824 ^ n10897 ^ 1'b0 ;
  assign n23826 = n23820 & n23825 ;
  assign n23827 = ( n8189 & ~n9922 ) | ( n8189 & n22186 ) | ( ~n9922 & n22186 ) ;
  assign n23828 = n6959 ^ n5948 ^ n3128 ;
  assign n23829 = n10465 ^ n3352 ^ n1233 ;
  assign n23834 = n19845 ^ n14744 ^ n2646 ;
  assign n23830 = n8707 ^ n420 ^ 1'b0 ;
  assign n23831 = ( n6230 & n8949 ) | ( n6230 & ~n23830 ) | ( n8949 & ~n23830 ) ;
  assign n23832 = n23831 ^ n10498 ^ n7554 ;
  assign n23833 = n6376 & n23832 ;
  assign n23835 = n23834 ^ n23833 ^ 1'b0 ;
  assign n23836 = n23835 ^ n12906 ^ 1'b0 ;
  assign n23837 = n23829 & ~n23836 ;
  assign n23838 = n23828 & n23837 ;
  assign n23839 = n23838 ^ n14505 ^ 1'b0 ;
  assign n23840 = n814 & ~n23839 ;
  assign n23841 = ( ~n13304 & n23827 ) | ( ~n13304 & n23840 ) | ( n23827 & n23840 ) ;
  assign n23843 = n5811 & n12391 ;
  assign n23842 = ~n15343 & n20082 ;
  assign n23844 = n23843 ^ n23842 ^ n13003 ;
  assign n23845 = ~n2649 & n7508 ;
  assign n23846 = ~n6635 & n23845 ;
  assign n23847 = n23846 ^ n21060 ^ n11624 ;
  assign n23848 = n19395 ^ n5162 ^ 1'b0 ;
  assign n23849 = n2888 | n23848 ;
  assign n23850 = n13869 ^ n10287 ^ n7298 ;
  assign n23851 = n23849 | n23850 ;
  assign n23852 = n23851 ^ n22615 ^ n5192 ;
  assign n23853 = ( x167 & ~n7740 ) | ( x167 & n12238 ) | ( ~n7740 & n12238 ) ;
  assign n23854 = n23853 ^ n9810 ^ n861 ;
  assign n23855 = n23854 ^ n7028 ^ n6189 ;
  assign n23856 = x222 & ~n7747 ;
  assign n23857 = n23856 ^ n1645 ^ 1'b0 ;
  assign n23858 = ( ~n724 & n14309 ) | ( ~n724 & n16066 ) | ( n14309 & n16066 ) ;
  assign n23861 = n4033 ^ n1406 ^ 1'b0 ;
  assign n23860 = ( n4295 & ~n13751 ) | ( n4295 & n22075 ) | ( ~n13751 & n22075 ) ;
  assign n23862 = n23861 ^ n23860 ^ 1'b0 ;
  assign n23863 = ~n4271 & n23862 ;
  assign n23859 = n11637 ^ n9815 ^ n7060 ;
  assign n23864 = n23863 ^ n23859 ^ 1'b0 ;
  assign n23865 = n7223 & n10204 ;
  assign n23866 = ( ~n6101 & n7240 ) | ( ~n6101 & n23865 ) | ( n7240 & n23865 ) ;
  assign n23868 = n4399 ^ n2214 ^ x65 ;
  assign n23867 = n17881 & ~n18670 ;
  assign n23869 = n23868 ^ n23867 ^ 1'b0 ;
  assign n23879 = n21172 ^ n914 ^ x144 ;
  assign n23875 = n11543 ^ n10826 ^ n3316 ;
  assign n23873 = n10305 ^ n5307 ^ n1198 ;
  assign n23874 = n423 & n23873 ;
  assign n23876 = n23875 ^ n23874 ^ 1'b0 ;
  assign n23877 = ( n4417 & n13355 ) | ( n4417 & n23876 ) | ( n13355 & n23876 ) ;
  assign n23878 = ( n1905 & n18920 ) | ( n1905 & ~n23877 ) | ( n18920 & ~n23877 ) ;
  assign n23870 = n2341 & n21577 ;
  assign n23871 = ~n7074 & n23870 ;
  assign n23872 = n23631 | n23871 ;
  assign n23880 = n23879 ^ n23878 ^ n23872 ;
  assign n23881 = n2083 ^ n1541 ^ n812 ;
  assign n23882 = n8035 | n23881 ;
  assign n23883 = ( ~n694 & n11299 ) | ( ~n694 & n23882 ) | ( n11299 & n23882 ) ;
  assign n23884 = n15772 ^ n8963 ^ n8383 ;
  assign n23885 = ~n7455 & n14091 ;
  assign n23888 = n17721 ^ n9120 ^ 1'b0 ;
  assign n23889 = ~n8569 & n23888 ;
  assign n23886 = ( n3899 & n16585 ) | ( n3899 & ~n19420 ) | ( n16585 & ~n19420 ) ;
  assign n23887 = n21271 & n23886 ;
  assign n23890 = n23889 ^ n23887 ^ 1'b0 ;
  assign n23891 = n18834 ^ n7776 ^ n1161 ;
  assign n23892 = n15687 ^ n4128 ^ x70 ;
  assign n23895 = n13688 ^ n2036 ^ 1'b0 ;
  assign n23896 = ~n8478 & n23895 ;
  assign n23897 = n17288 ^ n3072 ^ 1'b0 ;
  assign n23898 = n4718 | n23897 ;
  assign n23899 = ( ~n21359 & n23896 ) | ( ~n21359 & n23898 ) | ( n23896 & n23898 ) ;
  assign n23893 = n15642 ^ n8409 ^ 1'b0 ;
  assign n23894 = n1572 & n23893 ;
  assign n23900 = n23899 ^ n23894 ^ 1'b0 ;
  assign n23901 = ( ~n528 & n5085 ) | ( ~n528 & n17031 ) | ( n5085 & n17031 ) ;
  assign n23902 = n4554 & ~n23901 ;
  assign n23903 = n23663 ^ n12119 ^ 1'b0 ;
  assign n23904 = n3912 & ~n23903 ;
  assign n23905 = ( ~n476 & n1231 ) | ( ~n476 & n23904 ) | ( n1231 & n23904 ) ;
  assign n23906 = ( n20373 & n23902 ) | ( n20373 & ~n23905 ) | ( n23902 & ~n23905 ) ;
  assign n23908 = n18960 ^ n14766 ^ n446 ;
  assign n23907 = n10800 & n12646 ;
  assign n23909 = n23908 ^ n23907 ^ 1'b0 ;
  assign n23910 = n12889 & n15663 ;
  assign n23911 = n18127 & n23910 ;
  assign n23912 = n15797 ^ n11205 ^ n9719 ;
  assign n23915 = n1113 & ~n5918 ;
  assign n23913 = n6905 & ~n13949 ;
  assign n23914 = n23913 ^ n13200 ^ 1'b0 ;
  assign n23916 = n23915 ^ n23914 ^ 1'b0 ;
  assign n23917 = n10374 & n23916 ;
  assign n23918 = ( ~n17976 & n22245 ) | ( ~n17976 & n23057 ) | ( n22245 & n23057 ) ;
  assign n23919 = ~n1635 & n5817 ;
  assign n23920 = n23919 ^ n10066 ^ 1'b0 ;
  assign n23921 = n13219 | n21825 ;
  assign n23922 = ( n7830 & n8233 ) | ( n7830 & n22922 ) | ( n8233 & n22922 ) ;
  assign n23923 = n4452 | n10016 ;
  assign n23924 = n23922 & ~n23923 ;
  assign n23925 = n4757 & ~n9176 ;
  assign n23926 = n23925 ^ n8339 ^ 1'b0 ;
  assign n23927 = ( ~n4633 & n23924 ) | ( ~n4633 & n23926 ) | ( n23924 & n23926 ) ;
  assign n23928 = n9181 & ~n16171 ;
  assign n23929 = n23928 ^ n2763 ^ 1'b0 ;
  assign n23930 = n5851 & n23929 ;
  assign n23931 = ( ~n3793 & n9487 ) | ( ~n3793 & n10230 ) | ( n9487 & n10230 ) ;
  assign n23932 = n23931 ^ n9408 ^ n7292 ;
  assign n23933 = n9014 ^ n2298 ^ 1'b0 ;
  assign n23934 = n10342 ^ n2073 ^ 1'b0 ;
  assign n23935 = ( n3869 & n23933 ) | ( n3869 & n23934 ) | ( n23933 & n23934 ) ;
  assign n23936 = n23932 & ~n23935 ;
  assign n23937 = n8259 | n10739 ;
  assign n23938 = n2442 | n9829 ;
  assign n23939 = ( n7345 & n9189 ) | ( n7345 & ~n18321 ) | ( n9189 & ~n18321 ) ;
  assign n23940 = ( n467 & ~n6459 ) | ( n467 & n23939 ) | ( ~n6459 & n23939 ) ;
  assign n23941 = ( n2657 & ~n7397 ) | ( n2657 & n8065 ) | ( ~n7397 & n8065 ) ;
  assign n23942 = n23088 ^ n6745 ^ n6376 ;
  assign n23943 = ( n6111 & ~n15377 ) | ( n6111 & n23186 ) | ( ~n15377 & n23186 ) ;
  assign n23944 = ( n6623 & n14002 ) | ( n6623 & n23943 ) | ( n14002 & n23943 ) ;
  assign n23945 = ( n21729 & n23942 ) | ( n21729 & ~n23944 ) | ( n23942 & ~n23944 ) ;
  assign n23946 = ( n708 & ~n7908 ) | ( n708 & n18489 ) | ( ~n7908 & n18489 ) ;
  assign n23947 = n6999 ^ n3606 ^ 1'b0 ;
  assign n23948 = ( n2237 & n5838 ) | ( n2237 & ~n23947 ) | ( n5838 & ~n23947 ) ;
  assign n23949 = n23948 ^ n10921 ^ n4205 ;
  assign n23950 = n14432 ^ n8625 ^ 1'b0 ;
  assign n23951 = n19628 & n23950 ;
  assign n23952 = n23951 ^ n4476 ^ 1'b0 ;
  assign n23953 = n23949 & ~n23952 ;
  assign n23954 = n10998 & n23953 ;
  assign n23955 = n7687 ^ n3562 ^ 1'b0 ;
  assign n23956 = n1383 & n3701 ;
  assign n23957 = n17484 & n23956 ;
  assign n23958 = ( ~n8923 & n23955 ) | ( ~n8923 & n23957 ) | ( n23955 & n23957 ) ;
  assign n23959 = ~n5130 & n11936 ;
  assign n23970 = ( x105 & ~n5770 ) | ( x105 & n11878 ) | ( ~n5770 & n11878 ) ;
  assign n23968 = ( n2379 & n7766 ) | ( n2379 & ~n8152 ) | ( n7766 & ~n8152 ) ;
  assign n23969 = ( n617 & n16806 ) | ( n617 & ~n23968 ) | ( n16806 & ~n23968 ) ;
  assign n23960 = n6933 ^ n2164 ^ 1'b0 ;
  assign n23961 = n21318 ^ n17199 ^ n16918 ;
  assign n23962 = n23960 | n23961 ;
  assign n23963 = n19590 ^ n16573 ^ 1'b0 ;
  assign n23964 = ~n1635 & n23963 ;
  assign n23965 = n12861 & n23964 ;
  assign n23966 = ( n8178 & n23962 ) | ( n8178 & n23965 ) | ( n23962 & n23965 ) ;
  assign n23967 = n23966 ^ n18325 ^ n8436 ;
  assign n23971 = n23970 ^ n23969 ^ n23967 ;
  assign n23972 = ( n8654 & n15715 ) | ( n8654 & ~n16454 ) | ( n15715 & ~n16454 ) ;
  assign n23973 = n1158 & ~n14979 ;
  assign n23974 = n23973 ^ n8709 ^ 1'b0 ;
  assign n23975 = n23974 ^ n7338 ^ n845 ;
  assign n23976 = ( n16242 & n16322 ) | ( n16242 & n23975 ) | ( n16322 & n23975 ) ;
  assign n23977 = ( n8687 & ~n13726 ) | ( n8687 & n20330 ) | ( ~n13726 & n20330 ) ;
  assign n23978 = ~n8570 & n20077 ;
  assign n23979 = n23978 ^ n17330 ^ 1'b0 ;
  assign n23980 = n9767 & ~n23979 ;
  assign n23981 = n23980 ^ n22313 ^ 1'b0 ;
  assign n23994 = ( ~n1461 & n4608 ) | ( ~n1461 & n4992 ) | ( n4608 & n4992 ) ;
  assign n23995 = n23994 ^ n9807 ^ n6118 ;
  assign n23990 = ( n1104 & n5199 ) | ( n1104 & n6271 ) | ( n5199 & n6271 ) ;
  assign n23991 = n23990 ^ n7712 ^ 1'b0 ;
  assign n23992 = n5637 | n23991 ;
  assign n23993 = n23992 ^ n17383 ^ n8168 ;
  assign n23982 = n19739 ^ n5676 ^ n5425 ;
  assign n23983 = ( n8694 & n10960 ) | ( n8694 & n23982 ) | ( n10960 & n23982 ) ;
  assign n23984 = n7100 ^ n5463 ^ n4300 ;
  assign n23985 = n23984 ^ n14917 ^ 1'b0 ;
  assign n23986 = n23983 & ~n23985 ;
  assign n23987 = n3515 ^ n1694 ^ n1544 ;
  assign n23988 = n23987 ^ n21184 ^ 1'b0 ;
  assign n23989 = ( n4375 & ~n23986 ) | ( n4375 & n23988 ) | ( ~n23986 & n23988 ) ;
  assign n23996 = n23995 ^ n23993 ^ n23989 ;
  assign n23997 = n23411 ^ n8874 ^ n903 ;
  assign n23998 = n2540 | n4835 ;
  assign n23999 = n23998 ^ n1262 ^ 1'b0 ;
  assign n24000 = ( ~n9187 & n13974 ) | ( ~n9187 & n23999 ) | ( n13974 & n23999 ) ;
  assign n24001 = ( n11426 & n23997 ) | ( n11426 & n24000 ) | ( n23997 & n24000 ) ;
  assign n24002 = n17733 ^ n12860 ^ 1'b0 ;
  assign n24003 = ~n22877 & n24002 ;
  assign n24004 = n24003 ^ n19396 ^ n8949 ;
  assign n24005 = n12699 ^ n8586 ^ 1'b0 ;
  assign n24006 = n13793 & ~n24005 ;
  assign n24007 = n14146 ^ n9473 ^ n7181 ;
  assign n24008 = n24007 ^ n4647 ^ n740 ;
  assign n24009 = ( n11155 & n24006 ) | ( n11155 & ~n24008 ) | ( n24006 & ~n24008 ) ;
  assign n24010 = n9754 & n11186 ;
  assign n24011 = n6812 | n10369 ;
  assign n24012 = n24011 ^ n11631 ^ 1'b0 ;
  assign n24013 = ( n2661 & n24010 ) | ( n2661 & n24012 ) | ( n24010 & n24012 ) ;
  assign n24014 = ( n7273 & n14321 ) | ( n7273 & n24013 ) | ( n14321 & n24013 ) ;
  assign n24016 = ( n869 & n5236 ) | ( n869 & n11961 ) | ( n5236 & n11961 ) ;
  assign n24017 = ( n5774 & n5786 ) | ( n5774 & ~n24016 ) | ( n5786 & ~n24016 ) ;
  assign n24015 = n13053 ^ n9864 ^ n8775 ;
  assign n24018 = n24017 ^ n24015 ^ n7886 ;
  assign n24019 = n24018 ^ n16383 ^ n11000 ;
  assign n24020 = n3214 & ~n24019 ;
  assign n24021 = n8488 | n24020 ;
  assign n24022 = n903 & ~n24021 ;
  assign n24023 = n1006 & ~n21076 ;
  assign n24024 = ~n3027 & n24023 ;
  assign n24025 = n9477 ^ n6359 ^ 1'b0 ;
  assign n24026 = ( n4752 & n8673 ) | ( n4752 & ~n24024 ) | ( n8673 & ~n24024 ) ;
  assign n24027 = n7551 & ~n12473 ;
  assign n24028 = n7603 & n24027 ;
  assign n24029 = n19045 & ~n24028 ;
  assign n24030 = ~n24026 & n24029 ;
  assign n24031 = n24025 | n24030 ;
  assign n24032 = n2022 & ~n24031 ;
  assign n24033 = n24032 ^ n21851 ^ n4046 ;
  assign n24034 = n5948 & n24033 ;
  assign n24035 = n24034 ^ n12936 ^ 1'b0 ;
  assign n24036 = n24024 | n24035 ;
  assign n24037 = n2815 | n24036 ;
  assign n24038 = ~n10139 & n17915 ;
  assign n24039 = n16379 & n24038 ;
  assign n24040 = ( n9002 & n21032 ) | ( n9002 & n24039 ) | ( n21032 & n24039 ) ;
  assign n24041 = n24040 ^ n14679 ^ n6400 ;
  assign n24042 = ( n12857 & n15270 ) | ( n12857 & ~n23032 ) | ( n15270 & ~n23032 ) ;
  assign n24043 = n24042 ^ n10162 ^ 1'b0 ;
  assign n24044 = n8654 ^ n7601 ^ n2757 ;
  assign n24045 = n17091 | n24044 ;
  assign n24046 = n24045 ^ n3797 ^ 1'b0 ;
  assign n24047 = n21546 & ~n24046 ;
  assign n24048 = n17110 | n18127 ;
  assign n24049 = ( n791 & n2325 ) | ( n791 & n24048 ) | ( n2325 & n24048 ) ;
  assign n24050 = n6059 | n11271 ;
  assign n24051 = n2100 & ~n24050 ;
  assign n24052 = n5705 & n17262 ;
  assign n24053 = n5017 & n24052 ;
  assign n24054 = ~n12842 & n24053 ;
  assign n24055 = n6618 ^ n4519 ^ 1'b0 ;
  assign n24056 = ~n20947 & n24055 ;
  assign n24057 = ( ~n24051 & n24054 ) | ( ~n24051 & n24056 ) | ( n24054 & n24056 ) ;
  assign n24058 = n24057 ^ n19828 ^ n9697 ;
  assign n24059 = ( ~n4145 & n20105 ) | ( ~n4145 & n21110 ) | ( n20105 & n21110 ) ;
  assign n24063 = n13420 ^ n4519 ^ n2957 ;
  assign n24061 = ~n15845 & n16681 ;
  assign n24062 = n6341 | n24061 ;
  assign n24060 = n21522 ^ n19144 ^ n9362 ;
  assign n24064 = n24063 ^ n24062 ^ n24060 ;
  assign n24065 = ~n10721 & n16462 ;
  assign n24066 = n24065 ^ n18200 ^ 1'b0 ;
  assign n24068 = n1339 & ~n15741 ;
  assign n24069 = n24068 ^ n10640 ^ 1'b0 ;
  assign n24067 = n10989 ^ n7508 ^ n6655 ;
  assign n24070 = n24069 ^ n24067 ^ n1606 ;
  assign n24071 = ( n3410 & ~n23207 ) | ( n3410 & n24070 ) | ( ~n23207 & n24070 ) ;
  assign n24072 = n15911 ^ n1186 ^ 1'b0 ;
  assign n24073 = ( x70 & n2275 ) | ( x70 & n24072 ) | ( n2275 & n24072 ) ;
  assign n24074 = ( n1129 & n3715 ) | ( n1129 & ~n22286 ) | ( n3715 & ~n22286 ) ;
  assign n24075 = n1580 & n24074 ;
  assign n24076 = ( n2076 & ~n2893 ) | ( n2076 & n23853 ) | ( ~n2893 & n23853 ) ;
  assign n24077 = n6673 | n24076 ;
  assign n24078 = n24075 | n24077 ;
  assign n24079 = n24078 ^ n24037 ^ n16409 ;
  assign n24080 = n7217 & ~n11752 ;
  assign n24081 = n2069 | n24080 ;
  assign n24082 = n5382 ^ n4963 ^ 1'b0 ;
  assign n24083 = ~n9141 & n24082 ;
  assign n24084 = ~n1302 & n24083 ;
  assign n24087 = n11916 ^ n10174 ^ 1'b0 ;
  assign n24088 = n11029 & n24087 ;
  assign n24085 = n6414 ^ n3561 ^ n1422 ;
  assign n24086 = n24085 ^ n4124 ^ n1195 ;
  assign n24089 = n24088 ^ n24086 ^ 1'b0 ;
  assign n24090 = ( ~n9463 & n24084 ) | ( ~n9463 & n24089 ) | ( n24084 & n24089 ) ;
  assign n24093 = n9022 ^ n1067 ^ 1'b0 ;
  assign n24094 = ( n6988 & n21091 ) | ( n6988 & ~n24093 ) | ( n21091 & ~n24093 ) ;
  assign n24091 = n9066 ^ x247 ^ 1'b0 ;
  assign n24092 = n8614 & ~n24091 ;
  assign n24095 = n24094 ^ n24092 ^ n12122 ;
  assign n24096 = ( n10378 & n13012 ) | ( n10378 & ~n21988 ) | ( n13012 & ~n21988 ) ;
  assign n24099 = n16788 ^ n15288 ^ n5353 ;
  assign n24098 = ~n666 & n16862 ;
  assign n24100 = n24099 ^ n24098 ^ 1'b0 ;
  assign n24097 = n16054 | n21840 ;
  assign n24101 = n24100 ^ n24097 ^ 1'b0 ;
  assign n24102 = n3813 | n18532 ;
  assign n24103 = n2342 & n6745 ;
  assign n24104 = n24103 ^ n3474 ^ n1664 ;
  assign n24105 = n12158 | n16595 ;
  assign n24106 = n24105 ^ n13295 ^ n485 ;
  assign n24107 = ~n10082 & n24106 ;
  assign n24108 = n11040 & n24107 ;
  assign n24109 = ( n1391 & ~n4794 ) | ( n1391 & n5069 ) | ( ~n4794 & n5069 ) ;
  assign n24110 = n886 & n9714 ;
  assign n24111 = n24110 ^ n4135 ^ 1'b0 ;
  assign n24112 = ( n21189 & n21539 ) | ( n21189 & n24111 ) | ( n21539 & n24111 ) ;
  assign n24113 = n19748 & ~n24112 ;
  assign n24114 = n328 & n16389 ;
  assign n24115 = n19114 & n24114 ;
  assign n24116 = ( n686 & n7910 ) | ( n686 & ~n12957 ) | ( n7910 & ~n12957 ) ;
  assign n24117 = n14336 & n24116 ;
  assign n24118 = ( n3102 & n24115 ) | ( n3102 & n24117 ) | ( n24115 & n24117 ) ;
  assign n24119 = n24118 ^ n21265 ^ 1'b0 ;
  assign n24120 = ( ~n7373 & n9897 ) | ( ~n7373 & n10241 ) | ( n9897 & n10241 ) ;
  assign n24121 = n23289 ^ n3439 ^ 1'b0 ;
  assign n24122 = n2877 | n19341 ;
  assign n24123 = n3214 | n24122 ;
  assign n24124 = n24123 ^ n12066 ^ 1'b0 ;
  assign n24126 = n9402 ^ n2937 ^ n803 ;
  assign n24125 = ~n3101 & n3744 ;
  assign n24127 = n24126 ^ n24125 ^ 1'b0 ;
  assign n24128 = ~n3062 & n24127 ;
  assign n24129 = n24128 ^ n19603 ^ n827 ;
  assign n24130 = ~n5719 & n23737 ;
  assign n24131 = n6220 | n14016 ;
  assign n24132 = ( n5617 & n5996 ) | ( n5617 & n12695 ) | ( n5996 & n12695 ) ;
  assign n24133 = n24132 ^ n6728 ^ n586 ;
  assign n24134 = n5080 & n9277 ;
  assign n24135 = n10303 & n24134 ;
  assign n24136 = n7342 ^ n2043 ^ 1'b0 ;
  assign n24140 = n20521 ^ n8662 ^ n6857 ;
  assign n24137 = n10240 ^ n9002 ^ n4909 ;
  assign n24138 = n24137 ^ n15732 ^ n8492 ;
  assign n24139 = x28 & n24138 ;
  assign n24141 = n24140 ^ n24139 ^ n12702 ;
  assign n24142 = ( ~n4649 & n24136 ) | ( ~n4649 & n24141 ) | ( n24136 & n24141 ) ;
  assign n24143 = n24142 ^ n14513 ^ 1'b0 ;
  assign n24144 = n6130 & ~n24143 ;
  assign n24145 = n5576 & n24144 ;
  assign n24146 = ( n23762 & ~n24135 ) | ( n23762 & n24145 ) | ( ~n24135 & n24145 ) ;
  assign n24147 = n19979 ^ n1361 ^ 1'b0 ;
  assign n24148 = n2527 | n24147 ;
  assign n24149 = n17151 ^ n13847 ^ n788 ;
  assign n24150 = ( n2538 & n5292 ) | ( n2538 & ~n21189 ) | ( n5292 & ~n21189 ) ;
  assign n24151 = n24149 | n24150 ;
  assign n24152 = n24151 ^ n16345 ^ 1'b0 ;
  assign n24153 = ~n24148 & n24152 ;
  assign n24154 = ~n948 & n2648 ;
  assign n24155 = ~n1548 & n24154 ;
  assign n24156 = ~n5613 & n24155 ;
  assign n24157 = n11869 | n24156 ;
  assign n24158 = n24157 ^ n10684 ^ 1'b0 ;
  assign n24159 = n8257 & ~n8454 ;
  assign n24160 = ~n1637 & n24159 ;
  assign n24161 = n20205 ^ n19106 ^ n1626 ;
  assign n24162 = ( n8501 & n24160 ) | ( n8501 & ~n24161 ) | ( n24160 & ~n24161 ) ;
  assign n24163 = n24162 ^ n10587 ^ 1'b0 ;
  assign n24164 = n24163 ^ n19065 ^ 1'b0 ;
  assign n24165 = n11131 & n15776 ;
  assign n24170 = n7907 ^ n7759 ^ 1'b0 ;
  assign n24171 = n24170 ^ n7185 ^ n1514 ;
  assign n24168 = n15169 ^ n6442 ^ 1'b0 ;
  assign n24169 = n3949 & ~n24168 ;
  assign n24166 = n8126 | n13140 ;
  assign n24167 = ( n2657 & ~n16479 ) | ( n2657 & n24166 ) | ( ~n16479 & n24166 ) ;
  assign n24172 = n24171 ^ n24169 ^ n24167 ;
  assign n24173 = n19214 & ~n22630 ;
  assign n24174 = ~n9985 & n24173 ;
  assign n24175 = n11226 ^ n10152 ^ n9047 ;
  assign n24176 = ( n10801 & n10880 ) | ( n10801 & ~n24175 ) | ( n10880 & ~n24175 ) ;
  assign n24177 = n24176 ^ n8155 ^ 1'b0 ;
  assign n24178 = ( n2746 & ~n5359 ) | ( n2746 & n16174 ) | ( ~n5359 & n16174 ) ;
  assign n24179 = n24178 ^ n5906 ^ n460 ;
  assign n24180 = n5890 & n24179 ;
  assign n24181 = n21739 & n24180 ;
  assign n24182 = n11944 | n24181 ;
  assign n24183 = n18067 ^ n2206 ^ x242 ;
  assign n24184 = ~n21739 & n24183 ;
  assign n24185 = n5623 ^ n3111 ^ n2832 ;
  assign n24186 = n24185 ^ n20077 ^ n9501 ;
  assign n24187 = ( n3423 & n10028 ) | ( n3423 & n24186 ) | ( n10028 & n24186 ) ;
  assign n24188 = ( n18298 & n24184 ) | ( n18298 & ~n24187 ) | ( n24184 & ~n24187 ) ;
  assign n24189 = n1299 & ~n2288 ;
  assign n24190 = n24189 ^ n12243 ^ 1'b0 ;
  assign n24191 = n24190 ^ n9099 ^ 1'b0 ;
  assign n24192 = ( n1882 & n14750 ) | ( n1882 & n16365 ) | ( n14750 & n16365 ) ;
  assign n24193 = ( n1172 & n3351 ) | ( n1172 & ~n24192 ) | ( n3351 & ~n24192 ) ;
  assign n24194 = n8850 ^ x246 ^ 1'b0 ;
  assign n24195 = ( n3943 & n24193 ) | ( n3943 & ~n24194 ) | ( n24193 & ~n24194 ) ;
  assign n24196 = ~n9073 & n13132 ;
  assign n24197 = ( x134 & n6434 ) | ( x134 & n24196 ) | ( n6434 & n24196 ) ;
  assign n24198 = n24197 ^ n15868 ^ n7227 ;
  assign n24199 = n24198 ^ n4017 ^ x177 ;
  assign n24200 = n23425 ^ n10654 ^ 1'b0 ;
  assign n24205 = n8547 ^ n485 ^ 1'b0 ;
  assign n24206 = n5245 | n24205 ;
  assign n24207 = n8922 | n24206 ;
  assign n24208 = ( n13477 & n21365 ) | ( n13477 & n24207 ) | ( n21365 & n24207 ) ;
  assign n24202 = n2139 & ~n5253 ;
  assign n24203 = n18921 & ~n24202 ;
  assign n24201 = n653 & n14244 ;
  assign n24204 = n24203 ^ n24201 ^ 1'b0 ;
  assign n24209 = n24208 ^ n24204 ^ n15563 ;
  assign n24210 = n16771 ^ n1610 ^ x40 ;
  assign n24211 = n10270 ^ n7326 ^ n5235 ;
  assign n24212 = ( n16227 & ~n24210 ) | ( n16227 & n24211 ) | ( ~n24210 & n24211 ) ;
  assign n24213 = n24212 ^ n15573 ^ n10930 ;
  assign n24214 = ( n14398 & n23730 ) | ( n14398 & n24213 ) | ( n23730 & n24213 ) ;
  assign n24215 = n24214 ^ n10663 ^ 1'b0 ;
  assign n24216 = n24209 & ~n24215 ;
  assign n24221 = n17977 ^ n10112 ^ 1'b0 ;
  assign n24222 = n14449 | n24221 ;
  assign n24218 = n6396 ^ n3130 ^ n3102 ;
  assign n24217 = n3147 & n16307 ;
  assign n24219 = n24218 ^ n24217 ^ 1'b0 ;
  assign n24220 = n3929 | n24219 ;
  assign n24223 = n24222 ^ n24220 ^ 1'b0 ;
  assign n24224 = ( ~x24 & n12064 ) | ( ~x24 & n12475 ) | ( n12064 & n12475 ) ;
  assign n24225 = n15956 | n24224 ;
  assign n24226 = n23962 ^ n12128 ^ 1'b0 ;
  assign n24227 = ( n1647 & n4062 ) | ( n1647 & ~n6370 ) | ( n4062 & ~n6370 ) ;
  assign n24228 = n24227 ^ n8603 ^ n1507 ;
  assign n24229 = ~n6532 & n8614 ;
  assign n24230 = ~n2992 & n24229 ;
  assign n24231 = x67 & ~n24230 ;
  assign n24232 = ~n24228 & n24231 ;
  assign n24233 = n24232 ^ n10921 ^ 1'b0 ;
  assign n24234 = ~n1866 & n24233 ;
  assign n24235 = n24234 ^ n15784 ^ n13380 ;
  assign n24236 = n24235 ^ n15770 ^ n13008 ;
  assign n24237 = n24236 ^ n19718 ^ n5418 ;
  assign n24238 = n5233 & ~n20669 ;
  assign n24239 = n4262 & n24238 ;
  assign n24240 = n7655 ^ x140 ^ 1'b0 ;
  assign n24241 = ~n24239 & n24240 ;
  assign n24242 = n865 & n24241 ;
  assign n24243 = ~n6923 & n24242 ;
  assign n24247 = ~x4 & n19454 ;
  assign n24248 = n3433 & n24247 ;
  assign n24244 = n365 & n2086 ;
  assign n24245 = ( n3599 & ~n17559 ) | ( n3599 & n24244 ) | ( ~n17559 & n24244 ) ;
  assign n24246 = n24245 ^ n13652 ^ 1'b0 ;
  assign n24249 = n24248 ^ n24246 ^ 1'b0 ;
  assign n24250 = ~n4328 & n24249 ;
  assign n24251 = n8638 & ~n9101 ;
  assign n24252 = n24251 ^ n12413 ^ 1'b0 ;
  assign n24253 = ( n8364 & ~n13548 ) | ( n8364 & n24252 ) | ( ~n13548 & n24252 ) ;
  assign n24254 = n20314 ^ n18080 ^ n16443 ;
  assign n24255 = ( n6101 & n20997 ) | ( n6101 & n22501 ) | ( n20997 & n22501 ) ;
  assign n24256 = ( ~n563 & n2339 ) | ( ~n563 & n4044 ) | ( n2339 & n4044 ) ;
  assign n24257 = n24256 ^ n20894 ^ 1'b0 ;
  assign n24258 = n24257 ^ n1452 ^ 1'b0 ;
  assign n24259 = n3594 | n19946 ;
  assign n24260 = n4017 | n24259 ;
  assign n24261 = ( n905 & ~n13900 ) | ( n905 & n24260 ) | ( ~n13900 & n24260 ) ;
  assign n24262 = n17611 & n24261 ;
  assign n24263 = ( ~n9002 & n21762 ) | ( ~n9002 & n23880 ) | ( n21762 & n23880 ) ;
  assign n24264 = ( ~n717 & n3173 ) | ( ~n717 & n7768 ) | ( n3173 & n7768 ) ;
  assign n24265 = ( n7111 & n16447 ) | ( n7111 & ~n24264 ) | ( n16447 & ~n24264 ) ;
  assign n24266 = ( n5718 & ~n13869 ) | ( n5718 & n24265 ) | ( ~n13869 & n24265 ) ;
  assign n24267 = ( n3414 & n16573 ) | ( n3414 & n24266 ) | ( n16573 & n24266 ) ;
  assign n24268 = ( n16016 & ~n21142 ) | ( n16016 & n24267 ) | ( ~n21142 & n24267 ) ;
  assign n24269 = ~n2797 & n11882 ;
  assign n24270 = ~n5966 & n24269 ;
  assign n24271 = n5749 ^ n4357 ^ n2857 ;
  assign n24272 = ~n565 & n10057 ;
  assign n24273 = ~n16687 & n24272 ;
  assign n24274 = ( n24270 & ~n24271 ) | ( n24270 & n24273 ) | ( ~n24271 & n24273 ) ;
  assign n24275 = ( n4841 & ~n13378 ) | ( n4841 & n13737 ) | ( ~n13378 & n13737 ) ;
  assign n24276 = n7327 | n17790 ;
  assign n24277 = n24275 & ~n24276 ;
  assign n24279 = n6310 ^ n2221 ^ 1'b0 ;
  assign n24280 = n24279 ^ n19452 ^ n18045 ;
  assign n24281 = n24280 ^ n1330 ^ 1'b0 ;
  assign n24278 = n8547 ^ n3041 ^ n2016 ;
  assign n24282 = n24281 ^ n24278 ^ n20475 ;
  assign n24283 = ( n10853 & n13580 ) | ( n10853 & ~n17387 ) | ( n13580 & ~n17387 ) ;
  assign n24284 = n24283 ^ n18146 ^ 1'b0 ;
  assign n24285 = n4245 | n24284 ;
  assign n24286 = n10849 & ~n17721 ;
  assign n24287 = n5245 & n24286 ;
  assign n24288 = n16395 ^ n8499 ^ n4342 ;
  assign n24289 = ( n1957 & n11642 ) | ( n1957 & n24288 ) | ( n11642 & n24288 ) ;
  assign n24290 = ~n14100 & n23562 ;
  assign n24291 = n24290 ^ n20058 ^ 1'b0 ;
  assign n24292 = n23099 & ~n24291 ;
  assign n24293 = n3157 & ~n24292 ;
  assign n24294 = n12816 ^ n5290 ^ n1869 ;
  assign n24295 = n10485 ^ n3599 ^ 1'b0 ;
  assign n24296 = n24294 & n24295 ;
  assign n24298 = ( n7906 & ~n8790 ) | ( n7906 & n18484 ) | ( ~n8790 & n18484 ) ;
  assign n24297 = n19420 ^ n11782 ^ 1'b0 ;
  assign n24299 = n24298 ^ n24297 ^ n3384 ;
  assign n24300 = ( ~n4970 & n5479 ) | ( ~n4970 & n24299 ) | ( n5479 & n24299 ) ;
  assign n24301 = n8441 ^ n1799 ^ x49 ;
  assign n24302 = ( n13273 & ~n22218 ) | ( n13273 & n24301 ) | ( ~n22218 & n24301 ) ;
  assign n24303 = n7823 & n23270 ;
  assign n24304 = n18257 & n24303 ;
  assign n24305 = n24304 ^ x222 ^ 1'b0 ;
  assign n24306 = n24305 ^ n17557 ^ n2506 ;
  assign n24307 = ( n5818 & n16132 ) | ( n5818 & ~n24306 ) | ( n16132 & ~n24306 ) ;
  assign n24308 = n24307 ^ n21858 ^ n18762 ;
  assign n24309 = ( ~n7387 & n8021 ) | ( ~n7387 & n8882 ) | ( n8021 & n8882 ) ;
  assign n24313 = n2113 & ~n2931 ;
  assign n24310 = n23578 ^ n8790 ^ n2459 ;
  assign n24311 = ( n9795 & n10988 ) | ( n9795 & ~n24310 ) | ( n10988 & ~n24310 ) ;
  assign n24312 = n24311 ^ n8276 ^ 1'b0 ;
  assign n24314 = n24313 ^ n24312 ^ n14502 ;
  assign n24321 = n2433 ^ n1761 ^ 1'b0 ;
  assign n24317 = n10792 ^ n8017 ^ n6375 ;
  assign n24315 = x148 & ~n17783 ;
  assign n24316 = n9429 & n24315 ;
  assign n24318 = n24317 ^ n24316 ^ 1'b0 ;
  assign n24319 = ~n13674 & n24318 ;
  assign n24320 = n24319 ^ n14939 ^ 1'b0 ;
  assign n24322 = n24321 ^ n24320 ^ n10662 ;
  assign n24323 = n9729 & n10897 ;
  assign n24324 = n24323 ^ n18461 ^ n15191 ;
  assign n24325 = n5362 | n10036 ;
  assign n24326 = n5947 & ~n24325 ;
  assign n24327 = n5808 | n12341 ;
  assign n24328 = n24327 ^ n23987 ^ n22885 ;
  assign n24329 = n4824 & ~n10735 ;
  assign n24330 = n24329 ^ n23281 ^ n16645 ;
  assign n24331 = n12656 ^ n8616 ^ n788 ;
  assign n24332 = n5857 ^ n3738 ^ 1'b0 ;
  assign n24333 = n8240 ^ n6451 ^ n4442 ;
  assign n24334 = n1168 | n10360 ;
  assign n24335 = n24333 | n24334 ;
  assign n24336 = ( ~n15907 & n24332 ) | ( ~n15907 & n24335 ) | ( n24332 & n24335 ) ;
  assign n24337 = n17967 ^ n12762 ^ n376 ;
  assign n24338 = n24337 ^ n18128 ^ 1'b0 ;
  assign n24339 = ( n12056 & n18349 ) | ( n12056 & ~n24338 ) | ( n18349 & ~n24338 ) ;
  assign n24340 = n14625 ^ n14430 ^ 1'b0 ;
  assign n24342 = ( ~n8755 & n13084 ) | ( ~n8755 & n18895 ) | ( n13084 & n18895 ) ;
  assign n24343 = ( n2094 & n13205 ) | ( n2094 & ~n17940 ) | ( n13205 & ~n17940 ) ;
  assign n24344 = ( n18637 & ~n24342 ) | ( n18637 & n24343 ) | ( ~n24342 & n24343 ) ;
  assign n24345 = n12242 & ~n20222 ;
  assign n24346 = n9722 & n24345 ;
  assign n24347 = n24346 ^ n12635 ^ n1722 ;
  assign n24348 = n10940 ^ n4338 ^ n1762 ;
  assign n24349 = ( n1575 & n24347 ) | ( n1575 & ~n24348 ) | ( n24347 & ~n24348 ) ;
  assign n24350 = n24349 ^ n9228 ^ 1'b0 ;
  assign n24351 = ( n10863 & n24344 ) | ( n10863 & ~n24350 ) | ( n24344 & ~n24350 ) ;
  assign n24341 = n702 & n18551 ;
  assign n24352 = n24351 ^ n24341 ^ 1'b0 ;
  assign n24353 = ( ~n14725 & n15647 ) | ( ~n14725 & n24352 ) | ( n15647 & n24352 ) ;
  assign n24354 = n12095 ^ n1591 ^ 1'b0 ;
  assign n24355 = n2198 & ~n24354 ;
  assign n24356 = n24355 ^ n5849 ^ 1'b0 ;
  assign n24357 = n8818 ^ n3200 ^ n2026 ;
  assign n24358 = n24357 ^ n5890 ^ n4600 ;
  assign n24359 = n24358 ^ n8839 ^ 1'b0 ;
  assign n24360 = n4474 | n24359 ;
  assign n24361 = ( ~n2006 & n3438 ) | ( ~n2006 & n7432 ) | ( n3438 & n7432 ) ;
  assign n24362 = n5233 & n8339 ;
  assign n24363 = ~n24361 & n24362 ;
  assign n24364 = n24128 & ~n24363 ;
  assign n24365 = n19365 ^ n1716 ^ n1347 ;
  assign n24367 = n15414 ^ n14038 ^ 1'b0 ;
  assign n24366 = n11760 ^ n2170 ^ n956 ;
  assign n24368 = n24367 ^ n24366 ^ 1'b0 ;
  assign n24369 = n6949 ^ n4197 ^ 1'b0 ;
  assign n24370 = n24369 ^ n15736 ^ n478 ;
  assign n24371 = ( ~n6143 & n10718 ) | ( ~n6143 & n15302 ) | ( n10718 & n15302 ) ;
  assign n24372 = ~n18119 & n24371 ;
  assign n24373 = n24372 ^ n9033 ^ 1'b0 ;
  assign n24374 = n1843 | n5367 ;
  assign n24375 = n17877 & n24374 ;
  assign n24376 = n11587 & n24375 ;
  assign n24377 = n10118 | n11481 ;
  assign n24378 = n22573 ^ n1509 ^ 1'b0 ;
  assign n24379 = ( n24376 & n24377 ) | ( n24376 & ~n24378 ) | ( n24377 & ~n24378 ) ;
  assign n24389 = n10067 ^ n5562 ^ n1980 ;
  assign n24387 = ( n3130 & n4405 ) | ( n3130 & n6383 ) | ( n4405 & n6383 ) ;
  assign n24388 = n7236 & n24387 ;
  assign n24390 = n24389 ^ n24388 ^ 1'b0 ;
  assign n24380 = n10721 ^ n6918 ^ n5350 ;
  assign n24381 = ( n2163 & n5780 ) | ( n2163 & n8054 ) | ( n5780 & n8054 ) ;
  assign n24382 = ( n2842 & n4792 ) | ( n2842 & n7263 ) | ( n4792 & n7263 ) ;
  assign n24383 = n24381 & ~n24382 ;
  assign n24384 = n24383 ^ n21640 ^ 1'b0 ;
  assign n24385 = n24380 & ~n24384 ;
  assign n24386 = ( n7788 & n19970 ) | ( n7788 & ~n24385 ) | ( n19970 & ~n24385 ) ;
  assign n24391 = n24390 ^ n24386 ^ n3710 ;
  assign n24393 = n1001 & n3411 ;
  assign n24394 = n24393 ^ n11170 ^ 1'b0 ;
  assign n24395 = ( n2450 & ~n9678 ) | ( n2450 & n24394 ) | ( ~n9678 & n24394 ) ;
  assign n24392 = n17822 ^ n8672 ^ n6890 ;
  assign n24396 = n24395 ^ n24392 ^ n2442 ;
  assign n24397 = n24391 & n24396 ;
  assign n24398 = x247 & n4600 ;
  assign n24399 = n19102 ^ n14038 ^ n5910 ;
  assign n24400 = n12972 ^ n12150 ^ n6199 ;
  assign n24401 = ( n8525 & ~n10096 ) | ( n8525 & n14789 ) | ( ~n10096 & n14789 ) ;
  assign n24402 = n19646 ^ n6736 ^ n3026 ;
  assign n24403 = n5021 & n24402 ;
  assign n24404 = ( ~n20324 & n22941 ) | ( ~n20324 & n24403 ) | ( n22941 & n24403 ) ;
  assign n24405 = n9472 ^ n6103 ^ n1484 ;
  assign n24406 = n758 | n17914 ;
  assign n24407 = n2451 & ~n24406 ;
  assign n24408 = n24407 ^ n14155 ^ 1'b0 ;
  assign n24409 = ( x229 & n2222 ) | ( x229 & n24408 ) | ( n2222 & n24408 ) ;
  assign n24410 = ( n2926 & n10017 ) | ( n2926 & n24409 ) | ( n10017 & n24409 ) ;
  assign n24411 = n8107 ^ n6561 ^ n2527 ;
  assign n24412 = ( n8504 & n13425 ) | ( n8504 & n24411 ) | ( n13425 & n24411 ) ;
  assign n24413 = n24412 ^ n6582 ^ n3374 ;
  assign n24414 = ~n1363 & n24413 ;
  assign n24415 = n24414 ^ n7242 ^ 1'b0 ;
  assign n24416 = n14101 ^ n9881 ^ n6533 ;
  assign n24417 = ( n3591 & ~n4265 ) | ( n3591 & n4487 ) | ( ~n4265 & n4487 ) ;
  assign n24418 = n4267 & n24417 ;
  assign n24419 = ( n24415 & n24416 ) | ( n24415 & n24418 ) | ( n24416 & n24418 ) ;
  assign n24432 = n9668 | n21596 ;
  assign n24433 = n19465 | n24432 ;
  assign n24420 = n6097 ^ n4815 ^ n1844 ;
  assign n24421 = n24420 ^ n3643 ^ 1'b0 ;
  assign n24422 = n7168 & ~n24421 ;
  assign n24428 = n7661 ^ n4554 ^ n2333 ;
  assign n24423 = n17232 ^ n16240 ^ n3181 ;
  assign n24424 = n1237 & n8687 ;
  assign n24425 = n24424 ^ n10574 ^ 1'b0 ;
  assign n24426 = n2022 | n24425 ;
  assign n24427 = ( n7852 & n24423 ) | ( n7852 & n24426 ) | ( n24423 & n24426 ) ;
  assign n24429 = n24428 ^ n24427 ^ n16671 ;
  assign n24430 = n15911 | n24429 ;
  assign n24431 = n24422 | n24430 ;
  assign n24434 = n24433 ^ n24431 ^ n5901 ;
  assign n24435 = n11241 ^ n8058 ^ n3037 ;
  assign n24436 = n24435 ^ n1061 ^ 1'b0 ;
  assign n24437 = n24386 ^ n1032 ^ 1'b0 ;
  assign n24438 = n14239 & ~n24437 ;
  assign n24440 = ( n7965 & n12235 ) | ( n7965 & n13815 ) | ( n12235 & n13815 ) ;
  assign n24439 = n8822 & ~n18346 ;
  assign n24441 = n24440 ^ n24439 ^ 1'b0 ;
  assign n24442 = ( n9829 & ~n14649 ) | ( n9829 & n18687 ) | ( ~n14649 & n18687 ) ;
  assign n24443 = n12746 ^ n10752 ^ n1001 ;
  assign n24444 = n17334 & ~n24443 ;
  assign n24445 = ( n383 & ~n24442 ) | ( n383 & n24444 ) | ( ~n24442 & n24444 ) ;
  assign n24446 = n4801 & n11313 ;
  assign n24447 = n24446 ^ n7620 ^ 1'b0 ;
  assign n24448 = n24265 ^ n8877 ^ 1'b0 ;
  assign n24449 = ( n15999 & ~n24447 ) | ( n15999 & n24448 ) | ( ~n24447 & n24448 ) ;
  assign n24450 = ( n3012 & n8592 ) | ( n3012 & ~n9879 ) | ( n8592 & ~n9879 ) ;
  assign n24451 = n21223 ^ n15212 ^ n4873 ;
  assign n24452 = n24451 ^ n13585 ^ n12242 ;
  assign n24453 = ~n21606 & n24452 ;
  assign n24454 = n19786 & n24026 ;
  assign n24455 = n24454 ^ n7635 ^ 1'b0 ;
  assign n24456 = ( n9436 & ~n19660 ) | ( n9436 & n22811 ) | ( ~n19660 & n22811 ) ;
  assign n24457 = n24456 ^ n4035 ^ n1652 ;
  assign n24458 = ( n2427 & ~n7566 ) | ( n2427 & n18257 ) | ( ~n7566 & n18257 ) ;
  assign n24459 = n17335 ^ n9334 ^ 1'b0 ;
  assign n24460 = n24458 & n24459 ;
  assign n24461 = n24460 ^ n8730 ^ 1'b0 ;
  assign n24462 = ( n5261 & ~n11159 ) | ( n5261 & n24461 ) | ( ~n11159 & n24461 ) ;
  assign n24463 = ( n745 & n3196 ) | ( n745 & ~n7069 ) | ( n3196 & ~n7069 ) ;
  assign n24464 = n4182 & n24463 ;
  assign n24465 = n24464 ^ n20403 ^ 1'b0 ;
  assign n24466 = n16928 ^ n13066 ^ 1'b0 ;
  assign n24467 = n5504 | n24466 ;
  assign n24468 = n24467 ^ n372 ^ 1'b0 ;
  assign n24469 = n12743 & n24468 ;
  assign n24470 = n13381 & n14304 ;
  assign n24471 = n21991 ^ n16069 ^ n12953 ;
  assign n24472 = n8047 ^ n3907 ^ 1'b0 ;
  assign n24473 = n17293 ^ n5256 ^ n3120 ;
  assign n24478 = n18384 ^ n14038 ^ 1'b0 ;
  assign n24479 = ~n7060 & n24478 ;
  assign n24474 = n11653 ^ n10981 ^ n5197 ;
  assign n24475 = n15836 & ~n24474 ;
  assign n24476 = n24475 ^ n9716 ^ n6680 ;
  assign n24477 = n16227 & n24476 ;
  assign n24480 = n24479 ^ n24477 ^ n9639 ;
  assign n24481 = n15606 ^ n14727 ^ n13385 ;
  assign n24482 = n21970 ^ n8670 ^ 1'b0 ;
  assign n24483 = n7517 ^ n5709 ^ 1'b0 ;
  assign n24484 = ( n6478 & ~n6632 ) | ( n6478 & n10509 ) | ( ~n6632 & n10509 ) ;
  assign n24485 = n6555 ^ n4885 ^ n2899 ;
  assign n24486 = n24485 ^ n8096 ^ n1016 ;
  assign n24487 = n24486 ^ n16894 ^ n9345 ;
  assign n24488 = ( n9684 & n11704 ) | ( n9684 & n24487 ) | ( n11704 & n24487 ) ;
  assign n24489 = ( n24483 & ~n24484 ) | ( n24483 & n24488 ) | ( ~n24484 & n24488 ) ;
  assign n24490 = n9965 ^ n6378 ^ n3876 ;
  assign n24491 = n11126 ^ n5024 ^ 1'b0 ;
  assign n24492 = n24490 & ~n24491 ;
  assign n24493 = n24492 ^ n13930 ^ 1'b0 ;
  assign n24494 = n24493 ^ n17534 ^ 1'b0 ;
  assign n24495 = n20564 ^ n16134 ^ n10083 ;
  assign n24499 = n4935 ^ x61 ^ 1'b0 ;
  assign n24500 = n4971 & ~n24499 ;
  assign n24496 = n22138 ^ n21224 ^ 1'b0 ;
  assign n24497 = n1988 & n24496 ;
  assign n24498 = ~n10902 & n24497 ;
  assign n24501 = n24500 ^ n24498 ^ 1'b0 ;
  assign n24502 = n18439 ^ n16242 ^ 1'b0 ;
  assign n24503 = n9649 & ~n24502 ;
  assign n24504 = ~n10739 & n24503 ;
  assign n24505 = ( ~n1206 & n3234 ) | ( ~n1206 & n13279 ) | ( n3234 & n13279 ) ;
  assign n24506 = n24505 ^ n3870 ^ 1'b0 ;
  assign n24507 = n6103 | n24506 ;
  assign n24508 = n24507 ^ n16834 ^ n1200 ;
  assign n24509 = ( n8745 & ~n12992 ) | ( n8745 & n24508 ) | ( ~n12992 & n24508 ) ;
  assign n24510 = ( n5880 & n13105 ) | ( n5880 & ~n24509 ) | ( n13105 & ~n24509 ) ;
  assign n24511 = ( n5714 & n9929 ) | ( n5714 & n14677 ) | ( n9929 & n14677 ) ;
  assign n24512 = ( n1181 & ~n16066 ) | ( n1181 & n24511 ) | ( ~n16066 & n24511 ) ;
  assign n24513 = n20809 ^ n4873 ^ 1'b0 ;
  assign n24514 = ( n9944 & n22154 ) | ( n9944 & ~n24513 ) | ( n22154 & ~n24513 ) ;
  assign n24515 = n13078 | n14355 ;
  assign n24516 = n24514 & ~n24515 ;
  assign n24517 = n24516 ^ n5790 ^ n2139 ;
  assign n24518 = n834 & ~n5359 ;
  assign n24519 = ( ~n5717 & n16998 ) | ( ~n5717 & n24518 ) | ( n16998 & n24518 ) ;
  assign n24520 = n6220 & n9180 ;
  assign n24521 = ( n1502 & n3101 ) | ( n1502 & n24520 ) | ( n3101 & n24520 ) ;
  assign n24522 = n18558 ^ n14543 ^ 1'b0 ;
  assign n24523 = n24521 | n24522 ;
  assign n24524 = n3037 ^ n2105 ^ n948 ;
  assign n24525 = n24524 ^ n1562 ^ n1067 ;
  assign n24526 = n9438 & n24525 ;
  assign n24527 = n24523 | n24526 ;
  assign n24528 = n22137 | n24527 ;
  assign n24529 = n24519 & n24528 ;
  assign n24530 = n6111 ^ x136 ^ 1'b0 ;
  assign n24531 = n4450 & ~n7723 ;
  assign n24532 = ( ~n5350 & n24530 ) | ( ~n5350 & n24531 ) | ( n24530 & n24531 ) ;
  assign n24533 = n2437 & n20728 ;
  assign n24534 = n5157 & n24533 ;
  assign n24537 = ( ~n5598 & n13516 ) | ( ~n5598 & n24387 ) | ( n13516 & n24387 ) ;
  assign n24536 = ( n11259 & n13738 ) | ( n11259 & ~n19935 ) | ( n13738 & ~n19935 ) ;
  assign n24535 = n13757 ^ n4042 ^ 1'b0 ;
  assign n24538 = n24537 ^ n24536 ^ n24535 ;
  assign n24539 = n22756 ^ n8324 ^ n6558 ;
  assign n24540 = n655 & n2499 ;
  assign n24541 = n1095 & n24540 ;
  assign n24542 = n24541 ^ n17386 ^ n3763 ;
  assign n24543 = ( n1504 & n5917 ) | ( n1504 & ~n7827 ) | ( n5917 & ~n7827 ) ;
  assign n24544 = n24543 ^ n11914 ^ 1'b0 ;
  assign n24545 = ( ~n23574 & n24542 ) | ( ~n23574 & n24544 ) | ( n24542 & n24544 ) ;
  assign n24546 = ( ~n5212 & n6940 ) | ( ~n5212 & n20908 ) | ( n6940 & n20908 ) ;
  assign n24547 = ~n3257 & n5419 ;
  assign n24548 = ~n24546 & n24547 ;
  assign n24549 = n20169 ^ x193 ^ 1'b0 ;
  assign n24550 = n7758 & ~n24549 ;
  assign n24551 = n24550 ^ n21812 ^ 1'b0 ;
  assign n24552 = ~n24548 & n24551 ;
  assign n24553 = n24552 ^ n20751 ^ 1'b0 ;
  assign n24554 = n21767 ^ n14100 ^ n6901 ;
  assign n24555 = n24554 ^ n19736 ^ n14341 ;
  assign n24556 = ( n11879 & n16210 ) | ( n11879 & ~n24555 ) | ( n16210 & ~n24555 ) ;
  assign n24557 = ( ~n14410 & n20300 ) | ( ~n14410 & n24556 ) | ( n20300 & n24556 ) ;
  assign n24558 = n17686 ^ n2501 ^ 1'b0 ;
  assign n24559 = n21350 & ~n24558 ;
  assign n24560 = ( n6267 & ~n9475 ) | ( n6267 & n10007 ) | ( ~n9475 & n10007 ) ;
  assign n24561 = n24560 ^ n5444 ^ 1'b0 ;
  assign n24562 = n4248 & ~n24561 ;
  assign n24563 = n14537 ^ n3171 ^ n883 ;
  assign n24564 = ~n20233 & n24563 ;
  assign n24565 = ~n24562 & n24564 ;
  assign n24566 = n24559 & n24565 ;
  assign n24567 = n17658 & ~n21188 ;
  assign n24568 = n1500 & n24567 ;
  assign n24569 = n10321 ^ n4467 ^ n4466 ;
  assign n24570 = n24569 ^ n17738 ^ 1'b0 ;
  assign n24574 = ( ~n3814 & n5933 ) | ( ~n3814 & n8977 ) | ( n5933 & n8977 ) ;
  assign n24575 = ~n8231 & n13066 ;
  assign n24576 = ( n9641 & n24574 ) | ( n9641 & n24575 ) | ( n24574 & n24575 ) ;
  assign n24572 = n6204 ^ n5088 ^ n1456 ;
  assign n24571 = ( ~n2332 & n3767 ) | ( ~n2332 & n24030 ) | ( n3767 & n24030 ) ;
  assign n24573 = n24572 ^ n24571 ^ n3980 ;
  assign n24577 = n24576 ^ n24573 ^ n418 ;
  assign n24578 = n21252 ^ n17056 ^ n15421 ;
  assign n24579 = ( n14541 & n14960 ) | ( n14541 & n24578 ) | ( n14960 & n24578 ) ;
  assign n24586 = ~n5796 & n17254 ;
  assign n24587 = n24586 ^ n9243 ^ 1'b0 ;
  assign n24588 = ~n17244 & n24587 ;
  assign n24589 = n24588 ^ n11737 ^ 1'b0 ;
  assign n24580 = ~n9145 & n13536 ;
  assign n24581 = ~n3251 & n24580 ;
  assign n24582 = ( n2481 & n15567 ) | ( n2481 & ~n24581 ) | ( n15567 & ~n24581 ) ;
  assign n24583 = n16400 ^ n5327 ^ 1'b0 ;
  assign n24584 = n24582 & n24583 ;
  assign n24585 = ( ~n22506 & n22519 ) | ( ~n22506 & n24584 ) | ( n22519 & n24584 ) ;
  assign n24590 = n24589 ^ n24585 ^ n17509 ;
  assign n24591 = ( ~n2365 & n10577 ) | ( ~n2365 & n18916 ) | ( n10577 & n18916 ) ;
  assign n24592 = n4982 ^ n3651 ^ n713 ;
  assign n24593 = n3164 | n24592 ;
  assign n24594 = ( n1714 & ~n2216 ) | ( n1714 & n8635 ) | ( ~n2216 & n8635 ) ;
  assign n24595 = ~n12292 & n24594 ;
  assign n24596 = n15719 & ~n24595 ;
  assign n24597 = ( n3643 & ~n24593 ) | ( n3643 & n24596 ) | ( ~n24593 & n24596 ) ;
  assign n24598 = n24597 ^ n11479 ^ x178 ;
  assign n24599 = n8311 | n14773 ;
  assign n24600 = ( n5107 & n8570 ) | ( n5107 & n24599 ) | ( n8570 & n24599 ) ;
  assign n24601 = n24600 ^ n12156 ^ 1'b0 ;
  assign n24602 = n8431 & n24601 ;
  assign n24603 = n8493 ^ n7216 ^ 1'b0 ;
  assign n24604 = n2804 & n24603 ;
  assign n24605 = ~n4638 & n24604 ;
  assign n24606 = n24605 ^ n21491 ^ 1'b0 ;
  assign n24607 = ~n3312 & n24606 ;
  assign n24608 = n5819 ^ n5553 ^ 1'b0 ;
  assign n24609 = ( n4239 & n18409 ) | ( n4239 & ~n24608 ) | ( n18409 & ~n24608 ) ;
  assign n24611 = ( n3659 & n5428 ) | ( n3659 & n6901 ) | ( n5428 & n6901 ) ;
  assign n24610 = n7080 | n23584 ;
  assign n24612 = n24611 ^ n24610 ^ 1'b0 ;
  assign n24613 = ( n7296 & n7764 ) | ( n7296 & n17349 ) | ( n7764 & n17349 ) ;
  assign n24614 = ~n6065 & n24613 ;
  assign n24615 = ( n5877 & ~n9624 ) | ( n5877 & n19772 ) | ( ~n9624 & n19772 ) ;
  assign n24616 = n24615 ^ n17121 ^ n16612 ;
  assign n24617 = ~n8988 & n9641 ;
  assign n24618 = ~n7204 & n24617 ;
  assign n24619 = ( ~n6420 & n7859 ) | ( ~n6420 & n11673 ) | ( n7859 & n11673 ) ;
  assign n24620 = n17662 & ~n24619 ;
  assign n24621 = ( n17419 & n20064 ) | ( n17419 & ~n24620 ) | ( n20064 & ~n24620 ) ;
  assign n24622 = ~n24618 & n24621 ;
  assign n24623 = n24622 ^ n16624 ^ 1'b0 ;
  assign n24624 = n15321 ^ n6155 ^ 1'b0 ;
  assign n24627 = n21388 ^ n18308 ^ n15821 ;
  assign n24625 = n6091 | n8904 ;
  assign n24626 = n24625 ^ n10334 ^ 1'b0 ;
  assign n24628 = n24627 ^ n24626 ^ 1'b0 ;
  assign n24629 = ( ~n7375 & n24624 ) | ( ~n7375 & n24628 ) | ( n24624 & n24628 ) ;
  assign n24630 = ( n865 & n12453 ) | ( n865 & n15408 ) | ( n12453 & n15408 ) ;
  assign n24631 = ( ~n3506 & n8984 ) | ( ~n3506 & n11951 ) | ( n8984 & n11951 ) ;
  assign n24632 = n24026 ^ n13381 ^ n9993 ;
  assign n24633 = ( n14943 & n24631 ) | ( n14943 & n24632 ) | ( n24631 & n24632 ) ;
  assign n24634 = n24633 ^ n5253 ^ n3661 ;
  assign n24635 = n12454 ^ n3671 ^ 1'b0 ;
  assign n24636 = n983 & ~n24635 ;
  assign n24637 = n24636 ^ n1169 ^ 1'b0 ;
  assign n24638 = n24637 ^ n14568 ^ n8351 ;
  assign n24641 = n12007 ^ n2053 ^ 1'b0 ;
  assign n24642 = n24641 ^ n24156 ^ 1'b0 ;
  assign n24639 = n18768 ^ n571 ^ 1'b0 ;
  assign n24640 = n21699 | n24639 ;
  assign n24643 = n24642 ^ n24640 ^ n3645 ;
  assign n24646 = n9317 ^ n5838 ^ n3853 ;
  assign n24647 = ( n2851 & ~n5887 ) | ( n2851 & n24646 ) | ( ~n5887 & n24646 ) ;
  assign n24644 = ~n12037 & n14838 ;
  assign n24645 = n10538 & ~n24644 ;
  assign n24648 = n24647 ^ n24645 ^ 1'b0 ;
  assign n24649 = n24643 & ~n24648 ;
  assign n24650 = n24649 ^ n11772 ^ 1'b0 ;
  assign n24651 = ( ~n23053 & n24638 ) | ( ~n23053 & n24650 ) | ( n24638 & n24650 ) ;
  assign n24652 = ( n2865 & n4081 ) | ( n2865 & n5888 ) | ( n4081 & n5888 ) ;
  assign n24653 = n24652 ^ n14929 ^ n11255 ;
  assign n24654 = n24653 ^ n20035 ^ n9706 ;
  assign n24655 = n9602 ^ n6802 ^ n5382 ;
  assign n24656 = n21365 & n24655 ;
  assign n24657 = n11042 & n24656 ;
  assign n24658 = n24657 ^ n9033 ^ 1'b0 ;
  assign n24659 = n1717 & n5939 ;
  assign n24660 = n12743 & ~n24659 ;
  assign n24661 = n24660 ^ n14779 ^ 1'b0 ;
  assign n24662 = n24661 ^ n24548 ^ n8804 ;
  assign n24663 = ( n3757 & n3872 ) | ( n3757 & n24662 ) | ( n3872 & n24662 ) ;
  assign n24664 = ( n8387 & n9910 ) | ( n8387 & ~n18427 ) | ( n9910 & ~n18427 ) ;
  assign n24665 = n7135 ^ n861 ^ n558 ;
  assign n24666 = n24665 ^ n19550 ^ n6817 ;
  assign n24667 = n3459 & ~n24666 ;
  assign n24668 = ~n12340 & n24667 ;
  assign n24669 = ( ~n10808 & n24664 ) | ( ~n10808 & n24668 ) | ( n24664 & n24668 ) ;
  assign n24670 = n10298 ^ n7920 ^ 1'b0 ;
  assign n24671 = n24670 ^ n13364 ^ n3765 ;
  assign n24672 = ( x138 & n3715 ) | ( x138 & ~n15778 ) | ( n3715 & ~n15778 ) ;
  assign n24673 = n24671 & ~n24672 ;
  assign n24674 = ~n22886 & n24673 ;
  assign n24675 = n12528 ^ n10930 ^ 1'b0 ;
  assign n24676 = n24675 ^ n16073 ^ 1'b0 ;
  assign n24677 = n10498 | n24676 ;
  assign n24678 = n9846 ^ n1935 ^ 1'b0 ;
  assign n24679 = ( n18289 & ~n23006 ) | ( n18289 & n24678 ) | ( ~n23006 & n24678 ) ;
  assign n24681 = ~n3228 & n3405 ;
  assign n24682 = n24681 ^ n7209 ^ 1'b0 ;
  assign n24680 = n6326 & n8566 ;
  assign n24683 = n24682 ^ n24680 ^ n23521 ;
  assign n24687 = n7134 ^ n6887 ^ 1'b0 ;
  assign n24685 = n15599 ^ n14900 ^ n12917 ;
  assign n24684 = n7663 ^ n5829 ^ n2243 ;
  assign n24686 = n24685 ^ n24684 ^ n2472 ;
  assign n24688 = n24687 ^ n24686 ^ n11826 ;
  assign n24689 = n797 | n17813 ;
  assign n24690 = ( n10446 & ~n11729 ) | ( n10446 & n21483 ) | ( ~n11729 & n21483 ) ;
  assign n24691 = n23134 ^ n5523 ^ n4277 ;
  assign n24692 = n24691 ^ n8660 ^ 1'b0 ;
  assign n24693 = ( ~n12216 & n19226 ) | ( ~n12216 & n24692 ) | ( n19226 & n24692 ) ;
  assign n24694 = ( n4534 & ~n20467 ) | ( n4534 & n24693 ) | ( ~n20467 & n24693 ) ;
  assign n24695 = n24694 ^ n24348 ^ n19106 ;
  assign n24696 = x176 & n11784 ;
  assign n24698 = n8158 ^ n4705 ^ n2390 ;
  assign n24697 = ~n5956 & n8046 ;
  assign n24699 = n24698 ^ n24697 ^ n345 ;
  assign n24700 = ~n371 & n15232 ;
  assign n24701 = n21869 ^ n13556 ^ n7905 ;
  assign n24702 = n24701 ^ n16024 ^ 1'b0 ;
  assign n24703 = n19281 ^ n10852 ^ n9344 ;
  assign n24704 = ~n16154 & n24703 ;
  assign n24705 = ~n15724 & n24704 ;
  assign n24706 = n24702 & ~n24705 ;
  assign n24707 = n2311 & n24706 ;
  assign n24708 = ~n11241 & n15451 ;
  assign n24709 = n24707 & n24708 ;
  assign n24710 = ( ~n24699 & n24700 ) | ( ~n24699 & n24709 ) | ( n24700 & n24709 ) ;
  assign n24711 = n18489 ^ n12617 ^ n2756 ;
  assign n24712 = n24711 ^ n18536 ^ 1'b0 ;
  assign n24713 = n6582 & n24712 ;
  assign n24714 = n15498 ^ n2197 ^ n1404 ;
  assign n24715 = n23157 ^ n8495 ^ 1'b0 ;
  assign n24716 = n10590 & n24715 ;
  assign n24717 = n8842 & ~n9452 ;
  assign n24718 = n24717 ^ n7984 ^ 1'b0 ;
  assign n24719 = n14752 | n24718 ;
  assign n24720 = n24716 & n24719 ;
  assign n24721 = ( n1242 & ~n13932 ) | ( n1242 & n23664 ) | ( ~n13932 & n23664 ) ;
  assign n24724 = n6333 ^ n5033 ^ n2397 ;
  assign n24725 = n16791 & ~n24724 ;
  assign n24722 = n6386 ^ n2031 ^ 1'b0 ;
  assign n24723 = ( ~n7104 & n18185 ) | ( ~n7104 & n24722 ) | ( n18185 & n24722 ) ;
  assign n24726 = n24725 ^ n24723 ^ 1'b0 ;
  assign n24727 = n3181 & n24726 ;
  assign n24728 = n24452 ^ n8710 ^ 1'b0 ;
  assign n24729 = n21220 & n24728 ;
  assign n24730 = n9331 ^ n1526 ^ 1'b0 ;
  assign n24731 = n6428 | n24730 ;
  assign n24732 = n24731 ^ n9963 ^ n3254 ;
  assign n24733 = n5952 ^ n3279 ^ 1'b0 ;
  assign n24734 = n24733 ^ n11961 ^ 1'b0 ;
  assign n24735 = n6610 ^ n4138 ^ 1'b0 ;
  assign n24736 = n1210 | n24735 ;
  assign n24737 = n24736 ^ n9483 ^ n1575 ;
  assign n24738 = n19574 | n24737 ;
  assign n24739 = n20756 | n24738 ;
  assign n24740 = ( n1773 & ~n5566 ) | ( n1773 & n13220 ) | ( ~n5566 & n13220 ) ;
  assign n24741 = n10476 ^ n1936 ^ n484 ;
  assign n24742 = n24741 ^ n16254 ^ 1'b0 ;
  assign n24743 = n7673 | n24742 ;
  assign n24744 = ( n6375 & ~n24740 ) | ( n6375 & n24743 ) | ( ~n24740 & n24743 ) ;
  assign n24745 = n18439 ^ n7871 ^ 1'b0 ;
  assign n24746 = ~n786 & n24745 ;
  assign n24747 = n24746 ^ n16251 ^ n482 ;
  assign n24748 = ( n10314 & n22036 ) | ( n10314 & n24747 ) | ( n22036 & n24747 ) ;
  assign n24749 = ( ~n22418 & n24744 ) | ( ~n22418 & n24748 ) | ( n24744 & n24748 ) ;
  assign n24750 = ( n8067 & n18633 ) | ( n8067 & n20368 ) | ( n18633 & n20368 ) ;
  assign n24751 = n20856 ^ n9640 ^ n5690 ;
  assign n24752 = n24751 ^ n5296 ^ n4584 ;
  assign n24753 = n24752 ^ n18584 ^ 1'b0 ;
  assign n24754 = n2232 & n7020 ;
  assign n24755 = ~n24322 & n24754 ;
  assign n24756 = n16339 ^ n10389 ^ 1'b0 ;
  assign n24757 = n24756 ^ n13950 ^ n1093 ;
  assign n24764 = n20807 ^ n10787 ^ n9003 ;
  assign n24765 = ( ~n7727 & n14274 ) | ( ~n7727 & n24764 ) | ( n14274 & n24764 ) ;
  assign n24758 = n10318 ^ n1400 ^ x109 ;
  assign n24759 = n3009 ^ n2978 ^ 1'b0 ;
  assign n24760 = n8311 | n24759 ;
  assign n24761 = n10294 & n23726 ;
  assign n24762 = ( n24758 & n24760 ) | ( n24758 & n24761 ) | ( n24760 & n24761 ) ;
  assign n24763 = ( n7884 & n23465 ) | ( n7884 & n24762 ) | ( n23465 & n24762 ) ;
  assign n24766 = n24765 ^ n24763 ^ n5660 ;
  assign n24767 = ~n8390 & n10227 ;
  assign n24768 = ~n10444 & n24767 ;
  assign n24769 = n24768 ^ n7384 ^ n1675 ;
  assign n24770 = ( n945 & n9287 ) | ( n945 & n10974 ) | ( n9287 & n10974 ) ;
  assign n24771 = n24770 ^ n16373 ^ 1'b0 ;
  assign n24772 = ( ~n15310 & n24769 ) | ( ~n15310 & n24771 ) | ( n24769 & n24771 ) ;
  assign n24773 = n18455 & n24772 ;
  assign n24774 = n2545 ^ n931 ^ n599 ;
  assign n24775 = n24774 ^ n23802 ^ n16091 ;
  assign n24776 = ( n16930 & ~n19217 ) | ( n16930 & n19923 ) | ( ~n19217 & n19923 ) ;
  assign n24777 = ( n1167 & n9248 ) | ( n1167 & ~n11591 ) | ( n9248 & ~n11591 ) ;
  assign n24778 = ( n9103 & n10531 ) | ( n9103 & n24777 ) | ( n10531 & n24777 ) ;
  assign n24779 = n19842 ^ n14632 ^ n5648 ;
  assign n24780 = n2635 & n24779 ;
  assign n24781 = n24780 ^ n20878 ^ 1'b0 ;
  assign n24782 = ~n24509 & n24781 ;
  assign n24783 = n24486 & n24782 ;
  assign n24784 = n17133 & n17939 ;
  assign n24785 = n14255 ^ n12227 ^ n5689 ;
  assign n24786 = n8419 ^ n3006 ^ n1676 ;
  assign n24787 = n17279 ^ n9866 ^ n4152 ;
  assign n24788 = ( n677 & ~n8128 ) | ( n677 & n24787 ) | ( ~n8128 & n24787 ) ;
  assign n24789 = n9861 & ~n10124 ;
  assign n24790 = ~n20532 & n24789 ;
  assign n24791 = n5923 | n9625 ;
  assign n24792 = n24791 ^ n14749 ^ 1'b0 ;
  assign n24793 = n24792 ^ n17833 ^ n14795 ;
  assign n24794 = ( ~n4046 & n7222 ) | ( ~n4046 & n13407 ) | ( n7222 & n13407 ) ;
  assign n24795 = n14313 ^ n12776 ^ 1'b0 ;
  assign n24796 = n16769 & n24795 ;
  assign n24797 = ( n1433 & n24794 ) | ( n1433 & n24796 ) | ( n24794 & n24796 ) ;
  assign n24798 = n925 & n21839 ;
  assign n24799 = n24798 ^ n3448 ^ 1'b0 ;
  assign n24800 = n24799 ^ n7645 ^ n7644 ;
  assign n24801 = n4776 & n11982 ;
  assign n24802 = n7910 & n24801 ;
  assign n24803 = n11273 | n24802 ;
  assign n24804 = n24803 ^ n7605 ^ 1'b0 ;
  assign n24805 = n15947 ^ n3094 ^ 1'b0 ;
  assign n24816 = n22745 ^ n12432 ^ x174 ;
  assign n24815 = n7862 ^ n7188 ^ 1'b0 ;
  assign n24812 = ~n10935 & n12794 ;
  assign n24813 = n24812 ^ n15145 ^ 1'b0 ;
  assign n24807 = n10371 ^ n4529 ^ n2861 ;
  assign n24806 = ( ~n1963 & n8143 ) | ( ~n1963 & n10080 ) | ( n8143 & n10080 ) ;
  assign n24808 = n24807 ^ n24806 ^ n10217 ;
  assign n24809 = n24808 ^ n20698 ^ n3931 ;
  assign n24810 = n556 & ~n24809 ;
  assign n24811 = ~n9854 & n24810 ;
  assign n24814 = n24813 ^ n24811 ^ n5538 ;
  assign n24817 = n24816 ^ n24815 ^ n24814 ;
  assign n24818 = n12276 | n18578 ;
  assign n24819 = ( n11227 & n24560 ) | ( n11227 & ~n24818 ) | ( n24560 & ~n24818 ) ;
  assign n24820 = n15560 ^ n14550 ^ n6037 ;
  assign n24825 = ( n2728 & n11784 ) | ( n2728 & ~n12337 ) | ( n11784 & ~n12337 ) ;
  assign n24821 = n20675 ^ n17001 ^ 1'b0 ;
  assign n24822 = n12420 ^ n6755 ^ n291 ;
  assign n24823 = ( n11210 & n24821 ) | ( n11210 & n24822 ) | ( n24821 & n24822 ) ;
  assign n24824 = n9346 | n24823 ;
  assign n24826 = n24825 ^ n24824 ^ 1'b0 ;
  assign n24827 = ( n6713 & n12954 ) | ( n6713 & ~n13265 ) | ( n12954 & ~n13265 ) ;
  assign n24828 = n4333 ^ n1464 ^ 1'b0 ;
  assign n24829 = ~n5703 & n24828 ;
  assign n24830 = n24829 ^ n11339 ^ n2266 ;
  assign n24831 = n24827 & ~n24830 ;
  assign n24832 = ( n470 & n11781 ) | ( n470 & n22401 ) | ( n11781 & n22401 ) ;
  assign n24833 = ( n16060 & ~n20202 ) | ( n16060 & n24832 ) | ( ~n20202 & n24832 ) ;
  assign n24834 = n1108 & n4995 ;
  assign n24835 = ( n1078 & ~n4303 ) | ( n1078 & n17958 ) | ( ~n4303 & n17958 ) ;
  assign n24836 = n11209 ^ n9249 ^ n7022 ;
  assign n24837 = n24836 ^ n15261 ^ n5704 ;
  assign n24838 = n8736 & ~n16455 ;
  assign n24839 = ~n1048 & n24838 ;
  assign n24840 = ( n4329 & n7038 ) | ( n4329 & ~n8938 ) | ( n7038 & ~n8938 ) ;
  assign n24841 = n24840 ^ n18244 ^ n8947 ;
  assign n24842 = ~n24839 & n24841 ;
  assign n24843 = n24842 ^ n509 ^ 1'b0 ;
  assign n24844 = ( ~n13634 & n22276 ) | ( ~n13634 & n23435 ) | ( n22276 & n23435 ) ;
  assign n24845 = n24844 ^ n14448 ^ n6085 ;
  assign n24846 = n24845 ^ n21277 ^ 1'b0 ;
  assign n24847 = ( x82 & ~n14662 ) | ( x82 & n15155 ) | ( ~n14662 & n15155 ) ;
  assign n24848 = ( ~n10277 & n12437 ) | ( ~n10277 & n24847 ) | ( n12437 & n24847 ) ;
  assign n24849 = n24848 ^ n24063 ^ 1'b0 ;
  assign n24850 = n21888 ^ n14184 ^ n6480 ;
  assign n24851 = n21229 | n24850 ;
  assign n24852 = n24851 ^ n11208 ^ 1'b0 ;
  assign n24853 = n24852 ^ n15847 ^ n2948 ;
  assign n24857 = n14087 ^ n13027 ^ n10856 ;
  assign n24858 = n24857 ^ n21723 ^ 1'b0 ;
  assign n24859 = n8079 | n24858 ;
  assign n24854 = n12047 ^ n9959 ^ n8422 ;
  assign n24855 = n12491 | n18281 ;
  assign n24856 = n24854 & ~n24855 ;
  assign n24860 = n24859 ^ n24856 ^ 1'b0 ;
  assign n24861 = x70 & n10410 ;
  assign n24862 = n3051 & n24861 ;
  assign n24863 = n24862 ^ n11271 ^ n7437 ;
  assign n24864 = ( n3925 & n4126 ) | ( n3925 & ~n5501 ) | ( n4126 & ~n5501 ) ;
  assign n24865 = ~n5894 & n24864 ;
  assign n24866 = n24863 & n24865 ;
  assign n24867 = n14330 ^ n9660 ^ 1'b0 ;
  assign n24868 = n6028 | n24867 ;
  assign n24869 = n18540 ^ n3995 ^ 1'b0 ;
  assign n24870 = ( ~n4128 & n13944 ) | ( ~n4128 & n20105 ) | ( n13944 & n20105 ) ;
  assign n24871 = ( n2139 & n3221 ) | ( n2139 & n7483 ) | ( n3221 & n7483 ) ;
  assign n24872 = ( n418 & ~n7351 ) | ( n418 & n7377 ) | ( ~n7351 & n7377 ) ;
  assign n24873 = ( n14386 & n24871 ) | ( n14386 & ~n24872 ) | ( n24871 & ~n24872 ) ;
  assign n24874 = n23286 ^ n8089 ^ 1'b0 ;
  assign n24875 = ~n24873 & n24874 ;
  assign n24876 = ( n8034 & ~n8846 ) | ( n8034 & n21992 ) | ( ~n8846 & n21992 ) ;
  assign n24877 = ( ~n5343 & n6170 ) | ( ~n5343 & n24876 ) | ( n6170 & n24876 ) ;
  assign n24878 = n24877 ^ n11340 ^ 1'b0 ;
  assign n24884 = ( n13417 & n17542 ) | ( n13417 & ~n19119 ) | ( n17542 & ~n19119 ) ;
  assign n24883 = ~n649 & n1198 ;
  assign n24885 = n24884 ^ n24883 ^ 1'b0 ;
  assign n24879 = n938 & n2492 ;
  assign n24880 = n3619 ^ n3019 ^ n2425 ;
  assign n24881 = n5224 ^ n3956 ^ 1'b0 ;
  assign n24882 = ( n24879 & n24880 ) | ( n24879 & ~n24881 ) | ( n24880 & ~n24881 ) ;
  assign n24886 = n24885 ^ n24882 ^ n22164 ;
  assign n24887 = n20061 & n22931 ;
  assign n24888 = n1733 & n24887 ;
  assign n24889 = ( n4631 & ~n12708 ) | ( n4631 & n22507 ) | ( ~n12708 & n22507 ) ;
  assign n24890 = n24889 ^ n18269 ^ n3127 ;
  assign n24898 = n13523 ^ n13338 ^ n7526 ;
  assign n24893 = ~n2348 & n21101 ;
  assign n24894 = ~n2045 & n24893 ;
  assign n24892 = n22819 ^ n5018 ^ 1'b0 ;
  assign n24895 = n24894 ^ n24892 ^ n2753 ;
  assign n24891 = n6025 ^ n1577 ^ 1'b0 ;
  assign n24896 = n24895 ^ n24891 ^ 1'b0 ;
  assign n24897 = n2140 & n24896 ;
  assign n24899 = n24898 ^ n24897 ^ n18740 ;
  assign n24900 = ( ~n11756 & n18240 ) | ( ~n11756 & n21083 ) | ( n18240 & n21083 ) ;
  assign n24901 = n6732 ^ n3462 ^ n2659 ;
  assign n24902 = n13191 ^ n9102 ^ n2406 ;
  assign n24903 = n13719 ^ n2711 ^ n2403 ;
  assign n24904 = ~n17563 & n24903 ;
  assign n24905 = ~n3644 & n24904 ;
  assign n24906 = ~n5366 & n20107 ;
  assign n24907 = ~n5328 & n8201 ;
  assign n24908 = ~n18625 & n24907 ;
  assign n24909 = n24908 ^ n21274 ^ 1'b0 ;
  assign n24914 = n4163 | n18114 ;
  assign n24915 = n24914 ^ n3035 ^ 1'b0 ;
  assign n24910 = ( n1359 & n20902 ) | ( n1359 & ~n21248 ) | ( n20902 & ~n21248 ) ;
  assign n24911 = n15962 ^ x232 ^ 1'b0 ;
  assign n24912 = n8229 & ~n24911 ;
  assign n24913 = ( n21952 & n24910 ) | ( n21952 & n24912 ) | ( n24910 & n24912 ) ;
  assign n24916 = n24915 ^ n24913 ^ n6175 ;
  assign n24917 = n24916 ^ n20552 ^ n11418 ;
  assign n24918 = ( n4444 & n10363 ) | ( n4444 & ~n15935 ) | ( n10363 & ~n15935 ) ;
  assign n24919 = n24918 ^ n23299 ^ n18120 ;
  assign n24921 = n18791 ^ n7263 ^ 1'b0 ;
  assign n24922 = n7977 & ~n24921 ;
  assign n24920 = ( ~n15757 & n16198 ) | ( ~n15757 & n20540 ) | ( n16198 & n20540 ) ;
  assign n24923 = n24922 ^ n24920 ^ n10963 ;
  assign n24924 = n15270 ^ n9898 ^ n7448 ;
  assign n24925 = n24924 ^ n18428 ^ n12292 ;
  assign n24926 = n1626 | n3065 ;
  assign n24927 = n24926 ^ n399 ^ 1'b0 ;
  assign n24928 = ( x13 & n13286 ) | ( x13 & ~n24927 ) | ( n13286 & ~n24927 ) ;
  assign n24929 = ( n6524 & n24925 ) | ( n6524 & ~n24928 ) | ( n24925 & ~n24928 ) ;
  assign n24931 = x114 & n4954 ;
  assign n24932 = n24931 ^ n16749 ^ 1'b0 ;
  assign n24930 = ( n5185 & n9136 ) | ( n5185 & ~n13100 ) | ( n9136 & ~n13100 ) ;
  assign n24933 = n24932 ^ n24930 ^ n12592 ;
  assign n24934 = ~n17999 & n21410 ;
  assign n24935 = n19915 ^ n9017 ^ n7738 ;
  assign n24936 = n24935 ^ n13867 ^ n4512 ;
  assign n24937 = ( n10549 & n13746 ) | ( n10549 & n24936 ) | ( n13746 & n24936 ) ;
  assign n24938 = n5066 ^ n1658 ^ 1'b0 ;
  assign n24939 = n10603 & n20633 ;
  assign n24940 = n24939 ^ n22881 ^ 1'b0 ;
  assign n24941 = n20162 ^ n8659 ^ n3730 ;
  assign n24942 = n3063 & ~n5374 ;
  assign n24943 = n24942 ^ n8828 ^ 1'b0 ;
  assign n24944 = n7043 & ~n17149 ;
  assign n24945 = ~n24943 & n24944 ;
  assign n24946 = n24945 ^ n15833 ^ 1'b0 ;
  assign n24947 = n24941 & ~n24946 ;
  assign n24948 = n16267 ^ n7193 ^ 1'b0 ;
  assign n24949 = n20516 ^ n18164 ^ n717 ;
  assign n24950 = n15462 ^ n7986 ^ n5917 ;
  assign n24951 = n24950 ^ n11976 ^ n2379 ;
  assign n24952 = ~n5044 & n6592 ;
  assign n24953 = n4520 & n24952 ;
  assign n24954 = n18119 | n24028 ;
  assign n24955 = n4970 | n24954 ;
  assign n24956 = n6719 & n24955 ;
  assign n24957 = n24956 ^ n10485 ^ 1'b0 ;
  assign n24958 = n24957 ^ n8682 ^ x222 ;
  assign n24960 = ( ~n541 & n754 ) | ( ~n541 & n4015 ) | ( n754 & n4015 ) ;
  assign n24961 = ( n6392 & n12210 ) | ( n6392 & ~n24960 ) | ( n12210 & ~n24960 ) ;
  assign n24959 = n13738 ^ n4627 ^ n740 ;
  assign n24962 = n24961 ^ n24959 ^ n22154 ;
  assign n24963 = ( ~n2782 & n9000 ) | ( ~n2782 & n9679 ) | ( n9000 & n9679 ) ;
  assign n24964 = ( n5034 & ~n7247 ) | ( n5034 & n24963 ) | ( ~n7247 & n24963 ) ;
  assign n24968 = ( n534 & n18224 ) | ( n534 & n23970 ) | ( n18224 & n23970 ) ;
  assign n24965 = n12220 ^ n9496 ^ n1326 ;
  assign n24966 = n24965 ^ n16732 ^ n4954 ;
  assign n24967 = n11446 | n24966 ;
  assign n24969 = n24968 ^ n24967 ^ n21906 ;
  assign n24970 = ( n3064 & n7355 ) | ( n3064 & n22140 ) | ( n7355 & n22140 ) ;
  assign n24971 = ( n3118 & ~n6766 ) | ( n3118 & n14280 ) | ( ~n6766 & n14280 ) ;
  assign n24972 = n24971 ^ n7324 ^ 1'b0 ;
  assign n24973 = n13658 & ~n24972 ;
  assign n24974 = n20523 ^ n11537 ^ 1'b0 ;
  assign n24975 = n1304 & n24974 ;
  assign n24976 = ( n5567 & n14723 ) | ( n5567 & n24975 ) | ( n14723 & n24975 ) ;
  assign n24977 = n24976 ^ n3555 ^ n1125 ;
  assign n24978 = n24977 ^ x160 ^ 1'b0 ;
  assign n24979 = ( ~n4771 & n7495 ) | ( ~n4771 & n13538 ) | ( n7495 & n13538 ) ;
  assign n24981 = n7297 & ~n17747 ;
  assign n24980 = n5632 | n12810 ;
  assign n24982 = n24981 ^ n24980 ^ 1'b0 ;
  assign n24983 = n7845 | n24982 ;
  assign n24984 = ( n556 & n2262 ) | ( n556 & ~n4286 ) | ( n2262 & ~n4286 ) ;
  assign n24985 = n570 & ~n7022 ;
  assign n24986 = ( ~n24983 & n24984 ) | ( ~n24983 & n24985 ) | ( n24984 & n24985 ) ;
  assign n24987 = n355 & ~n11342 ;
  assign n24988 = n24987 ^ n12181 ^ n534 ;
  assign n24989 = ( n14805 & n15638 ) | ( n14805 & ~n24988 ) | ( n15638 & ~n24988 ) ;
  assign n24990 = ( ~n5149 & n8758 ) | ( ~n5149 & n19350 ) | ( n8758 & n19350 ) ;
  assign n24991 = n18184 | n20969 ;
  assign n24992 = n24991 ^ n20580 ^ 1'b0 ;
  assign n24993 = ~n5445 & n11223 ;
  assign n24994 = ~n13421 & n24993 ;
  assign n24995 = ( n3562 & ~n4070 ) | ( n3562 & n21966 ) | ( ~n4070 & n21966 ) ;
  assign n24996 = n24525 ^ n23421 ^ n5567 ;
  assign n24997 = n24995 & n24996 ;
  assign n24998 = ~n9424 & n24997 ;
  assign n24999 = ~n5626 & n19382 ;
  assign n25000 = n17955 & n19357 ;
  assign n25001 = n25000 ^ n1720 ^ 1'b0 ;
  assign n25002 = ( n17319 & n18580 ) | ( n17319 & ~n25001 ) | ( n18580 & ~n25001 ) ;
  assign n25003 = n17758 ^ n574 ^ 1'b0 ;
  assign n25004 = n25003 ^ n10998 ^ n7358 ;
  assign n25005 = n4627 ^ n4371 ^ 1'b0 ;
  assign n25006 = ~n25004 & n25005 ;
  assign n25008 = n6535 ^ n3672 ^ n2026 ;
  assign n25007 = ~n3014 & n12798 ;
  assign n25009 = n25008 ^ n25007 ^ 1'b0 ;
  assign n25010 = n1185 & ~n5391 ;
  assign n25011 = ~n10991 & n25010 ;
  assign n25012 = ( n1407 & n6627 ) | ( n1407 & ~n19904 ) | ( n6627 & ~n19904 ) ;
  assign n25013 = ~n6218 & n25012 ;
  assign n25014 = n20996 ^ n18830 ^ n6887 ;
  assign n25015 = n25014 ^ n3066 ^ 1'b0 ;
  assign n25016 = n7110 & n24958 ;
  assign n25017 = n12825 ^ n11580 ^ n9148 ;
  assign n25018 = ~n365 & n12716 ;
  assign n25019 = ~n12118 & n25018 ;
  assign n25020 = ( x218 & n25017 ) | ( x218 & n25019 ) | ( n25017 & n25019 ) ;
  assign n25021 = n4985 & n21656 ;
  assign n25022 = ~n12072 & n13550 ;
  assign n25023 = n8681 ^ n6619 ^ n1899 ;
  assign n25024 = n25022 & n25023 ;
  assign n25025 = n25024 ^ n14564 ^ 1'b0 ;
  assign n25026 = ( n6809 & n9621 ) | ( n6809 & n12250 ) | ( n9621 & n12250 ) ;
  assign n25027 = n25026 ^ n732 ^ 1'b0 ;
  assign n25028 = n25025 & ~n25027 ;
  assign n25029 = n25028 ^ n13687 ^ n6053 ;
  assign n25030 = ( ~n13742 & n25021 ) | ( ~n13742 & n25029 ) | ( n25021 & n25029 ) ;
  assign n25031 = n25030 ^ n7140 ^ 1'b0 ;
  assign n25032 = ( n6493 & ~n11080 ) | ( n6493 & n25031 ) | ( ~n11080 & n25031 ) ;
  assign n25033 = ( n15098 & n16624 ) | ( n15098 & ~n25032 ) | ( n16624 & ~n25032 ) ;
  assign n25034 = ( n1994 & ~n11053 ) | ( n1994 & n12160 ) | ( ~n11053 & n12160 ) ;
  assign n25035 = n15076 & n16418 ;
  assign n25036 = n23914 & n25035 ;
  assign n25037 = ( n17444 & ~n25034 ) | ( n17444 & n25036 ) | ( ~n25034 & n25036 ) ;
  assign n25043 = n3852 & ~n4939 ;
  assign n25044 = n25043 ^ n3522 ^ 1'b0 ;
  assign n25045 = n1104 & ~n25044 ;
  assign n25046 = n25045 ^ n17897 ^ n12695 ;
  assign n25038 = n5243 & ~n10895 ;
  assign n25039 = n25038 ^ n5051 ^ 1'b0 ;
  assign n25040 = n1339 | n11291 ;
  assign n25041 = n25039 | n25040 ;
  assign n25042 = n21653 & n25041 ;
  assign n25047 = n25046 ^ n25042 ^ 1'b0 ;
  assign n25048 = n4426 & ~n10266 ;
  assign n25049 = n5338 ^ n796 ^ 1'b0 ;
  assign n25050 = n25049 ^ n14152 ^ n11573 ;
  assign n25051 = n15087 ^ n5372 ^ 1'b0 ;
  assign n25052 = n25050 & n25051 ;
  assign n25053 = ( ~n4582 & n9451 ) | ( ~n4582 & n18416 ) | ( n9451 & n18416 ) ;
  assign n25054 = n10813 | n25053 ;
  assign n25055 = ( n2092 & n7110 ) | ( n2092 & n9949 ) | ( n7110 & n9949 ) ;
  assign n25056 = ( n8848 & n19955 ) | ( n8848 & ~n21687 ) | ( n19955 & ~n21687 ) ;
  assign n25057 = ( x7 & n3471 ) | ( x7 & n11183 ) | ( n3471 & n11183 ) ;
  assign n25058 = ( n14063 & ~n16552 ) | ( n14063 & n25057 ) | ( ~n16552 & n25057 ) ;
  assign n25059 = ~n15861 & n25058 ;
  assign n25060 = n25059 ^ n7020 ^ 1'b0 ;
  assign n25061 = ( n25055 & n25056 ) | ( n25055 & ~n25060 ) | ( n25056 & ~n25060 ) ;
  assign n25062 = ( n5485 & ~n8369 ) | ( n5485 & n16063 ) | ( ~n8369 & n16063 ) ;
  assign n25063 = n6706 | n25062 ;
  assign n25064 = n25063 ^ n20064 ^ 1'b0 ;
  assign n25065 = ( n9230 & ~n15025 ) | ( n9230 & n25064 ) | ( ~n15025 & n25064 ) ;
  assign n25066 = n9787 ^ n5428 ^ n2755 ;
  assign n25067 = n1582 | n5334 ;
  assign n25068 = n25067 ^ n1173 ^ 1'b0 ;
  assign n25069 = ~n433 & n24806 ;
  assign n25070 = ( n2707 & ~n20400 ) | ( n2707 & n25069 ) | ( ~n20400 & n25069 ) ;
  assign n25071 = n8068 ^ n1877 ^ n845 ;
  assign n25072 = ~n20011 & n25071 ;
  assign n25073 = n23265 ^ n2362 ^ 1'b0 ;
  assign n25074 = n3050 & n4216 ;
  assign n25075 = n721 & ~n9625 ;
  assign n25076 = ( n8038 & n8450 ) | ( n8038 & n25075 ) | ( n8450 & n25075 ) ;
  assign n25077 = ( ~n9424 & n12011 ) | ( ~n9424 & n25076 ) | ( n12011 & n25076 ) ;
  assign n25078 = ( n8602 & n17864 ) | ( n8602 & ~n23011 ) | ( n17864 & ~n23011 ) ;
  assign n25079 = ~n25077 & n25078 ;
  assign n25080 = n25079 ^ n19960 ^ n12388 ;
  assign n25081 = ( n3761 & ~n25074 ) | ( n3761 & n25080 ) | ( ~n25074 & n25080 ) ;
  assign n25082 = ( n891 & n5040 ) | ( n891 & n6076 ) | ( n5040 & n6076 ) ;
  assign n25083 = n25082 ^ n9930 ^ 1'b0 ;
  assign n25084 = n5748 | n25083 ;
  assign n25085 = ( n6112 & n12629 ) | ( n6112 & n19950 ) | ( n12629 & n19950 ) ;
  assign n25086 = n15627 ^ n6668 ^ n5693 ;
  assign n25087 = n21510 ^ n17605 ^ n11554 ;
  assign n25088 = ( n11816 & n12579 ) | ( n11816 & n15915 ) | ( n12579 & n15915 ) ;
  assign n25089 = ( n12518 & ~n16147 ) | ( n12518 & n20286 ) | ( ~n16147 & n20286 ) ;
  assign n25090 = n16625 ^ n3914 ^ n450 ;
  assign n25091 = ( n2181 & ~n25089 ) | ( n2181 & n25090 ) | ( ~n25089 & n25090 ) ;
  assign n25092 = n13613 | n25091 ;
  assign n25093 = n25088 & ~n25092 ;
  assign n25095 = ( n2175 & n6064 ) | ( n2175 & n6945 ) | ( n6064 & n6945 ) ;
  assign n25096 = ( ~x224 & n7425 ) | ( ~x224 & n7603 ) | ( n7425 & n7603 ) ;
  assign n25097 = n1029 & n25096 ;
  assign n25098 = ( n4109 & n25095 ) | ( n4109 & ~n25097 ) | ( n25095 & ~n25097 ) ;
  assign n25099 = ( n4673 & n8274 ) | ( n4673 & ~n25098 ) | ( n8274 & ~n25098 ) ;
  assign n25094 = n19098 | n22314 ;
  assign n25100 = n25099 ^ n25094 ^ 1'b0 ;
  assign n25101 = ~n2265 & n23398 ;
  assign n25102 = n25101 ^ n17784 ^ 1'b0 ;
  assign n25103 = ~n6525 & n11992 ;
  assign n25104 = ~n15980 & n25103 ;
  assign n25105 = ~n7908 & n17515 ;
  assign n25106 = n4910 & n25105 ;
  assign n25107 = n9163 & ~n13212 ;
  assign n25108 = n25107 ^ n14760 ^ 1'b0 ;
  assign n25109 = ( n8037 & n10784 ) | ( n8037 & ~n14296 ) | ( n10784 & ~n14296 ) ;
  assign n25110 = n9725 ^ n9573 ^ 1'b0 ;
  assign n25111 = n1002 & ~n25110 ;
  assign n25112 = n16855 & n25111 ;
  assign n25113 = n3008 & n25112 ;
  assign n25114 = ( ~n2605 & n15974 ) | ( ~n2605 & n23859 ) | ( n15974 & n23859 ) ;
  assign n25115 = ( n25109 & n25113 ) | ( n25109 & n25114 ) | ( n25113 & n25114 ) ;
  assign n25119 = n14721 ^ n14344 ^ 1'b0 ;
  assign n25120 = ( n560 & n5033 ) | ( n560 & n5674 ) | ( n5033 & n5674 ) ;
  assign n25121 = n25120 ^ n8372 ^ 1'b0 ;
  assign n25122 = n25119 | n25121 ;
  assign n25117 = n1344 & n3405 ;
  assign n25118 = ( n6026 & ~n15919 ) | ( n6026 & n25117 ) | ( ~n15919 & n25117 ) ;
  assign n25116 = ( n1068 & n1347 ) | ( n1068 & ~n6610 ) | ( n1347 & ~n6610 ) ;
  assign n25123 = n25122 ^ n25118 ^ n25116 ;
  assign n25124 = n25123 ^ n19582 ^ x231 ;
  assign n25125 = n12498 ^ n3716 ^ n2108 ;
  assign n25126 = n23065 ^ n18064 ^ n16615 ;
  assign n25129 = ~n934 & n3747 ;
  assign n25130 = n25129 ^ n6245 ^ 1'b0 ;
  assign n25131 = ( n1949 & n6051 ) | ( n1949 & n25130 ) | ( n6051 & n25130 ) ;
  assign n25132 = ( ~n10778 & n23662 ) | ( ~n10778 & n25131 ) | ( n23662 & n25131 ) ;
  assign n25127 = n12580 ^ n7445 ^ n2756 ;
  assign n25128 = ( n399 & ~n10924 ) | ( n399 & n25127 ) | ( ~n10924 & n25127 ) ;
  assign n25133 = n25132 ^ n25128 ^ x147 ;
  assign n25136 = n9335 ^ n8688 ^ n702 ;
  assign n25134 = ( n4030 & ~n4437 ) | ( n4030 & n21169 ) | ( ~n4437 & n21169 ) ;
  assign n25135 = n4263 | n25134 ;
  assign n25137 = n25136 ^ n25135 ^ 1'b0 ;
  assign n25138 = n16196 ^ n14037 ^ n5802 ;
  assign n25139 = ( n6012 & n25137 ) | ( n6012 & ~n25138 ) | ( n25137 & ~n25138 ) ;
  assign n25140 = ( n501 & n7371 ) | ( n501 & n14490 ) | ( n7371 & n14490 ) ;
  assign n25141 = n9635 | n25140 ;
  assign n25142 = n1818 | n25141 ;
  assign n25143 = ( n6910 & n25139 ) | ( n6910 & n25142 ) | ( n25139 & n25142 ) ;
  assign n25144 = ( n16168 & n20603 ) | ( n16168 & ~n24808 ) | ( n20603 & ~n24808 ) ;
  assign n25145 = n10635 | n16882 ;
  assign n25146 = n4902 & ~n25145 ;
  assign n25147 = ( n1606 & n2305 ) | ( n1606 & ~n5279 ) | ( n2305 & ~n5279 ) ;
  assign n25148 = ~n1982 & n25147 ;
  assign n25150 = n7503 ^ n5630 ^ n4723 ;
  assign n25149 = ~n10303 & n12118 ;
  assign n25151 = n25150 ^ n25149 ^ n17945 ;
  assign n25152 = ( n16010 & ~n25148 ) | ( n16010 & n25151 ) | ( ~n25148 & n25151 ) ;
  assign n25153 = n13002 & n25152 ;
  assign n25154 = ~n15501 & n25153 ;
  assign n25155 = n5985 & n25154 ;
  assign n25158 = n13663 ^ n13406 ^ n7845 ;
  assign n25156 = n9740 & n21113 ;
  assign n25157 = ~n21562 & n25156 ;
  assign n25159 = n25158 ^ n25157 ^ n5459 ;
  assign n25164 = x172 & ~n4178 ;
  assign n25160 = ( n3735 & ~n15113 ) | ( n3735 & n16393 ) | ( ~n15113 & n16393 ) ;
  assign n25161 = ( ~n1096 & n2084 ) | ( ~n1096 & n25160 ) | ( n2084 & n25160 ) ;
  assign n25162 = n25161 ^ n2931 ^ 1'b0 ;
  assign n25163 = n5243 & n25162 ;
  assign n25165 = n25164 ^ n25163 ^ n1173 ;
  assign n25166 = ~n4538 & n10174 ;
  assign n25167 = ~n18791 & n25166 ;
  assign n25168 = n25167 ^ n6441 ^ 1'b0 ;
  assign n25169 = ( n2797 & n15611 ) | ( n2797 & n25168 ) | ( n15611 & n25168 ) ;
  assign n25170 = n370 & ~n2016 ;
  assign n25171 = n25170 ^ n23081 ^ 1'b0 ;
  assign n25172 = ( n8967 & n16704 ) | ( n8967 & n25171 ) | ( n16704 & n25171 ) ;
  assign n25173 = ( n3951 & n4112 ) | ( n3951 & ~n18162 ) | ( n4112 & ~n18162 ) ;
  assign n25174 = ( ~n15371 & n23873 ) | ( ~n15371 & n25173 ) | ( n23873 & n25173 ) ;
  assign n25175 = ( n9444 & ~n10824 ) | ( n9444 & n25174 ) | ( ~n10824 & n25174 ) ;
  assign n25176 = n17557 ^ n6921 ^ n3993 ;
  assign n25177 = n25176 ^ n11679 ^ 1'b0 ;
  assign n25178 = n25177 ^ n13985 ^ 1'b0 ;
  assign n25179 = n1028 & ~n25178 ;
  assign n25180 = n25179 ^ n5836 ^ 1'b0 ;
  assign n25181 = n25175 & ~n25180 ;
  assign n25182 = ~n3997 & n7688 ;
  assign n25183 = n1718 | n25182 ;
  assign n25184 = n10851 & n25183 ;
  assign n25185 = n24930 ^ n18818 ^ 1'b0 ;
  assign n25186 = n6671 & ~n13930 ;
  assign n25187 = ~n2352 & n25186 ;
  assign n25188 = ( ~n3014 & n6111 ) | ( ~n3014 & n25187 ) | ( n6111 & n25187 ) ;
  assign n25189 = ( n18818 & n19262 ) | ( n18818 & ~n25188 ) | ( n19262 & ~n25188 ) ;
  assign n25190 = n2804 & n15356 ;
  assign n25191 = n17012 ^ n2485 ^ 1'b0 ;
  assign n25192 = ( n10133 & ~n12815 ) | ( n10133 & n13887 ) | ( ~n12815 & n13887 ) ;
  assign n25193 = n19326 ^ n1376 ^ 1'b0 ;
  assign n25194 = ( ~n13503 & n25192 ) | ( ~n13503 & n25193 ) | ( n25192 & n25193 ) ;
  assign n25195 = n25194 ^ n8289 ^ n4234 ;
  assign n25196 = n18116 ^ n17142 ^ n7876 ;
  assign n25197 = n1302 & n6178 ;
  assign n25198 = n25197 ^ n4982 ^ 1'b0 ;
  assign n25199 = n25198 ^ n4179 ^ 1'b0 ;
  assign n25200 = n25196 | n25199 ;
  assign n25201 = n25200 ^ n5736 ^ 1'b0 ;
  assign n25202 = n7466 & ~n25201 ;
  assign n25203 = n1422 & n8964 ;
  assign n25204 = n25203 ^ n1747 ^ 1'b0 ;
  assign n25208 = ~n12012 & n24716 ;
  assign n25209 = n5363 & n25208 ;
  assign n25205 = n17913 ^ x163 ^ 1'b0 ;
  assign n25206 = n16435 & n25205 ;
  assign n25207 = n11339 | n25206 ;
  assign n25210 = n25209 ^ n25207 ^ n9888 ;
  assign n25211 = n24306 ^ n23594 ^ 1'b0 ;
  assign n25212 = n6240 ^ n5704 ^ 1'b0 ;
  assign n25213 = ( n3773 & n13969 ) | ( n3773 & ~n20077 ) | ( n13969 & ~n20077 ) ;
  assign n25214 = n25212 & ~n25213 ;
  assign n25215 = n25211 & n25214 ;
  assign n25216 = ( ~n8976 & n13184 ) | ( ~n8976 & n25215 ) | ( n13184 & n25215 ) ;
  assign n25221 = n14303 ^ n2781 ^ n2026 ;
  assign n25219 = n14835 ^ n13434 ^ n3697 ;
  assign n25220 = n25219 ^ n21943 ^ n13410 ;
  assign n25217 = n19936 ^ n2353 ^ 1'b0 ;
  assign n25218 = n5928 & ~n25217 ;
  assign n25222 = n25221 ^ n25220 ^ n25218 ;
  assign n25223 = ( n11748 & ~n20189 ) | ( n11748 & n25222 ) | ( ~n20189 & n25222 ) ;
  assign n25224 = n25223 ^ n10855 ^ n5880 ;
  assign n25228 = n4399 ^ n2195 ^ 1'b0 ;
  assign n25225 = ~n4174 & n10169 ;
  assign n25226 = ~n6605 & n25225 ;
  assign n25227 = ( n2073 & n5189 ) | ( n2073 & ~n25226 ) | ( n5189 & ~n25226 ) ;
  assign n25229 = n25228 ^ n25227 ^ 1'b0 ;
  assign n25230 = n21775 & n25229 ;
  assign n25231 = n4933 & n5172 ;
  assign n25232 = n25231 ^ n7799 ^ 1'b0 ;
  assign n25233 = n15067 & ~n25232 ;
  assign n25234 = n25233 ^ n5907 ^ 1'b0 ;
  assign n25235 = n24044 ^ n10912 ^ n4485 ;
  assign n25236 = n25235 ^ n9772 ^ 1'b0 ;
  assign n25237 = n25234 & ~n25236 ;
  assign n25238 = n3242 & n15364 ;
  assign n25239 = n10948 & n25238 ;
  assign n25240 = n25239 ^ n11271 ^ 1'b0 ;
  assign n25241 = n8806 | n25240 ;
  assign n25250 = n3217 | n4331 ;
  assign n25251 = n14999 & ~n25250 ;
  assign n25243 = n20965 ^ n19699 ^ n3936 ;
  assign n25242 = ~n9122 & n10378 ;
  assign n25244 = n25243 ^ n25242 ^ n18123 ;
  assign n25245 = x108 & ~n25244 ;
  assign n25246 = ~n13050 & n25245 ;
  assign n25247 = ( n6861 & ~n15243 ) | ( n6861 & n25246 ) | ( ~n15243 & n25246 ) ;
  assign n25248 = n25247 ^ n22937 ^ 1'b0 ;
  assign n25249 = n3102 & ~n25248 ;
  assign n25252 = n25251 ^ n25249 ^ n8573 ;
  assign n25253 = ( ~n22472 & n25241 ) | ( ~n22472 & n25252 ) | ( n25241 & n25252 ) ;
  assign n25254 = n11828 ^ n10813 ^ 1'b0 ;
  assign n25255 = ( n2430 & n5163 ) | ( n2430 & ~n24178 ) | ( n5163 & ~n24178 ) ;
  assign n25256 = n12010 ^ n504 ^ 1'b0 ;
  assign n25257 = ( n6626 & n7425 ) | ( n6626 & n25256 ) | ( n7425 & n25256 ) ;
  assign n25258 = n7319 | n9602 ;
  assign n25259 = n25258 ^ n21966 ^ 1'b0 ;
  assign n25260 = n25257 & ~n25259 ;
  assign n25261 = n14106 ^ n9947 ^ n1459 ;
  assign n25262 = n25261 ^ n530 ^ 1'b0 ;
  assign n25263 = ( n678 & ~n4812 ) | ( n678 & n11592 ) | ( ~n4812 & n11592 ) ;
  assign n25264 = n25263 ^ n15222 ^ 1'b0 ;
  assign n25265 = ~n12963 & n25264 ;
  assign n25266 = ~n23686 & n25265 ;
  assign n25267 = n7793 ^ n5829 ^ 1'b0 ;
  assign n25268 = n25267 ^ n18361 ^ 1'b0 ;
  assign n25269 = ( ~n12254 & n17256 ) | ( ~n12254 & n24644 ) | ( n17256 & n24644 ) ;
  assign n25270 = n22423 ^ n12752 ^ n11652 ;
  assign n25271 = n25270 ^ n24280 ^ n8175 ;
  assign n25274 = ~n9684 & n10940 ;
  assign n25273 = n1490 | n4362 ;
  assign n25272 = ( ~n2302 & n3929 ) | ( ~n2302 & n23596 ) | ( n3929 & n23596 ) ;
  assign n25275 = n25274 ^ n25273 ^ n25272 ;
  assign n25276 = ~n4625 & n25275 ;
  assign n25277 = n10421 ^ n3352 ^ 1'b0 ;
  assign n25278 = n25277 ^ n23803 ^ n21712 ;
  assign n25279 = n8601 ^ n3889 ^ 1'b0 ;
  assign n25280 = n15024 & n25279 ;
  assign n25284 = ( n8203 & ~n21165 ) | ( n8203 & n21334 ) | ( ~n21165 & n21334 ) ;
  assign n25281 = n16230 ^ n3970 ^ 1'b0 ;
  assign n25282 = ~n21540 & n25281 ;
  assign n25283 = n13819 & n25282 ;
  assign n25285 = n25284 ^ n25283 ^ 1'b0 ;
  assign n25286 = n1649 & ~n12098 ;
  assign n25291 = n653 & ~n14927 ;
  assign n25292 = n25291 ^ n10403 ^ 1'b0 ;
  assign n25289 = n4888 & n7101 ;
  assign n25290 = n1870 & n25289 ;
  assign n25287 = ( ~n585 & n7260 ) | ( ~n585 & n16130 ) | ( n7260 & n16130 ) ;
  assign n25288 = n25287 ^ n12409 ^ 1'b0 ;
  assign n25293 = n25292 ^ n25290 ^ n25288 ;
  assign n25294 = n15115 ^ n13148 ^ n9835 ;
  assign n25295 = ( n12249 & n13875 ) | ( n12249 & ~n23653 ) | ( n13875 & ~n23653 ) ;
  assign n25297 = ( n2895 & n15845 ) | ( n2895 & n20150 ) | ( n15845 & n20150 ) ;
  assign n25296 = n7625 ^ n3222 ^ 1'b0 ;
  assign n25298 = n25297 ^ n25296 ^ n24350 ;
  assign n25299 = ( n4590 & n5153 ) | ( n4590 & n10550 ) | ( n5153 & n10550 ) ;
  assign n25300 = n5804 & n10797 ;
  assign n25301 = ~n1175 & n3720 ;
  assign n25302 = ( n14866 & n21163 ) | ( n14866 & ~n25301 ) | ( n21163 & ~n25301 ) ;
  assign n25303 = ~n393 & n5293 ;
  assign n25304 = ( ~n1513 & n4667 ) | ( ~n1513 & n23208 ) | ( n4667 & n23208 ) ;
  assign n25305 = ( n4584 & ~n25303 ) | ( n4584 & n25304 ) | ( ~n25303 & n25304 ) ;
  assign n25306 = n14270 & n25305 ;
  assign n25307 = ~n23772 & n25306 ;
  assign n25308 = ( ~n1444 & n3178 ) | ( ~n1444 & n7717 ) | ( n3178 & n7717 ) ;
  assign n25309 = ( ~n2285 & n15592 ) | ( ~n2285 & n17273 ) | ( n15592 & n17273 ) ;
  assign n25310 = n8022 & n13140 ;
  assign n25311 = ~n9173 & n25310 ;
  assign n25312 = n7527 & ~n25311 ;
  assign n25313 = n25312 ^ n19372 ^ n2867 ;
  assign n25314 = ( ~n7823 & n9285 ) | ( ~n7823 & n25313 ) | ( n9285 & n25313 ) ;
  assign n25315 = ( n25308 & n25309 ) | ( n25308 & ~n25314 ) | ( n25309 & ~n25314 ) ;
  assign n25316 = n9717 ^ n9174 ^ n1708 ;
  assign n25317 = n25316 ^ n9140 ^ n3223 ;
  assign n25320 = n15298 ^ n13936 ^ n11667 ;
  assign n25321 = ( n2120 & n15015 ) | ( n2120 & ~n25320 ) | ( n15015 & ~n25320 ) ;
  assign n25318 = n3030 & ~n15428 ;
  assign n25319 = n25318 ^ n18661 ^ 1'b0 ;
  assign n25322 = n25321 ^ n25319 ^ 1'b0 ;
  assign n25323 = n6670 | n25322 ;
  assign n25324 = n4279 ^ n401 ^ 1'b0 ;
  assign n25325 = n4342 & ~n25324 ;
  assign n25326 = n9745 | n13083 ;
  assign n25327 = n25326 ^ n16233 ^ 1'b0 ;
  assign n25328 = n9394 | n10849 ;
  assign n25329 = ( n9703 & ~n13618 ) | ( n9703 & n25328 ) | ( ~n13618 & n25328 ) ;
  assign n25330 = ( ~n1299 & n11725 ) | ( ~n1299 & n25329 ) | ( n11725 & n25329 ) ;
  assign n25331 = n10152 ^ n5992 ^ 1'b0 ;
  assign n25332 = n4630 & n25331 ;
  assign n25333 = ( n14231 & ~n14691 ) | ( n14231 & n25332 ) | ( ~n14691 & n25332 ) ;
  assign n25334 = ( ~n5405 & n10062 ) | ( ~n5405 & n10196 ) | ( n10062 & n10196 ) ;
  assign n25335 = ~n4792 & n16010 ;
  assign n25336 = n25335 ^ n9260 ^ n1921 ;
  assign n25337 = n25336 ^ n3268 ^ n1117 ;
  assign n25338 = n25334 & ~n25337 ;
  assign n25342 = n7270 ^ n4145 ^ x191 ;
  assign n25343 = ( ~n5782 & n22096 ) | ( ~n5782 & n25342 ) | ( n22096 & n25342 ) ;
  assign n25344 = ( ~n5710 & n14355 ) | ( ~n5710 & n25343 ) | ( n14355 & n25343 ) ;
  assign n25339 = ( ~n14630 & n18385 ) | ( ~n14630 & n22540 ) | ( n18385 & n22540 ) ;
  assign n25340 = ( ~n12802 & n20717 ) | ( ~n12802 & n25339 ) | ( n20717 & n25339 ) ;
  assign n25341 = n8319 | n25340 ;
  assign n25345 = n25344 ^ n25341 ^ 1'b0 ;
  assign n25346 = ~n4067 & n17121 ;
  assign n25347 = ~n14080 & n25346 ;
  assign n25348 = ( ~n10428 & n22250 ) | ( ~n10428 & n25347 ) | ( n22250 & n25347 ) ;
  assign n25350 = ( n1078 & n4879 ) | ( n1078 & ~n5871 ) | ( n4879 & ~n5871 ) ;
  assign n25351 = n22283 ^ n1606 ^ 1'b0 ;
  assign n25352 = n25350 | n25351 ;
  assign n25349 = ( n11947 & n11987 ) | ( n11947 & n20932 ) | ( n11987 & n20932 ) ;
  assign n25353 = n25352 ^ n25349 ^ n24461 ;
  assign n25355 = ( n6491 & ~n7727 ) | ( n6491 & n17418 ) | ( ~n7727 & n17418 ) ;
  assign n25356 = ~n11475 & n25355 ;
  assign n25357 = ~n6270 & n25356 ;
  assign n25354 = n8536 & ~n12013 ;
  assign n25358 = n25357 ^ n25354 ^ 1'b0 ;
  assign n25359 = ( ~n911 & n5035 ) | ( ~n911 & n16922 ) | ( n5035 & n16922 ) ;
  assign n25360 = n24521 | n25359 ;
  assign n25361 = n25358 | n25360 ;
  assign n25362 = n15784 ^ n12029 ^ 1'b0 ;
  assign n25363 = ~n15143 & n25362 ;
  assign n25364 = n10399 ^ n6561 ^ n1273 ;
  assign n25365 = n25364 ^ n343 ^ 1'b0 ;
  assign n25366 = n25365 ^ n17241 ^ n13452 ;
  assign n25367 = ( ~n3502 & n4540 ) | ( ~n3502 & n25366 ) | ( n4540 & n25366 ) ;
  assign n25368 = ( n2665 & ~n4418 ) | ( n2665 & n6320 ) | ( ~n4418 & n6320 ) ;
  assign n25369 = ( n6391 & n7322 ) | ( n6391 & ~n25368 ) | ( n7322 & ~n25368 ) ;
  assign n25370 = n25369 ^ n17411 ^ 1'b0 ;
  assign n25371 = ~n11448 & n25370 ;
  assign n25372 = ~n261 & n25371 ;
  assign n25373 = n25372 ^ n353 ^ 1'b0 ;
  assign n25374 = n12132 ^ n9528 ^ n7434 ;
  assign n25375 = n15866 ^ n5262 ^ n2984 ;
  assign n25376 = n10460 ^ n7706 ^ 1'b0 ;
  assign n25377 = n25376 ^ n13016 ^ 1'b0 ;
  assign n25378 = n5849 | n25377 ;
  assign n25379 = n25375 | n25378 ;
  assign n25380 = n25379 ^ n11178 ^ 1'b0 ;
  assign n25381 = n25380 ^ n12598 ^ 1'b0 ;
  assign n25382 = n2737 ^ n825 ^ 1'b0 ;
  assign n25383 = n25382 ^ n19952 ^ n3989 ;
  assign n25384 = ( n15553 & n25381 ) | ( n15553 & ~n25383 ) | ( n25381 & ~n25383 ) ;
  assign n25385 = n1711 & ~n25384 ;
  assign n25386 = n25374 & n25385 ;
  assign n25387 = n9301 ^ n8274 ^ n4524 ;
  assign n25388 = n13989 & n15170 ;
  assign n25389 = ~n25387 & n25388 ;
  assign n25390 = n328 & n5005 ;
  assign n25391 = n25390 ^ n18958 ^ 1'b0 ;
  assign n25392 = n25391 ^ n17100 ^ n9911 ;
  assign n25393 = ~n8305 & n25392 ;
  assign n25394 = ~n9073 & n25393 ;
  assign n25398 = n24574 ^ n9750 ^ 1'b0 ;
  assign n25399 = ( n17834 & ~n19123 ) | ( n17834 & n25398 ) | ( ~n19123 & n25398 ) ;
  assign n25400 = n25399 ^ n7577 ^ n790 ;
  assign n25396 = n24864 ^ n12089 ^ n4539 ;
  assign n25395 = n9956 ^ n989 ^ n306 ;
  assign n25397 = n25396 ^ n25395 ^ n2708 ;
  assign n25401 = n25400 ^ n25397 ^ n802 ;
  assign n25405 = ~x222 & n15556 ;
  assign n25403 = n16047 ^ n6936 ^ 1'b0 ;
  assign n25402 = n5184 ^ n2016 ^ 1'b0 ;
  assign n25404 = n25403 ^ n25402 ^ n16603 ;
  assign n25406 = n25405 ^ n25404 ^ 1'b0 ;
  assign n25407 = n6048 ^ n2393 ^ 1'b0 ;
  assign n25408 = n11328 & ~n25407 ;
  assign n25409 = n6730 & n8340 ;
  assign n25410 = ( ~n18994 & n25408 ) | ( ~n18994 & n25409 ) | ( n25408 & n25409 ) ;
  assign n25411 = n25410 ^ n3014 ^ 1'b0 ;
  assign n25412 = n19811 & ~n25411 ;
  assign n25413 = n16081 ^ n6997 ^ n3855 ;
  assign n25414 = n6117 & n11065 ;
  assign n25415 = n25413 & n25414 ;
  assign n25416 = ( n1665 & n5026 ) | ( n1665 & ~n25415 ) | ( n5026 & ~n25415 ) ;
  assign n25417 = ( n4328 & ~n13895 ) | ( n4328 & n25416 ) | ( ~n13895 & n25416 ) ;
  assign n25418 = n14602 ^ n8718 ^ 1'b0 ;
  assign n25421 = n12035 ^ n2357 ^ 1'b0 ;
  assign n25422 = n7754 & ~n25421 ;
  assign n25419 = ~n1473 & n15254 ;
  assign n25420 = n25419 ^ n11263 ^ 1'b0 ;
  assign n25423 = n25422 ^ n25420 ^ 1'b0 ;
  assign n25424 = ( ~n1378 & n12215 ) | ( ~n1378 & n25423 ) | ( n12215 & n25423 ) ;
  assign n25425 = ( n2486 & n8175 ) | ( n2486 & ~n10007 ) | ( n8175 & ~n10007 ) ;
  assign n25426 = n3910 & ~n11422 ;
  assign n25427 = n25425 & n25426 ;
  assign n25428 = n23998 ^ n9753 ^ n3504 ;
  assign n25429 = ~n4057 & n25428 ;
  assign n25430 = ~n14428 & n25429 ;
  assign n25431 = ( n1523 & n10360 ) | ( n1523 & ~n19843 ) | ( n10360 & ~n19843 ) ;
  assign n25432 = n21447 & n25431 ;
  assign n25433 = n25432 ^ n14455 ^ 1'b0 ;
  assign n25434 = ( ~n6687 & n25430 ) | ( ~n6687 & n25433 ) | ( n25430 & n25433 ) ;
  assign n25435 = n7454 & ~n21440 ;
  assign n25436 = n25435 ^ n21332 ^ 1'b0 ;
  assign n25437 = n25436 ^ n25292 ^ n14837 ;
  assign n25438 = ( n19059 & n19299 ) | ( n19059 & ~n22069 ) | ( n19299 & ~n22069 ) ;
  assign n25439 = n14223 ^ n7118 ^ 1'b0 ;
  assign n25440 = ~n17029 & n25439 ;
  assign n25441 = n20009 ^ x224 ^ 1'b0 ;
  assign n25442 = n24395 ^ n9591 ^ 1'b0 ;
  assign n25443 = ( n8145 & n14167 ) | ( n8145 & ~n25442 ) | ( n14167 & ~n25442 ) ;
  assign n25445 = n9167 ^ n4915 ^ n2141 ;
  assign n25446 = n13335 | n25445 ;
  assign n25447 = n14226 & ~n25446 ;
  assign n25444 = n18364 ^ n15997 ^ 1'b0 ;
  assign n25448 = n25447 ^ n25444 ^ n10849 ;
  assign n25449 = n4994 & ~n6604 ;
  assign n25450 = n25449 ^ n1376 ^ 1'b0 ;
  assign n25451 = ( ~n2427 & n6188 ) | ( ~n2427 & n19662 ) | ( n6188 & n19662 ) ;
  assign n25452 = ( n6295 & n20160 ) | ( n6295 & ~n20453 ) | ( n20160 & ~n20453 ) ;
  assign n25453 = ( n6282 & n14738 ) | ( n6282 & ~n25452 ) | ( n14738 & ~n25452 ) ;
  assign n25454 = ( n25450 & ~n25451 ) | ( n25450 & n25453 ) | ( ~n25451 & n25453 ) ;
  assign n25455 = ( ~n3964 & n12980 ) | ( ~n3964 & n15050 ) | ( n12980 & n15050 ) ;
  assign n25456 = n25455 ^ n11825 ^ n1265 ;
  assign n25457 = n14519 ^ n6547 ^ n5766 ;
  assign n25458 = ~n25456 & n25457 ;
  assign n25459 = ( n2178 & n3520 ) | ( n2178 & n19704 ) | ( n3520 & n19704 ) ;
  assign n25460 = n8854 & ~n9123 ;
  assign n25461 = n25459 & n25460 ;
  assign n25462 = n25461 ^ n460 ^ 1'b0 ;
  assign n25463 = n25458 | n25462 ;
  assign n25464 = n12322 ^ n11289 ^ 1'b0 ;
  assign n25465 = ~n1317 & n25464 ;
  assign n25466 = n25465 ^ n13959 ^ 1'b0 ;
  assign n25467 = ( n6234 & n19785 ) | ( n6234 & n25466 ) | ( n19785 & n25466 ) ;
  assign n25468 = n25467 ^ n6765 ^ n4810 ;
  assign n25469 = n25468 ^ n15657 ^ 1'b0 ;
  assign n25470 = ~n8928 & n18097 ;
  assign n25471 = ~n19810 & n25470 ;
  assign n25472 = n15530 ^ n6930 ^ n1507 ;
  assign n25473 = ( n15476 & n16102 ) | ( n15476 & n18671 ) | ( n16102 & n18671 ) ;
  assign n25474 = n16156 ^ n9032 ^ n8108 ;
  assign n25484 = n13921 ^ n10334 ^ n4931 ;
  assign n25475 = n14911 ^ n3673 ^ 1'b0 ;
  assign n25476 = n10523 ^ n3284 ^ 1'b0 ;
  assign n25477 = ~n16561 & n25476 ;
  assign n25478 = n7417 & ~n8315 ;
  assign n25479 = n3452 & ~n7922 ;
  assign n25480 = ( n1391 & n1413 ) | ( n1391 & n1897 ) | ( n1413 & n1897 ) ;
  assign n25481 = ( ~n19491 & n22259 ) | ( ~n19491 & n25480 ) | ( n22259 & n25480 ) ;
  assign n25482 = ( n25478 & ~n25479 ) | ( n25478 & n25481 ) | ( ~n25479 & n25481 ) ;
  assign n25483 = ( n25475 & ~n25477 ) | ( n25475 & n25482 ) | ( ~n25477 & n25482 ) ;
  assign n25485 = n25484 ^ n25483 ^ n16867 ;
  assign n25489 = n7018 ^ n874 ^ 1'b0 ;
  assign n25487 = ( n1898 & n6141 ) | ( n1898 & ~n7068 ) | ( n6141 & ~n7068 ) ;
  assign n25486 = ( n4925 & ~n5943 ) | ( n4925 & n22497 ) | ( ~n5943 & n22497 ) ;
  assign n25488 = n25487 ^ n25486 ^ 1'b0 ;
  assign n25490 = n25489 ^ n25488 ^ 1'b0 ;
  assign n25491 = ( n10495 & ~n22832 ) | ( n10495 & n25490 ) | ( ~n22832 & n25490 ) ;
  assign n25492 = n10991 ^ n3398 ^ n1911 ;
  assign n25493 = ( n11379 & n20527 ) | ( n11379 & ~n25492 ) | ( n20527 & ~n25492 ) ;
  assign n25494 = ( n6232 & ~n15980 ) | ( n6232 & n25493 ) | ( ~n15980 & n25493 ) ;
  assign n25495 = n6622 & n18444 ;
  assign n25496 = ~n11048 & n25495 ;
  assign n25497 = n16803 & n19648 ;
  assign n25498 = n25497 ^ n14938 ^ n14474 ;
  assign n25499 = n6041 & ~n25044 ;
  assign n25500 = n25499 ^ n21443 ^ 1'b0 ;
  assign n25501 = ( n8252 & ~n24170 ) | ( n8252 & n25500 ) | ( ~n24170 & n25500 ) ;
  assign n25502 = n2250 & n9289 ;
  assign n25503 = ( ~n1173 & n3673 ) | ( ~n1173 & n19240 ) | ( n3673 & n19240 ) ;
  assign n25504 = ( n10372 & n24733 ) | ( n10372 & ~n25503 ) | ( n24733 & ~n25503 ) ;
  assign n25505 = n5718 ^ n1951 ^ 1'b0 ;
  assign n25506 = n6376 & ~n11166 ;
  assign n25507 = n25506 ^ n24019 ^ 1'b0 ;
  assign n25508 = n25505 & ~n25507 ;
  assign n25509 = n18820 ^ n10438 ^ n2517 ;
  assign n25510 = n25509 ^ n17032 ^ 1'b0 ;
  assign n25511 = ( n22179 & n25508 ) | ( n22179 & ~n25510 ) | ( n25508 & ~n25510 ) ;
  assign n25512 = n24256 ^ n10449 ^ n8022 ;
  assign n25513 = ( ~n11328 & n23517 ) | ( ~n11328 & n25512 ) | ( n23517 & n25512 ) ;
  assign n25514 = n19368 ^ n12898 ^ 1'b0 ;
  assign n25515 = n12609 | n16500 ;
  assign n25516 = n25515 ^ n6841 ^ 1'b0 ;
  assign n25517 = ( ~n10151 & n25514 ) | ( ~n10151 & n25516 ) | ( n25514 & n25516 ) ;
  assign n25518 = n5675 & n8247 ;
  assign n25519 = n13231 ^ n10538 ^ n3452 ;
  assign n25520 = ( n7760 & n25518 ) | ( n7760 & ~n25519 ) | ( n25518 & ~n25519 ) ;
  assign n25521 = n16445 & ~n24224 ;
  assign n25522 = n25521 ^ n18905 ^ 1'b0 ;
  assign n25523 = n25520 & ~n25522 ;
  assign n25524 = n3900 & n25523 ;
  assign n25525 = ~n3713 & n11947 ;
  assign n25526 = n22801 ^ n11210 ^ 1'b0 ;
  assign n25527 = n25525 & n25526 ;
  assign n25528 = ( ~n10274 & n15172 ) | ( ~n10274 & n25527 ) | ( n15172 & n25527 ) ;
  assign n25529 = n22086 ^ n7861 ^ n6528 ;
  assign n25530 = n18680 & ~n20835 ;
  assign n25531 = n3025 | n10619 ;
  assign n25533 = n18385 ^ n14443 ^ 1'b0 ;
  assign n25534 = n25533 ^ n8316 ^ 1'b0 ;
  assign n25532 = n1202 | n4893 ;
  assign n25535 = n25534 ^ n25532 ^ n4485 ;
  assign n25536 = n637 | n25535 ;
  assign n25537 = n25536 ^ n24291 ^ n5192 ;
  assign n25538 = n21506 ^ n19875 ^ n7207 ;
  assign n25539 = n10628 & n25538 ;
  assign n25540 = n25539 ^ n25369 ^ n4911 ;
  assign n25541 = ( ~n459 & n1307 ) | ( ~n459 & n2974 ) | ( n1307 & n2974 ) ;
  assign n25542 = ( n4994 & n10327 ) | ( n4994 & n25541 ) | ( n10327 & n25541 ) ;
  assign n25543 = ( n7667 & n10017 ) | ( n7667 & ~n25542 ) | ( n10017 & ~n25542 ) ;
  assign n25544 = n5449 | n25543 ;
  assign n25545 = n2984 | n25544 ;
  assign n25546 = n12089 ^ n9477 ^ 1'b0 ;
  assign n25547 = n14544 & n25546 ;
  assign n25548 = n4297 ^ n650 ^ x173 ;
  assign n25549 = n25548 ^ n8751 ^ 1'b0 ;
  assign n25550 = n16332 | n22025 ;
  assign n25551 = ~n7207 & n25550 ;
  assign n25552 = n25549 & n25551 ;
  assign n25553 = n25036 ^ n21103 ^ n2197 ;
  assign n25554 = n8549 ^ n5980 ^ n1450 ;
  assign n25555 = ( ~n3614 & n4166 ) | ( ~n3614 & n25554 ) | ( n4166 & n25554 ) ;
  assign n25556 = ( ~n1588 & n4015 ) | ( ~n1588 & n20594 ) | ( n4015 & n20594 ) ;
  assign n25557 = ( n13632 & ~n25555 ) | ( n13632 & n25556 ) | ( ~n25555 & n25556 ) ;
  assign n25558 = n8889 ^ n8481 ^ 1'b0 ;
  assign n25559 = n25558 ^ n11533 ^ n7438 ;
  assign n25560 = n25559 ^ n14047 ^ 1'b0 ;
  assign n25561 = n25560 ^ n17781 ^ n11873 ;
  assign n25564 = ( n2655 & ~n6525 ) | ( n2655 & n8203 ) | ( ~n6525 & n8203 ) ;
  assign n25562 = ~n1705 & n8308 ;
  assign n25563 = ~n13840 & n25562 ;
  assign n25565 = n25564 ^ n25563 ^ n9707 ;
  assign n25566 = n25565 ^ n11556 ^ n5237 ;
  assign n25567 = n24511 ^ n9698 ^ n1402 ;
  assign n25569 = n19829 ^ n7237 ^ n2217 ;
  assign n25568 = n12371 & ~n19401 ;
  assign n25570 = n25569 ^ n25568 ^ 1'b0 ;
  assign n25571 = n25570 ^ n21754 ^ 1'b0 ;
  assign n25572 = n11219 & n25571 ;
  assign n25574 = n20423 ^ n7141 ^ 1'b0 ;
  assign n25575 = n7973 & ~n25574 ;
  assign n25573 = n18823 ^ n8262 ^ 1'b0 ;
  assign n25576 = n25575 ^ n25573 ^ 1'b0 ;
  assign n25577 = ( ~n9911 & n13481 ) | ( ~n9911 & n17038 ) | ( n13481 & n17038 ) ;
  assign n25578 = ( n7826 & n19452 ) | ( n7826 & ~n22337 ) | ( n19452 & ~n22337 ) ;
  assign n25579 = n16005 ^ n3528 ^ 1'b0 ;
  assign n25580 = n257 & ~n25579 ;
  assign n25581 = n25580 ^ n17413 ^ 1'b0 ;
  assign n25584 = ( ~n11498 & n11962 ) | ( ~n11498 & n16837 ) | ( n11962 & n16837 ) ;
  assign n25582 = n14205 ^ n8988 ^ n1278 ;
  assign n25583 = ~n3953 & n25582 ;
  assign n25585 = n25584 ^ n25583 ^ 1'b0 ;
  assign n25586 = n25303 ^ n15840 ^ n1321 ;
  assign n25587 = n7635 & n11160 ;
  assign n25588 = ~n25586 & n25587 ;
  assign n25589 = n6397 ^ n4591 ^ n3422 ;
  assign n25590 = n1123 & n25589 ;
  assign n25591 = ~n25588 & n25590 ;
  assign n25593 = n5637 ^ n2367 ^ n1535 ;
  assign n25594 = n13609 ^ n7209 ^ n7206 ;
  assign n25595 = n25594 ^ n6226 ^ 1'b0 ;
  assign n25596 = n8569 | n25595 ;
  assign n25597 = n22251 | n25596 ;
  assign n25598 = n6212 & ~n25597 ;
  assign n25599 = ( ~n18159 & n25593 ) | ( ~n18159 & n25598 ) | ( n25593 & n25598 ) ;
  assign n25600 = n14853 & ~n25599 ;
  assign n25601 = n9463 & n25600 ;
  assign n25592 = n5639 ^ n5533 ^ n1870 ;
  assign n25602 = n25601 ^ n25592 ^ n311 ;
  assign n25603 = n25602 ^ n3406 ^ 1'b0 ;
  assign n25604 = n3859 & n12884 ;
  assign n25605 = n25604 ^ n1257 ^ 1'b0 ;
  assign n25606 = x216 & n8800 ;
  assign n25607 = ~n20702 & n25606 ;
  assign n25608 = ~n2459 & n3674 ;
  assign n25609 = n4835 & n25608 ;
  assign n25610 = ( n8538 & ~n23473 ) | ( n8538 & n25609 ) | ( ~n23473 & n25609 ) ;
  assign n25611 = n25610 ^ n18620 ^ 1'b0 ;
  assign n25612 = n7517 ^ n699 ^ 1'b0 ;
  assign n25613 = ( n298 & ~n1108 ) | ( n298 & n5579 ) | ( ~n1108 & n5579 ) ;
  assign n25614 = n13994 & n22881 ;
  assign n25615 = n24279 | n25614 ;
  assign n25616 = n25615 ^ n11448 ^ 1'b0 ;
  assign n25617 = ~n5109 & n25616 ;
  assign n25618 = n10644 ^ n4433 ^ n779 ;
  assign n25623 = n19614 ^ n2454 ^ 1'b0 ;
  assign n25624 = n25623 ^ n8628 ^ 1'b0 ;
  assign n25619 = n2424 | n4329 ;
  assign n25620 = n25619 ^ n9557 ^ 1'b0 ;
  assign n25621 = n22100 ^ n12528 ^ n11227 ;
  assign n25622 = n25620 & n25621 ;
  assign n25625 = n25624 ^ n25622 ^ n11312 ;
  assign n25626 = ( n7145 & n10114 ) | ( n7145 & n13378 ) | ( n10114 & n13378 ) ;
  assign n25627 = ( n453 & ~n9212 ) | ( n453 & n11718 ) | ( ~n9212 & n11718 ) ;
  assign n25628 = n10287 | n10796 ;
  assign n25629 = n25628 ^ n6500 ^ 1'b0 ;
  assign n25630 = n25629 ^ n19445 ^ 1'b0 ;
  assign n25631 = ~n13634 & n25630 ;
  assign n25632 = n25631 ^ n19568 ^ x231 ;
  assign n25633 = ( ~n6063 & n6918 ) | ( ~n6063 & n25503 ) | ( n6918 & n25503 ) ;
  assign n25634 = ( n18699 & n25632 ) | ( n18699 & n25633 ) | ( n25632 & n25633 ) ;
  assign n25635 = ( n3325 & n4751 ) | ( n3325 & ~n24155 ) | ( n4751 & ~n24155 ) ;
  assign n25636 = n25635 ^ n12210 ^ 1'b0 ;
  assign n25640 = n15456 ^ x181 ^ 1'b0 ;
  assign n25638 = n5866 & ~n8889 ;
  assign n25639 = ~n2995 & n25638 ;
  assign n25637 = n23567 ^ n22003 ^ n973 ;
  assign n25641 = n25640 ^ n25639 ^ n25637 ;
  assign n25642 = ( n12097 & n23270 ) | ( n12097 & ~n25641 ) | ( n23270 & ~n25641 ) ;
  assign n25643 = n25636 | n25642 ;
  assign n25644 = n18684 ^ n5837 ^ n516 ;
  assign n25645 = n529 & ~n8223 ;
  assign n25646 = n25645 ^ n25222 ^ 1'b0 ;
  assign n25647 = ~n17937 & n25646 ;
  assign n25648 = n25647 ^ n4836 ^ 1'b0 ;
  assign n25649 = ( ~n4682 & n11692 ) | ( ~n4682 & n13333 ) | ( n11692 & n13333 ) ;
  assign n25650 = n25649 ^ n6898 ^ n1748 ;
  assign n25651 = n25650 ^ n19213 ^ n11969 ;
  assign n25652 = n10318 ^ n2004 ^ 1'b0 ;
  assign n25653 = n1345 | n25652 ;
  assign n25654 = n15721 & ~n25653 ;
  assign n25655 = n380 ^ x160 ^ 1'b0 ;
  assign n25656 = ( n16312 & n25654 ) | ( n16312 & ~n25655 ) | ( n25654 & ~n25655 ) ;
  assign n25657 = n16054 | n20870 ;
  assign n25658 = n25657 ^ n21040 ^ 1'b0 ;
  assign n25663 = ( n1109 & n2156 ) | ( n1109 & ~n4090 ) | ( n2156 & ~n4090 ) ;
  assign n25659 = n20949 & n24675 ;
  assign n25660 = n7954 & n25659 ;
  assign n25661 = n14336 & ~n25660 ;
  assign n25662 = n25661 ^ n837 ^ 1'b0 ;
  assign n25664 = n25663 ^ n25662 ^ 1'b0 ;
  assign n25665 = ( n2410 & n13756 ) | ( n2410 & ~n17902 ) | ( n13756 & ~n17902 ) ;
  assign n25666 = n25665 ^ n10766 ^ 1'b0 ;
  assign n25667 = n20138 ^ n13895 ^ n8599 ;
  assign n25668 = ( n1851 & n8648 ) | ( n1851 & n25667 ) | ( n8648 & n25667 ) ;
  assign n25669 = n1398 | n19027 ;
  assign n25670 = n11667 | n25669 ;
  assign n25671 = n9767 ^ n6394 ^ n2230 ;
  assign n25672 = ( n10127 & n11412 ) | ( n10127 & ~n25671 ) | ( n11412 & ~n25671 ) ;
  assign n25676 = n3942 & ~n4942 ;
  assign n25677 = n9904 & n25676 ;
  assign n25678 = ( n557 & n10155 ) | ( n557 & ~n25677 ) | ( n10155 & ~n25677 ) ;
  assign n25673 = n16057 ^ n9577 ^ 1'b0 ;
  assign n25674 = n20249 & n25673 ;
  assign n25675 = n12629 | n25674 ;
  assign n25679 = n25678 ^ n25675 ^ 1'b0 ;
  assign n25680 = n17591 ^ n13759 ^ n732 ;
  assign n25681 = ( n1554 & n10004 ) | ( n1554 & n11052 ) | ( n10004 & n11052 ) ;
  assign n25682 = ( ~n17346 & n22073 ) | ( ~n17346 & n25681 ) | ( n22073 & n25681 ) ;
  assign n25683 = n25682 ^ n7629 ^ 1'b0 ;
  assign n25684 = n3119 | n25683 ;
  assign n25685 = n20466 ^ n19190 ^ n8855 ;
  assign n25686 = ( n2704 & ~n21185 ) | ( n2704 & n23455 ) | ( ~n21185 & n23455 ) ;
  assign n25687 = n25686 ^ n7169 ^ 1'b0 ;
  assign n25688 = n25685 | n25687 ;
  assign n25689 = n13755 & ~n16081 ;
  assign n25690 = n25689 ^ n16595 ^ 1'b0 ;
  assign n25691 = ( n10620 & n20368 ) | ( n10620 & ~n25690 ) | ( n20368 & ~n25690 ) ;
  assign n25692 = n1422 ^ n1195 ^ 1'b0 ;
  assign n25693 = ( n2251 & n7222 ) | ( n2251 & n22233 ) | ( n7222 & n22233 ) ;
  assign n25694 = n10219 & n25693 ;
  assign n25695 = n10187 ^ n9663 ^ 1'b0 ;
  assign n25696 = ~n25694 & n25695 ;
  assign n25699 = n3280 ^ n687 ^ x47 ;
  assign n25698 = ( n3049 & n13617 ) | ( n3049 & ~n23069 ) | ( n13617 & ~n23069 ) ;
  assign n25700 = n25699 ^ n25698 ^ 1'b0 ;
  assign n25701 = ~n15280 & n25700 ;
  assign n25697 = n12526 ^ n2143 ^ 1'b0 ;
  assign n25702 = n25701 ^ n25697 ^ n4062 ;
  assign n25703 = n10604 ^ n3804 ^ 1'b0 ;
  assign n25704 = ~n9099 & n25703 ;
  assign n25705 = n23145 & n25704 ;
  assign n25706 = n20915 ^ n16119 ^ n12781 ;
  assign n25707 = n25706 ^ n23772 ^ n10996 ;
  assign n25708 = n7125 ^ n4703 ^ 1'b0 ;
  assign n25709 = ~n12848 & n25708 ;
  assign n25712 = n24357 ^ n11831 ^ n1830 ;
  assign n25713 = n8561 & ~n25712 ;
  assign n25711 = ( n3341 & n15358 ) | ( n3341 & ~n23452 ) | ( n15358 & ~n23452 ) ;
  assign n25710 = ( ~n9651 & n14095 ) | ( ~n9651 & n18684 ) | ( n14095 & n18684 ) ;
  assign n25714 = n25713 ^ n25711 ^ n25710 ;
  assign n25715 = n25709 & n25714 ;
  assign n25716 = ( n3164 & n13661 ) | ( n3164 & n16487 ) | ( n13661 & n16487 ) ;
  assign n25717 = n25716 ^ n18188 ^ n11390 ;
  assign n25718 = n21023 ^ n10394 ^ n4460 ;
  assign n25719 = n10040 ^ n6495 ^ n4320 ;
  assign n25720 = n18200 & ~n25719 ;
  assign n25721 = n25720 ^ n6249 ^ 1'b0 ;
  assign n25722 = ~n3630 & n25721 ;
  assign n25723 = n4802 & n25722 ;
  assign n25724 = n16828 & n18117 ;
  assign n25725 = n20630 ^ n3309 ^ x241 ;
  assign n25726 = n15615 ^ n1865 ^ 1'b0 ;
  assign n25727 = n3510 & n25726 ;
  assign n25728 = ( ~n6149 & n8544 ) | ( ~n6149 & n25727 ) | ( n8544 & n25727 ) ;
  assign n25729 = n25728 ^ n15025 ^ n1074 ;
  assign n25730 = n25729 ^ n13348 ^ n2064 ;
  assign n25731 = n25730 ^ n13867 ^ 1'b0 ;
  assign n25733 = n4744 & n9398 ;
  assign n25734 = n25733 ^ n12970 ^ 1'b0 ;
  assign n25732 = x127 & ~n12120 ;
  assign n25735 = n25734 ^ n25732 ^ 1'b0 ;
  assign n25736 = n1290 | n25735 ;
  assign n25737 = n22002 | n25736 ;
  assign n25738 = ~n6019 & n14209 ;
  assign n25739 = n19936 ^ n9873 ^ n3139 ;
  assign n25740 = n14160 ^ n12012 ^ n7191 ;
  assign n25741 = ( n25738 & n25739 ) | ( n25738 & n25740 ) | ( n25739 & n25740 ) ;
  assign n25742 = ( ~n2706 & n9067 ) | ( ~n2706 & n25741 ) | ( n9067 & n25741 ) ;
  assign n25743 = n5902 & ~n9103 ;
  assign n25744 = n25743 ^ n9775 ^ 1'b0 ;
  assign n25745 = n5552 & n21316 ;
  assign n25746 = ~n3285 & n25745 ;
  assign n25747 = ( n20927 & n25744 ) | ( n20927 & n25746 ) | ( n25744 & n25746 ) ;
  assign n25748 = n12646 ^ n6023 ^ n3738 ;
  assign n25749 = n5701 & ~n9864 ;
  assign n25750 = n25749 ^ n13078 ^ 1'b0 ;
  assign n25755 = n534 & n15204 ;
  assign n25756 = n25755 ^ n13304 ^ n3630 ;
  assign n25757 = n25756 ^ n7456 ^ n5374 ;
  assign n25751 = n16068 ^ n12035 ^ 1'b0 ;
  assign n25752 = ~n13691 & n25751 ;
  assign n25753 = n25752 ^ n10425 ^ 1'b0 ;
  assign n25754 = n16270 & n25753 ;
  assign n25758 = n25757 ^ n25754 ^ n14189 ;
  assign n25759 = n18909 ^ n18456 ^ n10093 ;
  assign n25760 = n3567 | n23622 ;
  assign n25761 = n23764 ^ n7739 ^ 1'b0 ;
  assign n25762 = n5416 | n25761 ;
  assign n25767 = n15424 ^ n7071 ^ n6285 ;
  assign n25763 = ~n3223 & n9808 ;
  assign n25764 = ~n13061 & n25763 ;
  assign n25765 = n25764 ^ n20597 ^ 1'b0 ;
  assign n25766 = n22134 | n25765 ;
  assign n25768 = n25767 ^ n25766 ^ 1'b0 ;
  assign n25769 = ( n6300 & ~n11384 ) | ( n6300 & n14116 ) | ( ~n11384 & n14116 ) ;
  assign n25770 = n25769 ^ n2981 ^ 1'b0 ;
  assign n25771 = n19205 ^ n14602 ^ n14340 ;
  assign n25772 = ( n9311 & ~n15025 ) | ( n9311 & n17902 ) | ( ~n15025 & n17902 ) ;
  assign n25773 = ( n12768 & n14478 ) | ( n12768 & ~n20244 ) | ( n14478 & ~n20244 ) ;
  assign n25774 = n25773 ^ n13086 ^ 1'b0 ;
  assign n25775 = n25772 & ~n25774 ;
  assign n25776 = n24108 & n25775 ;
  assign n25777 = n24849 ^ n10967 ^ n5335 ;
  assign n25778 = ( n12661 & n12876 ) | ( n12661 & n23375 ) | ( n12876 & n23375 ) ;
  assign n25779 = ( n2853 & n17868 ) | ( n2853 & n25778 ) | ( n17868 & n25778 ) ;
  assign n25780 = ( ~n1339 & n3301 ) | ( ~n1339 & n18982 ) | ( n3301 & n18982 ) ;
  assign n25781 = ( ~n8686 & n22130 ) | ( ~n8686 & n25780 ) | ( n22130 & n25780 ) ;
  assign n25782 = ~n3519 & n16598 ;
  assign n25783 = n4145 & n10801 ;
  assign n25785 = n17849 ^ n9000 ^ n6005 ;
  assign n25784 = n10611 | n15696 ;
  assign n25786 = n25785 ^ n25784 ^ 1'b0 ;
  assign n25787 = n11061 ^ n10726 ^ 1'b0 ;
  assign n25788 = n14001 ^ n6546 ^ n4926 ;
  assign n25789 = n25787 | n25788 ;
  assign n25790 = n25789 ^ n17265 ^ 1'b0 ;
  assign n25791 = n10766 ^ n9490 ^ 1'b0 ;
  assign n25792 = ~n7454 & n25791 ;
  assign n25793 = n9891 & ~n25792 ;
  assign n25794 = ~n23744 & n25420 ;
  assign n25795 = n6821 ^ n5792 ^ n4593 ;
  assign n25796 = ( n11916 & ~n23006 ) | ( n11916 & n25795 ) | ( ~n23006 & n25795 ) ;
  assign n25797 = n24920 ^ n7434 ^ 1'b0 ;
  assign n25798 = ~n22969 & n25797 ;
  assign n25799 = ( n1896 & n7679 ) | ( n1896 & n25798 ) | ( n7679 & n25798 ) ;
  assign n25803 = n17300 ^ n9074 ^ n5928 ;
  assign n25800 = n14598 & ~n23978 ;
  assign n25801 = n25800 ^ n22637 ^ 1'b0 ;
  assign n25802 = n5271 | n25801 ;
  assign n25804 = n25803 ^ n25802 ^ 1'b0 ;
  assign n25805 = n21048 ^ n4002 ^ 1'b0 ;
  assign n25806 = ( n7667 & n21772 ) | ( n7667 & n25805 ) | ( n21772 & n25805 ) ;
  assign n25807 = n14687 | n25806 ;
  assign n25808 = n11087 | n25807 ;
  assign n25813 = n12922 ^ n11745 ^ n4332 ;
  assign n25814 = ( x246 & n9601 ) | ( x246 & ~n25813 ) | ( n9601 & ~n25813 ) ;
  assign n25815 = x225 & n25814 ;
  assign n25816 = n19369 & n25815 ;
  assign n25811 = n12293 ^ n548 ^ 1'b0 ;
  assign n25809 = n23878 ^ n9428 ^ n7779 ;
  assign n25810 = ( n13999 & n21559 ) | ( n13999 & n25809 ) | ( n21559 & n25809 ) ;
  assign n25812 = n25811 ^ n25810 ^ n14348 ;
  assign n25817 = n25816 ^ n25812 ^ n6295 ;
  assign n25818 = n16701 ^ n11141 ^ n4729 ;
  assign n25819 = ( ~n10124 & n19104 ) | ( ~n10124 & n25818 ) | ( n19104 & n25818 ) ;
  assign n25820 = ( n6226 & n6850 ) | ( n6226 & n7692 ) | ( n6850 & n7692 ) ;
  assign n25821 = n4541 & n25820 ;
  assign n25822 = n25821 ^ n5189 ^ 1'b0 ;
  assign n25823 = n25819 & ~n25822 ;
  assign n25824 = ( n466 & n18584 ) | ( n466 & n25823 ) | ( n18584 & n25823 ) ;
  assign n25825 = n21198 ^ n7537 ^ n3345 ;
  assign n25826 = ( n7594 & ~n18994 ) | ( n7594 & n25825 ) | ( ~n18994 & n25825 ) ;
  assign n25830 = n5202 & n22287 ;
  assign n25831 = n25685 & n25830 ;
  assign n25827 = n13849 ^ n352 ^ 1'b0 ;
  assign n25828 = n6402 & ~n17552 ;
  assign n25829 = n25827 & n25828 ;
  assign n25832 = n25831 ^ n25829 ^ n7871 ;
  assign n25833 = n9526 ^ n7442 ^ x173 ;
  assign n25834 = n7659 & ~n20747 ;
  assign n25835 = ( n14657 & ~n18565 ) | ( n14657 & n25834 ) | ( ~n18565 & n25834 ) ;
  assign n25836 = n11286 | n25835 ;
  assign n25837 = ( n25832 & ~n25833 ) | ( n25832 & n25836 ) | ( ~n25833 & n25836 ) ;
  assign n25838 = n7780 ^ n7770 ^ n1507 ;
  assign n25839 = n1392 & n24070 ;
  assign n25840 = n25838 & n25839 ;
  assign n25841 = n2859 | n7761 ;
  assign n25842 = n25841 ^ n20083 ^ 1'b0 ;
  assign n25843 = ( ~n2644 & n8846 ) | ( ~n2644 & n16197 ) | ( n8846 & n16197 ) ;
  assign n25844 = n21319 ^ n20575 ^ n1949 ;
  assign n25845 = n7007 ^ n6759 ^ 1'b0 ;
  assign n25846 = ( ~n8804 & n14761 ) | ( ~n8804 & n25845 ) | ( n14761 & n25845 ) ;
  assign n25847 = ( ~n4102 & n9884 ) | ( ~n4102 & n12101 ) | ( n9884 & n12101 ) ;
  assign n25848 = n6480 ^ n6372 ^ x159 ;
  assign n25849 = ( ~n21713 & n25847 ) | ( ~n21713 & n25848 ) | ( n25847 & n25848 ) ;
  assign n25850 = ( ~n25844 & n25846 ) | ( ~n25844 & n25849 ) | ( n25846 & n25849 ) ;
  assign n25851 = n16970 ^ n13432 ^ 1'b0 ;
  assign n25852 = ~n4925 & n9252 ;
  assign n25853 = n25852 ^ n1550 ^ 1'b0 ;
  assign n25854 = n25853 ^ n15908 ^ n11892 ;
  assign n25855 = n25854 ^ n4512 ^ 1'b0 ;
  assign n25856 = n25855 ^ n5331 ^ 1'b0 ;
  assign n25857 = n24236 ^ n17082 ^ n6867 ;
  assign n25858 = ( n9062 & ~n11577 ) | ( n9062 & n25060 ) | ( ~n11577 & n25060 ) ;
  assign n25859 = n25858 ^ n24106 ^ n22561 ;
  assign n25860 = n2621 ^ n2447 ^ 1'b0 ;
  assign n25861 = ~n23995 & n25860 ;
  assign n25862 = n18660 & n25861 ;
  assign n25863 = ~n973 & n18269 ;
  assign n25864 = n25863 ^ n6901 ^ 1'b0 ;
  assign n25865 = ( n24043 & ~n25862 ) | ( n24043 & n25864 ) | ( ~n25862 & n25864 ) ;
  assign n25866 = n5503 & ~n7196 ;
  assign n25867 = ( n2515 & n9292 ) | ( n2515 & n10609 ) | ( n9292 & n10609 ) ;
  assign n25868 = n25867 ^ n13883 ^ n5489 ;
  assign n25869 = n8617 ^ n4705 ^ 1'b0 ;
  assign n25870 = n25869 ^ n21354 ^ n6017 ;
  assign n25871 = ~x14 & n4165 ;
  assign n25872 = ( ~n2819 & n6314 ) | ( ~n2819 & n25871 ) | ( n6314 & n25871 ) ;
  assign n25873 = ( n2348 & n12101 ) | ( n2348 & ~n14931 ) | ( n12101 & ~n14931 ) ;
  assign n25874 = ( n25870 & n25872 ) | ( n25870 & ~n25873 ) | ( n25872 & ~n25873 ) ;
  assign n25876 = n22230 ^ n15804 ^ n7450 ;
  assign n25875 = n9295 & n16397 ;
  assign n25877 = n25876 ^ n25875 ^ 1'b0 ;
  assign n25878 = ( n4895 & n16712 ) | ( n4895 & n25877 ) | ( n16712 & n25877 ) ;
  assign n25879 = n1085 & n25878 ;
  assign n25880 = n10698 ^ n315 ^ 1'b0 ;
  assign n25881 = ~n25879 & n25880 ;
  assign n25882 = ( n1087 & n4319 ) | ( n1087 & n8961 ) | ( n4319 & n8961 ) ;
  assign n25883 = ( n2176 & n5383 ) | ( n2176 & ~n25882 ) | ( n5383 & ~n25882 ) ;
  assign n25884 = n25883 ^ n13305 ^ 1'b0 ;
  assign n25885 = n4363 | n25884 ;
  assign n25892 = ~n13732 & n15251 ;
  assign n25889 = ( n5833 & n10691 ) | ( n5833 & n14420 ) | ( n10691 & n14420 ) ;
  assign n25890 = n25889 ^ n10870 ^ 1'b0 ;
  assign n25891 = n3781 | n25890 ;
  assign n25886 = ( n6581 & n10460 ) | ( n6581 & ~n17476 ) | ( n10460 & ~n17476 ) ;
  assign n25887 = n3089 & ~n25886 ;
  assign n25888 = n25887 ^ n22756 ^ n9296 ;
  assign n25893 = n25892 ^ n25891 ^ n25888 ;
  assign n25894 = n12992 & ~n16111 ;
  assign n25895 = ( ~n5159 & n15419 ) | ( ~n5159 & n25894 ) | ( n15419 & n25894 ) ;
  assign n25896 = n7292 | n19448 ;
  assign n25897 = ( ~n7180 & n14410 ) | ( ~n7180 & n20870 ) | ( n14410 & n20870 ) ;
  assign n25898 = ~n25896 & n25897 ;
  assign n25899 = n8541 & ~n15301 ;
  assign n25900 = ( n2916 & n9123 ) | ( n2916 & n9369 ) | ( n9123 & n9369 ) ;
  assign n25901 = n2980 | n3019 ;
  assign n25902 = ~n25900 & n25901 ;
  assign n25903 = n25902 ^ n14062 ^ 1'b0 ;
  assign n25905 = ~n11318 & n13504 ;
  assign n25906 = ~n8878 & n25905 ;
  assign n25904 = n1604 & n4282 ;
  assign n25907 = n25906 ^ n25904 ^ 1'b0 ;
  assign n25908 = ( ~n2182 & n2747 ) | ( ~n2182 & n7100 ) | ( n2747 & n7100 ) ;
  assign n25909 = n20045 | n25908 ;
  assign n25910 = n9765 ^ n4764 ^ n2473 ;
  assign n25911 = n5418 | n24850 ;
  assign n25912 = ( ~n10267 & n14657 ) | ( ~n10267 & n18477 ) | ( n14657 & n18477 ) ;
  assign n25913 = n25912 ^ n3108 ^ n1694 ;
  assign n25914 = n7905 | n14558 ;
  assign n25915 = ( n2913 & n9947 ) | ( n2913 & n19130 ) | ( n9947 & n19130 ) ;
  assign n25916 = ( n22328 & ~n25914 ) | ( n22328 & n25915 ) | ( ~n25914 & n25915 ) ;
  assign n25917 = ~n4026 & n13722 ;
  assign n25918 = n25917 ^ n17756 ^ n6760 ;
  assign n25919 = ( n16732 & ~n25916 ) | ( n16732 & n25918 ) | ( ~n25916 & n25918 ) ;
  assign n25920 = n12414 ^ n12368 ^ 1'b0 ;
  assign n25921 = ~n22972 & n25920 ;
  assign n25922 = n25921 ^ n9951 ^ 1'b0 ;
  assign n25923 = ~n24502 & n24936 ;
  assign n25924 = n25923 ^ n2547 ^ 1'b0 ;
  assign n25925 = ( n7926 & n18101 ) | ( n7926 & n19345 ) | ( n18101 & n19345 ) ;
  assign n25926 = n25925 ^ n11959 ^ 1'b0 ;
  assign n25927 = n7722 | n25926 ;
  assign n25928 = n15313 ^ n607 ^ 1'b0 ;
  assign n25929 = n16230 & ~n25928 ;
  assign n25930 = n25929 ^ n20285 ^ 1'b0 ;
  assign n25931 = n15300 ^ n8683 ^ n6030 ;
  assign n25932 = ( ~n14488 & n25930 ) | ( ~n14488 & n25931 ) | ( n25930 & n25931 ) ;
  assign n25933 = n20047 ^ n8232 ^ n5224 ;
  assign n25934 = ( ~n11060 & n14878 ) | ( ~n11060 & n25933 ) | ( n14878 & n25933 ) ;
  assign n25935 = n4265 | n22416 ;
  assign n25936 = n25935 ^ n11301 ^ 1'b0 ;
  assign n25937 = ( n3920 & n5014 ) | ( n3920 & ~n25936 ) | ( n5014 & ~n25936 ) ;
  assign n25938 = ( n13170 & ~n25787 ) | ( n13170 & n25937 ) | ( ~n25787 & n25937 ) ;
  assign n25940 = ( ~n3937 & n5407 ) | ( ~n3937 & n15457 ) | ( n5407 & n15457 ) ;
  assign n25939 = n13759 ^ n11957 ^ n11351 ;
  assign n25941 = n25940 ^ n25939 ^ 1'b0 ;
  assign n25942 = n2835 ^ n2502 ^ 1'b0 ;
  assign n25943 = ~x23 & n25942 ;
  assign n25947 = n5411 & ~n10502 ;
  assign n25948 = ~n10841 & n25947 ;
  assign n25944 = ~n5917 & n18790 ;
  assign n25945 = n14437 & n25944 ;
  assign n25946 = n25945 ^ n17256 ^ n6343 ;
  assign n25949 = n25948 ^ n25946 ^ 1'b0 ;
  assign n25950 = ( ~n16839 & n25943 ) | ( ~n16839 & n25949 ) | ( n25943 & n25949 ) ;
  assign n25951 = ( ~n20042 & n25941 ) | ( ~n20042 & n25950 ) | ( n25941 & n25950 ) ;
  assign n25952 = x251 & ~n20566 ;
  assign n25953 = n25952 ^ n10339 ^ 1'b0 ;
  assign n25956 = n11385 ^ n9851 ^ 1'b0 ;
  assign n25957 = ( ~n834 & n19536 ) | ( ~n834 & n25956 ) | ( n19536 & n25956 ) ;
  assign n25954 = ( n1170 & ~n11817 ) | ( n1170 & n22461 ) | ( ~n11817 & n22461 ) ;
  assign n25955 = n25954 ^ n11965 ^ n5149 ;
  assign n25958 = n25957 ^ n25955 ^ n2774 ;
  assign n25959 = n6628 ^ n2724 ^ n2649 ;
  assign n25960 = n4502 & n5888 ;
  assign n25961 = n3800 & ~n4578 ;
  assign n25962 = n25961 ^ n6859 ^ n3669 ;
  assign n25963 = n25960 & ~n25962 ;
  assign n25964 = n15196 ^ x49 ^ 1'b0 ;
  assign n25965 = ~n25963 & n25964 ;
  assign n25966 = ~n22532 & n25965 ;
  assign n25967 = n25959 & n25966 ;
  assign n25968 = n25967 ^ n20726 ^ 1'b0 ;
  assign n25969 = ~n11524 & n17395 ;
  assign n25970 = n25969 ^ n20782 ^ n5216 ;
  assign n25971 = n17986 ^ n5368 ^ n727 ;
  assign n25972 = ( n9333 & n12812 ) | ( n9333 & n16400 ) | ( n12812 & n16400 ) ;
  assign n25973 = ( n8047 & ~n18198 ) | ( n8047 & n25972 ) | ( ~n18198 & n25972 ) ;
  assign n25974 = n8379 ^ n4665 ^ 1'b0 ;
  assign n25975 = n25974 ^ n10065 ^ 1'b0 ;
  assign n25976 = n8992 | n25975 ;
  assign n25977 = n25976 ^ n15154 ^ n14512 ;
  assign n25978 = n3581 ^ n1928 ^ n1813 ;
  assign n25979 = n8628 & n25978 ;
  assign n25980 = n1883 & ~n8267 ;
  assign n25981 = ~n10574 & n25980 ;
  assign n25982 = n25981 ^ n3925 ^ n1610 ;
  assign n25983 = ( ~n7736 & n10530 ) | ( ~n7736 & n14611 ) | ( n10530 & n14611 ) ;
  assign n25984 = ( n1025 & n3781 ) | ( n1025 & n9825 ) | ( n3781 & n9825 ) ;
  assign n25985 = n11427 ^ n6702 ^ n6126 ;
  assign n25986 = ( ~n25983 & n25984 ) | ( ~n25983 & n25985 ) | ( n25984 & n25985 ) ;
  assign n25987 = n25986 ^ n10477 ^ n5710 ;
  assign n25988 = n17431 ^ n9899 ^ n6459 ;
  assign n25989 = n11189 | n25988 ;
  assign n25990 = ( n22932 & ~n25861 ) | ( n22932 & n25989 ) | ( ~n25861 & n25989 ) ;
  assign n25992 = ~n2687 & n7285 ;
  assign n25993 = n25992 ^ n5633 ^ 1'b0 ;
  assign n25994 = n25993 ^ n2203 ^ 1'b0 ;
  assign n25995 = n15056 & n25994 ;
  assign n25996 = n2759 & n25995 ;
  assign n25991 = n12697 & ~n14696 ;
  assign n25997 = n25996 ^ n25991 ^ n6470 ;
  assign n25998 = n6982 ^ n1768 ^ n801 ;
  assign n25999 = ( ~n22515 & n23388 ) | ( ~n22515 & n25998 ) | ( n23388 & n25998 ) ;
  assign n26005 = ( n4072 & n4598 ) | ( n4072 & n7264 ) | ( n4598 & n7264 ) ;
  assign n26000 = n24028 ^ n16278 ^ n5657 ;
  assign n26001 = n13712 | n26000 ;
  assign n26002 = ~n9518 & n26001 ;
  assign n26003 = n26002 ^ n263 ^ 1'b0 ;
  assign n26004 = n7094 & ~n26003 ;
  assign n26006 = n26005 ^ n26004 ^ 1'b0 ;
  assign n26007 = ( ~n4826 & n6054 ) | ( ~n4826 & n7989 ) | ( n6054 & n7989 ) ;
  assign n26008 = n19110 ^ n4247 ^ 1'b0 ;
  assign n26009 = ~n26007 & n26008 ;
  assign n26013 = n7220 ^ n6579 ^ n1111 ;
  assign n26014 = ( n3999 & ~n23679 ) | ( n3999 & n26013 ) | ( ~n23679 & n26013 ) ;
  assign n26010 = n16184 ^ n15600 ^ 1'b0 ;
  assign n26011 = n14943 & ~n26010 ;
  assign n26012 = n26011 ^ n12085 ^ 1'b0 ;
  assign n26015 = n26014 ^ n26012 ^ n18167 ;
  assign n26016 = ( n25134 & n26009 ) | ( n25134 & n26015 ) | ( n26009 & n26015 ) ;
  assign n26017 = n18848 | n23633 ;
  assign n26018 = n26017 ^ n7586 ^ 1'b0 ;
  assign n26019 = n26018 ^ n5434 ^ 1'b0 ;
  assign n26020 = n10498 ^ n8641 ^ 1'b0 ;
  assign n26021 = ~n2129 & n26020 ;
  assign n26022 = n9820 & n26021 ;
  assign n26023 = n11074 & ~n26022 ;
  assign n26024 = n26023 ^ n12453 ^ n4472 ;
  assign n26025 = n12554 ^ n4492 ^ 1'b0 ;
  assign n26026 = ~n16540 & n26025 ;
  assign n26027 = ( n6447 & n15337 ) | ( n6447 & ~n26026 ) | ( n15337 & ~n26026 ) ;
  assign n26028 = n26027 ^ n18865 ^ n17144 ;
  assign n26029 = ( n6784 & ~n13730 ) | ( n6784 & n25867 ) | ( ~n13730 & n25867 ) ;
  assign n26032 = ( ~n1588 & n18922 ) | ( ~n1588 & n22725 ) | ( n18922 & n22725 ) ;
  assign n26030 = n4138 & n23157 ;
  assign n26031 = n1222 & n26030 ;
  assign n26033 = n26032 ^ n26031 ^ n2504 ;
  assign n26037 = n2380 | n13420 ;
  assign n26038 = n26037 ^ n11492 ^ 1'b0 ;
  assign n26034 = n5707 ^ n4754 ^ n1413 ;
  assign n26035 = ( n586 & ~n1633 ) | ( n586 & n25481 ) | ( ~n1633 & n25481 ) ;
  assign n26036 = n26034 & n26035 ;
  assign n26039 = n26038 ^ n26036 ^ 1'b0 ;
  assign n26040 = n5757 | n10913 ;
  assign n26041 = n7229 & n15444 ;
  assign n26042 = ( ~n5812 & n12860 ) | ( ~n5812 & n26041 ) | ( n12860 & n26041 ) ;
  assign n26043 = n15361 | n23125 ;
  assign n26044 = n26043 ^ n11410 ^ 1'b0 ;
  assign n26045 = ( n21247 & n26042 ) | ( n21247 & ~n26044 ) | ( n26042 & ~n26044 ) ;
  assign n26046 = ( n14487 & ~n19420 ) | ( n14487 & n20148 ) | ( ~n19420 & n20148 ) ;
  assign n26047 = ( n3290 & ~n9501 ) | ( n3290 & n26046 ) | ( ~n9501 & n26046 ) ;
  assign n26048 = n26047 ^ n22899 ^ 1'b0 ;
  assign n26049 = ( ~n4201 & n23979 ) | ( ~n4201 & n26048 ) | ( n23979 & n26048 ) ;
  assign n26050 = n8877 ^ n8731 ^ 1'b0 ;
  assign n26051 = n5403 & ~n26050 ;
  assign n26052 = ~n1797 & n26051 ;
  assign n26053 = n26052 ^ n20479 ^ 1'b0 ;
  assign n26055 = n6648 ^ n3223 ^ 1'b0 ;
  assign n26056 = n26055 ^ n3758 ^ 1'b0 ;
  assign n26054 = n480 & ~n674 ;
  assign n26057 = n26056 ^ n26054 ^ 1'b0 ;
  assign n26058 = n18518 & n26057 ;
  assign n26059 = n5567 & n26058 ;
  assign n26060 = n26059 ^ n11693 ^ 1'b0 ;
  assign n26061 = n6615 | n26060 ;
  assign n26062 = n12915 ^ n5216 ^ 1'b0 ;
  assign n26063 = n2174 | n14240 ;
  assign n26064 = n9879 | n26063 ;
  assign n26065 = ( n7573 & n26062 ) | ( n7573 & ~n26064 ) | ( n26062 & ~n26064 ) ;
  assign n26066 = n23657 ^ n9363 ^ n8769 ;
  assign n26067 = ( n6106 & n9570 ) | ( n6106 & ~n26066 ) | ( n9570 & ~n26066 ) ;
  assign n26068 = ( ~n5249 & n13144 ) | ( ~n5249 & n26067 ) | ( n13144 & n26067 ) ;
  assign n26072 = n9170 ^ n658 ^ x81 ;
  assign n26069 = n4011 ^ n524 ^ 1'b0 ;
  assign n26070 = n10790 & ~n11586 ;
  assign n26071 = ( n347 & ~n26069 ) | ( n347 & n26070 ) | ( ~n26069 & n26070 ) ;
  assign n26073 = n26072 ^ n26071 ^ 1'b0 ;
  assign n26074 = n4384 & n26073 ;
  assign n26075 = ( n1124 & n10134 ) | ( n1124 & n26074 ) | ( n10134 & n26074 ) ;
  assign n26078 = n4817 & ~n6112 ;
  assign n26079 = ~n17509 & n26078 ;
  assign n26076 = n16448 ^ n10850 ^ 1'b0 ;
  assign n26077 = n26076 ^ n10656 ^ n4457 ;
  assign n26080 = n26079 ^ n26077 ^ n23239 ;
  assign n26081 = n10346 ^ n10316 ^ 1'b0 ;
  assign n26082 = n26081 ^ n16561 ^ 1'b0 ;
  assign n26083 = n4872 & n15161 ;
  assign n26084 = ~n12717 & n26083 ;
  assign n26085 = ( n4306 & ~n7730 ) | ( n4306 & n26084 ) | ( ~n7730 & n26084 ) ;
  assign n26086 = ~n16158 & n19660 ;
  assign n26087 = n26086 ^ n18839 ^ 1'b0 ;
  assign n26088 = ( n6340 & n13065 ) | ( n6340 & n26087 ) | ( n13065 & n26087 ) ;
  assign n26089 = ~n26085 & n26088 ;
  assign n26090 = n26082 & n26089 ;
  assign n26091 = n19829 ^ n5383 ^ 1'b0 ;
  assign n26092 = n25993 ^ n13738 ^ 1'b0 ;
  assign n26093 = ~n19814 & n26092 ;
  assign n26094 = n26093 ^ n16925 ^ n2214 ;
  assign n26097 = ~n2657 & n14278 ;
  assign n26098 = ( n4692 & n9344 ) | ( n4692 & n26097 ) | ( n9344 & n26097 ) ;
  assign n26095 = ~n583 & n3889 ;
  assign n26096 = n26095 ^ n13986 ^ n5044 ;
  assign n26099 = n26098 ^ n26096 ^ n18686 ;
  assign n26100 = n6461 ^ n548 ^ 1'b0 ;
  assign n26101 = n26100 ^ n16834 ^ n4781 ;
  assign n26102 = ~n17452 & n17520 ;
  assign n26103 = n26101 & n26102 ;
  assign n26104 = n26103 ^ n1920 ^ 1'b0 ;
  assign n26105 = ( n2976 & n5695 ) | ( n2976 & ~n13023 ) | ( n5695 & ~n13023 ) ;
  assign n26106 = ~n22730 & n26105 ;
  assign n26107 = ( n11093 & n26104 ) | ( n11093 & n26106 ) | ( n26104 & n26106 ) ;
  assign n26110 = n20580 & n21298 ;
  assign n26108 = ( n3936 & n13665 ) | ( n3936 & n18757 ) | ( n13665 & n18757 ) ;
  assign n26109 = ( n9658 & n22401 ) | ( n9658 & ~n26108 ) | ( n22401 & ~n26108 ) ;
  assign n26111 = n26110 ^ n26109 ^ n10825 ;
  assign n26112 = n11819 & ~n26111 ;
  assign n26113 = n26112 ^ n20029 ^ 1'b0 ;
  assign n26119 = n11051 ^ n7428 ^ n5202 ;
  assign n26114 = n17737 | n25582 ;
  assign n26115 = n19023 | n26114 ;
  assign n26116 = n11633 ^ n9067 ^ n2443 ;
  assign n26117 = ( ~n9177 & n26115 ) | ( ~n9177 & n26116 ) | ( n26115 & n26116 ) ;
  assign n26118 = ~n21463 & n26117 ;
  assign n26120 = n26119 ^ n26118 ^ 1'b0 ;
  assign n26121 = n15351 & n19723 ;
  assign n26122 = ( ~n427 & n1170 ) | ( ~n427 & n25139 ) | ( n1170 & n25139 ) ;
  assign n26123 = ~n24283 & n26122 ;
  assign n26124 = n26121 & n26123 ;
  assign n26125 = n25529 ^ n5930 ^ 1'b0 ;
  assign n26126 = n379 | n26125 ;
  assign n26129 = n10432 ^ n3198 ^ 1'b0 ;
  assign n26130 = ~n989 & n26129 ;
  assign n26131 = ( ~n5037 & n18625 ) | ( ~n5037 & n26130 ) | ( n18625 & n26130 ) ;
  assign n26132 = n1224 ^ n422 ^ 1'b0 ;
  assign n26133 = ( ~n970 & n26131 ) | ( ~n970 & n26132 ) | ( n26131 & n26132 ) ;
  assign n26134 = n26133 ^ n10525 ^ n10230 ;
  assign n26127 = n10722 ^ n6218 ^ n1366 ;
  assign n26128 = ( n10343 & n12801 ) | ( n10343 & ~n26127 ) | ( n12801 & ~n26127 ) ;
  assign n26135 = n26134 ^ n26128 ^ n21411 ;
  assign n26136 = n13410 ^ n8682 ^ 1'b0 ;
  assign n26137 = n26136 ^ n18836 ^ n8911 ;
  assign n26138 = n7585 & n26137 ;
  assign n26139 = ( n5394 & ~n6841 ) | ( n5394 & n26138 ) | ( ~n6841 & n26138 ) ;
  assign n26140 = n8860 & ~n26139 ;
  assign n26141 = n540 & ~n2479 ;
  assign n26142 = n26141 ^ n5096 ^ 1'b0 ;
  assign n26143 = n26142 ^ n14010 ^ 1'b0 ;
  assign n26144 = n1614 & n26143 ;
  assign n26145 = n1751 | n3488 ;
  assign n26146 = n10316 | n26145 ;
  assign n26147 = ( n4469 & ~n12212 ) | ( n4469 & n26146 ) | ( ~n12212 & n26146 ) ;
  assign n26148 = ( n10334 & n12535 ) | ( n10334 & ~n24241 ) | ( n12535 & ~n24241 ) ;
  assign n26149 = n19906 ^ n6624 ^ x53 ;
  assign n26150 = ( n5864 & n9429 ) | ( n5864 & n26149 ) | ( n9429 & n26149 ) ;
  assign n26151 = ( n3707 & n12855 ) | ( n3707 & ~n26150 ) | ( n12855 & ~n26150 ) ;
  assign n26152 = ~n16763 & n26151 ;
  assign n26153 = ( n6422 & n19070 ) | ( n6422 & ~n26152 ) | ( n19070 & ~n26152 ) ;
  assign n26154 = n12143 ^ n6325 ^ n4880 ;
  assign n26155 = n14595 ^ n11975 ^ n3877 ;
  assign n26156 = n5897 & n26155 ;
  assign n26157 = ~n993 & n26156 ;
  assign n26158 = n589 | n1968 ;
  assign n26159 = n2256 & ~n26158 ;
  assign n26160 = n5153 & ~n26159 ;
  assign n26161 = n7242 | n8020 ;
  assign n26162 = n26160 | n26161 ;
  assign n26163 = ~n3369 & n12864 ;
  assign n26164 = ( n5249 & n20001 ) | ( n5249 & n26163 ) | ( n20001 & n26163 ) ;
  assign n26165 = ( n7625 & n13007 ) | ( n7625 & ~n15805 ) | ( n13007 & ~n15805 ) ;
  assign n26166 = ~n24760 & n26165 ;
  assign n26167 = n486 | n20575 ;
  assign n26168 = n20612 & ~n26167 ;
  assign n26169 = ~n16188 & n24162 ;
  assign n26170 = n26168 | n26169 ;
  assign n26171 = ( x23 & n3573 ) | ( x23 & n5848 ) | ( n3573 & n5848 ) ;
  assign n26172 = n14929 | n22356 ;
  assign n26173 = n21031 | n26172 ;
  assign n26174 = ( n12550 & n26171 ) | ( n12550 & n26173 ) | ( n26171 & n26173 ) ;
  assign n26175 = ( ~n9535 & n21348 ) | ( ~n9535 & n26174 ) | ( n21348 & n26174 ) ;
  assign n26178 = n2768 & n15153 ;
  assign n26176 = n9815 ^ n7736 ^ n3384 ;
  assign n26177 = n6838 | n26176 ;
  assign n26179 = n26178 ^ n26177 ^ 1'b0 ;
  assign n26180 = n26179 ^ n12539 ^ 1'b0 ;
  assign n26181 = n6062 | n26180 ;
  assign n26182 = n3738 | n9148 ;
  assign n26183 = n26182 ^ n11085 ^ 1'b0 ;
  assign n26184 = ( n5827 & ~n6277 ) | ( n5827 & n7169 ) | ( ~n6277 & n7169 ) ;
  assign n26195 = n8571 ^ n6059 ^ 1'b0 ;
  assign n26196 = n24205 ^ n17643 ^ n13070 ;
  assign n26197 = n2336 & n26196 ;
  assign n26198 = ~n26195 & n26197 ;
  assign n26185 = n2227 ^ x10 ^ 1'b0 ;
  assign n26186 = n4582 & n26185 ;
  assign n26187 = ( ~x116 & n3072 ) | ( ~x116 & n12019 ) | ( n3072 & n12019 ) ;
  assign n26188 = ( n7086 & n22137 ) | ( n7086 & n26187 ) | ( n22137 & n26187 ) ;
  assign n26189 = n26188 ^ n24280 ^ 1'b0 ;
  assign n26190 = n16435 & n26189 ;
  assign n26191 = ( ~n1668 & n12176 ) | ( ~n1668 & n26190 ) | ( n12176 & n26190 ) ;
  assign n26192 = ( n11577 & n12581 ) | ( n11577 & n26191 ) | ( n12581 & n26191 ) ;
  assign n26193 = ( n24385 & n26186 ) | ( n24385 & n26192 ) | ( n26186 & n26192 ) ;
  assign n26194 = n26193 ^ n6073 ^ 1'b0 ;
  assign n26199 = n26198 ^ n26194 ^ 1'b0 ;
  assign n26200 = n14235 & n26199 ;
  assign n26201 = n20234 & n26200 ;
  assign n26202 = ~n26184 & n26201 ;
  assign n26203 = n9334 ^ n2113 ^ 1'b0 ;
  assign n26204 = ( ~n9496 & n11199 ) | ( ~n9496 & n26203 ) | ( n11199 & n26203 ) ;
  assign n26205 = n9473 ^ n1775 ^ 1'b0 ;
  assign n26206 = x78 & n26205 ;
  assign n26207 = n18828 ^ n2570 ^ 1'b0 ;
  assign n26208 = n26206 & ~n26207 ;
  assign n26209 = n6651 ^ n1855 ^ 1'b0 ;
  assign n26210 = n18947 & ~n26209 ;
  assign n26211 = n6808 | n26210 ;
  assign n26212 = ( n2777 & n4790 ) | ( n2777 & n19782 ) | ( n4790 & n19782 ) ;
  assign n26213 = n10712 & n21878 ;
  assign n26214 = ( n26211 & n26212 ) | ( n26211 & ~n26213 ) | ( n26212 & ~n26213 ) ;
  assign n26215 = ( n1702 & ~n17288 ) | ( n1702 & n22062 ) | ( ~n17288 & n22062 ) ;
  assign n26216 = ~n3142 & n11944 ;
  assign n26217 = n5658 & n13074 ;
  assign n26218 = n16265 & n26217 ;
  assign n26219 = ( n20651 & n26216 ) | ( n20651 & n26218 ) | ( n26216 & n26218 ) ;
  assign n26220 = ( n16296 & n23665 ) | ( n16296 & ~n26219 ) | ( n23665 & ~n26219 ) ;
  assign n26221 = n26220 ^ n8598 ^ n3605 ;
  assign n26222 = n3309 | n13303 ;
  assign n26223 = n26222 ^ n21887 ^ 1'b0 ;
  assign n26224 = n22964 ^ n17175 ^ n1175 ;
  assign n26225 = n582 & ~n21229 ;
  assign n26226 = n15634 & n26225 ;
  assign n26227 = n16065 ^ n7270 ^ n5820 ;
  assign n26229 = n7256 ^ n3027 ^ 1'b0 ;
  assign n26230 = n17262 & n26229 ;
  assign n26231 = n26230 ^ n12362 ^ 1'b0 ;
  assign n26228 = n21130 ^ n14197 ^ n4000 ;
  assign n26232 = n26231 ^ n26228 ^ n11696 ;
  assign n26233 = x113 & ~n1386 ;
  assign n26234 = n26233 ^ n1795 ^ 1'b0 ;
  assign n26235 = n24856 | n26234 ;
  assign n26236 = n10048 ^ n7926 ^ 1'b0 ;
  assign n26237 = n5475 & n26236 ;
  assign n26238 = ( ~n16795 & n22034 ) | ( ~n16795 & n26237 ) | ( n22034 & n26237 ) ;
  assign n26239 = ( ~n4380 & n11107 ) | ( ~n4380 & n24278 ) | ( n11107 & n24278 ) ;
  assign n26241 = n5637 | n7414 ;
  assign n26242 = ( n12741 & n14302 ) | ( n12741 & ~n26241 ) | ( n14302 & ~n26241 ) ;
  assign n26240 = ( ~n3196 & n17645 ) | ( ~n3196 & n24115 ) | ( n17645 & n24115 ) ;
  assign n26243 = n26242 ^ n26240 ^ n5423 ;
  assign n26244 = n13261 & n13414 ;
  assign n26245 = n26244 ^ n2552 ^ 1'b0 ;
  assign n26246 = n26245 ^ n9217 ^ n2654 ;
  assign n26247 = ( n7374 & n7671 ) | ( n7374 & ~n26246 ) | ( n7671 & ~n26246 ) ;
  assign n26248 = n7868 & ~n22369 ;
  assign n26249 = n26248 ^ n12128 ^ 1'b0 ;
  assign n26250 = ( ~x19 & n5520 ) | ( ~x19 & n13138 ) | ( n5520 & n13138 ) ;
  assign n26255 = ( n5953 & ~n12915 ) | ( n5953 & n14257 ) | ( ~n12915 & n14257 ) ;
  assign n26251 = n3444 | n4493 ;
  assign n26252 = n26251 ^ n2586 ^ 1'b0 ;
  assign n26253 = ~n22871 & n26252 ;
  assign n26254 = ~n6397 & n26253 ;
  assign n26256 = n26255 ^ n26254 ^ n25744 ;
  assign n26257 = ( n7172 & n20515 ) | ( n7172 & ~n22981 ) | ( n20515 & ~n22981 ) ;
  assign n26259 = n3397 ^ n3044 ^ n2964 ;
  assign n26260 = n26259 ^ n668 ^ 1'b0 ;
  assign n26261 = n310 | n26260 ;
  assign n26258 = n3042 & ~n17750 ;
  assign n26262 = n26261 ^ n26258 ^ 1'b0 ;
  assign n26263 = ( ~x163 & n2760 ) | ( ~x163 & n12168 ) | ( n2760 & n12168 ) ;
  assign n26264 = n17096 ^ n2832 ^ 1'b0 ;
  assign n26265 = n10915 ^ n6820 ^ n4748 ;
  assign n26267 = ( n2565 & n3663 ) | ( n2565 & ~n16168 ) | ( n3663 & ~n16168 ) ;
  assign n26266 = ( ~n1741 & n7092 ) | ( ~n1741 & n8050 ) | ( n7092 & n8050 ) ;
  assign n26268 = n26267 ^ n26266 ^ 1'b0 ;
  assign n26269 = n2452 & ~n5106 ;
  assign n26270 = ~n26268 & n26269 ;
  assign n26271 = n9839 ^ n6840 ^ 1'b0 ;
  assign n26273 = ( n787 & ~n13016 ) | ( n787 & n13080 ) | ( ~n13016 & n13080 ) ;
  assign n26272 = n18664 & n23651 ;
  assign n26274 = n26273 ^ n26272 ^ 1'b0 ;
  assign n26275 = n18963 | n26274 ;
  assign n26276 = n26275 ^ n6896 ^ 1'b0 ;
  assign n26277 = ( ~n7863 & n10307 ) | ( ~n7863 & n10880 ) | ( n10307 & n10880 ) ;
  assign n26278 = n3874 & n3890 ;
  assign n26279 = ( x105 & ~n17899 ) | ( x105 & n25077 ) | ( ~n17899 & n25077 ) ;
  assign n26280 = n26279 ^ n21543 ^ n4120 ;
  assign n26281 = n2334 & n3540 ;
  assign n26282 = n6075 & ~n26281 ;
  assign n26284 = n7544 & n7625 ;
  assign n26285 = n26284 ^ n1730 ^ 1'b0 ;
  assign n26286 = n26285 ^ n8990 ^ n1061 ;
  assign n26287 = ( n13347 & n13709 ) | ( n13347 & n26286 ) | ( n13709 & n26286 ) ;
  assign n26288 = ( ~n15240 & n21461 ) | ( ~n15240 & n26287 ) | ( n21461 & n26287 ) ;
  assign n26283 = n20886 | n24389 ;
  assign n26289 = n26288 ^ n26283 ^ 1'b0 ;
  assign n26290 = n18755 ^ n12209 ^ 1'b0 ;
  assign n26291 = ( n3332 & ~n24127 ) | ( n3332 & n26290 ) | ( ~n24127 & n26290 ) ;
  assign n26292 = n2937 & ~n8241 ;
  assign n26293 = ( n9123 & n16301 ) | ( n9123 & ~n26292 ) | ( n16301 & ~n26292 ) ;
  assign n26294 = ( ~n10658 & n26291 ) | ( ~n10658 & n26293 ) | ( n26291 & n26293 ) ;
  assign n26295 = n1883 & ~n11822 ;
  assign n26296 = n14721 ^ n5462 ^ n3191 ;
  assign n26297 = ~n1918 & n11709 ;
  assign n26298 = n10285 & ~n26297 ;
  assign n26299 = n26296 & ~n26298 ;
  assign n26300 = ~n10940 & n26299 ;
  assign n26301 = n9349 ^ n9092 ^ n7630 ;
  assign n26302 = n26301 ^ n15761 ^ n10935 ;
  assign n26303 = n25222 ^ n21342 ^ n15229 ;
  assign n26304 = n22490 ^ n16863 ^ x105 ;
  assign n26305 = n26304 ^ n9844 ^ 1'b0 ;
  assign n26306 = ( n2929 & n4314 ) | ( n2929 & ~n4923 ) | ( n4314 & ~n4923 ) ;
  assign n26307 = ( n2693 & n10672 ) | ( n2693 & ~n26306 ) | ( n10672 & ~n26306 ) ;
  assign n26308 = ( ~n645 & n3572 ) | ( ~n645 & n13244 ) | ( n3572 & n13244 ) ;
  assign n26309 = n10651 ^ n3064 ^ x240 ;
  assign n26310 = n6005 | n15207 ;
  assign n26311 = n8429 & ~n26310 ;
  assign n26312 = ( n8274 & n26309 ) | ( n8274 & n26311 ) | ( n26309 & n26311 ) ;
  assign n26313 = ( n5162 & ~n11418 ) | ( n5162 & n26312 ) | ( ~n11418 & n26312 ) ;
  assign n26314 = ( ~n26307 & n26308 ) | ( ~n26307 & n26313 ) | ( n26308 & n26313 ) ;
  assign n26315 = n12173 ^ n11626 ^ 1'b0 ;
  assign n26317 = ( n2545 & n2949 ) | ( n2545 & ~n6907 ) | ( n2949 & ~n6907 ) ;
  assign n26318 = ( n8685 & ~n20890 ) | ( n8685 & n24170 ) | ( ~n20890 & n24170 ) ;
  assign n26319 = n22515 ^ n2753 ^ 1'b0 ;
  assign n26320 = ~n26318 & n26319 ;
  assign n26321 = n26320 ^ n13162 ^ 1'b0 ;
  assign n26322 = ( n13444 & n26317 ) | ( n13444 & ~n26321 ) | ( n26317 & ~n26321 ) ;
  assign n26316 = n17861 ^ n11159 ^ 1'b0 ;
  assign n26323 = n26322 ^ n26316 ^ n676 ;
  assign n26324 = n8800 ^ n5955 ^ n2536 ;
  assign n26325 = n16635 ^ n12763 ^ n933 ;
  assign n26326 = ~n2305 & n10690 ;
  assign n26327 = n12823 ^ n4101 ^ 1'b0 ;
  assign n26328 = n26327 ^ n995 ^ 1'b0 ;
  assign n26329 = n23335 ^ n22317 ^ n15180 ;
  assign n26330 = ( n14095 & ~n26328 ) | ( n14095 & n26329 ) | ( ~n26328 & n26329 ) ;
  assign n26332 = ~n2888 & n3103 ;
  assign n26331 = ( n6666 & n6676 ) | ( n6666 & n12200 ) | ( n6676 & n12200 ) ;
  assign n26333 = n26332 ^ n26331 ^ n2106 ;
  assign n26334 = n3270 | n26333 ;
  assign n26335 = n8201 & ~n10853 ;
  assign n26336 = n4205 & ~n26335 ;
  assign n26337 = ~n16581 & n26336 ;
  assign n26338 = n8496 & ~n26337 ;
  assign n26339 = n26338 ^ n13528 ^ 1'b0 ;
  assign n26340 = ( ~n2339 & n4474 ) | ( ~n2339 & n16846 ) | ( n4474 & n16846 ) ;
  assign n26344 = ~n4059 & n6997 ;
  assign n26345 = n26344 ^ n7641 ^ 1'b0 ;
  assign n26341 = n11622 ^ n5565 ^ n2315 ;
  assign n26342 = n26341 ^ n23499 ^ 1'b0 ;
  assign n26343 = n4684 & ~n26342 ;
  assign n26346 = n26345 ^ n26343 ^ n6195 ;
  assign n26347 = ( n523 & n6208 ) | ( n523 & n18322 ) | ( n6208 & n18322 ) ;
  assign n26348 = ( n4326 & ~n13577 ) | ( n4326 & n25219 ) | ( ~n13577 & n25219 ) ;
  assign n26349 = n26348 ^ n7549 ^ n4479 ;
  assign n26350 = ( n15228 & n26347 ) | ( n15228 & n26349 ) | ( n26347 & n26349 ) ;
  assign n26351 = n12707 ^ n3207 ^ n2971 ;
  assign n26352 = ~n19596 & n26351 ;
  assign n26353 = ~n26350 & n26352 ;
  assign n26354 = ( ~n7645 & n23722 ) | ( ~n7645 & n26353 ) | ( n23722 & n26353 ) ;
  assign n26358 = n14590 ^ n13969 ^ n5988 ;
  assign n26356 = n4895 & ~n10080 ;
  assign n26357 = ~n11442 & n26356 ;
  assign n26359 = n26358 ^ n26357 ^ 1'b0 ;
  assign n26355 = n18775 ^ n15368 ^ 1'b0 ;
  assign n26360 = n26359 ^ n26355 ^ n20036 ;
  assign n26362 = n357 & n5418 ;
  assign n26363 = n2667 & n26362 ;
  assign n26361 = ( n4154 & n4249 ) | ( n4154 & n25391 ) | ( n4249 & n25391 ) ;
  assign n26364 = n26363 ^ n26361 ^ n7888 ;
  assign n26365 = n26364 ^ n14887 ^ n13774 ;
  assign n26366 = n26365 ^ n14219 ^ 1'b0 ;
  assign n26367 = n2130 & ~n26366 ;
  assign n26368 = n26367 ^ n13257 ^ n6486 ;
  assign n26376 = ~n4030 & n17058 ;
  assign n26377 = n26376 ^ n4881 ^ 1'b0 ;
  assign n26369 = n2514 ^ n2250 ^ n2145 ;
  assign n26370 = ( n1578 & n15491 ) | ( n1578 & ~n26369 ) | ( n15491 & ~n26369 ) ;
  assign n26371 = n18416 ^ n10650 ^ n3204 ;
  assign n26372 = ~n26370 & n26371 ;
  assign n26373 = n26372 ^ n8830 ^ 1'b0 ;
  assign n26374 = n21836 & n26373 ;
  assign n26375 = n26374 ^ n17142 ^ 1'b0 ;
  assign n26378 = n26377 ^ n26375 ^ n18244 ;
  assign n26379 = ~n6995 & n10574 ;
  assign n26380 = ( n2345 & n5608 ) | ( n2345 & ~n26379 ) | ( n5608 & ~n26379 ) ;
  assign n26381 = ( x83 & ~n7132 ) | ( x83 & n8965 ) | ( ~n7132 & n8965 ) ;
  assign n26382 = ~n26380 & n26381 ;
  assign n26383 = n8013 ^ n4957 ^ 1'b0 ;
  assign n26384 = n13220 & ~n26383 ;
  assign n26385 = x158 & n26384 ;
  assign n26386 = n22921 ^ n860 ^ 1'b0 ;
  assign n26387 = n8842 ^ n2867 ^ n699 ;
  assign n26388 = ( n545 & n600 ) | ( n545 & ~n12123 ) | ( n600 & ~n12123 ) ;
  assign n26389 = ~n5151 & n8242 ;
  assign n26390 = ( ~n15452 & n26388 ) | ( ~n15452 & n26389 ) | ( n26388 & n26389 ) ;
  assign n26391 = n9105 ^ n2139 ^ 1'b0 ;
  assign n26392 = n13787 ^ n5952 ^ n3571 ;
  assign n26393 = n6479 & n10335 ;
  assign n26394 = n26393 ^ n3223 ^ 1'b0 ;
  assign n26395 = n26394 ^ n16277 ^ 1'b0 ;
  assign n26396 = n16931 | n26395 ;
  assign n26397 = n11894 & ~n18820 ;
  assign n26398 = n23380 ^ n11262 ^ n10842 ;
  assign n26399 = n18242 ^ n6469 ^ 1'b0 ;
  assign n26400 = n26399 ^ n25455 ^ n2960 ;
  assign n26401 = n23140 ^ n18587 ^ n2932 ;
  assign n26402 = n22925 | n26401 ;
  assign n26403 = n2956 & n6586 ;
  assign n26404 = ~n9666 & n26403 ;
  assign n26405 = n26404 ^ n22025 ^ n12719 ;
  assign n26408 = n11341 | n11354 ;
  assign n26409 = n3096 | n26408 ;
  assign n26406 = ( n1848 & ~n5968 ) | ( n1848 & n8771 ) | ( ~n5968 & n8771 ) ;
  assign n26407 = n26406 ^ n23275 ^ n5829 ;
  assign n26410 = n26409 ^ n26407 ^ n6210 ;
  assign n26412 = n14098 ^ n6437 ^ n1823 ;
  assign n26413 = ( ~n11964 & n20449 ) | ( ~n11964 & n26412 ) | ( n20449 & n26412 ) ;
  assign n26411 = n21803 & ~n23375 ;
  assign n26414 = n26413 ^ n26411 ^ 1'b0 ;
  assign n26415 = ~n1011 & n20107 ;
  assign n26416 = n5974 ^ n2141 ^ 1'b0 ;
  assign n26417 = n3232 & n26416 ;
  assign n26418 = n26417 ^ n6982 ^ 1'b0 ;
  assign n26419 = n8607 & ~n22693 ;
  assign n26420 = ~n25509 & n26419 ;
  assign n26421 = n3362 & n7454 ;
  assign n26422 = n26421 ^ n7808 ^ 1'b0 ;
  assign n26423 = ( n11462 & ~n25492 ) | ( n11462 & n26422 ) | ( ~n25492 & n26422 ) ;
  assign n26424 = ~n1440 & n6330 ;
  assign n26425 = ~n3626 & n26424 ;
  assign n26426 = n25375 ^ n16899 ^ 1'b0 ;
  assign n26427 = n26425 | n26426 ;
  assign n26428 = ( ~n12471 & n24894 ) | ( ~n12471 & n26427 ) | ( n24894 & n26427 ) ;
  assign n26429 = n1962 | n4113 ;
  assign n26430 = n26429 ^ n11873 ^ n8915 ;
  assign n26431 = ( ~n3363 & n13736 ) | ( ~n3363 & n16795 ) | ( n13736 & n16795 ) ;
  assign n26432 = n26431 ^ n19404 ^ 1'b0 ;
  assign n26433 = n26430 & n26432 ;
  assign n26434 = ( ~n13369 & n17835 ) | ( ~n13369 & n17966 ) | ( n17835 & n17966 ) ;
  assign n26435 = ( n10189 & n14818 ) | ( n10189 & ~n26434 ) | ( n14818 & ~n26434 ) ;
  assign n26436 = n15496 ^ n12284 ^ 1'b0 ;
  assign n26437 = ~n9775 & n11924 ;
  assign n26438 = n26437 ^ n1821 ^ 1'b0 ;
  assign n26439 = ( n7034 & n26436 ) | ( n7034 & n26438 ) | ( n26436 & n26438 ) ;
  assign n26440 = n4202 ^ n3674 ^ n3398 ;
  assign n26441 = ( n1158 & n14145 ) | ( n1158 & n18917 ) | ( n14145 & n18917 ) ;
  assign n26442 = n23535 ^ n2491 ^ 1'b0 ;
  assign n26443 = n19957 & ~n26442 ;
  assign n26444 = n2666 & ~n26443 ;
  assign n26445 = ( ~n2961 & n16845 ) | ( ~n2961 & n26444 ) | ( n16845 & n26444 ) ;
  assign n26446 = n10985 | n12725 ;
  assign n26447 = n14762 ^ n12013 ^ n9063 ;
  assign n26448 = n26447 ^ n4225 ^ n2585 ;
  assign n26449 = n4524 ^ n1753 ^ n1381 ;
  assign n26450 = ~n10045 & n26449 ;
  assign n26451 = ~n8827 & n26450 ;
  assign n26452 = ( ~n395 & n5512 ) | ( ~n395 & n19158 ) | ( n5512 & n19158 ) ;
  assign n26453 = n4584 | n5277 ;
  assign n26454 = n26452 | n26453 ;
  assign n26455 = n26454 ^ n8258 ^ 1'b0 ;
  assign n26456 = ( ~n1843 & n26451 ) | ( ~n1843 & n26455 ) | ( n26451 & n26455 ) ;
  assign n26457 = ( n2704 & n11339 ) | ( n2704 & ~n26456 ) | ( n11339 & ~n26456 ) ;
  assign n26461 = ( n1137 & n1711 ) | ( n1137 & n9166 ) | ( n1711 & n9166 ) ;
  assign n26458 = n23707 ^ n6990 ^ n914 ;
  assign n26459 = ( n5248 & n7357 ) | ( n5248 & n26458 ) | ( n7357 & n26458 ) ;
  assign n26460 = n20751 | n26459 ;
  assign n26462 = n26461 ^ n26460 ^ 1'b0 ;
  assign n26463 = ( n17983 & ~n26457 ) | ( n17983 & n26462 ) | ( ~n26457 & n26462 ) ;
  assign n26464 = n26463 ^ n13001 ^ n11975 ;
  assign n26465 = n23068 ^ n3806 ^ 1'b0 ;
  assign n26466 = ( ~n5335 & n20336 ) | ( ~n5335 & n26465 ) | ( n20336 & n26465 ) ;
  assign n26467 = n3459 ^ n3290 ^ 1'b0 ;
  assign n26468 = n14552 | n26467 ;
  assign n26469 = n26468 ^ n1572 ^ 1'b0 ;
  assign n26470 = n5224 & ~n26469 ;
  assign n26471 = n7991 | n19831 ;
  assign n26472 = ~n14618 & n26471 ;
  assign n26473 = n26472 ^ n17301 ^ 1'b0 ;
  assign n26474 = n24741 ^ n15315 ^ n3961 ;
  assign n26475 = n18924 ^ n12608 ^ n8649 ;
  assign n26476 = ( n26473 & n26474 ) | ( n26473 & ~n26475 ) | ( n26474 & ~n26475 ) ;
  assign n26477 = ~n2527 & n13232 ;
  assign n26478 = n26477 ^ n15238 ^ 1'b0 ;
  assign n26479 = n16503 & ~n26478 ;
  assign n26480 = ~n19274 & n26479 ;
  assign n26481 = ( n3042 & ~n7491 ) | ( n3042 & n26480 ) | ( ~n7491 & n26480 ) ;
  assign n26482 = ( n3738 & ~n6053 ) | ( n3738 & n15033 ) | ( ~n6053 & n15033 ) ;
  assign n26483 = n26482 ^ n7357 ^ n2580 ;
  assign n26488 = n11518 ^ n3789 ^ n3661 ;
  assign n26489 = ~n11025 & n26488 ;
  assign n26490 = ~n8210 & n26489 ;
  assign n26485 = n8322 & ~n13191 ;
  assign n26486 = n26485 ^ n9794 ^ 1'b0 ;
  assign n26487 = ( n16760 & ~n17728 ) | ( n16760 & n26486 ) | ( ~n17728 & n26486 ) ;
  assign n26484 = ( n1014 & n3414 ) | ( n1014 & n9380 ) | ( n3414 & n9380 ) ;
  assign n26491 = n26490 ^ n26487 ^ n26484 ;
  assign n26492 = ( n1294 & n12961 ) | ( n1294 & ~n13459 ) | ( n12961 & ~n13459 ) ;
  assign n26493 = ( n12902 & n25118 ) | ( n12902 & n26492 ) | ( n25118 & n26492 ) ;
  assign n26494 = n8241 ^ n7601 ^ 1'b0 ;
  assign n26495 = n26494 ^ n20606 ^ n6829 ;
  assign n26496 = n10976 ^ n5122 ^ n2090 ;
  assign n26497 = n16398 ^ n4192 ^ n2489 ;
  assign n26498 = n26497 ^ n13362 ^ n4777 ;
  assign n26499 = n14890 & ~n26286 ;
  assign n26500 = n26499 ^ n18720 ^ 1'b0 ;
  assign n26501 = n17012 ^ n13465 ^ 1'b0 ;
  assign n26502 = n2651 & n2722 ;
  assign n26503 = n26502 ^ n7600 ^ n1918 ;
  assign n26504 = ( n8561 & ~n26501 ) | ( n8561 & n26503 ) | ( ~n26501 & n26503 ) ;
  assign n26505 = ( n3959 & n13473 ) | ( n3959 & n14263 ) | ( n13473 & n14263 ) ;
  assign n26506 = n26505 ^ n24239 ^ 1'b0 ;
  assign n26507 = n10605 & ~n26506 ;
  assign n26510 = n11942 & n13131 ;
  assign n26511 = n26510 ^ n2334 ^ 1'b0 ;
  assign n26512 = n26511 ^ n2445 ^ 1'b0 ;
  assign n26513 = n9372 & ~n26512 ;
  assign n26508 = n15450 ^ n8749 ^ 1'b0 ;
  assign n26509 = n17918 & ~n26508 ;
  assign n26514 = n26513 ^ n26509 ^ n14390 ;
  assign n26515 = n26514 ^ n6505 ^ 1'b0 ;
  assign n26516 = n11780 | n26515 ;
  assign n26517 = n11205 ^ n10389 ^ 1'b0 ;
  assign n26518 = ( ~n1408 & n7357 ) | ( ~n1408 & n26517 ) | ( n7357 & n26517 ) ;
  assign n26519 = n7065 ^ n7056 ^ n4673 ;
  assign n26520 = ( n1191 & n26518 ) | ( n1191 & n26519 ) | ( n26518 & n26519 ) ;
  assign n26521 = n26520 ^ n23199 ^ 1'b0 ;
  assign n26522 = n12166 & ~n12222 ;
  assign n26523 = ( n2198 & ~n15543 ) | ( n2198 & n26522 ) | ( ~n15543 & n26522 ) ;
  assign n26524 = n8982 & ~n10389 ;
  assign n26525 = n26524 ^ n13016 ^ 1'b0 ;
  assign n26526 = ( n1085 & n12725 ) | ( n1085 & ~n26525 ) | ( n12725 & ~n26525 ) ;
  assign n26527 = n7197 | n14516 ;
  assign n26528 = n26527 ^ n12040 ^ 1'b0 ;
  assign n26531 = n20163 ^ n6205 ^ 1'b0 ;
  assign n26529 = n19297 & ~n24813 ;
  assign n26530 = n26529 ^ n12202 ^ 1'b0 ;
  assign n26532 = n26531 ^ n26530 ^ 1'b0 ;
  assign n26533 = ~n18919 & n26532 ;
  assign n26534 = n1634 | n25943 ;
  assign n26535 = n12246 | n26534 ;
  assign n26536 = n8195 & n26535 ;
  assign n26537 = n26105 & n26536 ;
  assign n26538 = n23510 ^ n9716 ^ n1459 ;
  assign n26539 = n24196 ^ n17680 ^ n7721 ;
  assign n26540 = ( ~n6127 & n14279 ) | ( ~n6127 & n14580 ) | ( n14279 & n14580 ) ;
  assign n26541 = ( ~n5074 & n8053 ) | ( ~n5074 & n26540 ) | ( n8053 & n26540 ) ;
  assign n26542 = ~n11468 & n15672 ;
  assign n26543 = n5269 & ~n24762 ;
  assign n26544 = ~n26542 & n26543 ;
  assign n26545 = n18027 ^ n15847 ^ 1'b0 ;
  assign n26546 = n26544 | n26545 ;
  assign n26550 = ( n1433 & n12622 ) | ( n1433 & ~n17514 ) | ( n12622 & ~n17514 ) ;
  assign n26549 = n16368 ^ n11487 ^ 1'b0 ;
  assign n26551 = n26550 ^ n26549 ^ n760 ;
  assign n26547 = n23248 ^ n8607 ^ n5009 ;
  assign n26548 = n10332 | n26547 ;
  assign n26552 = n26551 ^ n26548 ^ 1'b0 ;
  assign n26556 = ( n12241 & n13665 ) | ( n12241 & ~n14590 ) | ( n13665 & ~n14590 ) ;
  assign n26553 = ( ~n1728 & n15897 ) | ( ~n1728 & n21076 ) | ( n15897 & n21076 ) ;
  assign n26554 = ~n7928 & n11305 ;
  assign n26555 = ~n26553 & n26554 ;
  assign n26557 = n26556 ^ n26555 ^ 1'b0 ;
  assign n26558 = n26557 ^ n13413 ^ n4908 ;
  assign n26562 = ( n5858 & n12776 ) | ( n5858 & ~n22397 ) | ( n12776 & ~n22397 ) ;
  assign n26560 = n5077 & ~n5833 ;
  assign n26559 = n374 & ~n20663 ;
  assign n26561 = n26560 ^ n26559 ^ 1'b0 ;
  assign n26563 = n26562 ^ n26561 ^ n6067 ;
  assign n26564 = n13581 & ~n24074 ;
  assign n26568 = ( n2403 & n2706 ) | ( n2403 & n25120 ) | ( n2706 & n25120 ) ;
  assign n26565 = n8822 & n9741 ;
  assign n26566 = n26565 ^ n1127 ^ 1'b0 ;
  assign n26567 = n23508 & n26566 ;
  assign n26569 = n26568 ^ n26567 ^ 1'b0 ;
  assign n26570 = x92 & n5662 ;
  assign n26571 = n9105 & n26570 ;
  assign n26572 = n26571 ^ n3961 ^ n1340 ;
  assign n26573 = n26572 ^ n12906 ^ n1297 ;
  assign n26574 = n17244 | n25945 ;
  assign n26575 = n26574 ^ n21039 ^ 1'b0 ;
  assign n26576 = n26573 | n26575 ;
  assign n26577 = n25660 ^ n7562 ^ 1'b0 ;
  assign n26578 = x239 & n1227 ;
  assign n26579 = n12750 ^ n4447 ^ 1'b0 ;
  assign n26580 = n7353 & n26579 ;
  assign n26581 = ( n2881 & ~n6970 ) | ( n2881 & n26580 ) | ( ~n6970 & n26580 ) ;
  assign n26582 = ~n26578 & n26581 ;
  assign n26583 = n26582 ^ n19491 ^ n632 ;
  assign n26584 = n12086 ^ n4795 ^ 1'b0 ;
  assign n26585 = n14678 ^ x38 ^ 1'b0 ;
  assign n26586 = n12673 ^ n4497 ^ n3680 ;
  assign n26587 = n10525 | n26586 ;
  assign n26588 = n26478 & n26587 ;
  assign n26589 = ( n12851 & n16016 ) | ( n12851 & n17861 ) | ( n16016 & n17861 ) ;
  assign n26590 = n13844 ^ n12847 ^ n12644 ;
  assign n26591 = n26590 ^ n10585 ^ 1'b0 ;
  assign n26592 = n26589 & n26591 ;
  assign n26593 = n11424 ^ n1457 ^ n407 ;
  assign n26594 = n11863 ^ n872 ^ 1'b0 ;
  assign n26595 = n7641 & ~n26594 ;
  assign n26596 = n26593 & n26595 ;
  assign n26597 = n26596 ^ n11161 ^ 1'b0 ;
  assign n26598 = n26597 ^ n402 ^ 1'b0 ;
  assign n26599 = n5213 | n20216 ;
  assign n26600 = n7077 | n26599 ;
  assign n26601 = x161 & ~n6583 ;
  assign n26602 = n26601 ^ n5920 ^ 1'b0 ;
  assign n26603 = ( n8044 & n26047 ) | ( n8044 & n26602 ) | ( n26047 & n26602 ) ;
  assign n26604 = ( n2108 & n3671 ) | ( n2108 & n11489 ) | ( n3671 & n11489 ) ;
  assign n26605 = ( n4024 & ~n8010 ) | ( n4024 & n13884 ) | ( ~n8010 & n13884 ) ;
  assign n26606 = n26605 ^ n22092 ^ 1'b0 ;
  assign n26607 = n502 & ~n26606 ;
  assign n26608 = n26607 ^ n15193 ^ n11356 ;
  assign n26609 = n6681 & ~n16240 ;
  assign n26610 = ~n1113 & n26609 ;
  assign n26611 = n26610 ^ n15429 ^ 1'b0 ;
  assign n26612 = n16739 ^ x24 ^ 1'b0 ;
  assign n26613 = ( n1170 & n1197 ) | ( n1170 & n10259 ) | ( n1197 & n10259 ) ;
  assign n26614 = ( n927 & n21832 ) | ( n927 & n26613 ) | ( n21832 & n26613 ) ;
  assign n26615 = ( n5630 & n26612 ) | ( n5630 & ~n26614 ) | ( n26612 & ~n26614 ) ;
  assign n26616 = n15993 ^ n8840 ^ n7910 ;
  assign n26617 = ~n12818 & n22675 ;
  assign n26618 = n26617 ^ n2603 ^ 1'b0 ;
  assign n26619 = n4585 & n22878 ;
  assign n26621 = n16963 | n22898 ;
  assign n26622 = n12213 | n26621 ;
  assign n26620 = n15993 ^ n7977 ^ 1'b0 ;
  assign n26623 = n26622 ^ n26620 ^ n2871 ;
  assign n26624 = ( n4295 & ~n12739 ) | ( n4295 & n19946 ) | ( ~n12739 & n19946 ) ;
  assign n26625 = ( ~n1401 & n18798 ) | ( ~n1401 & n26624 ) | ( n18798 & n26624 ) ;
  assign n26626 = n26625 ^ n8048 ^ n6664 ;
  assign n26627 = ( n919 & ~n1960 ) | ( n919 & n12212 ) | ( ~n1960 & n12212 ) ;
  assign n26628 = n11920 ^ n2645 ^ 1'b0 ;
  assign n26629 = n11516 & ~n26628 ;
  assign n26630 = ~n26627 & n26629 ;
  assign n26631 = n10331 | n11110 ;
  assign n26632 = n19358 | n26631 ;
  assign n26633 = n17998 ^ n13263 ^ n10345 ;
  assign n26634 = ( n9390 & n12152 ) | ( n9390 & ~n26633 ) | ( n12152 & ~n26633 ) ;
  assign n26635 = n15914 ^ n8887 ^ 1'b0 ;
  assign n26636 = n26635 ^ n24975 ^ n18808 ;
  assign n26637 = n10067 ^ n5351 ^ n2016 ;
  assign n26638 = n5656 & n12029 ;
  assign n26639 = n10091 ^ n444 ^ 1'b0 ;
  assign n26640 = ( n12894 & n26638 ) | ( n12894 & n26639 ) | ( n26638 & n26639 ) ;
  assign n26641 = n16888 ^ n453 ^ 1'b0 ;
  assign n26642 = ( ~x109 & n1473 ) | ( ~x109 & n8772 ) | ( n1473 & n8772 ) ;
  assign n26643 = n4521 ^ n1454 ^ 1'b0 ;
  assign n26644 = n8526 ^ n3902 ^ 1'b0 ;
  assign n26645 = ~n9988 & n26644 ;
  assign n26646 = ( n11386 & ~n26643 ) | ( n11386 & n26645 ) | ( ~n26643 & n26645 ) ;
  assign n26647 = ( n26641 & n26642 ) | ( n26641 & ~n26646 ) | ( n26642 & ~n26646 ) ;
  assign n26648 = ( n26637 & n26640 ) | ( n26637 & ~n26647 ) | ( n26640 & ~n26647 ) ;
  assign n26649 = n15251 ^ n11601 ^ 1'b0 ;
  assign n26650 = ( n20380 & n21927 ) | ( n20380 & n26649 ) | ( n21927 & n26649 ) ;
  assign n26651 = n13066 ^ n5638 ^ n4334 ;
  assign n26652 = ~n6775 & n11837 ;
  assign n26653 = n26651 & n26652 ;
  assign n26654 = n26653 ^ n21377 ^ 1'b0 ;
  assign n26655 = ( n9225 & n26650 ) | ( n9225 & n26654 ) | ( n26650 & n26654 ) ;
  assign n26656 = n22811 ^ n7713 ^ 1'b0 ;
  assign n26657 = n15208 | n26656 ;
  assign n26658 = n26553 ^ n13224 ^ 1'b0 ;
  assign n26659 = ( ~n4172 & n13380 ) | ( ~n4172 & n26658 ) | ( n13380 & n26658 ) ;
  assign n26662 = n12281 | n14498 ;
  assign n26663 = n4452 & ~n26662 ;
  assign n26660 = n7738 & ~n8494 ;
  assign n26661 = n26660 ^ n19523 ^ n15520 ;
  assign n26664 = n26663 ^ n26661 ^ n15491 ;
  assign n26665 = n1299 | n21158 ;
  assign n26666 = ( ~n10137 & n15222 ) | ( ~n10137 & n26665 ) | ( n15222 & n26665 ) ;
  assign n26667 = ~n3245 & n22186 ;
  assign n26668 = ( ~n845 & n7327 ) | ( ~n845 & n16569 ) | ( n7327 & n16569 ) ;
  assign n26669 = n26668 ^ n17234 ^ n14760 ;
  assign n26670 = n26669 ^ n5075 ^ 1'b0 ;
  assign n26671 = ~n25755 & n26670 ;
  assign n26672 = n9706 ^ n6622 ^ n2019 ;
  assign n26673 = n1663 & n2045 ;
  assign n26674 = ( n10352 & n26672 ) | ( n10352 & n26673 ) | ( n26672 & n26673 ) ;
  assign n26675 = ( ~n8250 & n16741 ) | ( ~n8250 & n23272 ) | ( n16741 & n23272 ) ;
  assign n26676 = n4361 | n26675 ;
  assign n26677 = n6703 | n26676 ;
  assign n26678 = ~n9491 & n26677 ;
  assign n26679 = n26678 ^ n1301 ^ 1'b0 ;
  assign n26680 = n26679 ^ n24943 ^ 1'b0 ;
  assign n26681 = n657 & ~n9703 ;
  assign n26682 = ( ~n3043 & n5230 ) | ( ~n3043 & n13821 ) | ( n5230 & n13821 ) ;
  assign n26683 = ( n26680 & n26681 ) | ( n26680 & n26682 ) | ( n26681 & n26682 ) ;
  assign n26684 = ( n11401 & ~n22785 ) | ( n11401 & n25028 ) | ( ~n22785 & n25028 ) ;
  assign n26685 = n26684 ^ n23974 ^ n2912 ;
  assign n26686 = n1363 | n18763 ;
  assign n26687 = ~n2594 & n26637 ;
  assign n26688 = n15407 ^ n5890 ^ n4396 ;
  assign n26689 = n26688 ^ n21839 ^ n12481 ;
  assign n26691 = ( n5421 & n5904 ) | ( n5421 & n14993 ) | ( n5904 & n14993 ) ;
  assign n26690 = n8910 & ~n12943 ;
  assign n26692 = n26691 ^ n26690 ^ n17198 ;
  assign n26693 = ( n1461 & n4304 ) | ( n1461 & ~n6994 ) | ( n4304 & ~n6994 ) ;
  assign n26694 = ~n5520 & n13891 ;
  assign n26695 = n26693 & n26694 ;
  assign n26696 = n3085 & n6222 ;
  assign n26697 = ~n18666 & n26696 ;
  assign n26698 = n26697 ^ n25691 ^ 1'b0 ;
  assign n26699 = n26695 | n26698 ;
  assign n26701 = n12741 ^ n5907 ^ x67 ;
  assign n26702 = n4592 | n26701 ;
  assign n26703 = ~n1541 & n26702 ;
  assign n26704 = n26703 ^ n3962 ^ 1'b0 ;
  assign n26700 = n6383 & ~n13303 ;
  assign n26705 = n26704 ^ n26700 ^ 1'b0 ;
  assign n26706 = n26705 ^ n15930 ^ n1949 ;
  assign n26707 = ( n4342 & n10114 ) | ( n4342 & ~n18857 ) | ( n10114 & ~n18857 ) ;
  assign n26708 = n19101 ^ n16470 ^ n3514 ;
  assign n26709 = n26708 ^ n12108 ^ n6850 ;
  assign n26711 = ( ~n4590 & n6434 ) | ( ~n4590 & n7556 ) | ( n6434 & n7556 ) ;
  assign n26710 = n14765 ^ n6460 ^ x33 ;
  assign n26712 = n26711 ^ n26710 ^ n5856 ;
  assign n26713 = n12644 ^ n7321 ^ n4548 ;
  assign n26714 = ~n25510 & n26713 ;
  assign n26715 = n15114 | n18589 ;
  assign n26716 = ( ~n412 & n2417 ) | ( ~n412 & n2609 ) | ( n2417 & n2609 ) ;
  assign n26717 = n8762 ^ n6523 ^ 1'b0 ;
  assign n26718 = n4810 & n26717 ;
  assign n26719 = ( n21652 & ~n26716 ) | ( n21652 & n26718 ) | ( ~n26716 & n26718 ) ;
  assign n26720 = n26425 ^ n20687 ^ n11942 ;
  assign n26721 = n20990 ^ n9521 ^ 1'b0 ;
  assign n26722 = n26720 | n26721 ;
  assign n26723 = n18293 & ~n25877 ;
  assign n26724 = n6103 & n26723 ;
  assign n26725 = n1777 & n8752 ;
  assign n26729 = ~n1675 & n8574 ;
  assign n26730 = n4876 | n9154 ;
  assign n26731 = n26729 | n26730 ;
  assign n26728 = n6622 ^ n4463 ^ n1818 ;
  assign n26726 = n20609 ^ n11730 ^ 1'b0 ;
  assign n26727 = ~n3811 & n26726 ;
  assign n26732 = n26731 ^ n26728 ^ n26727 ;
  assign n26733 = ( n5844 & n8421 ) | ( n5844 & n15116 ) | ( n8421 & n15116 ) ;
  assign n26734 = n8405 ^ n2521 ^ n1650 ;
  assign n26735 = n11084 & n26734 ;
  assign n26736 = ~n26733 & n26735 ;
  assign n26737 = ~n15123 & n15932 ;
  assign n26738 = n26737 ^ n9866 ^ 1'b0 ;
  assign n26739 = n26738 ^ n8979 ^ 1'b0 ;
  assign n26740 = n23949 & ~n26739 ;
  assign n26741 = n11990 ^ n11274 ^ n5670 ;
  assign n26742 = n20293 ^ n13862 ^ n4090 ;
  assign n26743 = ( ~x81 & n26741 ) | ( ~x81 & n26742 ) | ( n26741 & n26742 ) ;
  assign n26744 = n26743 ^ n21664 ^ n10061 ;
  assign n26745 = n13047 & n21319 ;
  assign n26746 = ( n21165 & ~n26744 ) | ( n21165 & n26745 ) | ( ~n26744 & n26745 ) ;
  assign n26747 = n21245 ^ n10233 ^ 1'b0 ;
  assign n26748 = n22115 | n26747 ;
  assign n26749 = ( ~n7285 & n12509 ) | ( ~n7285 & n26748 ) | ( n12509 & n26748 ) ;
  assign n26750 = n23899 ^ n7252 ^ n914 ;
  assign n26751 = ( ~x167 & n7770 ) | ( ~x167 & n26750 ) | ( n7770 & n26750 ) ;
  assign n26752 = ( n8289 & ~n13369 ) | ( n8289 & n24329 ) | ( ~n13369 & n24329 ) ;
  assign n26753 = n26751 | n26752 ;
  assign n26754 = n26753 ^ n2413 ^ 1'b0 ;
  assign n26756 = n8909 ^ n1440 ^ n1320 ;
  assign n26755 = n24768 ^ n7184 ^ n1416 ;
  assign n26757 = n26756 ^ n26755 ^ 1'b0 ;
  assign n26758 = n18580 ^ n15765 ^ n15109 ;
  assign n26759 = n26758 ^ n21431 ^ 1'b0 ;
  assign n26760 = n8318 | n26759 ;
  assign n26761 = n2641 & n9027 ;
  assign n26762 = n22092 ^ n18834 ^ n16815 ;
  assign n26763 = n22603 ^ n6637 ^ n578 ;
  assign n26764 = n26763 ^ n23088 ^ 1'b0 ;
  assign n26765 = ~n7142 & n7708 ;
  assign n26766 = ~n26174 & n26765 ;
  assign n26767 = ( n20534 & n20833 ) | ( n20534 & n26766 ) | ( n20833 & n26766 ) ;
  assign n26768 = ( ~n7654 & n13598 ) | ( ~n7654 & n26767 ) | ( n13598 & n26767 ) ;
  assign n26769 = n10741 ^ n5153 ^ n4764 ;
  assign n26770 = n19967 ^ n13933 ^ n4049 ;
  assign n26771 = n850 & n26770 ;
  assign n26772 = n26769 & ~n26771 ;
  assign n26773 = n8504 | n26351 ;
  assign n26774 = n20337 ^ n1510 ^ 1'b0 ;
  assign n26775 = n26773 | n26774 ;
  assign n26776 = n26775 ^ n13607 ^ 1'b0 ;
  assign n26777 = n26772 | n26776 ;
  assign n26778 = n12339 ^ n4447 ^ n1517 ;
  assign n26779 = n26778 ^ n11468 ^ 1'b0 ;
  assign n26780 = ( n6293 & n10106 ) | ( n6293 & ~n26779 ) | ( n10106 & ~n26779 ) ;
  assign n26782 = n25077 ^ n9792 ^ n568 ;
  assign n26781 = ~n7318 & n15173 ;
  assign n26783 = n26782 ^ n26781 ^ 1'b0 ;
  assign n26784 = n10150 & n19554 ;
  assign n26785 = n26784 ^ n4494 ^ 1'b0 ;
  assign n26787 = ~n11899 & n12861 ;
  assign n26788 = ~n16650 & n26787 ;
  assign n26789 = ( n1799 & n7285 ) | ( n1799 & ~n19136 ) | ( n7285 & ~n19136 ) ;
  assign n26790 = n26788 | n26789 ;
  assign n26791 = n26790 ^ n24025 ^ 1'b0 ;
  assign n26786 = n18479 ^ n11422 ^ n10348 ;
  assign n26792 = n26791 ^ n26786 ^ n1079 ;
  assign n26793 = n25974 ^ n16722 ^ n12029 ;
  assign n26794 = n12454 & n13689 ;
  assign n26795 = ( n22859 & n26793 ) | ( n22859 & n26794 ) | ( n26793 & n26794 ) ;
  assign n26796 = n18566 ^ n13538 ^ n8839 ;
  assign n26797 = n7220 & n10283 ;
  assign n26798 = ~n26796 & n26797 ;
  assign n26799 = ( n8155 & ~n22433 ) | ( n8155 & n26798 ) | ( ~n22433 & n26798 ) ;
  assign n26801 = ( n6687 & n7295 ) | ( n6687 & n10291 ) | ( n7295 & n10291 ) ;
  assign n26800 = ~n4224 & n9695 ;
  assign n26802 = n26801 ^ n26800 ^ n23124 ;
  assign n26803 = n25641 ^ n12574 ^ n1315 ;
  assign n26804 = ~n6885 & n26803 ;
  assign n26805 = n10705 & n25179 ;
  assign n26806 = n19227 & n26805 ;
  assign n26807 = n25050 ^ n17384 ^ 1'b0 ;
  assign n26808 = n24306 & n26807 ;
  assign n26809 = n15870 ^ n12914 ^ n8335 ;
  assign n26810 = ( n8861 & n17239 ) | ( n8861 & ~n17667 ) | ( n17239 & ~n17667 ) ;
  assign n26811 = n5800 & n9052 ;
  assign n26812 = ( n7758 & ~n17020 ) | ( n7758 & n25949 ) | ( ~n17020 & n25949 ) ;
  assign n26813 = ( n2708 & n9767 ) | ( n2708 & ~n12529 ) | ( n9767 & ~n12529 ) ;
  assign n26815 = n1421 & n6977 ;
  assign n26816 = n26815 ^ n26018 ^ n16985 ;
  assign n26817 = n5515 & ~n19670 ;
  assign n26818 = ~n5421 & n6914 ;
  assign n26819 = n777 | n26818 ;
  assign n26820 = n26817 & ~n26819 ;
  assign n26821 = ( n6928 & n26816 ) | ( n6928 & n26820 ) | ( n26816 & n26820 ) ;
  assign n26814 = ( n2020 & n3925 ) | ( n2020 & ~n8239 ) | ( n3925 & ~n8239 ) ;
  assign n26822 = n26821 ^ n26814 ^ 1'b0 ;
  assign n26829 = n3369 & ~n25134 ;
  assign n26823 = n14610 ^ n5662 ^ n4464 ;
  assign n26824 = n13924 & n26823 ;
  assign n26826 = n19883 ^ n9324 ^ n5374 ;
  assign n26825 = n18601 ^ n15377 ^ n3950 ;
  assign n26827 = n26826 ^ n26825 ^ n10778 ;
  assign n26828 = ( n3119 & n26824 ) | ( n3119 & ~n26827 ) | ( n26824 & ~n26827 ) ;
  assign n26830 = n26829 ^ n26828 ^ n12398 ;
  assign n26831 = ( n15535 & ~n23609 ) | ( n15535 & n26607 ) | ( ~n23609 & n26607 ) ;
  assign n26832 = ~n3622 & n4922 ;
  assign n26833 = n16377 & n26832 ;
  assign n26834 = ( n2075 & ~n5147 ) | ( n2075 & n13691 ) | ( ~n5147 & n13691 ) ;
  assign n26835 = ( n8854 & ~n15134 ) | ( n8854 & n26834 ) | ( ~n15134 & n26834 ) ;
  assign n26836 = n26835 ^ n11361 ^ n2688 ;
  assign n26837 = ~n10247 & n21911 ;
  assign n26838 = n13567 ^ n13117 ^ n8729 ;
  assign n26839 = n26838 ^ n18056 ^ 1'b0 ;
  assign n26840 = n26549 & n26682 ;
  assign n26841 = n2674 & ~n22494 ;
  assign n26842 = n8472 | n24071 ;
  assign n26843 = n26842 ^ n11688 ^ 1'b0 ;
  assign n26844 = n14029 & n17754 ;
  assign n26845 = n6976 ^ x173 ^ 1'b0 ;
  assign n26846 = ~n26844 & n26845 ;
  assign n26847 = n26846 ^ n11608 ^ 1'b0 ;
  assign n26848 = n26847 ^ n25877 ^ 1'b0 ;
  assign n26849 = ( ~n8337 & n17513 ) | ( ~n8337 & n18596 ) | ( n17513 & n18596 ) ;
  assign n26850 = ( ~n5118 & n5687 ) | ( ~n5118 & n26849 ) | ( n5687 & n26849 ) ;
  assign n26851 = n16507 ^ n15881 ^ n576 ;
  assign n26852 = n1158 & n20727 ;
  assign n26853 = n9042 & n26852 ;
  assign n26854 = ( n4190 & n23990 ) | ( n4190 & ~n26853 ) | ( n23990 & ~n26853 ) ;
  assign n26855 = n11552 ^ x4 ^ 1'b0 ;
  assign n26856 = ( n12592 & n17121 ) | ( n12592 & n18651 ) | ( n17121 & n18651 ) ;
  assign n26857 = ( n10201 & n15425 ) | ( n10201 & n26856 ) | ( n15425 & n26856 ) ;
  assign n26858 = ( ~n7840 & n9114 ) | ( ~n7840 & n26857 ) | ( n9114 & n26857 ) ;
  assign n26859 = n17420 ^ n2918 ^ 1'b0 ;
  assign n26860 = n942 | n26859 ;
  assign n26861 = n11271 ^ n1790 ^ 1'b0 ;
  assign n26862 = ( n18631 & ~n25148 ) | ( n18631 & n26861 ) | ( ~n25148 & n26861 ) ;
  assign n26863 = n6047 ^ n3204 ^ 1'b0 ;
  assign n26864 = n4400 & n26863 ;
  assign n26865 = n1927 | n5302 ;
  assign n26866 = n26865 ^ n9501 ^ n3254 ;
  assign n26867 = ( ~n18830 & n26864 ) | ( ~n18830 & n26866 ) | ( n26864 & n26866 ) ;
  assign n26868 = n25823 ^ n13598 ^ n486 ;
  assign n26869 = ( ~n20131 & n26867 ) | ( ~n20131 & n26868 ) | ( n26867 & n26868 ) ;
  assign n26870 = n5522 ^ n1009 ^ 1'b0 ;
  assign n26871 = ( n3659 & n5864 ) | ( n3659 & ~n26870 ) | ( n5864 & ~n26870 ) ;
  assign n26872 = n11831 ^ n5744 ^ 1'b0 ;
  assign n26874 = n1611 & ~n4790 ;
  assign n26873 = n5366 | n13418 ;
  assign n26875 = n26874 ^ n26873 ^ n10277 ;
  assign n26876 = n18643 & ~n26875 ;
  assign n26877 = n26876 ^ n19807 ^ 1'b0 ;
  assign n26878 = n15110 ^ n13385 ^ n3849 ;
  assign n26879 = ~n21104 & n23804 ;
  assign n26880 = n26878 & n26879 ;
  assign n26881 = n26877 | n26880 ;
  assign n26882 = n6810 | n26881 ;
  assign n26883 = ( n1019 & ~n15414 ) | ( n1019 & n15644 ) | ( ~n15414 & n15644 ) ;
  assign n26884 = n17903 & ~n26883 ;
  assign n26885 = n26884 ^ n17974 ^ n11414 ;
  assign n26886 = ( n5212 & n5870 ) | ( n5212 & n12940 ) | ( n5870 & n12940 ) ;
  assign n26887 = ( ~n6240 & n11106 ) | ( ~n6240 & n26886 ) | ( n11106 & n26886 ) ;
  assign n26889 = n4749 ^ n3126 ^ 1'b0 ;
  assign n26888 = n1365 & ~n12093 ;
  assign n26890 = n26889 ^ n26888 ^ 1'b0 ;
  assign n26891 = x84 & ~n26890 ;
  assign n26892 = ( n5405 & ~n10422 ) | ( n5405 & n26891 ) | ( ~n10422 & n26891 ) ;
  assign n26893 = ~n26887 & n26892 ;
  assign n26894 = ( n4349 & n4417 ) | ( n4349 & ~n24026 ) | ( n4417 & ~n24026 ) ;
  assign n26895 = n19048 ^ n12789 ^ 1'b0 ;
  assign n26896 = n2350 | n26895 ;
  assign n26897 = n25398 ^ n11144 ^ n1681 ;
  assign n26898 = ( n13544 & n26896 ) | ( n13544 & ~n26897 ) | ( n26896 & ~n26897 ) ;
  assign n26899 = ( n10473 & n26894 ) | ( n10473 & ~n26898 ) | ( n26894 & ~n26898 ) ;
  assign n26903 = n14153 ^ n8169 ^ n4043 ;
  assign n26900 = n5674 ^ n2173 ^ 1'b0 ;
  assign n26901 = n1851 & ~n26900 ;
  assign n26902 = n26901 ^ n14474 ^ n14208 ;
  assign n26904 = n26903 ^ n26902 ^ 1'b0 ;
  assign n26905 = n17191 ^ n10814 ^ 1'b0 ;
  assign n26906 = n26905 ^ n15504 ^ 1'b0 ;
  assign n26907 = ( n11582 & ~n22096 ) | ( n11582 & n22490 ) | ( ~n22096 & n22490 ) ;
  assign n26908 = n26907 ^ n12744 ^ 1'b0 ;
  assign n26909 = n3287 & n26908 ;
  assign n26910 = n10840 ^ n8475 ^ 1'b0 ;
  assign n26911 = n7331 & n26910 ;
  assign n26912 = n8269 ^ n4197 ^ 1'b0 ;
  assign n26913 = ~n5755 & n26912 ;
  assign n26914 = n2154 & ~n26913 ;
  assign n26915 = ~n26911 & n26914 ;
  assign n26916 = ~n3862 & n18772 ;
  assign n26917 = ~n604 & n26907 ;
  assign n26918 = n12808 & ~n19427 ;
  assign n26919 = n19705 ^ n15155 ^ n6735 ;
  assign n26920 = n25986 ^ n11102 ^ 1'b0 ;
  assign n26921 = ~n26919 & n26920 ;
  assign n26922 = ~n5908 & n6045 ;
  assign n26923 = n11652 & n26922 ;
  assign n26924 = ( n4211 & ~n6357 ) | ( n4211 & n15158 ) | ( ~n6357 & n15158 ) ;
  assign n26925 = ( ~n6555 & n9897 ) | ( ~n6555 & n26924 ) | ( n9897 & n26924 ) ;
  assign n26926 = n4884 & ~n24894 ;
  assign n26927 = ~n6992 & n26926 ;
  assign n26928 = ( n17885 & n26925 ) | ( n17885 & ~n26927 ) | ( n26925 & ~n26927 ) ;
  assign n26929 = ( n3917 & n26923 ) | ( n3917 & n26928 ) | ( n26923 & n26928 ) ;
  assign n26930 = n16982 ^ n6385 ^ n3158 ;
  assign n26931 = n10602 ^ n8426 ^ n3322 ;
  assign n26932 = n26931 ^ n3900 ^ 1'b0 ;
  assign n26933 = ( n13875 & ~n21729 ) | ( n13875 & n22876 ) | ( ~n21729 & n22876 ) ;
  assign n26934 = n14688 & ~n26933 ;
  assign n26935 = n12742 & n26934 ;
  assign n26936 = n6377 ^ n5456 ^ n777 ;
  assign n26937 = ( ~n6252 & n7711 ) | ( ~n6252 & n26936 ) | ( n7711 & n26936 ) ;
  assign n26938 = n26937 ^ n21975 ^ n10743 ;
  assign n26939 = x85 | n26938 ;
  assign n26940 = n15203 ^ n13688 ^ n7778 ;
  assign n26941 = n26940 ^ n22487 ^ 1'b0 ;
  assign n26942 = n26941 ^ n24493 ^ n15950 ;
  assign n26943 = n20257 ^ n6639 ^ n5701 ;
  assign n26944 = n13894 ^ n2782 ^ 1'b0 ;
  assign n26945 = n13903 & ~n26944 ;
  assign n26946 = n1755 & n22122 ;
  assign n26947 = n3873 & n26946 ;
  assign n26948 = n26947 ^ n20312 ^ 1'b0 ;
  assign n26953 = n3826 ^ n3657 ^ n3391 ;
  assign n26949 = n9737 ^ n7566 ^ n7324 ;
  assign n26950 = n26949 ^ n9542 ^ n6703 ;
  assign n26951 = ( n14282 & n16594 ) | ( n14282 & n26950 ) | ( n16594 & n26950 ) ;
  assign n26952 = ( n13540 & n17630 ) | ( n13540 & ~n26951 ) | ( n17630 & ~n26951 ) ;
  assign n26954 = n26953 ^ n26952 ^ n24758 ;
  assign n26955 = ~n7569 & n17855 ;
  assign n26956 = n26955 ^ n18476 ^ n9958 ;
  assign n26957 = ( ~x15 & n26356 ) | ( ~x15 & n26956 ) | ( n26356 & n26956 ) ;
  assign n26958 = n26957 ^ n15293 ^ n1931 ;
  assign n26959 = n3989 & ~n22397 ;
  assign n26960 = n26959 ^ n18659 ^ n9152 ;
  assign n26961 = ( n11208 & n26958 ) | ( n11208 & n26960 ) | ( n26958 & n26960 ) ;
  assign n26962 = n10961 & n26961 ;
  assign n26963 = n26954 & n26962 ;
  assign n26964 = n20004 ^ n5479 ^ n4889 ;
  assign n26965 = ( ~n6849 & n8417 ) | ( ~n6849 & n20175 ) | ( n8417 & n20175 ) ;
  assign n26966 = ( n11453 & ~n26964 ) | ( n11453 & n26965 ) | ( ~n26964 & n26965 ) ;
  assign n26967 = ( n4808 & n7525 ) | ( n4808 & ~n23526 ) | ( n7525 & ~n23526 ) ;
  assign n26968 = ~n10185 & n26967 ;
  assign n26969 = n26968 ^ n6987 ^ 1'b0 ;
  assign n26970 = n20065 ^ n12054 ^ 1'b0 ;
  assign n26971 = n26969 & ~n26970 ;
  assign n26972 = ( ~n1084 & n9238 ) | ( ~n1084 & n21352 ) | ( n9238 & n21352 ) ;
  assign n26973 = n14524 | n17833 ;
  assign n26974 = ~n19845 & n22168 ;
  assign n26975 = n26974 ^ n9484 ^ n8790 ;
  assign n26976 = ( n1317 & n4767 ) | ( n1317 & ~n19550 ) | ( n4767 & ~n19550 ) ;
  assign n26977 = n26976 ^ n7693 ^ 1'b0 ;
  assign n26978 = n5548 & n26977 ;
  assign n26979 = n10223 ^ n1833 ^ 1'b0 ;
  assign n26980 = ~n23506 & n26979 ;
  assign n26981 = n26980 ^ n11076 ^ 1'b0 ;
  assign n26983 = ~n6878 & n8800 ;
  assign n26984 = n3998 & n26983 ;
  assign n26982 = ~n1486 & n6590 ;
  assign n26985 = n26984 ^ n26982 ^ 1'b0 ;
  assign n26986 = ( ~n4380 & n20044 ) | ( ~n4380 & n26985 ) | ( n20044 & n26985 ) ;
  assign n26990 = ( n1579 & ~n5241 ) | ( n1579 & n23041 ) | ( ~n5241 & n23041 ) ;
  assign n26987 = ( ~n4751 & n16111 ) | ( ~n4751 & n19473 ) | ( n16111 & n19473 ) ;
  assign n26988 = n26987 ^ n14828 ^ n8817 ;
  assign n26989 = ( n7035 & ~n11858 ) | ( n7035 & n26988 ) | ( ~n11858 & n26988 ) ;
  assign n26991 = n26990 ^ n26989 ^ n11591 ;
  assign n26992 = n6652 & ~n15772 ;
  assign n26993 = ~n11158 & n26992 ;
  assign n26994 = n17802 | n26993 ;
  assign n26995 = ( n6699 & n9169 ) | ( n6699 & ~n26994 ) | ( n9169 & ~n26994 ) ;
  assign n26996 = n20871 ^ n5611 ^ n3178 ;
  assign n26997 = n26996 ^ n23151 ^ n22462 ;
  assign n26998 = ( n2453 & n2880 ) | ( n2453 & n5083 ) | ( n2880 & n5083 ) ;
  assign n26999 = ( n700 & n6092 ) | ( n700 & n26998 ) | ( n6092 & n26998 ) ;
  assign n27000 = n26999 ^ n26653 ^ 1'b0 ;
  assign n27001 = n19532 ^ n10161 ^ 1'b0 ;
  assign n27003 = n2856 & ~n5527 ;
  assign n27004 = n1634 & n27003 ;
  assign n27002 = n1288 ^ n545 ^ 1'b0 ;
  assign n27005 = n27004 ^ n27002 ^ n12150 ;
  assign n27006 = n2819 ^ n2412 ^ n662 ;
  assign n27007 = n27006 ^ n16201 ^ n6609 ;
  assign n27008 = n16064 ^ n9086 ^ 1'b0 ;
  assign n27009 = n7070 & n27008 ;
  assign n27010 = n22615 ^ n840 ^ 1'b0 ;
  assign n27011 = n27010 ^ n22484 ^ n15196 ;
  assign n27013 = n5637 ^ n1007 ^ 1'b0 ;
  assign n27014 = n27013 ^ n17754 ^ n6540 ;
  assign n27012 = n4769 | n12035 ;
  assign n27015 = n27014 ^ n27012 ^ 1'b0 ;
  assign n27016 = ( n10455 & n17037 ) | ( n10455 & n25847 ) | ( n17037 & n25847 ) ;
  assign n27017 = n1400 & n24578 ;
  assign n27018 = n27017 ^ n8746 ^ 1'b0 ;
  assign n27019 = n1110 & ~n11360 ;
  assign n27020 = n4969 & n27019 ;
  assign n27021 = n2742 & ~n9874 ;
  assign n27022 = ~n15943 & n27021 ;
  assign n27023 = n14535 ^ n7821 ^ n2492 ;
  assign n27024 = ( n3270 & n21762 ) | ( n3270 & ~n27023 ) | ( n21762 & ~n27023 ) ;
  assign n27025 = ( ~n2722 & n18115 ) | ( ~n2722 & n27024 ) | ( n18115 & n27024 ) ;
  assign n27026 = ( n15457 & n16675 ) | ( n15457 & n27025 ) | ( n16675 & n27025 ) ;
  assign n27027 = n1352 & ~n9580 ;
  assign n27028 = n27027 ^ n17631 ^ 1'b0 ;
  assign n27029 = n27028 ^ n24608 ^ n1212 ;
  assign n27030 = n26668 ^ n23934 ^ n8480 ;
  assign n27031 = ( n10307 & n15657 ) | ( n10307 & ~n27030 ) | ( n15657 & ~n27030 ) ;
  assign n27032 = n25623 ^ n8880 ^ 1'b0 ;
  assign n27033 = ~n2435 & n9955 ;
  assign n27034 = n27033 ^ n8458 ^ 1'b0 ;
  assign n27035 = n2007 & n27034 ;
  assign n27036 = n7642 ^ n1410 ^ x15 ;
  assign n27037 = n27035 & ~n27036 ;
  assign n27038 = n13466 ^ n7659 ^ 1'b0 ;
  assign n27039 = n27037 & n27038 ;
  assign n27040 = n27039 ^ n20910 ^ 1'b0 ;
  assign n27041 = n1906 | n11226 ;
  assign n27042 = n27041 ^ n3813 ^ 1'b0 ;
  assign n27043 = n4155 & n11356 ;
  assign n27044 = n27043 ^ n16446 ^ 1'b0 ;
  assign n27045 = ( n13799 & n27042 ) | ( n13799 & ~n27044 ) | ( n27042 & ~n27044 ) ;
  assign n27046 = ( n267 & ~n5232 ) | ( n267 & n14535 ) | ( ~n5232 & n14535 ) ;
  assign n27047 = n3319 | n27046 ;
  assign n27048 = n27047 ^ n11816 ^ n2725 ;
  assign n27049 = n11904 & n27048 ;
  assign n27050 = ( n6880 & n27045 ) | ( n6880 & ~n27049 ) | ( n27045 & ~n27049 ) ;
  assign n27051 = n19459 ^ n4878 ^ n2797 ;
  assign n27052 = n22885 ^ n10808 ^ n4069 ;
  assign n27053 = ( n12089 & n20933 ) | ( n12089 & ~n27052 ) | ( n20933 & ~n27052 ) ;
  assign n27054 = ( n2999 & n14755 ) | ( n2999 & n15446 ) | ( n14755 & n15446 ) ;
  assign n27055 = n27054 ^ n15905 ^ n1276 ;
  assign n27058 = n14684 ^ n1626 ^ 1'b0 ;
  assign n27059 = n2406 | n27058 ;
  assign n27060 = ( n2627 & n8061 ) | ( n2627 & ~n27059 ) | ( n8061 & ~n27059 ) ;
  assign n27057 = ( n1757 & ~n4597 ) | ( n1757 & n16168 ) | ( ~n4597 & n16168 ) ;
  assign n27061 = n27060 ^ n27057 ^ n2652 ;
  assign n27056 = n8709 & n14332 ;
  assign n27062 = n27061 ^ n27056 ^ 1'b0 ;
  assign n27063 = ( n5376 & n20274 ) | ( n5376 & n20331 ) | ( n20274 & n20331 ) ;
  assign n27064 = n17188 ^ n726 ^ 1'b0 ;
  assign n27065 = n8339 & n27064 ;
  assign n27066 = n27065 ^ n11663 ^ n1860 ;
  assign n27067 = n27066 ^ n15362 ^ 1'b0 ;
  assign n27068 = n16542 & n27067 ;
  assign n27069 = ( ~n25559 & n27063 ) | ( ~n25559 & n27068 ) | ( n27063 & n27068 ) ;
  assign n27070 = ( n7228 & n10259 ) | ( n7228 & ~n16963 ) | ( n10259 & ~n16963 ) ;
  assign n27071 = ~n1061 & n1538 ;
  assign n27072 = n27071 ^ n7952 ^ 1'b0 ;
  assign n27073 = ( ~n4880 & n12995 ) | ( ~n4880 & n27072 ) | ( n12995 & n27072 ) ;
  assign n27074 = ( n7050 & ~n27070 ) | ( n7050 & n27073 ) | ( ~n27070 & n27073 ) ;
  assign n27075 = ( ~n11428 & n24638 ) | ( ~n11428 & n27074 ) | ( n24638 & n27074 ) ;
  assign n27076 = n8066 & n8922 ;
  assign n27077 = n27076 ^ n24731 ^ x50 ;
  assign n27078 = n26234 ^ n17128 ^ 1'b0 ;
  assign n27079 = ( n9866 & n13114 ) | ( n9866 & ~n13497 ) | ( n13114 & ~n13497 ) ;
  assign n27080 = n27079 ^ n20391 ^ n12953 ;
  assign n27081 = ~n23473 & n27080 ;
  assign n27082 = n15632 ^ n4694 ^ n2740 ;
  assign n27083 = n6608 & n13988 ;
  assign n27084 = ( n1708 & n12414 ) | ( n1708 & ~n27083 ) | ( n12414 & ~n27083 ) ;
  assign n27085 = n2942 & n27084 ;
  assign n27086 = ( n2070 & n6981 ) | ( n2070 & ~n20062 ) | ( n6981 & ~n20062 ) ;
  assign n27087 = n27086 ^ n23427 ^ n4507 ;
  assign n27089 = n23801 ^ n3350 ^ 1'b0 ;
  assign n27090 = n10219 | n27089 ;
  assign n27088 = n12443 & n16093 ;
  assign n27091 = n27090 ^ n27088 ^ 1'b0 ;
  assign n27092 = ( n14543 & n23334 ) | ( n14543 & n27091 ) | ( n23334 & n27091 ) ;
  assign n27093 = ( n12264 & n17183 ) | ( n12264 & n27092 ) | ( n17183 & n27092 ) ;
  assign n27094 = n15889 ^ n13134 ^ n9364 ;
  assign n27095 = n4135 & ~n27094 ;
  assign n27096 = ~n16401 & n27095 ;
  assign n27097 = ( n1997 & n9502 ) | ( n1997 & n27096 ) | ( n9502 & n27096 ) ;
  assign n27098 = n9694 & ~n23351 ;
  assign n27099 = ~n815 & n27098 ;
  assign n27100 = n16222 | n27099 ;
  assign n27101 = n15034 | n27100 ;
  assign n27102 = n14613 ^ n12646 ^ n6457 ;
  assign n27103 = ( n2579 & n19941 ) | ( n2579 & ~n21169 ) | ( n19941 & ~n21169 ) ;
  assign n27104 = ( n5917 & ~n7842 ) | ( n5917 & n21920 ) | ( ~n7842 & n21920 ) ;
  assign n27105 = ~n27103 & n27104 ;
  assign n27106 = n11299 | n13674 ;
  assign n27107 = n27106 ^ n2897 ^ 1'b0 ;
  assign n27108 = n14964 ^ n9408 ^ n890 ;
  assign n27109 = ( n1682 & n2752 ) | ( n1682 & ~n27108 ) | ( n2752 & ~n27108 ) ;
  assign n27110 = n22358 ^ n14233 ^ n1272 ;
  assign n27111 = ( ~n3694 & n10658 ) | ( ~n3694 & n27110 ) | ( n10658 & n27110 ) ;
  assign n27112 = n16559 ^ n5966 ^ 1'b0 ;
  assign n27113 = ~n4026 & n18044 ;
  assign n27114 = ~n3350 & n27113 ;
  assign n27115 = n27112 & ~n27114 ;
  assign n27116 = n27115 ^ n7527 ^ 1'b0 ;
  assign n27121 = n19969 ^ n13076 ^ n8777 ;
  assign n27120 = n14813 ^ n6840 ^ n557 ;
  assign n27122 = n27121 ^ n27120 ^ n14742 ;
  assign n27118 = n21388 ^ n16083 ^ n11605 ;
  assign n27117 = n7386 & ~n17500 ;
  assign n27119 = n27118 ^ n27117 ^ n11959 ;
  assign n27123 = n27122 ^ n27119 ^ n10477 ;
  assign n27124 = n11429 & ~n22489 ;
  assign n27125 = n2892 & n6732 ;
  assign n27126 = ( n12711 & n19496 ) | ( n12711 & ~n27125 ) | ( n19496 & ~n27125 ) ;
  assign n27127 = n3038 & ~n9017 ;
  assign n27128 = ~n19793 & n27127 ;
  assign n27129 = n895 & ~n27128 ;
  assign n27130 = n27129 ^ n1229 ^ 1'b0 ;
  assign n27131 = n8660 & ~n27130 ;
  assign n27132 = n16485 ^ n13076 ^ 1'b0 ;
  assign n27133 = n11306 & n27132 ;
  assign n27134 = ( n766 & n2859 ) | ( n766 & n22092 ) | ( n2859 & n22092 ) ;
  assign n27135 = ( n5675 & n22770 ) | ( n5675 & n27134 ) | ( n22770 & n27134 ) ;
  assign n27136 = n4110 ^ n3229 ^ x212 ;
  assign n27137 = n3161 | n27136 ;
  assign n27138 = n27135 | n27137 ;
  assign n27143 = n20255 ^ n7290 ^ n1101 ;
  assign n27139 = n12403 ^ n7093 ^ 1'b0 ;
  assign n27140 = n9027 & n27139 ;
  assign n27141 = n27140 ^ n18348 ^ n3021 ;
  assign n27142 = n14155 & ~n27141 ;
  assign n27144 = n27143 ^ n27142 ^ n8096 ;
  assign n27145 = n10578 & n18268 ;
  assign n27147 = n1791 | n18838 ;
  assign n27146 = n9105 & ~n18258 ;
  assign n27148 = n27147 ^ n27146 ^ n25996 ;
  assign n27149 = ( n3766 & n3804 ) | ( n3766 & ~n7774 ) | ( n3804 & ~n7774 ) ;
  assign n27150 = n4916 & ~n27149 ;
  assign n27151 = n24990 ^ n1194 ^ 1'b0 ;
  assign n27152 = ~n27150 & n27151 ;
  assign n27153 = ~n412 & n2195 ;
  assign n27154 = n27153 ^ n6971 ^ 1'b0 ;
  assign n27155 = n24389 ^ n12340 ^ n710 ;
  assign n27156 = n7957 & n27155 ;
  assign n27157 = ~n19355 & n27156 ;
  assign n27158 = ( n6857 & ~n10928 ) | ( n6857 & n27157 ) | ( ~n10928 & n27157 ) ;
  assign n27159 = ( n4025 & ~n5113 ) | ( n4025 & n24701 ) | ( ~n5113 & n24701 ) ;
  assign n27160 = n3287 & ~n6272 ;
  assign n27161 = ~n8488 & n27160 ;
  assign n27162 = ( n760 & ~n27159 ) | ( n760 & n27161 ) | ( ~n27159 & n27161 ) ;
  assign n27163 = ( ~n4241 & n14406 ) | ( ~n4241 & n17760 ) | ( n14406 & n17760 ) ;
  assign n27164 = n27163 ^ n19671 ^ n13794 ;
  assign n27165 = n3369 | n12095 ;
  assign n27166 = n27165 ^ n16653 ^ 1'b0 ;
  assign n27167 = n27164 | n27166 ;
  assign n27168 = n4563 | n16474 ;
  assign n27169 = n27168 ^ n16420 ^ 1'b0 ;
  assign n27170 = ~n2865 & n3424 ;
  assign n27171 = n27169 & n27170 ;
  assign n27172 = n16894 ^ n5703 ^ 1'b0 ;
  assign n27174 = n9477 ^ n9105 ^ n7067 ;
  assign n27173 = n5983 & ~n10430 ;
  assign n27175 = n27174 ^ n27173 ^ 1'b0 ;
  assign n27176 = ( ~n10914 & n27172 ) | ( ~n10914 & n27175 ) | ( n27172 & n27175 ) ;
  assign n27177 = ( ~n14588 & n27171 ) | ( ~n14588 & n27176 ) | ( n27171 & n27176 ) ;
  assign n27178 = n4800 & n24829 ;
  assign n27179 = n27178 ^ n3171 ^ 1'b0 ;
  assign n27180 = n27179 ^ n22526 ^ n3813 ;
  assign n27181 = n27180 ^ n21950 ^ 1'b0 ;
  assign n27182 = ~n9608 & n25334 ;
  assign n27183 = n1461 | n27182 ;
  assign n27184 = n23663 | n27183 ;
  assign n27185 = ( n1869 & n19713 ) | ( n1869 & n20244 ) | ( n19713 & n20244 ) ;
  assign n27186 = ( n1316 & ~n6494 ) | ( n1316 & n11840 ) | ( ~n6494 & n11840 ) ;
  assign n27187 = n27186 ^ n3740 ^ n1768 ;
  assign n27188 = n15462 ^ n13962 ^ 1'b0 ;
  assign n27189 = n27188 ^ n3971 ^ n1357 ;
  assign n27190 = n24469 ^ n9370 ^ n5100 ;
  assign n27191 = n10617 | n15300 ;
  assign n27192 = n18767 & ~n27191 ;
  assign n27193 = n27192 ^ n14343 ^ n1147 ;
  assign n27194 = ( ~n5680 & n18156 ) | ( ~n5680 & n27193 ) | ( n18156 & n27193 ) ;
  assign n27195 = n22092 ^ n1726 ^ 1'b0 ;
  assign n27196 = n27195 ^ n19831 ^ n4175 ;
  assign n27197 = n18772 & n26549 ;
  assign n27198 = n27196 & n27197 ;
  assign n27199 = n14723 ^ n8984 ^ x72 ;
  assign n27200 = n708 & n27199 ;
  assign n27201 = n27198 & n27200 ;
  assign n27202 = ( n3053 & ~n4906 ) | ( n3053 & n5462 ) | ( ~n4906 & n5462 ) ;
  assign n27203 = n10762 ^ n6207 ^ 1'b0 ;
  assign n27204 = n5686 & ~n27203 ;
  assign n27205 = n27204 ^ n13354 ^ n817 ;
  assign n27206 = n22487 ^ n2967 ^ 1'b0 ;
  assign n27207 = n2995 & ~n27206 ;
  assign n27208 = ~n27205 & n27207 ;
  assign n27209 = n27208 ^ n12999 ^ 1'b0 ;
  assign n27210 = n27209 ^ n1056 ^ 1'b0 ;
  assign n27211 = n3993 & n7882 ;
  assign n27212 = n8946 & n9755 ;
  assign n27213 = ~n19845 & n27212 ;
  assign n27216 = n8694 & ~n14745 ;
  assign n27214 = x55 & n9829 ;
  assign n27215 = ( ~n9634 & n23547 ) | ( ~n9634 & n27214 ) | ( n23547 & n27214 ) ;
  assign n27217 = n27216 ^ n27215 ^ 1'b0 ;
  assign n27218 = n22714 ^ n18797 ^ n17189 ;
  assign n27219 = n27218 ^ n25272 ^ n6653 ;
  assign n27220 = ( n925 & ~n16338 ) | ( n925 & n16495 ) | ( ~n16338 & n16495 ) ;
  assign n27221 = n27220 ^ n21552 ^ n3694 ;
  assign n27222 = n27221 ^ n935 ^ n667 ;
  assign n27223 = n1720 ^ n967 ^ 1'b0 ;
  assign n27224 = ( n877 & n4537 ) | ( n877 & ~n10082 ) | ( n4537 & ~n10082 ) ;
  assign n27225 = n17925 ^ n4567 ^ 1'b0 ;
  assign n27226 = ~n18384 & n27225 ;
  assign n27227 = n27226 ^ n8077 ^ 1'b0 ;
  assign n27228 = n4802 | n27227 ;
  assign n27229 = n17918 ^ n8903 ^ 1'b0 ;
  assign n27230 = n27229 ^ n19838 ^ n934 ;
  assign n27231 = n15684 ^ n8405 ^ 1'b0 ;
  assign n27232 = ( ~n1507 & n4226 ) | ( ~n1507 & n27231 ) | ( n4226 & n27231 ) ;
  assign n27233 = n27232 ^ n9328 ^ n3040 ;
  assign n27234 = n4292 | n10407 ;
  assign n27235 = n4023 | n27234 ;
  assign n27236 = ~n24329 & n27235 ;
  assign n27237 = n2365 | n9561 ;
  assign n27238 = n27237 ^ n26987 ^ n14455 ;
  assign n27239 = n25639 ^ n8184 ^ n3360 ;
  assign n27240 = n27239 ^ n16794 ^ n498 ;
  assign n27241 = n1022 | n10303 ;
  assign n27242 = n883 | n27241 ;
  assign n27243 = n10100 ^ n1278 ^ x62 ;
  assign n27244 = n12949 & n27243 ;
  assign n27245 = n17747 ^ n8714 ^ n3648 ;
  assign n27246 = ( n907 & n21992 ) | ( n907 & n27245 ) | ( n21992 & n27245 ) ;
  assign n27247 = ( ~n27242 & n27244 ) | ( ~n27242 & n27246 ) | ( n27244 & n27246 ) ;
  assign n27248 = n12609 ^ n9886 ^ n9103 ;
  assign n27249 = n19406 & n27248 ;
  assign n27250 = n14195 ^ n10743 ^ n4399 ;
  assign n27251 = n27250 ^ n1060 ^ 1'b0 ;
  assign n27252 = n27111 ^ n18255 ^ 1'b0 ;
  assign n27253 = n27251 | n27252 ;
  assign n27254 = n1728 & n9709 ;
  assign n27255 = n27254 ^ n3167 ^ 1'b0 ;
  assign n27256 = ( ~n2142 & n7123 ) | ( ~n2142 & n27255 ) | ( n7123 & n27255 ) ;
  assign n27257 = n27256 ^ n5302 ^ n2806 ;
  assign n27258 = n27257 ^ n1830 ^ 1'b0 ;
  assign n27262 = n4056 & n13351 ;
  assign n27263 = n27262 ^ n4311 ^ 1'b0 ;
  assign n27264 = ( n947 & n17752 ) | ( n947 & n27263 ) | ( n17752 & n27263 ) ;
  assign n27260 = n10690 & n11219 ;
  assign n27259 = n15213 ^ n11529 ^ n10075 ;
  assign n27261 = n27260 ^ n27259 ^ n3899 ;
  assign n27265 = n27264 ^ n27261 ^ n13394 ;
  assign n27269 = ( n8177 & n10922 ) | ( n8177 & n11621 ) | ( n10922 & n11621 ) ;
  assign n27266 = ~n5654 & n9264 ;
  assign n27267 = n27266 ^ n12790 ^ 1'b0 ;
  assign n27268 = ~n1074 & n27267 ;
  assign n27270 = n27269 ^ n27268 ^ 1'b0 ;
  assign n27271 = ( n910 & n1151 ) | ( n910 & ~n20164 ) | ( n1151 & ~n20164 ) ;
  assign n27272 = n27271 ^ n17470 ^ n6626 ;
  assign n27273 = n27272 ^ n12900 ^ 1'b0 ;
  assign n27278 = n7748 & n7883 ;
  assign n27279 = n27278 ^ n18707 ^ 1'b0 ;
  assign n27274 = n13609 ^ n1505 ^ n1029 ;
  assign n27275 = n24513 & n27274 ;
  assign n27276 = n13777 ^ n3223 ^ n2872 ;
  assign n27277 = ( n3214 & n27275 ) | ( n3214 & n27276 ) | ( n27275 & n27276 ) ;
  assign n27280 = n27279 ^ n27277 ^ n14981 ;
  assign n27281 = ( n1961 & n8335 ) | ( n1961 & n27280 ) | ( n8335 & n27280 ) ;
  assign n27282 = n24104 ^ n3948 ^ 1'b0 ;
  assign n27283 = n1406 ^ n1196 ^ 1'b0 ;
  assign n27284 = n27283 ^ n13851 ^ n13226 ;
  assign n27285 = ( n431 & n6325 ) | ( n431 & ~n21479 ) | ( n6325 & ~n21479 ) ;
  assign n27286 = n11631 | n27285 ;
  assign n27287 = ( n13194 & ~n27284 ) | ( n13194 & n27286 ) | ( ~n27284 & n27286 ) ;
  assign n27288 = ( n10091 & n10822 ) | ( n10091 & n14777 ) | ( n10822 & n14777 ) ;
  assign n27289 = ( n17821 & n24198 ) | ( n17821 & n27288 ) | ( n24198 & n27288 ) ;
  assign n27290 = ( n4631 & n25152 ) | ( n4631 & n27289 ) | ( n25152 & n27289 ) ;
  assign n27291 = n2105 | n27290 ;
  assign n27292 = n3594 | n7809 ;
  assign n27293 = n9097 & ~n27292 ;
  assign n27294 = n27293 ^ n21606 ^ 1'b0 ;
  assign n27295 = n18018 | n27294 ;
  assign n27300 = n2979 & n10739 ;
  assign n27301 = n27300 ^ n12073 ^ 1'b0 ;
  assign n27296 = n10836 ^ n3948 ^ 1'b0 ;
  assign n27297 = n27296 ^ n15838 ^ 1'b0 ;
  assign n27298 = n7672 & n27297 ;
  assign n27299 = n27298 ^ n574 ^ 1'b0 ;
  assign n27302 = n27301 ^ n27299 ^ n7605 ;
  assign n27303 = n27302 ^ n20596 ^ 1'b0 ;
  assign n27304 = n5411 & ~n27303 ;
  assign n27305 = n27304 ^ n18253 ^ n12207 ;
  assign n27306 = ( n6489 & n13533 ) | ( n6489 & n27305 ) | ( n13533 & n27305 ) ;
  assign n27307 = n13094 ^ n3322 ^ 1'b0 ;
  assign n27308 = n2797 ^ n1098 ^ 1'b0 ;
  assign n27309 = n16420 | n27308 ;
  assign n27310 = n9995 | n12694 ;
  assign n27311 = n20127 & ~n27310 ;
  assign n27312 = n1546 ^ x143 ^ 1'b0 ;
  assign n27313 = n27312 ^ n13969 ^ n8297 ;
  assign n27314 = n10794 & ~n24389 ;
  assign n27315 = ( n15002 & n26820 ) | ( n15002 & ~n27314 ) | ( n26820 & ~n27314 ) ;
  assign n27316 = ( ~n478 & n14443 ) | ( ~n478 & n21355 ) | ( n14443 & n21355 ) ;
  assign n27317 = ~n13747 & n20681 ;
  assign n27318 = ( n1916 & n27316 ) | ( n1916 & ~n27317 ) | ( n27316 & ~n27317 ) ;
  assign n27319 = ( n6033 & ~n9326 ) | ( n6033 & n20678 ) | ( ~n9326 & n20678 ) ;
  assign n27320 = n15999 & ~n16250 ;
  assign n27321 = n27320 ^ n9980 ^ 1'b0 ;
  assign n27322 = n23265 ^ n7911 ^ n1457 ;
  assign n27323 = n27322 ^ n23761 ^ n4269 ;
  assign n27324 = n23225 & n27323 ;
  assign n27325 = n27321 & n27324 ;
  assign n27326 = n2302 & n27325 ;
  assign n27327 = n27326 ^ n8342 ^ 1'b0 ;
  assign n27328 = n19645 & ~n27018 ;
  assign n27329 = n27328 ^ n3525 ^ 1'b0 ;
  assign n27330 = n20226 ^ n19158 ^ n7058 ;
  assign n27331 = n3963 ^ n1871 ^ 1'b0 ;
  assign n27332 = n27330 & ~n27331 ;
  assign n27333 = n10939 ^ n10391 ^ n10352 ;
  assign n27334 = n27333 ^ n25914 ^ n8923 ;
  assign n27335 = n27334 ^ n14610 ^ n3505 ;
  assign n27336 = n27335 ^ n2995 ^ 1'b0 ;
  assign n27337 = n19370 ^ n13639 ^ 1'b0 ;
  assign n27338 = n10087 ^ n8371 ^ n6500 ;
  assign n27339 = ~n2432 & n27338 ;
  assign n27340 = n27339 ^ n2199 ^ n1139 ;
  assign n27342 = n25263 ^ n23156 ^ 1'b0 ;
  assign n27343 = n2548 & ~n27342 ;
  assign n27341 = ( n8598 & ~n16831 ) | ( n8598 & n25978 ) | ( ~n16831 & n25978 ) ;
  assign n27344 = n27343 ^ n27341 ^ n19139 ;
  assign n27345 = n19969 ^ n3098 ^ 1'b0 ;
  assign n27346 = ~n19930 & n27345 ;
  assign n27347 = n959 & ~n6241 ;
  assign n27348 = ~n11021 & n27347 ;
  assign n27349 = n4211 | n24751 ;
  assign n27350 = n9689 | n27349 ;
  assign n27351 = n18219 ^ n12977 ^ 1'b0 ;
  assign n27352 = ~n5173 & n27351 ;
  assign n27353 = n27352 ^ n25039 ^ n1002 ;
  assign n27354 = ( ~n8791 & n27350 ) | ( ~n8791 & n27353 ) | ( n27350 & n27353 ) ;
  assign n27355 = ( n7257 & ~n27348 ) | ( n7257 & n27354 ) | ( ~n27348 & n27354 ) ;
  assign n27356 = n27355 ^ n3624 ^ 1'b0 ;
  assign n27357 = n27356 ^ n21109 ^ 1'b0 ;
  assign n27358 = n11626 ^ n10037 ^ n2931 ;
  assign n27359 = ( ~n2110 & n8549 ) | ( ~n2110 & n27358 ) | ( n8549 & n27358 ) ;
  assign n27360 = n12310 ^ n1745 ^ 1'b0 ;
  assign n27362 = ~n2311 & n11051 ;
  assign n27363 = n6771 & n27362 ;
  assign n27361 = n23717 ^ n11220 ^ n7780 ;
  assign n27364 = n27363 ^ n27361 ^ n5596 ;
  assign n27365 = n27364 ^ n3617 ^ 1'b0 ;
  assign n27366 = n9675 | n27365 ;
  assign n27367 = n27366 ^ n7995 ^ 1'b0 ;
  assign n27368 = ~n22142 & n27367 ;
  assign n27369 = n15507 ^ n3107 ^ n2826 ;
  assign n27370 = n27369 ^ n21461 ^ n6049 ;
  assign n27371 = n7395 ^ n3262 ^ n381 ;
  assign n27372 = n27371 ^ n11908 ^ n708 ;
  assign n27373 = ( ~n8889 & n22168 ) | ( ~n8889 & n23184 ) | ( n22168 & n23184 ) ;
  assign n27374 = n19255 ^ n18649 ^ n12394 ;
  assign n27375 = ( n3587 & ~n5959 ) | ( n3587 & n27374 ) | ( ~n5959 & n27374 ) ;
  assign n27376 = n27375 ^ n21262 ^ n9002 ;
  assign n27377 = n22887 ^ n16485 ^ 1'b0 ;
  assign n27378 = n24346 & ~n27377 ;
  assign n27379 = ~n27376 & n27378 ;
  assign n27380 = ~n27373 & n27379 ;
  assign n27381 = ( n7270 & n11710 ) | ( n7270 & n22092 ) | ( n11710 & n22092 ) ;
  assign n27382 = n27381 ^ n12322 ^ 1'b0 ;
  assign n27383 = n27380 | n27382 ;
  assign n27384 = n16882 ^ n10481 ^ n10167 ;
  assign n27385 = n4543 ^ n3890 ^ 1'b0 ;
  assign n27386 = ( n6164 & n10004 ) | ( n6164 & ~n27385 ) | ( n10004 & ~n27385 ) ;
  assign n27387 = n25036 ^ n20651 ^ n17212 ;
  assign n27395 = n10514 & ~n11097 ;
  assign n27393 = n904 & n12360 ;
  assign n27394 = n27393 ^ n3872 ^ 1'b0 ;
  assign n27396 = n27395 ^ n27394 ^ 1'b0 ;
  assign n27388 = n3211 & ~n4155 ;
  assign n27389 = ~n10081 & n27388 ;
  assign n27390 = n22787 ^ n8933 ^ n2753 ;
  assign n27391 = ( n11153 & n27389 ) | ( n11153 & ~n27390 ) | ( n27389 & ~n27390 ) ;
  assign n27392 = n3230 | n27391 ;
  assign n27397 = n27396 ^ n27392 ^ 1'b0 ;
  assign n27398 = n27397 ^ n24626 ^ n12853 ;
  assign n27399 = n10085 ^ n8395 ^ 1'b0 ;
  assign n27400 = n11697 ^ n8980 ^ n8501 ;
  assign n27401 = n27400 ^ n15957 ^ 1'b0 ;
  assign n27402 = n21528 & n27401 ;
  assign n27403 = ~n27399 & n27402 ;
  assign n27404 = ( n4316 & n8363 ) | ( n4316 & n10389 ) | ( n8363 & n10389 ) ;
  assign n27405 = n11067 & ~n17476 ;
  assign n27406 = n27405 ^ n13862 ^ n5381 ;
  assign n27407 = ( n1066 & ~n27404 ) | ( n1066 & n27406 ) | ( ~n27404 & n27406 ) ;
  assign n27408 = n9477 | n27407 ;
  assign n27409 = n7420 | n27408 ;
  assign n27410 = n21369 ^ n9111 ^ 1'b0 ;
  assign n27413 = n3235 & n13913 ;
  assign n27414 = ~n1828 & n27413 ;
  assign n27415 = n27414 ^ n8397 ^ n8233 ;
  assign n27416 = n27415 ^ n20022 ^ 1'b0 ;
  assign n27412 = n8601 & ~n13186 ;
  assign n27417 = n27416 ^ n27412 ^ 1'b0 ;
  assign n27411 = n3764 & n25050 ;
  assign n27418 = n27417 ^ n27411 ^ 1'b0 ;
  assign n27419 = n18491 & n27348 ;
  assign n27420 = n27419 ^ n5396 ^ 1'b0 ;
  assign n27421 = ( ~n12997 & n17182 ) | ( ~n12997 & n19677 ) | ( n17182 & n19677 ) ;
  assign n27422 = n27421 ^ n5065 ^ 1'b0 ;
  assign n27423 = n711 & n27422 ;
  assign n27424 = n10784 & n27423 ;
  assign n27425 = ( n2736 & n7792 ) | ( n2736 & ~n16254 ) | ( n7792 & ~n16254 ) ;
  assign n27426 = n18971 ^ n17470 ^ 1'b0 ;
  assign n27427 = n27425 | n27426 ;
  assign n27428 = ( n6972 & n27424 ) | ( n6972 & n27427 ) | ( n27424 & n27427 ) ;
  assign n27429 = n22562 & n27428 ;
  assign n27430 = n13212 ^ n2101 ^ n1002 ;
  assign n27431 = n25413 ^ n11759 ^ n3629 ;
  assign n27432 = ( ~n18665 & n27430 ) | ( ~n18665 & n27431 ) | ( n27430 & n27431 ) ;
  assign n27433 = n27432 ^ n24849 ^ n10352 ;
  assign n27434 = n15038 ^ n8904 ^ 1'b0 ;
  assign n27435 = n25374 ^ n3611 ^ 1'b0 ;
  assign n27436 = n2139 & n27435 ;
  assign n27437 = n27434 & n27436 ;
  assign n27439 = n10507 & ~n20776 ;
  assign n27440 = ~n8220 & n27439 ;
  assign n27438 = n7333 ^ n1459 ^ 1'b0 ;
  assign n27441 = n27440 ^ n27438 ^ n7415 ;
  assign n27442 = n6730 & n15047 ;
  assign n27443 = ~n15449 & n27442 ;
  assign n27444 = ( n4886 & n13725 ) | ( n4886 & n18923 ) | ( n13725 & n18923 ) ;
  assign n27445 = n27444 ^ n13011 ^ 1'b0 ;
  assign n27446 = n23571 & n27445 ;
  assign n27447 = n27446 ^ n10227 ^ n8703 ;
  assign n27448 = n19561 & n27447 ;
  assign n27449 = ( n1680 & n27443 ) | ( n1680 & ~n27448 ) | ( n27443 & ~n27448 ) ;
  assign n27451 = ( n5196 & n9763 ) | ( n5196 & ~n19159 ) | ( n9763 & ~n19159 ) ;
  assign n27450 = n15515 & ~n20540 ;
  assign n27452 = n27451 ^ n27450 ^ 1'b0 ;
  assign n27454 = n13516 ^ n8889 ^ n7715 ;
  assign n27455 = n27454 ^ n8193 ^ 1'b0 ;
  assign n27453 = n23601 ^ n4438 ^ 1'b0 ;
  assign n27456 = n27455 ^ n27453 ^ x103 ;
  assign n27457 = ( n1126 & n2271 ) | ( n1126 & ~n13554 ) | ( n2271 & ~n13554 ) ;
  assign n27458 = n27457 ^ n14383 ^ n10189 ;
  assign n27459 = n27456 & ~n27458 ;
  assign n27460 = ( ~n4563 & n17550 ) | ( ~n4563 & n22095 ) | ( n17550 & n22095 ) ;
  assign n27461 = n27460 ^ n715 ^ 1'b0 ;
  assign n27462 = ( n768 & n4054 ) | ( n768 & ~n16354 ) | ( n4054 & ~n16354 ) ;
  assign n27463 = ( n2472 & ~n8573 ) | ( n2472 & n27462 ) | ( ~n8573 & n27462 ) ;
  assign n27464 = ( ~n570 & n668 ) | ( ~n570 & n3017 ) | ( n668 & n3017 ) ;
  assign n27465 = n1112 & ~n27464 ;
  assign n27466 = n2926 ^ n834 ^ 1'b0 ;
  assign n27467 = ( ~n23099 & n24903 ) | ( ~n23099 & n27466 ) | ( n24903 & n27466 ) ;
  assign n27468 = ( ~n3890 & n6945 ) | ( ~n3890 & n7920 ) | ( n6945 & n7920 ) ;
  assign n27469 = n3704 & ~n27468 ;
  assign n27470 = n18633 & n27469 ;
  assign n27471 = n18643 ^ n13878 ^ x178 ;
  assign n27472 = n27471 ^ n3170 ^ 1'b0 ;
  assign n27473 = n10444 & ~n21143 ;
  assign n27474 = ~n13450 & n27473 ;
  assign n27475 = n21477 ^ n2750 ^ 1'b0 ;
  assign n27476 = n27474 | n27475 ;
  assign n27477 = n27476 ^ n12596 ^ n3824 ;
  assign n27478 = ( n12456 & n20022 ) | ( n12456 & ~n21102 ) | ( n20022 & ~n21102 ) ;
  assign n27479 = n27478 ^ n17138 ^ 1'b0 ;
  assign n27480 = n15651 ^ n8990 ^ n271 ;
  assign n27481 = n26027 ^ n18298 ^ n15293 ;
  assign n27482 = n27481 ^ n14946 ^ n393 ;
  assign n27483 = ( n2638 & n27480 ) | ( n2638 & n27482 ) | ( n27480 & n27482 ) ;
  assign n27484 = n12611 & ~n16680 ;
  assign n27485 = n27484 ^ n23067 ^ n10373 ;
  assign n27486 = n27485 ^ n25653 ^ n22250 ;
  assign n27487 = n9712 & ~n27486 ;
  assign n27488 = ~n5203 & n27487 ;
  assign n27489 = n16083 & n21584 ;
  assign n27490 = n27489 ^ n13900 ^ 1'b0 ;
  assign n27491 = ( n622 & n7939 ) | ( n622 & n22039 ) | ( n7939 & n22039 ) ;
  assign n27492 = ( ~n7497 & n20606 ) | ( ~n7497 & n27491 ) | ( n20606 & n27491 ) ;
  assign n27493 = n16990 ^ n15178 ^ n11587 ;
  assign n27494 = n3399 | n27493 ;
  assign n27495 = n8688 | n10694 ;
  assign n27496 = n8072 & ~n27495 ;
  assign n27497 = n27496 ^ n12876 ^ 1'b0 ;
  assign n27498 = n27494 & n27497 ;
  assign n27499 = ( ~n2152 & n12802 ) | ( ~n2152 & n27498 ) | ( n12802 & n27498 ) ;
  assign n27500 = ( x197 & n18856 ) | ( x197 & n27499 ) | ( n18856 & n27499 ) ;
  assign n27501 = ( n12107 & n16990 ) | ( n12107 & n17608 ) | ( n16990 & n17608 ) ;
  assign n27502 = n27501 ^ n13548 ^ n781 ;
  assign n27503 = ( n2987 & ~n5080 ) | ( n2987 & n15491 ) | ( ~n5080 & n15491 ) ;
  assign n27504 = ( n6378 & n15017 ) | ( n6378 & ~n27503 ) | ( n15017 & ~n27503 ) ;
  assign n27505 = n27504 ^ n22969 ^ n14684 ;
  assign n27506 = ( n8226 & n18406 ) | ( n8226 & n27505 ) | ( n18406 & n27505 ) ;
  assign n27507 = n15980 ^ n6461 ^ 1'b0 ;
  assign n27508 = ~n20744 & n27507 ;
  assign n27509 = ~n24572 & n27508 ;
  assign n27510 = ~n27506 & n27509 ;
  assign n27512 = ( ~n2214 & n5722 ) | ( ~n2214 & n27047 ) | ( n5722 & n27047 ) ;
  assign n27511 = ~n13969 & n22485 ;
  assign n27513 = n27512 ^ n27511 ^ n18642 ;
  assign n27514 = n27513 ^ n17112 ^ 1'b0 ;
  assign n27515 = n11873 & n23091 ;
  assign n27516 = ( x56 & n3104 ) | ( x56 & n27515 ) | ( n3104 & n27515 ) ;
  assign n27517 = n8444 | n9312 ;
  assign n27518 = n27517 ^ n14127 ^ 1'b0 ;
  assign n27519 = n805 & n5196 ;
  assign n27520 = n27519 ^ n9780 ^ 1'b0 ;
  assign n27521 = n27520 ^ n25847 ^ 1'b0 ;
  assign n27522 = n27518 | n27521 ;
  assign n27523 = n20448 ^ n18374 ^ n6883 ;
  assign n27524 = ( n975 & ~n27522 ) | ( n975 & n27523 ) | ( ~n27522 & n27523 ) ;
  assign n27525 = n14844 ^ n2031 ^ 1'b0 ;
  assign n27526 = n10836 ^ n2622 ^ 1'b0 ;
  assign n27527 = n27526 ^ n16752 ^ 1'b0 ;
  assign n27528 = n27527 ^ n9084 ^ 1'b0 ;
  assign n27529 = ~n4608 & n27528 ;
  assign n27530 = n27394 ^ n26096 ^ n12900 ;
  assign n27531 = n19319 | n23707 ;
  assign n27532 = n27531 ^ n11472 ^ n407 ;
  assign n27533 = n25554 ^ n14137 ^ n8781 ;
  assign n27534 = n27533 ^ n18349 ^ n1499 ;
  assign n27535 = n1258 | n9164 ;
  assign n27536 = n27535 ^ n25049 ^ 1'b0 ;
  assign n27537 = n3259 & ~n6976 ;
  assign n27541 = n10501 ^ n9180 ^ 1'b0 ;
  assign n27542 = ~n16782 & n27541 ;
  assign n27543 = n9600 | n27542 ;
  assign n27538 = n22363 ^ n13436 ^ n8730 ;
  assign n27539 = n21787 ^ n19124 ^ 1'b0 ;
  assign n27540 = n27538 | n27539 ;
  assign n27544 = n27543 ^ n27540 ^ n11417 ;
  assign n27545 = n6997 ^ n942 ^ 1'b0 ;
  assign n27546 = n10521 & ~n27545 ;
  assign n27547 = n27546 ^ n13104 ^ n9128 ;
  assign n27548 = ( n11356 & n11955 ) | ( n11356 & n27547 ) | ( n11955 & n27547 ) ;
  assign n27549 = n27548 ^ n14152 ^ n13763 ;
  assign n27550 = n17081 & ~n20735 ;
  assign n27553 = n14081 ^ n12675 ^ n1091 ;
  assign n27551 = n24777 ^ n6477 ^ n5576 ;
  assign n27552 = ( n1643 & n23815 ) | ( n1643 & ~n27551 ) | ( n23815 & ~n27551 ) ;
  assign n27554 = n27553 ^ n27552 ^ n9852 ;
  assign n27555 = ( n12857 & ~n17604 ) | ( n12857 & n27554 ) | ( ~n17604 & n27554 ) ;
  assign n27556 = n27550 & ~n27555 ;
  assign n27557 = ~n8564 & n20924 ;
  assign n27558 = n27557 ^ n13471 ^ 1'b0 ;
  assign n27559 = n19267 ^ n10507 ^ n10142 ;
  assign n27560 = n27559 ^ n14685 ^ n7432 ;
  assign n27561 = n27558 & ~n27560 ;
  assign n27562 = n13444 & n27561 ;
  assign n27563 = n15371 & ~n23669 ;
  assign n27564 = n18670 & n27563 ;
  assign n27565 = n10762 & ~n27564 ;
  assign n27566 = n10698 ^ n7911 ^ n4250 ;
  assign n27567 = n27206 ^ n6042 ^ n3902 ;
  assign n27568 = n18626 | n27567 ;
  assign n27569 = n27566 & ~n27568 ;
  assign n27571 = n10635 | n24516 ;
  assign n27572 = n27571 ^ n23806 ^ 1'b0 ;
  assign n27570 = n8105 | n20497 ;
  assign n27573 = n27572 ^ n27570 ^ 1'b0 ;
  assign n27574 = ( x100 & n2584 ) | ( x100 & n5888 ) | ( n2584 & n5888 ) ;
  assign n27575 = n8462 & n9359 ;
  assign n27576 = n27575 ^ x104 ^ 1'b0 ;
  assign n27577 = ( ~n19050 & n24486 ) | ( ~n19050 & n27576 ) | ( n24486 & n27576 ) ;
  assign n27578 = n27574 | n27577 ;
  assign n27579 = ( x3 & n22790 ) | ( x3 & n27578 ) | ( n22790 & n27578 ) ;
  assign n27580 = n20985 ^ n6101 ^ 1'b0 ;
  assign n27588 = ( x56 & n2194 ) | ( x56 & n9271 ) | ( n2194 & n9271 ) ;
  assign n27581 = n3180 ^ n2036 ^ n859 ;
  assign n27582 = ~n18778 & n27581 ;
  assign n27583 = n27582 ^ n6888 ^ n6300 ;
  assign n27584 = n7611 ^ n3949 ^ n2143 ;
  assign n27585 = ( n2688 & n5813 ) | ( n2688 & n27584 ) | ( n5813 & n27584 ) ;
  assign n27586 = n27583 | n27585 ;
  assign n27587 = n1316 | n27586 ;
  assign n27589 = n27588 ^ n27587 ^ n4077 ;
  assign n27593 = n13496 ^ n11868 ^ n8246 ;
  assign n27592 = n10525 ^ n9898 ^ n3914 ;
  assign n27590 = n25023 ^ n18946 ^ n11404 ;
  assign n27591 = n27590 ^ n11232 ^ n1735 ;
  assign n27594 = n27593 ^ n27592 ^ n27591 ;
  assign n27595 = ( ~n1169 & n4923 ) | ( ~n1169 & n7415 ) | ( n4923 & n7415 ) ;
  assign n27596 = n27595 ^ n18772 ^ n14537 ;
  assign n27604 = ( n7120 & ~n7867 ) | ( n7120 & n27243 ) | ( ~n7867 & n27243 ) ;
  assign n27599 = n18506 ^ n12438 ^ n6609 ;
  assign n27600 = ( n6368 & ~n7057 ) | ( n6368 & n12852 ) | ( ~n7057 & n12852 ) ;
  assign n27601 = n27599 & ~n27600 ;
  assign n27602 = n15768 & n27601 ;
  assign n27597 = n20523 ^ n12719 ^ 1'b0 ;
  assign n27598 = n10411 & ~n27597 ;
  assign n27603 = n27602 ^ n27598 ^ 1'b0 ;
  assign n27605 = n27604 ^ n27603 ^ 1'b0 ;
  assign n27606 = n6843 | n24407 ;
  assign n27607 = n14526 & ~n27606 ;
  assign n27608 = n12989 & ~n27607 ;
  assign n27609 = n27608 ^ n5164 ^ 1'b0 ;
  assign n27610 = n9237 ^ n406 ^ 1'b0 ;
  assign n27611 = n1530 | n27610 ;
  assign n27612 = ( ~n408 & n8315 ) | ( ~n408 & n27515 ) | ( n8315 & n27515 ) ;
  assign n27613 = ( n26298 & n26633 ) | ( n26298 & ~n27612 ) | ( n26633 & ~n27612 ) ;
  assign n27614 = n26637 ^ n15728 ^ n9105 ;
  assign n27615 = n27614 ^ n23965 ^ n1659 ;
  assign n27616 = x91 & ~n7197 ;
  assign n27617 = n12696 ^ n5526 ^ 1'b0 ;
  assign n27618 = n27617 ^ n15515 ^ n9272 ;
  assign n27619 = n10434 & n27618 ;
  assign n27620 = ~n9185 & n10571 ;
  assign n27621 = n27620 ^ n8235 ^ 1'b0 ;
  assign n27622 = ( ~n715 & n27619 ) | ( ~n715 & n27621 ) | ( n27619 & n27621 ) ;
  assign n27623 = n27622 ^ n2717 ^ 1'b0 ;
  assign n27624 = n17845 | n27623 ;
  assign n27625 = n3812 & n6205 ;
  assign n27626 = n27625 ^ n10900 ^ n3182 ;
  assign n27627 = ~n21412 & n27626 ;
  assign n27628 = n27627 ^ n1645 ^ 1'b0 ;
  assign n27629 = ( ~n11913 & n15553 ) | ( ~n11913 & n23635 ) | ( n15553 & n23635 ) ;
  assign n27636 = n18920 ^ n13634 ^ n903 ;
  assign n27631 = n897 | n2523 ;
  assign n27632 = n27631 ^ n5098 ^ 1'b0 ;
  assign n27633 = n2310 ^ n1156 ^ 1'b0 ;
  assign n27634 = n5437 & ~n27633 ;
  assign n27635 = ( n20256 & n27632 ) | ( n20256 & ~n27634 ) | ( n27632 & ~n27634 ) ;
  assign n27637 = n27636 ^ n27635 ^ n19401 ;
  assign n27638 = ( n13356 & ~n24019 ) | ( n13356 & n27637 ) | ( ~n24019 & n27637 ) ;
  assign n27630 = ( n2164 & ~n14268 ) | ( n2164 & n16882 ) | ( ~n14268 & n16882 ) ;
  assign n27639 = n27638 ^ n27630 ^ n11859 ;
  assign n27640 = n17740 ^ n7351 ^ n3077 ;
  assign n27641 = n27640 ^ n8984 ^ n6481 ;
  assign n27642 = ( n2257 & ~n6007 ) | ( n2257 & n16517 ) | ( ~n6007 & n16517 ) ;
  assign n27643 = n5232 & n15405 ;
  assign n27644 = n27643 ^ n19893 ^ 1'b0 ;
  assign n27645 = n27644 ^ n19040 ^ n12859 ;
  assign n27646 = ~n22795 & n27645 ;
  assign n27647 = n4116 & n27646 ;
  assign n27648 = n14332 ^ n12818 ^ 1'b0 ;
  assign n27649 = n9391 ^ x132 ^ 1'b0 ;
  assign n27650 = ( ~x45 & n3983 ) | ( ~x45 & n16170 ) | ( n3983 & n16170 ) ;
  assign n27651 = n6980 ^ n2758 ^ 1'b0 ;
  assign n27652 = n2280 & n27651 ;
  assign n27653 = ( n4331 & ~n18110 ) | ( n4331 & n27652 ) | ( ~n18110 & n27652 ) ;
  assign n27654 = n18944 ^ n7378 ^ n4670 ;
  assign n27655 = ( n23250 & ~n27653 ) | ( n23250 & n27654 ) | ( ~n27653 & n27654 ) ;
  assign n27656 = n18972 & n27655 ;
  assign n27657 = ~n27650 & n27656 ;
  assign n27658 = ( n1979 & ~n5124 ) | ( n1979 & n9907 ) | ( ~n5124 & n9907 ) ;
  assign n27659 = ~n2157 & n27658 ;
  assign n27660 = ~n1879 & n27659 ;
  assign n27661 = n27660 ^ n25097 ^ 1'b0 ;
  assign n27662 = ( n11470 & n11576 ) | ( n11470 & ~n26718 ) | ( n11576 & ~n26718 ) ;
  assign n27663 = n9418 & ~n27662 ;
  assign n27664 = n4879 & n27663 ;
  assign n27665 = ( n18337 & ~n20891 ) | ( n18337 & n27664 ) | ( ~n20891 & n27664 ) ;
  assign n27666 = ~n14193 & n21306 ;
  assign n27667 = ( ~n11409 & n15065 ) | ( ~n11409 & n24562 ) | ( n15065 & n24562 ) ;
  assign n27668 = ( n2501 & n24546 ) | ( n2501 & ~n27667 ) | ( n24546 & ~n27667 ) ;
  assign n27669 = n14544 ^ n1057 ^ n628 ;
  assign n27670 = n25030 & ~n27669 ;
  assign n27671 = ~n6260 & n27670 ;
  assign n27672 = ( n799 & n12926 ) | ( n799 & n14687 ) | ( n12926 & n14687 ) ;
  assign n27673 = n24487 & n27672 ;
  assign n27674 = ( n683 & n27671 ) | ( n683 & n27673 ) | ( n27671 & n27673 ) ;
  assign n27675 = n17718 ^ n6981 ^ n4904 ;
  assign n27676 = ( n306 & n9047 ) | ( n306 & n20293 ) | ( n9047 & n20293 ) ;
  assign n27677 = n24234 ^ n6951 ^ n3487 ;
  assign n27678 = ( n1942 & n27676 ) | ( n1942 & n27677 ) | ( n27676 & n27677 ) ;
  assign n27679 = n27678 ^ n22886 ^ 1'b0 ;
  assign n27680 = ~n18203 & n18711 ;
  assign n27681 = ~n13012 & n27680 ;
  assign n27685 = n23192 ^ n20687 ^ 1'b0 ;
  assign n27682 = ~n2958 & n4605 ;
  assign n27683 = n27682 ^ n1539 ^ 1'b0 ;
  assign n27684 = n27683 ^ n5313 ^ 1'b0 ;
  assign n27686 = n27685 ^ n27684 ^ n10853 ;
  assign n27691 = ( ~n10584 & n13744 ) | ( ~n10584 & n26889 ) | ( n13744 & n26889 ) ;
  assign n27692 = n27691 ^ n4447 ^ 1'b0 ;
  assign n27687 = n7848 ^ n7353 ^ x188 ;
  assign n27688 = ( n2324 & n15507 ) | ( n2324 & ~n27687 ) | ( n15507 & ~n27687 ) ;
  assign n27689 = n27688 ^ n14470 ^ n4639 ;
  assign n27690 = ( n15978 & n25128 ) | ( n15978 & ~n27689 ) | ( n25128 & ~n27689 ) ;
  assign n27693 = n27692 ^ n27690 ^ n27496 ;
  assign n27694 = n15096 ^ n6495 ^ 1'b0 ;
  assign n27695 = n11206 | n27694 ;
  assign n27696 = n18467 ^ n8254 ^ 1'b0 ;
  assign n27697 = ~n27695 & n27696 ;
  assign n27698 = n27697 ^ n23237 ^ n15875 ;
  assign n27699 = n17232 ^ n2379 ^ n1942 ;
  assign n27700 = ~n2081 & n27699 ;
  assign n27701 = n27700 ^ n12468 ^ 1'b0 ;
  assign n27707 = n9706 & n14197 ;
  assign n27708 = n9335 & n27707 ;
  assign n27706 = n17835 ^ n1957 ^ 1'b0 ;
  assign n27709 = n27708 ^ n27706 ^ n25368 ;
  assign n27702 = n14364 ^ n5494 ^ n4605 ;
  assign n27703 = n15919 ^ n6801 ^ n639 ;
  assign n27704 = ( n19002 & n27702 ) | ( n19002 & ~n27703 ) | ( n27702 & ~n27703 ) ;
  assign n27705 = ( n2470 & n18056 ) | ( n2470 & n27704 ) | ( n18056 & n27704 ) ;
  assign n27710 = n27709 ^ n27705 ^ n21407 ;
  assign n27711 = n16054 | n26712 ;
  assign n27712 = n27711 ^ n3445 ^ 1'b0 ;
  assign n27713 = ( n1646 & ~n2888 ) | ( n1646 & n10574 ) | ( ~n2888 & n10574 ) ;
  assign n27714 = ~n3024 & n4407 ;
  assign n27715 = ( n9403 & n13000 ) | ( n9403 & ~n27714 ) | ( n13000 & ~n27714 ) ;
  assign n27716 = ( n16689 & n24317 ) | ( n16689 & n27715 ) | ( n24317 & n27715 ) ;
  assign n27717 = ( n1477 & n6575 ) | ( n1477 & ~n27716 ) | ( n6575 & ~n27716 ) ;
  assign n27718 = n783 | n3551 ;
  assign n27720 = n17908 ^ n12764 ^ n8061 ;
  assign n27719 = ( n9338 & n9668 ) | ( n9338 & ~n23987 ) | ( n9668 & ~n23987 ) ;
  assign n27721 = n27720 ^ n27719 ^ 1'b0 ;
  assign n27722 = ( n22174 & n27718 ) | ( n22174 & n27721 ) | ( n27718 & n27721 ) ;
  assign n27723 = n681 ^ n441 ^ x152 ;
  assign n27724 = ~n11969 & n27723 ;
  assign n27725 = ~n11140 & n27724 ;
  assign n27726 = ( n4852 & ~n10880 ) | ( n4852 & n27725 ) | ( ~n10880 & n27725 ) ;
  assign n27727 = ( n1856 & ~n7297 ) | ( n1856 & n27726 ) | ( ~n7297 & n27726 ) ;
  assign n27728 = n13878 ^ n7924 ^ n1496 ;
  assign n27729 = ( n10745 & n13336 ) | ( n10745 & ~n27728 ) | ( n13336 & ~n27728 ) ;
  assign n27730 = n27729 ^ n7062 ^ n2857 ;
  assign n27731 = n9274 & ~n13361 ;
  assign n27732 = ( n502 & n4136 ) | ( n502 & n7238 ) | ( n4136 & n7238 ) ;
  assign n27733 = ( ~n6587 & n27731 ) | ( ~n6587 & n27732 ) | ( n27731 & n27732 ) ;
  assign n27734 = n27733 ^ n14030 ^ n12015 ;
  assign n27735 = ( n25329 & n27730 ) | ( n25329 & ~n27734 ) | ( n27730 & ~n27734 ) ;
  assign n27736 = n8780 ^ n423 ^ n376 ;
  assign n27737 = n27736 ^ n17482 ^ n5465 ;
  assign n27738 = n27737 ^ n25119 ^ n6910 ;
  assign n27742 = n20763 ^ n15575 ^ n9765 ;
  assign n27739 = n593 & n11202 ;
  assign n27740 = n27739 ^ n15303 ^ n7208 ;
  assign n27741 = n1598 | n27740 ;
  assign n27743 = n27742 ^ n27741 ^ 1'b0 ;
  assign n27744 = n23053 ^ n18032 ^ 1'b0 ;
  assign n27746 = ( n1252 & n4498 ) | ( n1252 & n23680 ) | ( n4498 & n23680 ) ;
  assign n27745 = n15112 | n24126 ;
  assign n27747 = n27746 ^ n27745 ^ 1'b0 ;
  assign n27748 = n11144 & ~n27747 ;
  assign n27749 = n27748 ^ n7643 ^ 1'b0 ;
  assign n27752 = n20485 & ~n26052 ;
  assign n27753 = n9239 & n27752 ;
  assign n27750 = n16432 ^ n11300 ^ 1'b0 ;
  assign n27751 = n6968 & ~n27750 ;
  assign n27754 = n27753 ^ n27751 ^ 1'b0 ;
  assign n27755 = n1144 | n2347 ;
  assign n27756 = n27755 ^ n13547 ^ n5707 ;
  assign n27757 = ( n5933 & n8064 ) | ( n5933 & n27756 ) | ( n8064 & n27756 ) ;
  assign n27758 = n5407 ^ n4000 ^ n1423 ;
  assign n27759 = n14195 ^ n13073 ^ n2494 ;
  assign n27760 = ( n7176 & n27758 ) | ( n7176 & ~n27759 ) | ( n27758 & ~n27759 ) ;
  assign n27761 = n10581 ^ n5304 ^ n4506 ;
  assign n27762 = n27761 ^ n8527 ^ 1'b0 ;
  assign n27763 = ( n9243 & n22374 ) | ( n9243 & ~n27762 ) | ( n22374 & ~n27762 ) ;
  assign n27764 = n11137 ^ n9152 ^ n5961 ;
  assign n27765 = ~n18573 & n27764 ;
  assign n27766 = n27765 ^ n25503 ^ n833 ;
  assign n27767 = n19989 ^ n13335 ^ 1'b0 ;
  assign n27768 = n13279 ^ n11354 ^ n6400 ;
  assign n27769 = ( n13689 & ~n27767 ) | ( n13689 & n27768 ) | ( ~n27767 & n27768 ) ;
  assign n27770 = n27769 ^ n4038 ^ 1'b0 ;
  assign n27771 = n4472 & ~n27770 ;
  assign n27772 = n2791 & n27771 ;
  assign n27773 = n17641 & n27772 ;
  assign n27774 = n15229 ^ n6786 ^ 1'b0 ;
  assign n27779 = n20512 ^ n15537 ^ n15208 ;
  assign n27775 = n8506 & n9489 ;
  assign n27776 = n22726 ^ n3213 ^ 1'b0 ;
  assign n27777 = n9223 | n27776 ;
  assign n27778 = ( ~n7346 & n27775 ) | ( ~n7346 & n27777 ) | ( n27775 & n27777 ) ;
  assign n27780 = n27779 ^ n27778 ^ n4145 ;
  assign n27781 = n27780 ^ n5013 ^ 1'b0 ;
  assign n27782 = ~n27774 & n27781 ;
  assign n27783 = ( n5182 & n12966 ) | ( n5182 & ~n17262 ) | ( n12966 & ~n17262 ) ;
  assign n27784 = ( n11917 & n14678 ) | ( n11917 & ~n27783 ) | ( n14678 & ~n27783 ) ;
  assign n27785 = ( n1651 & n5562 ) | ( n1651 & ~n22899 ) | ( n5562 & ~n22899 ) ;
  assign n27786 = n27785 ^ n15936 ^ n2613 ;
  assign n27787 = n14872 ^ n5177 ^ 1'b0 ;
  assign n27788 = ~n21628 & n27787 ;
  assign n27789 = n19509 ^ n10663 ^ 1'b0 ;
  assign n27790 = n24871 ^ n4562 ^ n1132 ;
  assign n27791 = ( ~x226 & n3303 ) | ( ~x226 & n9097 ) | ( n3303 & n9097 ) ;
  assign n27792 = n27790 & ~n27791 ;
  assign n27793 = n27792 ^ n4623 ^ 1'b0 ;
  assign n27794 = n27789 | n27793 ;
  assign n27795 = n27794 ^ n26169 ^ 1'b0 ;
  assign n27796 = ~n27788 & n27795 ;
  assign n27797 = ( n1153 & ~n7968 ) | ( n1153 & n13434 ) | ( ~n7968 & n13434 ) ;
  assign n27798 = ( ~n13605 & n19309 ) | ( ~n13605 & n20112 ) | ( n19309 & n20112 ) ;
  assign n27799 = n5649 & ~n27798 ;
  assign n27800 = n27799 ^ n4767 ^ 1'b0 ;
  assign n27801 = n402 | n27800 ;
  assign n27802 = n7974 | n27801 ;
  assign n27803 = n27797 | n27802 ;
  assign n27804 = n15622 & ~n17810 ;
  assign n27805 = n7784 & ~n24053 ;
  assign n27806 = ~n3918 & n27805 ;
  assign n27807 = n19386 ^ n2895 ^ 1'b0 ;
  assign n27808 = ( ~n16453 & n21199 ) | ( ~n16453 & n27807 ) | ( n21199 & n27807 ) ;
  assign n27809 = n16134 ^ n14934 ^ 1'b0 ;
  assign n27810 = ~n8790 & n27809 ;
  assign n27811 = n27810 ^ n13058 ^ n7340 ;
  assign n27814 = ( n5877 & n13625 ) | ( n5877 & ~n25945 ) | ( n13625 & ~n25945 ) ;
  assign n27812 = n15560 ^ n14720 ^ 1'b0 ;
  assign n27813 = n27812 ^ n19044 ^ 1'b0 ;
  assign n27815 = n27814 ^ n27813 ^ n5901 ;
  assign n27816 = n19144 ^ n14599 ^ x33 ;
  assign n27817 = n27816 ^ n26488 ^ n9612 ;
  assign n27818 = ( n3724 & n8882 ) | ( n3724 & ~n11899 ) | ( n8882 & ~n11899 ) ;
  assign n27819 = n10507 & ~n27818 ;
  assign n27820 = ~n12837 & n27819 ;
  assign n27821 = n13339 ^ n7909 ^ 1'b0 ;
  assign n27822 = n16290 ^ n4120 ^ n2957 ;
  assign n27823 = n27822 ^ n13291 ^ 1'b0 ;
  assign n27825 = n4260 ^ n2273 ^ 1'b0 ;
  assign n27826 = n27825 ^ n21061 ^ n2258 ;
  assign n27824 = n11683 & ~n27635 ;
  assign n27827 = n27826 ^ n27824 ^ 1'b0 ;
  assign n27828 = ~n8921 & n21445 ;
  assign n27829 = ~n13972 & n27828 ;
  assign n27830 = ( n672 & ~n15078 ) | ( n672 & n21323 ) | ( ~n15078 & n21323 ) ;
  assign n27831 = ( ~n3045 & n23300 ) | ( ~n3045 & n27830 ) | ( n23300 & n27830 ) ;
  assign n27832 = n3330 | n6834 ;
  assign n27833 = n18255 ^ n5307 ^ 1'b0 ;
  assign n27834 = n7914 & ~n27833 ;
  assign n27835 = ( n11180 & n19758 ) | ( n11180 & n27834 ) | ( n19758 & n27834 ) ;
  assign n27836 = n27835 ^ n16970 ^ 1'b0 ;
  assign n27837 = ( n24573 & n27832 ) | ( n24573 & n27836 ) | ( n27832 & n27836 ) ;
  assign n27838 = n23965 ^ n6050 ^ 1'b0 ;
  assign n27839 = n7183 ^ n3588 ^ n713 ;
  assign n27840 = n27839 ^ n13468 ^ n1530 ;
  assign n27841 = ( ~n14870 & n23275 ) | ( ~n14870 & n27840 ) | ( n23275 & n27840 ) ;
  assign n27842 = n1109 | n27841 ;
  assign n27843 = n8770 | n27842 ;
  assign n27844 = ( ~n4928 & n5285 ) | ( ~n4928 & n7417 ) | ( n5285 & n7417 ) ;
  assign n27845 = n18397 ^ n729 ^ 1'b0 ;
  assign n27846 = n27844 & ~n27845 ;
  assign n27847 = n27846 ^ n6069 ^ 1'b0 ;
  assign n27848 = n20094 ^ n11345 ^ n10155 ;
  assign n27849 = n27848 ^ n21726 ^ n12902 ;
  assign n27850 = n27849 ^ n15384 ^ n15114 ;
  assign n27851 = ( n2096 & ~n10031 ) | ( n2096 & n13196 ) | ( ~n10031 & n13196 ) ;
  assign n27852 = n19378 | n27851 ;
  assign n27853 = n14830 | n27852 ;
  assign n27854 = ( n11920 & ~n22062 ) | ( n11920 & n23364 ) | ( ~n22062 & n23364 ) ;
  assign n27855 = n7826 ^ n3595 ^ 1'b0 ;
  assign n27859 = n8313 ^ n2905 ^ n1633 ;
  assign n27856 = n721 | n6316 ;
  assign n27857 = n27856 ^ n1297 ^ 1'b0 ;
  assign n27858 = ( ~n15335 & n21079 ) | ( ~n15335 & n27857 ) | ( n21079 & n27857 ) ;
  assign n27860 = n27859 ^ n27858 ^ n344 ;
  assign n27861 = n7775 | n27860 ;
  assign n27862 = ( n14619 & n27855 ) | ( n14619 & n27861 ) | ( n27855 & n27861 ) ;
  assign n27863 = n26121 ^ n22440 ^ n7867 ;
  assign n27864 = n11651 ^ n3298 ^ x119 ;
  assign n27865 = n9478 ^ n4850 ^ 1'b0 ;
  assign n27866 = n8653 & n27865 ;
  assign n27867 = n27864 & ~n27866 ;
  assign n27868 = ( n2747 & n13059 ) | ( n2747 & ~n27867 ) | ( n13059 & ~n27867 ) ;
  assign n27869 = n9312 | n19259 ;
  assign n27870 = n7525 & ~n27869 ;
  assign n27871 = n27870 ^ n10292 ^ n2455 ;
  assign n27872 = n19288 ^ n5294 ^ 1'b0 ;
  assign n27873 = ( n6124 & ~n8760 ) | ( n6124 & n10362 ) | ( ~n8760 & n10362 ) ;
  assign n27874 = ~n8750 & n27873 ;
  assign n27875 = n27872 & n27874 ;
  assign n27877 = n4554 & ~n12497 ;
  assign n27878 = n27877 ^ n20589 ^ n12263 ;
  assign n27876 = n6048 & ~n27245 ;
  assign n27879 = n27878 ^ n27876 ^ n1755 ;
  assign n27880 = ~n14941 & n27879 ;
  assign n27881 = ( n2199 & ~n17557 ) | ( n2199 & n18571 ) | ( ~n17557 & n18571 ) ;
  assign n27882 = n25888 ^ n6858 ^ 1'b0 ;
  assign n27883 = n27881 | n27882 ;
  assign n27888 = n14357 ^ n4225 ^ 1'b0 ;
  assign n27889 = n6763 & n27888 ;
  assign n27887 = n22244 ^ n10466 ^ n5471 ;
  assign n27890 = n27889 ^ n27887 ^ n27425 ;
  assign n27884 = n7615 | n7653 ;
  assign n27885 = n27884 ^ n15949 ^ 1'b0 ;
  assign n27886 = n27885 ^ n17332 ^ n5848 ;
  assign n27891 = n27890 ^ n27886 ^ n7694 ;
  assign n27892 = n9573 & ~n12456 ;
  assign n27893 = ~n393 & n468 ;
  assign n27894 = n15164 & n27893 ;
  assign n27895 = n8448 | n27894 ;
  assign n27896 = n17127 ^ n2762 ^ 1'b0 ;
  assign n27897 = ~n16702 & n27896 ;
  assign n27898 = n14146 ^ n5049 ^ 1'b0 ;
  assign n27899 = n4911 | n27898 ;
  assign n27900 = n6375 ^ n549 ^ 1'b0 ;
  assign n27901 = n3925 | n27900 ;
  assign n27902 = ( n4792 & ~n23966 ) | ( n4792 & n27901 ) | ( ~n23966 & n27901 ) ;
  assign n27903 = n19503 ^ n18840 ^ n5326 ;
  assign n27904 = ( n9064 & n19444 ) | ( n9064 & n23783 ) | ( n19444 & n23783 ) ;
  assign n27905 = n5796 ^ n5409 ^ 1'b0 ;
  assign n27906 = n7167 & ~n27905 ;
  assign n27907 = n27906 ^ n25594 ^ n24187 ;
  assign n27908 = n10419 ^ n7830 ^ n898 ;
  assign n27909 = ( ~n3228 & n4860 ) | ( ~n3228 & n13800 ) | ( n4860 & n13800 ) ;
  assign n27910 = ( n8521 & n27908 ) | ( n8521 & n27909 ) | ( n27908 & n27909 ) ;
  assign n27911 = ( ~n4873 & n12834 ) | ( ~n4873 & n17215 ) | ( n12834 & n17215 ) ;
  assign n27912 = n27911 ^ n23687 ^ n15298 ;
  assign n27918 = n16606 & ~n19573 ;
  assign n27917 = ~n12893 & n22389 ;
  assign n27913 = n4159 & ~n9927 ;
  assign n27914 = n26623 ^ n25697 ^ n23984 ;
  assign n27915 = n12695 & n27914 ;
  assign n27916 = ~n27913 & n27915 ;
  assign n27919 = n27918 ^ n27917 ^ n27916 ;
  assign n27921 = n3395 & n4444 ;
  assign n27920 = ~n993 & n7262 ;
  assign n27922 = n27921 ^ n27920 ^ 1'b0 ;
  assign n27925 = n14992 ^ n7633 ^ n6764 ;
  assign n27926 = ( n6671 & n19179 ) | ( n6671 & n27925 ) | ( n19179 & n27925 ) ;
  assign n27923 = ~n7261 & n9802 ;
  assign n27924 = n27923 ^ n13711 ^ 1'b0 ;
  assign n27927 = n27926 ^ n27924 ^ 1'b0 ;
  assign n27928 = n5344 & n27927 ;
  assign n27929 = n17626 & n27928 ;
  assign n27930 = ~n27922 & n27929 ;
  assign n27936 = ( n7110 & n17840 ) | ( n7110 & n18351 ) | ( n17840 & n18351 ) ;
  assign n27935 = n3482 & n16694 ;
  assign n27937 = n27936 ^ n27935 ^ 1'b0 ;
  assign n27938 = ( n801 & n22164 ) | ( n801 & ~n27937 ) | ( n22164 & ~n27937 ) ;
  assign n27931 = ( n762 & ~n10092 ) | ( n762 & n25263 ) | ( ~n10092 & n25263 ) ;
  assign n27932 = n16901 ^ n6578 ^ 1'b0 ;
  assign n27933 = n12732 & ~n27932 ;
  assign n27934 = ~n27931 & n27933 ;
  assign n27939 = n27938 ^ n27934 ^ 1'b0 ;
  assign n27940 = ( n2526 & n14480 ) | ( n2526 & n18920 ) | ( n14480 & n18920 ) ;
  assign n27941 = n27940 ^ n16189 ^ n501 ;
  assign n27942 = n5536 ^ n3950 ^ 1'b0 ;
  assign n27943 = n27941 | n27942 ;
  assign n27947 = ( n446 & n8769 ) | ( n446 & n17887 ) | ( n8769 & n17887 ) ;
  assign n27944 = ~n13728 & n23215 ;
  assign n27945 = ~n12133 & n27944 ;
  assign n27946 = n10423 & ~n27945 ;
  assign n27948 = n27947 ^ n27946 ^ 1'b0 ;
  assign n27949 = ( ~n5941 & n10763 ) | ( ~n5941 & n15302 ) | ( n10763 & n15302 ) ;
  assign n27950 = ( n16420 & n22615 ) | ( n16420 & n22925 ) | ( n22615 & n22925 ) ;
  assign n27951 = n11611 ^ n2043 ^ 1'b0 ;
  assign n27952 = ( n27949 & ~n27950 ) | ( n27949 & n27951 ) | ( ~n27950 & n27951 ) ;
  assign n27953 = n6667 ^ n903 ^ 1'b0 ;
  assign n27954 = n13481 ^ n8677 ^ 1'b0 ;
  assign n27955 = ( n8357 & n27953 ) | ( n8357 & ~n27954 ) | ( n27953 & ~n27954 ) ;
  assign n27956 = n27955 ^ n19937 ^ x230 ;
  assign n27957 = ( n6841 & n15778 ) | ( n6841 & n27956 ) | ( n15778 & n27956 ) ;
  assign n27958 = ~n5707 & n15393 ;
  assign n27959 = n27958 ^ n27121 ^ 1'b0 ;
  assign n27960 = ( n8878 & ~n21583 ) | ( n8878 & n27959 ) | ( ~n21583 & n27959 ) ;
  assign n27961 = ( ~n20508 & n23724 ) | ( ~n20508 & n27960 ) | ( n23724 & n27960 ) ;
  assign n27962 = n19233 ^ n4174 ^ 1'b0 ;
  assign n27963 = n7032 & ~n9042 ;
  assign n27964 = n27963 ^ n4051 ^ 1'b0 ;
  assign n27965 = ( n8884 & ~n27962 ) | ( n8884 & n27964 ) | ( ~n27962 & n27964 ) ;
  assign n27966 = n1245 & n27965 ;
  assign n27967 = n27966 ^ n9046 ^ 1'b0 ;
  assign n27968 = ~n12150 & n18542 ;
  assign n27969 = n27968 ^ n10566 ^ n8148 ;
  assign n27970 = n8001 & n15506 ;
  assign n27971 = n27970 ^ n6849 ^ 1'b0 ;
  assign n27972 = n27971 ^ n19047 ^ n401 ;
  assign n27973 = n15813 ^ n13875 ^ n5231 ;
  assign n27974 = n19949 & n27973 ;
  assign n27975 = ( n3801 & ~n14549 ) | ( n3801 & n27974 ) | ( ~n14549 & n27974 ) ;
  assign n27976 = n15184 ^ n9339 ^ 1'b0 ;
  assign n27977 = ( n5682 & n18729 ) | ( n5682 & n27976 ) | ( n18729 & n27976 ) ;
  assign n27978 = n25960 ^ n18308 ^ n7028 ;
  assign n27979 = n27978 ^ n17319 ^ 1'b0 ;
  assign n27980 = ~n23264 & n27979 ;
  assign n27981 = n27980 ^ n26522 ^ n13899 ;
  assign n27982 = n20912 & n27981 ;
  assign n27984 = n5498 ^ n4768 ^ n1822 ;
  assign n27983 = n1755 & ~n23568 ;
  assign n27985 = n27984 ^ n27983 ^ 1'b0 ;
  assign n27986 = n966 | n27985 ;
  assign n27988 = n9863 ^ n5248 ^ 1'b0 ;
  assign n27989 = n1340 & ~n27988 ;
  assign n27990 = n27989 ^ n3415 ^ 1'b0 ;
  assign n27987 = n6493 ^ n1995 ^ 1'b0 ;
  assign n27991 = n27990 ^ n27987 ^ n22107 ;
  assign n27992 = n5614 & n6463 ;
  assign n27993 = ~n25117 & n27992 ;
  assign n27994 = ( ~n17576 & n19163 ) | ( ~n17576 & n27993 ) | ( n19163 & n27993 ) ;
  assign n27998 = ( x231 & n10979 ) | ( x231 & n19260 ) | ( n10979 & n19260 ) ;
  assign n27995 = n5154 & ~n17577 ;
  assign n27996 = ~n20398 & n27995 ;
  assign n27997 = ( n6985 & n19891 ) | ( n6985 & n27996 ) | ( n19891 & n27996 ) ;
  assign n27999 = n27998 ^ n27997 ^ 1'b0 ;
  assign n28000 = n16500 ^ n14584 ^ 1'b0 ;
  assign n28001 = n19599 ^ n12094 ^ n5629 ;
  assign n28002 = ( ~n10498 & n13906 ) | ( ~n10498 & n28001 ) | ( n13906 & n28001 ) ;
  assign n28003 = n25312 ^ n8965 ^ 1'b0 ;
  assign n28004 = ( n5688 & n19767 ) | ( n5688 & ~n28003 ) | ( n19767 & ~n28003 ) ;
  assign n28005 = n21966 ^ n6557 ^ n4229 ;
  assign n28006 = n24541 ^ n10727 ^ 1'b0 ;
  assign n28007 = ~n28005 & n28006 ;
  assign n28009 = n27669 ^ n10091 ^ n534 ;
  assign n28008 = n23619 ^ n8938 ^ n5755 ;
  assign n28010 = n28009 ^ n28008 ^ 1'b0 ;
  assign n28011 = n1604 & ~n23501 ;
  assign n28012 = ~n21365 & n28011 ;
  assign n28013 = n13255 ^ n1670 ^ 1'b0 ;
  assign n28014 = n3171 & ~n28013 ;
  assign n28015 = ~n5923 & n28014 ;
  assign n28016 = ~n1376 & n28015 ;
  assign n28017 = ( n22034 & n28012 ) | ( n22034 & ~n28016 ) | ( n28012 & ~n28016 ) ;
  assign n28018 = n12208 | n16377 ;
  assign n28019 = n28017 & ~n28018 ;
  assign n28020 = n10649 ^ n5890 ^ n1805 ;
  assign n28021 = n5506 ^ n1674 ^ 1'b0 ;
  assign n28022 = n28020 & ~n28021 ;
  assign n28023 = ~n27543 & n28022 ;
  assign n28024 = ( n1873 & n10885 ) | ( n1873 & n11471 ) | ( n10885 & n11471 ) ;
  assign n28025 = n17593 ^ n3833 ^ n1017 ;
  assign n28026 = ( ~n18388 & n21373 ) | ( ~n18388 & n28025 ) | ( n21373 & n28025 ) ;
  assign n28027 = ( n1926 & n28024 ) | ( n1926 & n28026 ) | ( n28024 & n28026 ) ;
  assign n28030 = ~n11035 & n25876 ;
  assign n28031 = n15868 & n28030 ;
  assign n28029 = ( n3759 & n5929 ) | ( n3759 & n24241 ) | ( n5929 & n24241 ) ;
  assign n28028 = ~n1739 & n4991 ;
  assign n28032 = n28031 ^ n28029 ^ n28028 ;
  assign n28033 = ( ~n19743 & n24366 ) | ( ~n19743 & n28032 ) | ( n24366 & n28032 ) ;
  assign n28034 = ~n23510 & n27024 ;
  assign n28035 = n9750 ^ n3429 ^ n696 ;
  assign n28036 = n12166 ^ n8905 ^ n8430 ;
  assign n28037 = n22261 | n28036 ;
  assign n28038 = ~n11093 & n28037 ;
  assign n28039 = ~n20858 & n28038 ;
  assign n28040 = ( n28034 & n28035 ) | ( n28034 & n28039 ) | ( n28035 & n28039 ) ;
  assign n28041 = n9838 & ~n27072 ;
  assign n28042 = ~n1821 & n28041 ;
  assign n28043 = n16973 | n28042 ;
  assign n28044 = n28040 | n28043 ;
  assign n28045 = n28044 ^ n24746 ^ n1599 ;
  assign n28046 = n16281 ^ n6604 ^ 1'b0 ;
  assign n28047 = n28046 ^ n13392 ^ n4172 ;
  assign n28049 = n12622 ^ n1491 ^ n500 ;
  assign n28050 = ~n1005 & n28049 ;
  assign n28048 = n15268 ^ n8418 ^ n431 ;
  assign n28051 = n28050 ^ n28048 ^ n5305 ;
  assign n28053 = n5324 ^ n2962 ^ n1850 ;
  assign n28052 = ( ~n20047 & n20405 ) | ( ~n20047 & n20708 ) | ( n20405 & n20708 ) ;
  assign n28054 = n28053 ^ n28052 ^ n3117 ;
  assign n28055 = n28054 ^ n23662 ^ n13183 ;
  assign n28056 = n10401 | n28055 ;
  assign n28057 = n28051 | n28056 ;
  assign n28058 = n17927 & ~n22527 ;
  assign n28059 = n28058 ^ x66 ^ 1'b0 ;
  assign n28060 = ( n7421 & n14545 ) | ( n7421 & n27341 ) | ( n14545 & n27341 ) ;
  assign n28063 = n18835 ^ n5084 ^ n4078 ;
  assign n28061 = n19508 ^ n7813 ^ n7668 ;
  assign n28062 = n4888 & n28061 ;
  assign n28064 = n28063 ^ n28062 ^ 1'b0 ;
  assign n28065 = n22401 ^ n4855 ^ n1774 ;
  assign n28066 = n28065 ^ n14649 ^ n9673 ;
  assign n28067 = n28066 ^ n22398 ^ n2240 ;
  assign n28068 = n28067 ^ n11106 ^ 1'b0 ;
  assign n28069 = n14495 & n21712 ;
  assign n28070 = ~n25484 & n28069 ;
  assign n28071 = n11168 | n25378 ;
  assign n28072 = n21206 | n28071 ;
  assign n28074 = n4980 ^ n4603 ^ 1'b0 ;
  assign n28075 = n818 & n28074 ;
  assign n28076 = ( n3535 & n10092 ) | ( n3535 & ~n28075 ) | ( n10092 & ~n28075 ) ;
  assign n28077 = n28076 ^ n6461 ^ n6214 ;
  assign n28078 = n2085 | n4060 ;
  assign n28079 = n26708 ^ n22725 ^ n15757 ;
  assign n28080 = ( n13121 & n28078 ) | ( n13121 & ~n28079 ) | ( n28078 & ~n28079 ) ;
  assign n28081 = n15887 & n28080 ;
  assign n28082 = ( n21552 & ~n28077 ) | ( n21552 & n28081 ) | ( ~n28077 & n28081 ) ;
  assign n28083 = ( n2232 & n20086 ) | ( n2232 & ~n28082 ) | ( n20086 & ~n28082 ) ;
  assign n28073 = ( n2673 & ~n3143 ) | ( n2673 & n5876 ) | ( ~n3143 & n5876 ) ;
  assign n28084 = n28083 ^ n28073 ^ 1'b0 ;
  assign n28085 = ( n7012 & ~n16094 ) | ( n7012 & n16753 ) | ( ~n16094 & n16753 ) ;
  assign n28086 = n18738 ^ n8973 ^ 1'b0 ;
  assign n28087 = ( ~n1191 & n24492 ) | ( ~n1191 & n24523 ) | ( n24492 & n24523 ) ;
  assign n28088 = n28087 ^ n25056 ^ n19573 ;
  assign n28089 = n28088 ^ n20796 ^ n6176 ;
  assign n28090 = n15356 ^ n6855 ^ 1'b0 ;
  assign n28091 = n22646 & ~n28090 ;
  assign n28092 = n28091 ^ n9305 ^ n3747 ;
  assign n28093 = n20515 ^ n15222 ^ n3387 ;
  assign n28094 = n28093 ^ n25130 ^ n11406 ;
  assign n28095 = n20534 & ~n28094 ;
  assign n28096 = n26192 & n28095 ;
  assign n28097 = ~n870 & n7368 ;
  assign n28098 = ( ~n13524 & n20979 ) | ( ~n13524 & n28097 ) | ( n20979 & n28097 ) ;
  assign n28099 = ( n756 & n18167 ) | ( n756 & ~n23121 ) | ( n18167 & ~n23121 ) ;
  assign n28100 = ( n26915 & n28098 ) | ( n26915 & ~n28099 ) | ( n28098 & ~n28099 ) ;
  assign n28101 = n19908 ^ n17215 ^ n11897 ;
  assign n28102 = ( n2355 & n13972 ) | ( n2355 & n22046 ) | ( n13972 & n22046 ) ;
  assign n28103 = n28102 ^ n25853 ^ n5830 ;
  assign n28104 = n547 & n6068 ;
  assign n28105 = n28104 ^ n25671 ^ 1'b0 ;
  assign n28106 = n23830 | n28105 ;
  assign n28107 = ( n6946 & n22417 ) | ( n6946 & n28106 ) | ( n22417 & n28106 ) ;
  assign n28108 = n3985 & n20560 ;
  assign n28109 = n28108 ^ n8971 ^ 1'b0 ;
  assign n28110 = n28109 ^ n10804 ^ n10084 ;
  assign n28111 = n6640 | n28082 ;
  assign n28112 = ( n2765 & n13687 ) | ( n2765 & ~n16756 ) | ( n13687 & ~n16756 ) ;
  assign n28113 = ( n3260 & n11580 ) | ( n3260 & ~n28112 ) | ( n11580 & ~n28112 ) ;
  assign n28114 = n28113 ^ n19844 ^ n1087 ;
  assign n28115 = n9366 & n11280 ;
  assign n28116 = n28115 ^ n25337 ^ 1'b0 ;
  assign n28117 = n27913 ^ n16601 ^ n4586 ;
  assign n28118 = n18848 ^ n3078 ^ 1'b0 ;
  assign n28121 = ( n4653 & ~n6355 ) | ( n4653 & n9248 ) | ( ~n6355 & n9248 ) ;
  assign n28119 = n12600 & n18847 ;
  assign n28120 = n28119 ^ n15931 ^ 1'b0 ;
  assign n28122 = n28121 ^ n28120 ^ 1'b0 ;
  assign n28123 = n17595 ^ n14771 ^ n4080 ;
  assign n28124 = n8313 & ~n27616 ;
  assign n28125 = n28124 ^ n14305 ^ 1'b0 ;
  assign n28128 = n27658 ^ n20198 ^ 1'b0 ;
  assign n28129 = ~n4555 & n28128 ;
  assign n28126 = n14795 ^ n9941 ^ 1'b0 ;
  assign n28127 = n4326 & ~n28126 ;
  assign n28130 = n28129 ^ n28127 ^ n20960 ;
  assign n28133 = ( n2033 & n2948 ) | ( n2033 & n12299 ) | ( n2948 & n12299 ) ;
  assign n28132 = ( n4540 & ~n8428 ) | ( n4540 & n17578 ) | ( ~n8428 & n17578 ) ;
  assign n28131 = n18337 ^ n9170 ^ 1'b0 ;
  assign n28134 = n28133 ^ n28132 ^ n28131 ;
  assign n28136 = n23010 ^ n4122 ^ 1'b0 ;
  assign n28137 = ( ~n7156 & n14996 ) | ( ~n7156 & n17404 ) | ( n14996 & n17404 ) ;
  assign n28138 = n28137 ^ n3539 ^ 1'b0 ;
  assign n28139 = n4459 | n28138 ;
  assign n28140 = ( n835 & n7202 ) | ( n835 & ~n28139 ) | ( n7202 & ~n28139 ) ;
  assign n28141 = n28136 & ~n28140 ;
  assign n28135 = n2345 & n20711 ;
  assign n28142 = n28141 ^ n28135 ^ 1'b0 ;
  assign n28143 = x70 & ~n3046 ;
  assign n28144 = n18820 & n28143 ;
  assign n28145 = n2569 | n26266 ;
  assign n28146 = n28145 ^ n7549 ^ 1'b0 ;
  assign n28147 = n1221 & ~n14628 ;
  assign n28156 = n4489 & n5622 ;
  assign n28157 = n28156 ^ n1399 ^ 1'b0 ;
  assign n28150 = n6749 | n10797 ;
  assign n28151 = n28150 ^ n20800 ^ 1'b0 ;
  assign n28152 = ~n5172 & n11450 ;
  assign n28153 = n28151 & n28152 ;
  assign n28154 = ~n19649 & n28153 ;
  assign n28155 = n28154 ^ n17754 ^ n1381 ;
  assign n28148 = ( n2610 & n20239 ) | ( n2610 & n25029 ) | ( n20239 & n25029 ) ;
  assign n28149 = n28148 ^ n26738 ^ n23657 ;
  assign n28158 = n28157 ^ n28155 ^ n28149 ;
  assign n28159 = n17845 ^ n9135 ^ n8377 ;
  assign n28163 = n9344 & ~n25026 ;
  assign n28164 = n28163 ^ n22765 ^ 1'b0 ;
  assign n28165 = n22512 ^ n2559 ^ 1'b0 ;
  assign n28166 = n28164 & ~n28165 ;
  assign n28160 = n21951 ^ n20766 ^ n2018 ;
  assign n28161 = n28160 ^ n18072 ^ n8881 ;
  assign n28162 = n28161 ^ n13758 ^ n5740 ;
  assign n28167 = n28166 ^ n28162 ^ n16597 ;
  assign n28169 = ~n2786 & n6601 ;
  assign n28170 = n28169 ^ n5705 ^ n5311 ;
  assign n28168 = n17494 ^ n12542 ^ 1'b0 ;
  assign n28171 = n28170 ^ n28168 ^ n20409 ;
  assign n28172 = n4862 ^ n3952 ^ 1'b0 ;
  assign n28173 = n1720 | n18485 ;
  assign n28174 = n28173 ^ n11974 ^ 1'b0 ;
  assign n28175 = ~n7954 & n16519 ;
  assign n28176 = n28175 ^ n20895 ^ 1'b0 ;
  assign n28177 = ( n1097 & ~n4047 ) | ( n1097 & n10835 ) | ( ~n4047 & n10835 ) ;
  assign n28178 = n28176 | n28177 ;
  assign n28179 = ( x134 & ~n11886 ) | ( x134 & n15041 ) | ( ~n11886 & n15041 ) ;
  assign n28180 = n8656 ^ n7150 ^ n598 ;
  assign n28181 = ( n11470 & n13073 ) | ( n11470 & n28180 ) | ( n13073 & n28180 ) ;
  assign n28182 = ( n7891 & ~n21125 ) | ( n7891 & n28181 ) | ( ~n21125 & n28181 ) ;
  assign n28183 = ( ~n5370 & n11363 ) | ( ~n5370 & n15214 ) | ( n11363 & n15214 ) ;
  assign n28184 = ~n903 & n19625 ;
  assign n28185 = n14206 & n28184 ;
  assign n28186 = n7247 ^ n5739 ^ n2747 ;
  assign n28187 = n28186 ^ n13016 ^ 1'b0 ;
  assign n28188 = n28187 ^ n24046 ^ n9866 ;
  assign n28189 = n17323 | n19395 ;
  assign n28190 = n28189 ^ x60 ^ 1'b0 ;
  assign n28191 = n2302 | n14240 ;
  assign n28192 = n23473 ^ n10700 ^ 1'b0 ;
  assign n28193 = n28191 & ~n28192 ;
  assign n28194 = ( ~n747 & n13003 ) | ( ~n747 & n28193 ) | ( n13003 & n28193 ) ;
  assign n28195 = ~n16373 & n27319 ;
  assign n28196 = ~n28194 & n28195 ;
  assign n28197 = n5743 ^ n1451 ^ 1'b0 ;
  assign n28198 = n3083 | n28197 ;
  assign n28199 = n4245 | n4406 ;
  assign n28200 = n28198 | n28199 ;
  assign n28201 = n2876 & ~n28200 ;
  assign n28204 = n325 & n10583 ;
  assign n28205 = ( n7021 & n13967 ) | ( n7021 & ~n28204 ) | ( n13967 & ~n28204 ) ;
  assign n28206 = n28205 ^ n14623 ^ n9639 ;
  assign n28207 = n11730 & ~n20751 ;
  assign n28208 = ~n28206 & n28207 ;
  assign n28202 = n4281 ^ n1420 ^ 1'b0 ;
  assign n28203 = n15071 | n28202 ;
  assign n28209 = n28208 ^ n28203 ^ 1'b0 ;
  assign n28213 = n6956 | n28065 ;
  assign n28214 = n14057 & ~n28213 ;
  assign n28210 = ( ~n1988 & n3621 ) | ( ~n1988 & n17976 ) | ( n3621 & n17976 ) ;
  assign n28211 = ( n10603 & n13933 ) | ( n10603 & n28210 ) | ( n13933 & n28210 ) ;
  assign n28212 = ( n10370 & ~n16161 ) | ( n10370 & n28211 ) | ( ~n16161 & n28211 ) ;
  assign n28215 = n28214 ^ n28212 ^ n6873 ;
  assign n28216 = ( n7110 & n21848 ) | ( n7110 & ~n27024 ) | ( n21848 & ~n27024 ) ;
  assign n28217 = ( n19101 & n24456 ) | ( n19101 & ~n24879 ) | ( n24456 & ~n24879 ) ;
  assign n28218 = n20697 ^ n8555 ^ n5556 ;
  assign n28219 = n22336 & n28218 ;
  assign n28220 = ~n14343 & n28219 ;
  assign n28221 = n4100 & n19156 ;
  assign n28222 = ( n8755 & ~n10840 ) | ( n8755 & n28221 ) | ( ~n10840 & n28221 ) ;
  assign n28223 = n23068 ^ n436 ^ 1'b0 ;
  assign n28224 = n4086 & ~n14133 ;
  assign n28225 = n16019 ^ n1706 ^ 1'b0 ;
  assign n28226 = ( n6444 & n8616 ) | ( n6444 & ~n22862 ) | ( n8616 & ~n22862 ) ;
  assign n28227 = n28226 ^ n5275 ^ n1627 ;
  assign n28228 = ( n12343 & ~n28225 ) | ( n12343 & n28227 ) | ( ~n28225 & n28227 ) ;
  assign n28229 = n19326 ^ n18152 ^ x70 ;
  assign n28230 = n22979 ^ n20463 ^ 1'b0 ;
  assign n28231 = n6555 & ~n28230 ;
  assign n28232 = n28231 ^ n14698 ^ n10727 ;
  assign n28233 = ( ~n12247 & n25308 ) | ( ~n12247 & n28112 ) | ( n25308 & n28112 ) ;
  assign n28234 = ( n8086 & n17687 ) | ( n8086 & n22401 ) | ( n17687 & n22401 ) ;
  assign n28235 = ( n817 & n15174 ) | ( n817 & n28234 ) | ( n15174 & n28234 ) ;
  assign n28236 = n28235 ^ n14912 ^ 1'b0 ;
  assign n28237 = n26013 ^ n16321 ^ 1'b0 ;
  assign n28238 = ~n19920 & n28237 ;
  assign n28239 = n9054 ^ n3091 ^ n2797 ;
  assign n28240 = n28239 ^ n5475 ^ 1'b0 ;
  assign n28241 = n28238 & ~n28240 ;
  assign n28242 = n23914 ^ n20504 ^ n14426 ;
  assign n28245 = n11777 ^ n11180 ^ n9895 ;
  assign n28243 = n11526 ^ n1447 ^ 1'b0 ;
  assign n28244 = n12271 & ~n28243 ;
  assign n28246 = n28245 ^ n28244 ^ 1'b0 ;
  assign n28247 = n18253 ^ n17398 ^ 1'b0 ;
  assign n28248 = ( n10420 & n15358 ) | ( n10420 & n28247 ) | ( n15358 & n28247 ) ;
  assign n28249 = ( n8917 & n27692 ) | ( n8917 & n28248 ) | ( n27692 & n28248 ) ;
  assign n28250 = ( n28242 & ~n28246 ) | ( n28242 & n28249 ) | ( ~n28246 & n28249 ) ;
  assign n28251 = n18653 & n23088 ;
  assign n28252 = n15882 & n28251 ;
  assign n28253 = n22876 | n28252 ;
  assign n28254 = n28250 & ~n28253 ;
  assign n28255 = n13082 ^ n10089 ^ n1400 ;
  assign n28256 = n8784 ^ n6623 ^ 1'b0 ;
  assign n28257 = ~n28255 & n28256 ;
  assign n28258 = ( n2862 & n7432 ) | ( n2862 & ~n28257 ) | ( n7432 & ~n28257 ) ;
  assign n28259 = n20205 ^ n14545 ^ n6667 ;
  assign n28260 = n12340 ^ n6735 ^ 1'b0 ;
  assign n28261 = n2239 | n28260 ;
  assign n28262 = n28261 ^ n17835 ^ 1'b0 ;
  assign n28263 = n5660 & n28262 ;
  assign n28265 = n11348 ^ x123 ^ 1'b0 ;
  assign n28264 = n19821 ^ n5761 ^ n3006 ;
  assign n28266 = n28265 ^ n28264 ^ 1'b0 ;
  assign n28267 = n28263 & ~n28266 ;
  assign n28268 = ~n28259 & n28267 ;
  assign n28269 = n9146 & n28268 ;
  assign n28270 = n28269 ^ n8670 ^ n496 ;
  assign n28271 = ( ~n5058 & n14859 ) | ( ~n5058 & n26675 ) | ( n14859 & n26675 ) ;
  assign n28272 = n24020 ^ n14339 ^ 1'b0 ;
  assign n28273 = n12630 | n21866 ;
  assign n28274 = n22140 ^ n16312 ^ n11995 ;
  assign n28275 = ~n9296 & n28274 ;
  assign n28276 = n28275 ^ n21671 ^ 1'b0 ;
  assign n28281 = ( n2315 & ~n12012 ) | ( n2315 & n20584 ) | ( ~n12012 & n20584 ) ;
  assign n28279 = ( ~n3268 & n4619 ) | ( ~n3268 & n7919 ) | ( n4619 & n7919 ) ;
  assign n28280 = n28279 ^ n3383 ^ n2911 ;
  assign n28282 = n28281 ^ n28280 ^ x137 ;
  assign n28277 = ( n7352 & n10915 ) | ( n7352 & n14054 ) | ( n10915 & n14054 ) ;
  assign n28278 = n28277 ^ n5340 ^ 1'b0 ;
  assign n28283 = n28282 ^ n28278 ^ n17605 ;
  assign n28284 = n26285 ^ n12215 ^ n4362 ;
  assign n28285 = n28284 ^ n14375 ^ 1'b0 ;
  assign n28286 = n28285 ^ n27717 ^ n6346 ;
  assign n28287 = n25883 ^ n16573 ^ n5074 ;
  assign n28288 = n28287 ^ n7896 ^ 1'b0 ;
  assign n28293 = n8378 ^ n5477 ^ n3916 ;
  assign n28294 = n28293 ^ n24960 ^ n13675 ;
  assign n28295 = n6317 & ~n28294 ;
  assign n28290 = n15853 ^ n10762 ^ 1'b0 ;
  assign n28291 = n28290 ^ n21617 ^ n2810 ;
  assign n28292 = n28291 ^ n20666 ^ n13628 ;
  assign n28289 = n13558 ^ n11042 ^ x83 ;
  assign n28296 = n28295 ^ n28292 ^ n28289 ;
  assign n28297 = n14467 ^ n1981 ^ 1'b0 ;
  assign n28298 = n9235 ^ n3423 ^ 1'b0 ;
  assign n28299 = ~n26984 & n28298 ;
  assign n28300 = n28299 ^ n21032 ^ n2961 ;
  assign n28301 = ( n21683 & n28297 ) | ( n21683 & n28300 ) | ( n28297 & n28300 ) ;
  assign n28302 = n9687 ^ n2842 ^ 1'b0 ;
  assign n28303 = n28302 ^ n10483 ^ n4619 ;
  assign n28304 = ( n5951 & n19922 ) | ( n5951 & ~n23493 ) | ( n19922 & ~n23493 ) ;
  assign n28305 = n28303 & n28304 ;
  assign n28306 = n10367 & n28305 ;
  assign n28307 = ~n7246 & n19029 ;
  assign n28308 = n28307 ^ n4005 ^ 1'b0 ;
  assign n28309 = n12027 & n28308 ;
  assign n28310 = n28309 ^ n28206 ^ 1'b0 ;
  assign n28311 = n28310 ^ n18044 ^ 1'b0 ;
  assign n28312 = n28311 ^ n19067 ^ n9796 ;
  assign n28313 = ~n12316 & n12840 ;
  assign n28317 = n23119 ^ n19338 ^ n7605 ;
  assign n28318 = n8638 ^ n550 ^ 1'b0 ;
  assign n28319 = n28317 & ~n28318 ;
  assign n28320 = n28319 ^ n8993 ^ n1315 ;
  assign n28316 = ( n6658 & n9468 ) | ( n6658 & n19385 ) | ( n9468 & n19385 ) ;
  assign n28314 = n4790 & ~n6500 ;
  assign n28315 = ( n1515 & ~n9343 ) | ( n1515 & n28314 ) | ( ~n9343 & n28314 ) ;
  assign n28321 = n28320 ^ n28316 ^ n28315 ;
  assign n28322 = ( ~n744 & n6425 ) | ( ~n744 & n8418 ) | ( n6425 & n8418 ) ;
  assign n28323 = n28322 ^ n24985 ^ n13070 ;
  assign n28324 = n11669 ^ n8605 ^ n7992 ;
  assign n28325 = ~n9114 & n28324 ;
  assign n28326 = n28325 ^ n11064 ^ n8613 ;
  assign n28327 = n3154 | n11703 ;
  assign n28328 = n28327 ^ n22505 ^ 1'b0 ;
  assign n28329 = ( n16688 & ~n28326 ) | ( n16688 & n28328 ) | ( ~n28326 & n28328 ) ;
  assign n28330 = ~n6083 & n25095 ;
  assign n28331 = ( ~n5235 & n8464 ) | ( ~n5235 & n13020 ) | ( n8464 & n13020 ) ;
  assign n28332 = ~n2920 & n11949 ;
  assign n28333 = ( n10414 & n28331 ) | ( n10414 & n28332 ) | ( n28331 & n28332 ) ;
  assign n28334 = n28333 ^ n24535 ^ 1'b0 ;
  assign n28335 = n28330 | n28334 ;
  assign n28336 = n8683 | n28335 ;
  assign n28337 = n23978 & ~n28336 ;
  assign n28340 = n9712 ^ n872 ^ 1'b0 ;
  assign n28338 = n24779 ^ n5080 ^ 1'b0 ;
  assign n28339 = n16429 & n28338 ;
  assign n28341 = n28340 ^ n28339 ^ 1'b0 ;
  assign n28342 = ~n12238 & n28341 ;
  assign n28343 = n28342 ^ n17332 ^ 1'b0 ;
  assign n28344 = n28343 ^ n19592 ^ n11334 ;
  assign n28345 = ( n1023 & n11934 ) | ( n1023 & ~n25641 ) | ( n11934 & ~n25641 ) ;
  assign n28346 = n16967 | n18707 ;
  assign n28347 = n28346 ^ n16714 ^ 1'b0 ;
  assign n28348 = n26911 ^ n17163 ^ n5142 ;
  assign n28349 = n28348 ^ n18722 ^ 1'b0 ;
  assign n28350 = ( ~x166 & n5599 ) | ( ~x166 & n8193 ) | ( n5599 & n8193 ) ;
  assign n28351 = n4526 ^ n4083 ^ x34 ;
  assign n28352 = n28351 ^ n25232 ^ 1'b0 ;
  assign n28353 = n18651 | n28352 ;
  assign n28354 = n3335 | n3937 ;
  assign n28355 = n28354 ^ n7730 ^ 1'b0 ;
  assign n28356 = ( n4748 & n18116 ) | ( n4748 & ~n28355 ) | ( n18116 & ~n28355 ) ;
  assign n28357 = n1018 & n15196 ;
  assign n28358 = ( n22582 & n28356 ) | ( n22582 & ~n28357 ) | ( n28356 & ~n28357 ) ;
  assign n28359 = n22714 ^ n20148 ^ n3471 ;
  assign n28360 = ( n3934 & n6463 ) | ( n3934 & n15109 ) | ( n6463 & n15109 ) ;
  assign n28361 = ~n28359 & n28360 ;
  assign n28362 = n364 | n11291 ;
  assign n28363 = n28362 ^ n12637 ^ n12589 ;
  assign n28364 = ( n6439 & n23379 ) | ( n6439 & ~n25198 ) | ( n23379 & ~n25198 ) ;
  assign n28368 = n12320 & ~n21481 ;
  assign n28365 = n13916 ^ n5609 ^ 1'b0 ;
  assign n28366 = n7114 & n28365 ;
  assign n28367 = ( n3878 & n17953 ) | ( n3878 & ~n28366 ) | ( n17953 & ~n28366 ) ;
  assign n28369 = n28368 ^ n28367 ^ 1'b0 ;
  assign n28370 = n20140 ^ n19548 ^ n5145 ;
  assign n28374 = n10880 ^ n945 ^ 1'b0 ;
  assign n28371 = ~n1866 & n6340 ;
  assign n28372 = n1509 & n28371 ;
  assign n28373 = n28372 ^ n7551 ^ n4540 ;
  assign n28375 = n28374 ^ n28373 ^ 1'b0 ;
  assign n28376 = n11774 ^ n5655 ^ n2425 ;
  assign n28377 = ( n13651 & n28375 ) | ( n13651 & ~n28376 ) | ( n28375 & ~n28376 ) ;
  assign n28378 = ( n8717 & ~n22807 ) | ( n8717 & n28377 ) | ( ~n22807 & n28377 ) ;
  assign n28379 = n11673 ^ n3808 ^ 1'b0 ;
  assign n28380 = n10584 & ~n28379 ;
  assign n28381 = ( n5052 & n22568 ) | ( n5052 & ~n28380 ) | ( n22568 & ~n28380 ) ;
  assign n28382 = n2021 & n12614 ;
  assign n28383 = n28382 ^ n1694 ^ 1'b0 ;
  assign n28384 = n28383 ^ n19762 ^ n1355 ;
  assign n28385 = ( n5311 & n24831 ) | ( n5311 & ~n28384 ) | ( n24831 & ~n28384 ) ;
  assign n28386 = ~n919 & n3337 ;
  assign n28387 = n28386 ^ n13712 ^ 1'b0 ;
  assign n28388 = n28387 ^ n20427 ^ 1'b0 ;
  assign n28389 = n15911 ^ n9370 ^ 1'b0 ;
  assign n28390 = x77 & n26138 ;
  assign n28391 = n17501 ^ n14458 ^ 1'b0 ;
  assign n28392 = ( n16485 & n19120 ) | ( n16485 & n26951 ) | ( n19120 & n26951 ) ;
  assign n28393 = ( ~n14613 & n17218 ) | ( ~n14613 & n21604 ) | ( n17218 & n21604 ) ;
  assign n28394 = ( n2527 & n15309 ) | ( n2527 & ~n27023 ) | ( n15309 & ~n27023 ) ;
  assign n28395 = n28394 ^ n22399 ^ n18453 ;
  assign n28396 = ( n17358 & ~n24936 ) | ( n17358 & n28395 ) | ( ~n24936 & n28395 ) ;
  assign n28397 = n8967 & n17166 ;
  assign n28398 = n3374 & ~n17283 ;
  assign n28399 = ~n28397 & n28398 ;
  assign n28400 = n28399 ^ n10371 ^ 1'b0 ;
  assign n28401 = n1347 | n4196 ;
  assign n28402 = n24518 | n28401 ;
  assign n28403 = ( n1979 & n16735 ) | ( n1979 & n28402 ) | ( n16735 & n28402 ) ;
  assign n28404 = ( ~n3733 & n10399 ) | ( ~n3733 & n10501 ) | ( n10399 & n10501 ) ;
  assign n28408 = ~n3113 & n27993 ;
  assign n28405 = ( n1920 & n4349 ) | ( n1920 & ~n7151 ) | ( n4349 & ~n7151 ) ;
  assign n28406 = ( ~n9597 & n14731 ) | ( ~n9597 & n28405 ) | ( n14731 & n28405 ) ;
  assign n28407 = n7031 & n28406 ;
  assign n28409 = n28408 ^ n28407 ^ 1'b0 ;
  assign n28410 = n6386 ^ n5488 ^ n770 ;
  assign n28411 = n28410 ^ n15545 ^ 1'b0 ;
  assign n28412 = ~n27028 & n28411 ;
  assign n28413 = n27689 & n28412 ;
  assign n28414 = n28413 ^ n12998 ^ 1'b0 ;
  assign n28418 = n7733 & ~n26889 ;
  assign n28419 = n28418 ^ n6460 ^ 1'b0 ;
  assign n28415 = n586 & n1434 ;
  assign n28416 = n10066 & n28415 ;
  assign n28417 = n14586 & ~n28416 ;
  assign n28420 = n28419 ^ n28417 ^ 1'b0 ;
  assign n28421 = x209 & ~n9866 ;
  assign n28422 = ~n2358 & n28421 ;
  assign n28423 = ( n8383 & n28420 ) | ( n8383 & ~n28422 ) | ( n28420 & ~n28422 ) ;
  assign n28427 = n12000 | n12927 ;
  assign n28424 = n1003 & n20597 ;
  assign n28425 = ( n8756 & n21769 ) | ( n8756 & ~n28424 ) | ( n21769 & ~n28424 ) ;
  assign n28426 = n24470 | n28425 ;
  assign n28428 = n28427 ^ n28426 ^ 1'b0 ;
  assign n28429 = n21116 ^ n15663 ^ n15496 ;
  assign n28430 = n28429 ^ n13883 ^ n2977 ;
  assign n28431 = ( n653 & n1349 ) | ( n653 & ~n24965 ) | ( n1349 & ~n24965 ) ;
  assign n28432 = n1367 & ~n6538 ;
  assign n28433 = n28432 ^ n12715 ^ 1'b0 ;
  assign n28434 = n28433 ^ n19357 ^ 1'b0 ;
  assign n28435 = n26743 ^ n25078 ^ n12019 ;
  assign n28440 = n6615 ^ n1645 ^ 1'b0 ;
  assign n28438 = n11891 ^ n11221 ^ n841 ;
  assign n28436 = n26087 ^ n5686 ^ 1'b0 ;
  assign n28437 = n23773 & n28436 ;
  assign n28439 = n28438 ^ n28437 ^ n16256 ;
  assign n28441 = n28440 ^ n28439 ^ n9360 ;
  assign n28448 = n18917 | n19419 ;
  assign n28449 = n17677 | n27159 ;
  assign n28450 = n28448 | n28449 ;
  assign n28442 = n2311 | n3487 ;
  assign n28443 = n18324 | n28442 ;
  assign n28444 = ( n2550 & ~n14179 ) | ( n2550 & n28443 ) | ( ~n14179 & n28443 ) ;
  assign n28445 = n16294 ^ n3209 ^ 1'b0 ;
  assign n28446 = n28444 & n28445 ;
  assign n28447 = ~n16488 & n28446 ;
  assign n28451 = n28450 ^ n28447 ^ 1'b0 ;
  assign n28458 = n24053 ^ n3228 ^ n642 ;
  assign n28452 = n3557 | n3775 ;
  assign n28453 = n18191 | n28452 ;
  assign n28454 = n2463 & n4754 ;
  assign n28455 = n3366 & n28454 ;
  assign n28456 = n28455 ^ n6188 ^ 1'b0 ;
  assign n28457 = n28453 & n28456 ;
  assign n28459 = n28458 ^ n28457 ^ n11991 ;
  assign n28460 = ( n3083 & ~n11137 ) | ( n3083 & n15952 ) | ( ~n11137 & n15952 ) ;
  assign n28461 = n13075 & ~n22089 ;
  assign n28462 = x191 & ~n580 ;
  assign n28463 = n28462 ^ n12663 ^ n11924 ;
  assign n28464 = n4316 | n28463 ;
  assign n28465 = n25123 ^ n19672 ^ n15664 ;
  assign n28466 = n28465 ^ n10495 ^ n4676 ;
  assign n28467 = n17850 ^ n12818 ^ n9313 ;
  assign n28468 = n10955 ^ n7754 ^ n3291 ;
  assign n28469 = n14232 ^ n1433 ^ 1'b0 ;
  assign n28470 = n4592 & n16379 ;
  assign n28471 = n28470 ^ x49 ^ 1'b0 ;
  assign n28472 = n10936 | n28471 ;
  assign n28473 = x237 | n28472 ;
  assign n28474 = ( n336 & ~n24338 ) | ( n336 & n25882 ) | ( ~n24338 & n25882 ) ;
  assign n28475 = n1592 | n28474 ;
  assign n28476 = n28473 | n28475 ;
  assign n28477 = n2515 | n7107 ;
  assign n28478 = n28477 ^ n2222 ^ 1'b0 ;
  assign n28479 = ( n2402 & ~n16925 ) | ( n2402 & n28478 ) | ( ~n16925 & n28478 ) ;
  assign n28480 = n14921 ^ n3628 ^ 1'b0 ;
  assign n28483 = n25096 ^ n20330 ^ 1'b0 ;
  assign n28481 = n6480 & ~n22310 ;
  assign n28482 = ( ~n17032 & n20623 ) | ( ~n17032 & n28481 ) | ( n20623 & n28481 ) ;
  assign n28484 = n28483 ^ n28482 ^ n2463 ;
  assign n28485 = n3701 ^ n1006 ^ 1'b0 ;
  assign n28486 = n1511 & n28485 ;
  assign n28487 = n28486 ^ n9020 ^ x49 ;
  assign n28488 = ( n14136 & ~n18843 ) | ( n14136 & n28487 ) | ( ~n18843 & n28487 ) ;
  assign n28489 = n9318 ^ n4805 ^ 1'b0 ;
  assign n28490 = ~n1200 & n28489 ;
  assign n28491 = n25681 ^ n21710 ^ n21442 ;
  assign n28492 = n23802 & ~n27785 ;
  assign n28493 = ~x129 & n28492 ;
  assign n28494 = n11516 ^ n3841 ^ n1789 ;
  assign n28495 = n28494 ^ n21532 ^ 1'b0 ;
  assign n28496 = n11540 ^ n8166 ^ n7659 ;
  assign n28498 = n12406 ^ n9550 ^ x218 ;
  assign n28497 = n20553 & n21778 ;
  assign n28499 = n28498 ^ n28497 ^ 1'b0 ;
  assign n28500 = n25160 ^ n7743 ^ n3601 ;
  assign n28501 = ( n4726 & ~n9949 ) | ( n4726 & n28500 ) | ( ~n9949 & n28500 ) ;
  assign n28502 = n28501 ^ n26806 ^ 1'b0 ;
  assign n28503 = n14497 ^ n7292 ^ n1809 ;
  assign n28504 = x134 & ~n28503 ;
  assign n28505 = n28504 ^ n3597 ^ 1'b0 ;
  assign n28506 = n28505 ^ n26514 ^ n22017 ;
  assign n28507 = n10235 & ~n22184 ;
  assign n28508 = n28507 ^ n9209 ^ n8635 ;
  assign n28509 = n28508 ^ n5929 ^ 1'b0 ;
  assign n28510 = n6673 & n22028 ;
  assign n28511 = ( n14887 & ~n15386 ) | ( n14887 & n28510 ) | ( ~n15386 & n28510 ) ;
  assign n28512 = n28511 ^ n26705 ^ n24703 ;
  assign n28513 = n22553 ^ n8432 ^ n7037 ;
  assign n28514 = ( n1121 & ~n1554 ) | ( n1121 & n28513 ) | ( ~n1554 & n28513 ) ;
  assign n28515 = n28514 ^ n3258 ^ 1'b0 ;
  assign n28516 = n8508 & n18905 ;
  assign n28517 = n25489 & n28516 ;
  assign n28518 = n18448 | n28517 ;
  assign n28519 = n28518 ^ n20835 ^ 1'b0 ;
  assign n28522 = ( ~n7204 & n8697 ) | ( ~n7204 & n19911 ) | ( n8697 & n19911 ) ;
  assign n28523 = ( ~n4540 & n10543 ) | ( ~n4540 & n28522 ) | ( n10543 & n28522 ) ;
  assign n28520 = n8571 | n8954 ;
  assign n28521 = n28520 ^ n19241 ^ 1'b0 ;
  assign n28524 = n28523 ^ n28521 ^ n3214 ;
  assign n28525 = n28524 ^ n9782 ^ n7565 ;
  assign n28526 = ( ~n6735 & n28519 ) | ( ~n6735 & n28525 ) | ( n28519 & n28525 ) ;
  assign n28527 = ( n868 & ~n17587 ) | ( n868 & n21015 ) | ( ~n17587 & n21015 ) ;
  assign n28528 = n28527 ^ n1641 ^ 1'b0 ;
  assign n28531 = n6490 ^ n3315 ^ 1'b0 ;
  assign n28529 = n9412 ^ n6402 ^ 1'b0 ;
  assign n28530 = n14515 & n28529 ;
  assign n28532 = n28531 ^ n28530 ^ 1'b0 ;
  assign n28533 = ~n8701 & n26607 ;
  assign n28536 = n21172 ^ n478 ^ 1'b0 ;
  assign n28537 = n895 | n1124 ;
  assign n28538 = n28537 ^ n8311 ^ n5829 ;
  assign n28539 = ( n581 & n7984 ) | ( n581 & ~n28538 ) | ( n7984 & ~n28538 ) ;
  assign n28540 = ( n27272 & n28536 ) | ( n27272 & n28539 ) | ( n28536 & n28539 ) ;
  assign n28534 = n26228 ^ n25138 ^ n19469 ;
  assign n28535 = n28534 ^ n19015 ^ 1'b0 ;
  assign n28541 = n28540 ^ n28535 ^ n6701 ;
  assign n28542 = n22578 ^ n8934 ^ n6138 ;
  assign n28543 = ( n1777 & n8692 ) | ( n1777 & n8818 ) | ( n8692 & n8818 ) ;
  assign n28544 = n22882 ^ n13779 ^ n6944 ;
  assign n28545 = ( n2552 & n28543 ) | ( n2552 & ~n28544 ) | ( n28543 & ~n28544 ) ;
  assign n28546 = n6954 ^ n6490 ^ 1'b0 ;
  assign n28547 = n1268 | n28546 ;
  assign n28548 = n22167 & ~n28547 ;
  assign n28549 = ~n594 & n28548 ;
  assign n28550 = n28549 ^ n480 ^ 1'b0 ;
  assign n28551 = n10088 | n28550 ;
  assign n28552 = n6913 | n13148 ;
  assign n28553 = n28552 ^ n26961 ^ 1'b0 ;
  assign n28554 = n21259 ^ n7374 ^ x106 ;
  assign n28555 = n12230 | n24256 ;
  assign n28556 = n13398 | n28555 ;
  assign n28557 = n28554 & ~n28556 ;
  assign n28558 = ( n4978 & n19729 ) | ( n4978 & n22485 ) | ( n19729 & n22485 ) ;
  assign n28559 = n17272 ^ n14631 ^ 1'b0 ;
  assign n28560 = n28558 | n28559 ;
  assign n28561 = n28560 ^ n9499 ^ n3572 ;
  assign n28562 = n15995 & n28561 ;
  assign n28563 = ~x212 & n28562 ;
  assign n28564 = n16039 ^ n9484 ^ n9200 ;
  assign n28565 = ( n23612 & n27848 ) | ( n23612 & n28564 ) | ( n27848 & n28564 ) ;
  assign n28566 = n8905 ^ n1088 ^ 1'b0 ;
  assign n28567 = ~n325 & n661 ;
  assign n28568 = ~n28566 & n28567 ;
  assign n28569 = n19282 | n28568 ;
  assign n28570 = n28565 & ~n28569 ;
  assign n28572 = n7061 & n7670 ;
  assign n28573 = ( n8881 & ~n11781 ) | ( n8881 & n28572 ) | ( ~n11781 & n28572 ) ;
  assign n28574 = n6745 & n28573 ;
  assign n28575 = n28574 ^ n1194 ^ 1'b0 ;
  assign n28571 = n10519 ^ n8526 ^ n7348 ;
  assign n28576 = n28575 ^ n28571 ^ n10756 ;
  assign n28577 = n28576 ^ n14292 ^ 1'b0 ;
  assign n28578 = n9579 & ~n28577 ;
  assign n28580 = n6776 ^ n6649 ^ n3591 ;
  assign n28581 = ~n5638 & n28580 ;
  assign n28579 = n12502 ^ n11645 ^ n3358 ;
  assign n28582 = n28581 ^ n28579 ^ n14749 ;
  assign n28583 = n12310 ^ n5296 ^ 1'b0 ;
  assign n28586 = n16917 ^ n4229 ^ n1003 ;
  assign n28584 = n22356 ^ n2766 ^ 1'b0 ;
  assign n28585 = n16503 & ~n28584 ;
  assign n28587 = n28586 ^ n28585 ^ 1'b0 ;
  assign n28588 = n1227 | n28587 ;
  assign n28589 = ( n15115 & n20095 ) | ( n15115 & n28588 ) | ( n20095 & n28588 ) ;
  assign n28590 = n5199 | n5538 ;
  assign n28591 = ( n17036 & n20576 ) | ( n17036 & ~n28590 ) | ( n20576 & ~n28590 ) ;
  assign n28592 = n17090 ^ n12004 ^ 1'b0 ;
  assign n28593 = n28592 ^ n13226 ^ n6095 ;
  assign n28594 = ~n27851 & n28593 ;
  assign n28595 = ( n3645 & n28591 ) | ( n3645 & n28594 ) | ( n28591 & n28594 ) ;
  assign n28596 = ( n6136 & n8475 ) | ( n6136 & n10067 ) | ( n8475 & n10067 ) ;
  assign n28597 = ( n15067 & ~n19142 ) | ( n15067 & n25026 ) | ( ~n19142 & n25026 ) ;
  assign n28600 = ~n13084 & n15840 ;
  assign n28598 = n23931 ^ n5976 ^ 1'b0 ;
  assign n28599 = n5340 & ~n28598 ;
  assign n28601 = n28600 ^ n28599 ^ n15760 ;
  assign n28602 = n2876 | n4916 ;
  assign n28603 = n28602 ^ n20580 ^ 1'b0 ;
  assign n28604 = n16515 | n28603 ;
  assign n28605 = n28604 ^ n11750 ^ n3369 ;
  assign n28606 = ( n4529 & n6033 ) | ( n4529 & ~n27839 ) | ( n6033 & ~n27839 ) ;
  assign n28607 = n8104 | n28606 ;
  assign n28608 = n26905 ^ n5076 ^ 1'b0 ;
  assign n28609 = n27940 & ~n28608 ;
  assign n28610 = n1915 | n27431 ;
  assign n28611 = ( n6955 & n12227 ) | ( n6955 & ~n15214 ) | ( n12227 & ~n15214 ) ;
  assign n28612 = ( ~n16839 & n17731 ) | ( ~n16839 & n23947 ) | ( n17731 & n23947 ) ;
  assign n28613 = n12455 ^ n906 ^ n370 ;
  assign n28614 = n5415 & n18152 ;
  assign n28615 = ( ~n3643 & n14023 ) | ( ~n3643 & n28614 ) | ( n14023 & n28614 ) ;
  assign n28616 = ( n14836 & n23561 ) | ( n14836 & n28615 ) | ( n23561 & n28615 ) ;
  assign n28618 = n12394 | n13488 ;
  assign n28617 = n8522 | n24852 ;
  assign n28619 = n28618 ^ n28617 ^ 1'b0 ;
  assign n28621 = n2142 & ~n13880 ;
  assign n28620 = ( n3841 & n18285 ) | ( n3841 & ~n20336 ) | ( n18285 & ~n20336 ) ;
  assign n28622 = n28621 ^ n28620 ^ n11747 ;
  assign n28623 = n331 & n12010 ;
  assign n28624 = n28623 ^ n3384 ^ 1'b0 ;
  assign n28625 = ~n3572 & n6618 ;
  assign n28626 = n863 & n1979 ;
  assign n28627 = n28626 ^ n28498 ^ 1'b0 ;
  assign n28628 = n28625 | n28627 ;
  assign n28629 = n23263 ^ n18201 ^ 1'b0 ;
  assign n28630 = n12420 & ~n28629 ;
  assign n28631 = ( n7036 & n28628 ) | ( n7036 & ~n28630 ) | ( n28628 & ~n28630 ) ;
  assign n28632 = n6669 & n20405 ;
  assign n28633 = ~n10541 & n28632 ;
  assign n28636 = n531 & ~n15278 ;
  assign n28634 = n7144 | n14782 ;
  assign n28635 = n28634 ^ n24770 ^ 1'b0 ;
  assign n28637 = n28636 ^ n28635 ^ n4858 ;
  assign n28638 = ~n2128 & n3255 ;
  assign n28639 = n15023 ^ n7727 ^ 1'b0 ;
  assign n28640 = n28638 | n28639 ;
  assign n28641 = ( n17045 & n28637 ) | ( n17045 & ~n28640 ) | ( n28637 & ~n28640 ) ;
  assign n28642 = n12379 | n17588 ;
  assign n28643 = n13827 & ~n28642 ;
  assign n28644 = n2015 & ~n28643 ;
  assign n28645 = n6899 & n12665 ;
  assign n28646 = ( n15434 & n26989 ) | ( n15434 & ~n28645 ) | ( n26989 & ~n28645 ) ;
  assign n28647 = n4339 ^ n4245 ^ n642 ;
  assign n28648 = n28647 ^ n22518 ^ n6592 ;
  assign n28654 = n19338 ^ n16023 ^ n11725 ;
  assign n28652 = n13210 & n18397 ;
  assign n28653 = n28652 ^ n19445 ^ 1'b0 ;
  assign n28650 = n10394 ^ n3617 ^ 1'b0 ;
  assign n28649 = x183 & n19257 ;
  assign n28651 = n28650 ^ n28649 ^ n7799 ;
  assign n28655 = n28654 ^ n28653 ^ n28651 ;
  assign n28656 = n18821 ^ n11811 ^ n5224 ;
  assign n28657 = n14402 & n28656 ;
  assign n28658 = ~n4039 & n4967 ;
  assign n28659 = n28658 ^ n13478 ^ n5176 ;
  assign n28662 = ( n3399 & n13661 ) | ( n3399 & ~n17188 ) | ( n13661 & ~n17188 ) ;
  assign n28660 = n13803 & ~n20067 ;
  assign n28661 = n14696 & n28660 ;
  assign n28663 = n28662 ^ n28661 ^ n17026 ;
  assign n28667 = n24502 ^ n22512 ^ n14619 ;
  assign n28664 = ( n5376 & n5711 ) | ( n5376 & n8156 ) | ( n5711 & n8156 ) ;
  assign n28665 = ( ~n10615 & n22319 ) | ( ~n10615 & n28664 ) | ( n22319 & n28664 ) ;
  assign n28666 = n28665 ^ n18530 ^ 1'b0 ;
  assign n28668 = n28667 ^ n28666 ^ x4 ;
  assign n28669 = n16565 ^ n10848 ^ n487 ;
  assign n28670 = n18760 ^ n4625 ^ 1'b0 ;
  assign n28671 = n23187 ^ n2336 ^ 1'b0 ;
  assign n28672 = n28670 & ~n28671 ;
  assign n28673 = n14792 ^ n1565 ^ 1'b0 ;
  assign n28674 = n28673 ^ n8165 ^ n7330 ;
  assign n28675 = ( n14186 & ~n27140 ) | ( n14186 & n28674 ) | ( ~n27140 & n28674 ) ;
  assign n28676 = ( n28669 & n28672 ) | ( n28669 & n28675 ) | ( n28672 & n28675 ) ;
  assign n28677 = n14944 ^ n11507 ^ n5766 ;
  assign n28678 = n28677 ^ n3250 ^ n2601 ;
  assign n28679 = ( ~n3887 & n14595 ) | ( ~n3887 & n28678 ) | ( n14595 & n28678 ) ;
  assign n28680 = ( n7253 & n14963 ) | ( n7253 & ~n23187 ) | ( n14963 & ~n23187 ) ;
  assign n28681 = n28680 ^ n4942 ^ 1'b0 ;
  assign n28682 = n3402 | n14672 ;
  assign n28685 = n15816 ^ n6690 ^ n2815 ;
  assign n28683 = n23410 ^ n19945 ^ 1'b0 ;
  assign n28684 = n7832 & ~n28683 ;
  assign n28686 = n28685 ^ n28684 ^ n22328 ;
  assign n28696 = n28180 ^ n434 ^ 1'b0 ;
  assign n28687 = n2864 & n13651 ;
  assign n28688 = ~n16671 & n28687 ;
  assign n28689 = n10656 | n28688 ;
  assign n28690 = n28689 ^ n6985 ^ 1'b0 ;
  assign n28691 = n21185 ^ n17339 ^ n11534 ;
  assign n28692 = n28691 ^ x57 ^ 1'b0 ;
  assign n28693 = ~n25614 & n28692 ;
  assign n28694 = n28693 ^ n19045 ^ 1'b0 ;
  assign n28695 = n28690 & n28694 ;
  assign n28697 = n28696 ^ n28695 ^ n13957 ;
  assign n28698 = n9350 | n15096 ;
  assign n28699 = ~n2638 & n10595 ;
  assign n28700 = ~n16405 & n28699 ;
  assign n28701 = ( n9011 & ~n28698 ) | ( n9011 & n28700 ) | ( ~n28698 & n28700 ) ;
  assign n28702 = n11923 ^ n3617 ^ 1'b0 ;
  assign n28703 = ( ~n2598 & n8199 ) | ( ~n2598 & n12211 ) | ( n8199 & n12211 ) ;
  assign n28704 = n11998 | n28703 ;
  assign n28705 = ~n8345 & n28704 ;
  assign n28707 = n8475 | n15905 ;
  assign n28706 = n15930 ^ n14296 ^ n11073 ;
  assign n28708 = n28707 ^ n28706 ^ n14879 ;
  assign n28715 = n27363 ^ n21615 ^ x73 ;
  assign n28709 = n6450 ^ n3722 ^ 1'b0 ;
  assign n28710 = n7983 & ~n28709 ;
  assign n28711 = ( ~n6325 & n12493 ) | ( ~n6325 & n28556 ) | ( n12493 & n28556 ) ;
  assign n28712 = n28711 ^ n28621 ^ 1'b0 ;
  assign n28713 = n16492 & ~n28712 ;
  assign n28714 = ( n12366 & n28710 ) | ( n12366 & ~n28713 ) | ( n28710 & ~n28713 ) ;
  assign n28716 = n28715 ^ n28714 ^ 1'b0 ;
  assign n28717 = n10582 & ~n28716 ;
  assign n28718 = ~n6197 & n13460 ;
  assign n28719 = n28718 ^ n805 ^ 1'b0 ;
  assign n28720 = n11651 ^ x111 ^ 1'b0 ;
  assign n28721 = n22716 & ~n28720 ;
  assign n28722 = n28721 ^ n11573 ^ n3538 ;
  assign n28723 = n28719 | n28722 ;
  assign n28724 = n28723 ^ n23388 ^ 1'b0 ;
  assign n28725 = n11930 | n28724 ;
  assign n28726 = n22589 & ~n28725 ;
  assign n28727 = n26005 ^ n11603 ^ n3062 ;
  assign n28728 = n28727 ^ n18848 ^ 1'b0 ;
  assign n28729 = n28728 ^ n28684 ^ n17945 ;
  assign n28730 = n28729 ^ n25349 ^ n21742 ;
  assign n28731 = n26169 ^ n10912 ^ 1'b0 ;
  assign n28732 = ( ~n6678 & n19000 ) | ( ~n6678 & n21290 ) | ( n19000 & n21290 ) ;
  assign n28733 = n11768 ^ n1233 ^ 1'b0 ;
  assign n28734 = ~n18687 & n28733 ;
  assign n28735 = n28734 ^ n11602 ^ 1'b0 ;
  assign n28736 = n6473 & ~n14438 ;
  assign n28737 = n7120 & n28736 ;
  assign n28738 = n9962 & n16322 ;
  assign n28739 = ( n21866 & n25008 ) | ( n21866 & n28738 ) | ( n25008 & n28738 ) ;
  assign n28740 = ( n9863 & n10399 ) | ( n9863 & n12334 ) | ( n10399 & n12334 ) ;
  assign n28741 = ( n1385 & ~n18115 ) | ( n1385 & n18638 ) | ( ~n18115 & n18638 ) ;
  assign n28742 = ( ~n1631 & n6046 ) | ( ~n1631 & n19098 ) | ( n6046 & n19098 ) ;
  assign n28743 = n12195 ^ n6706 ^ n5056 ;
  assign n28744 = n28743 ^ n26349 ^ 1'b0 ;
  assign n28745 = n28744 ^ n21609 ^ 1'b0 ;
  assign n28746 = n6511 & ~n28745 ;
  assign n28747 = ( ~n7854 & n23474 ) | ( ~n7854 & n26898 ) | ( n23474 & n26898 ) ;
  assign n28748 = ~n11899 & n19352 ;
  assign n28749 = n2840 | n17153 ;
  assign n28750 = n28749 ^ n20504 ^ 1'b0 ;
  assign n28751 = n28750 ^ n27083 ^ n9531 ;
  assign n28752 = n22213 ^ n2995 ^ 1'b0 ;
  assign n28754 = ( n4801 & ~n5659 ) | ( n4801 & n18935 ) | ( ~n5659 & n18935 ) ;
  assign n28753 = n13761 ^ n10339 ^ 1'b0 ;
  assign n28755 = n28754 ^ n28753 ^ n28448 ;
  assign n28756 = ( n3275 & ~n4424 ) | ( n3275 & n28755 ) | ( ~n4424 & n28755 ) ;
  assign n28757 = ( n6841 & n28752 ) | ( n6841 & ~n28756 ) | ( n28752 & ~n28756 ) ;
  assign n28758 = n17299 ^ n8738 ^ n2974 ;
  assign n28759 = n8573 | n21790 ;
  assign n28760 = ~n405 & n20510 ;
  assign n28761 = ( ~n6460 & n25654 ) | ( ~n6460 & n28760 ) | ( n25654 & n28760 ) ;
  assign n28762 = ( n14591 & ~n26014 ) | ( n14591 & n26878 ) | ( ~n26014 & n26878 ) ;
  assign n28763 = n1279 & ~n11572 ;
  assign n28764 = n7428 & n28763 ;
  assign n28765 = ( n3180 & n10377 ) | ( n3180 & n12699 ) | ( n10377 & n12699 ) ;
  assign n28766 = ( n27558 & n28764 ) | ( n27558 & ~n28765 ) | ( n28764 & ~n28765 ) ;
  assign n28767 = ( n4499 & n4886 ) | ( n4499 & ~n13097 ) | ( n4886 & ~n13097 ) ;
  assign n28768 = ( ~n10380 & n15038 ) | ( ~n10380 & n26175 ) | ( n15038 & n26175 ) ;
  assign n28769 = n25791 ^ n3111 ^ n1783 ;
  assign n28770 = ( n286 & n429 ) | ( n286 & ~n447 ) | ( n429 & ~n447 ) ;
  assign n28771 = n23809 & n28770 ;
  assign n28772 = n28771 ^ n27518 ^ 1'b0 ;
  assign n28773 = ( n2408 & n28440 ) | ( n2408 & n28772 ) | ( n28440 & n28772 ) ;
  assign n28774 = n26685 ^ n4562 ^ 1'b0 ;
  assign n28775 = n28774 ^ x122 ^ 1'b0 ;
  assign n28776 = n3715 & n4677 ;
  assign n28777 = n28776 ^ n4160 ^ 1'b0 ;
  assign n28778 = ( ~n550 & n15784 ) | ( ~n550 & n28777 ) | ( n15784 & n28777 ) ;
  assign n28779 = n16870 ^ n6703 ^ n5511 ;
  assign n28780 = n28779 ^ n11414 ^ 1'b0 ;
  assign n28781 = ( n2980 & ~n14653 ) | ( n2980 & n19441 ) | ( ~n14653 & n19441 ) ;
  assign n28782 = ( n8711 & n10852 ) | ( n8711 & ~n28781 ) | ( n10852 & ~n28781 ) ;
  assign n28783 = n16206 ^ n15032 ^ n8871 ;
  assign n28784 = ( ~n3927 & n8909 ) | ( ~n3927 & n28783 ) | ( n8909 & n28783 ) ;
  assign n28785 = n555 & n14861 ;
  assign n28786 = n10196 & n28785 ;
  assign n28787 = n28786 ^ n16607 ^ n3669 ;
  assign n28788 = ( n21313 & ~n22752 ) | ( n21313 & n28787 ) | ( ~n22752 & n28787 ) ;
  assign n28789 = ( n12673 & n12793 ) | ( n12673 & n20123 ) | ( n12793 & n20123 ) ;
  assign n28790 = n19725 ^ n12875 ^ n7436 ;
  assign n28791 = n12528 ^ n12039 ^ n2474 ;
  assign n28792 = n28791 ^ n25614 ^ n24581 ;
  assign n28793 = ( n21552 & ~n28790 ) | ( n21552 & n28792 ) | ( ~n28790 & n28792 ) ;
  assign n28794 = ( n498 & ~n9347 ) | ( n498 & n28793 ) | ( ~n9347 & n28793 ) ;
  assign n28795 = n28794 ^ n17605 ^ 1'b0 ;
  assign n28796 = n28789 | n28795 ;
  assign n28797 = n1332 & ~n7268 ;
  assign n28798 = ( ~n3304 & n7645 ) | ( ~n3304 & n27301 ) | ( n7645 & n27301 ) ;
  assign n28799 = n15805 ^ n3208 ^ 1'b0 ;
  assign n28800 = ~n28798 & n28799 ;
  assign n28801 = ( n6841 & n28797 ) | ( n6841 & n28800 ) | ( n28797 & n28800 ) ;
  assign n28802 = n1777 ^ x100 ^ 1'b0 ;
  assign n28803 = n28801 & ~n28802 ;
  assign n28804 = n21903 ^ n9692 ^ n1315 ;
  assign n28808 = ( ~n3391 & n4154 ) | ( ~n3391 & n4723 ) | ( n4154 & n4723 ) ;
  assign n28805 = n27799 ^ n5243 ^ n2230 ;
  assign n28806 = n28805 ^ n13744 ^ 1'b0 ;
  assign n28807 = n2625 & ~n28806 ;
  assign n28809 = n28808 ^ n28807 ^ n22299 ;
  assign n28810 = n3977 & n18124 ;
  assign n28811 = ~n18584 & n28810 ;
  assign n28814 = n8683 ^ n3774 ^ n1626 ;
  assign n28812 = ( n8681 & n12674 ) | ( n8681 & n16838 ) | ( n12674 & n16838 ) ;
  assign n28813 = ( n4636 & n11522 ) | ( n4636 & ~n28812 ) | ( n11522 & ~n28812 ) ;
  assign n28815 = n28814 ^ n28813 ^ n17877 ;
  assign n28816 = ( n15296 & ~n16615 ) | ( n15296 & n24487 ) | ( ~n16615 & n24487 ) ;
  assign n28817 = n28816 ^ n14004 ^ 1'b0 ;
  assign n28818 = ( ~n5079 & n28815 ) | ( ~n5079 & n28817 ) | ( n28815 & n28817 ) ;
  assign n28819 = ( ~n4099 & n7515 ) | ( ~n4099 & n28444 ) | ( n7515 & n28444 ) ;
  assign n28820 = n3860 ^ n2226 ^ n2019 ;
  assign n28821 = ( n5242 & n13580 ) | ( n5242 & ~n28820 ) | ( n13580 & ~n28820 ) ;
  assign n28822 = ( n19184 & ~n21179 ) | ( n19184 & n28821 ) | ( ~n21179 & n28821 ) ;
  assign n28823 = n25136 ^ n10170 ^ 1'b0 ;
  assign n28824 = n2485 | n28823 ;
  assign n28825 = n17962 & n20816 ;
  assign n28826 = n28825 ^ n27652 ^ 1'b0 ;
  assign n28827 = n5035 ^ n1459 ^ 1'b0 ;
  assign n28828 = n5502 & ~n8188 ;
  assign n28829 = n28828 ^ n7741 ^ 1'b0 ;
  assign n28830 = n15635 ^ n5732 ^ 1'b0 ;
  assign n28831 = n28830 ^ n8712 ^ 1'b0 ;
  assign n28832 = n6781 | n28831 ;
  assign n28833 = n12471 ^ n9919 ^ n861 ;
  assign n28834 = n18855 ^ n2845 ^ 1'b0 ;
  assign n28835 = n3071 | n28834 ;
  assign n28836 = ( ~n10738 & n14581 ) | ( ~n10738 & n15287 ) | ( n14581 & n15287 ) ;
  assign n28837 = n28836 ^ n12523 ^ n12217 ;
  assign n28838 = ( n6640 & n25432 ) | ( n6640 & n28837 ) | ( n25432 & n28837 ) ;
  assign n28839 = n7912 & n22433 ;
  assign n28840 = n28838 & n28839 ;
  assign n28841 = ( n28833 & ~n28835 ) | ( n28833 & n28840 ) | ( ~n28835 & n28840 ) ;
  assign n28842 = ( n8586 & ~n11811 ) | ( n8586 & n17423 ) | ( ~n11811 & n17423 ) ;
  assign n28843 = n23342 & ~n28842 ;
  assign n28844 = n25596 ^ n18818 ^ n17485 ;
  assign n28845 = n28844 ^ n24716 ^ n5487 ;
  assign n28846 = ( n1383 & n14242 ) | ( n1383 & n24323 ) | ( n14242 & n24323 ) ;
  assign n28847 = n28846 ^ n2962 ^ 1'b0 ;
  assign n28848 = n24635 ^ n5565 ^ n4481 ;
  assign n28849 = ( n1511 & n16610 ) | ( n1511 & ~n28848 ) | ( n16610 & ~n28848 ) ;
  assign n28850 = n600 & ~n14319 ;
  assign n28851 = n28850 ^ n28093 ^ 1'b0 ;
  assign n28852 = ( ~n28847 & n28849 ) | ( ~n28847 & n28851 ) | ( n28849 & n28851 ) ;
  assign n28853 = n27354 ^ n10969 ^ n3725 ;
  assign n28854 = n13292 ^ n5463 ^ 1'b0 ;
  assign n28855 = n7282 ^ n2848 ^ 1'b0 ;
  assign n28856 = ~n28854 & n28855 ;
  assign n28857 = n28856 ^ n5174 ^ n1544 ;
  assign n28858 = n22646 ^ n4156 ^ n2987 ;
  assign n28863 = ( n571 & n8418 ) | ( n571 & n10458 ) | ( n8418 & n10458 ) ;
  assign n28864 = ( n10330 & n16978 ) | ( n10330 & ~n28863 ) | ( n16978 & ~n28863 ) ;
  assign n28859 = n21483 ^ n19943 ^ n261 ;
  assign n28860 = n4874 | n20805 ;
  assign n28861 = n6817 | n28860 ;
  assign n28862 = ~n28859 & n28861 ;
  assign n28865 = n28864 ^ n28862 ^ 1'b0 ;
  assign n28866 = ( n28857 & n28858 ) | ( n28857 & ~n28865 ) | ( n28858 & ~n28865 ) ;
  assign n28867 = ( n12759 & n15629 ) | ( n12759 & n27471 ) | ( n15629 & n27471 ) ;
  assign n28868 = ( x1 & ~n6436 ) | ( x1 & n15099 ) | ( ~n6436 & n15099 ) ;
  assign n28869 = n14470 ^ n7435 ^ 1'b0 ;
  assign n28870 = n12237 ^ n6403 ^ n2670 ;
  assign n28871 = ( n2010 & ~n3774 ) | ( n2010 & n26593 ) | ( ~n3774 & n26593 ) ;
  assign n28872 = ( n1409 & n28870 ) | ( n1409 & n28871 ) | ( n28870 & n28871 ) ;
  assign n28873 = n1217 | n8687 ;
  assign n28874 = n3881 | n28873 ;
  assign n28875 = n28874 ^ n5928 ^ n1383 ;
  assign n28876 = n28875 ^ n13536 ^ n5248 ;
  assign n28877 = n13462 | n24545 ;
  assign n28878 = n20765 ^ n5520 ^ n1871 ;
  assign n28879 = n28878 ^ n6285 ^ x41 ;
  assign n28880 = n3734 | n11798 ;
  assign n28881 = n28880 ^ n8031 ^ 1'b0 ;
  assign n28882 = n28881 ^ n4000 ^ n406 ;
  assign n28883 = ( n9625 & ~n28879 ) | ( n9625 & n28882 ) | ( ~n28879 & n28882 ) ;
  assign n28884 = n20132 & n28883 ;
  assign n28885 = n19027 & n28884 ;
  assign n28886 = n15020 ^ n3515 ^ 1'b0 ;
  assign n28887 = n28886 ^ n14135 ^ 1'b0 ;
  assign n28888 = ~n5002 & n28887 ;
  assign n28889 = n9004 ^ n4493 ^ n4414 ;
  assign n28890 = n28889 ^ n27474 ^ 1'b0 ;
  assign n28891 = n28888 & ~n28890 ;
  assign n28892 = n15330 & ~n27636 ;
  assign n28893 = n28892 ^ n1910 ^ 1'b0 ;
  assign n28894 = ~n16201 & n28893 ;
  assign n28895 = n23731 ^ n12314 ^ n11892 ;
  assign n28896 = ( n1191 & ~n5037 ) | ( n1191 & n28895 ) | ( ~n5037 & n28895 ) ;
  assign n28897 = n23863 & ~n26954 ;
  assign n28898 = n28897 ^ n18058 ^ 1'b0 ;
  assign n28906 = ( ~n1747 & n10399 ) | ( ~n1747 & n14225 ) | ( n10399 & n14225 ) ;
  assign n28904 = n5937 & n12088 ;
  assign n28905 = n28904 ^ n5346 ^ 1'b0 ;
  assign n28899 = n16594 ^ n5366 ^ n1790 ;
  assign n28900 = n28899 ^ n16166 ^ 1'b0 ;
  assign n28901 = ~n19688 & n28900 ;
  assign n28902 = n21553 ^ n12823 ^ 1'b0 ;
  assign n28903 = n28901 & ~n28902 ;
  assign n28907 = n28906 ^ n28905 ^ n28903 ;
  assign n28912 = ( n2348 & n7099 ) | ( n2348 & n8512 ) | ( n7099 & n8512 ) ;
  assign n28913 = ( n3405 & ~n6240 ) | ( n3405 & n6716 ) | ( ~n6240 & n6716 ) ;
  assign n28914 = ( n408 & n2751 ) | ( n408 & ~n28913 ) | ( n2751 & ~n28913 ) ;
  assign n28915 = n28914 ^ n6164 ^ n2216 ;
  assign n28916 = ( n15883 & ~n28912 ) | ( n15883 & n28915 ) | ( ~n28912 & n28915 ) ;
  assign n28917 = n27790 ^ n12092 ^ n11636 ;
  assign n28918 = n28917 ^ n11029 ^ n6994 ;
  assign n28919 = ( n19406 & n28916 ) | ( n19406 & n28918 ) | ( n28916 & n28918 ) ;
  assign n28909 = ~n2960 & n9279 ;
  assign n28910 = n23455 & n28909 ;
  assign n28908 = ( n2285 & n13006 ) | ( n2285 & n16615 ) | ( n13006 & n16615 ) ;
  assign n28911 = n28910 ^ n28908 ^ n20704 ;
  assign n28920 = n28919 ^ n28911 ^ 1'b0 ;
  assign n28921 = n12321 | n26254 ;
  assign n28922 = n28921 ^ n19482 ^ 1'b0 ;
  assign n28923 = n4855 & ~n7006 ;
  assign n28924 = n2871 & n28923 ;
  assign n28925 = ~x112 & n28924 ;
  assign n28926 = n28925 ^ n14080 ^ 1'b0 ;
  assign n28927 = ( n919 & n9412 ) | ( n919 & n28926 ) | ( n9412 & n28926 ) ;
  assign n28928 = n12687 ^ n5623 ^ n4122 ;
  assign n28929 = n22777 ^ n13403 ^ 1'b0 ;
  assign n28930 = n8346 | n28929 ;
  assign n28931 = ~n349 & n17867 ;
  assign n28932 = n1716 & n28931 ;
  assign n28933 = n22363 ^ n2785 ^ 1'b0 ;
  assign n28934 = ( n18924 & n19736 ) | ( n18924 & ~n28933 ) | ( n19736 & ~n28933 ) ;
  assign n28935 = n1169 & ~n11071 ;
  assign n28936 = n28935 ^ n21936 ^ n10815 ;
  assign n28937 = n28936 ^ n12188 ^ 1'b0 ;
  assign n28938 = n26984 ^ n6029 ^ 1'b0 ;
  assign n28939 = n4045 & n28938 ;
  assign n28940 = n7623 & n28939 ;
  assign n28941 = n16551 ^ n14767 ^ n11962 ;
  assign n28942 = n14226 ^ n13189 ^ n11792 ;
  assign n28943 = n28942 ^ n14452 ^ 1'b0 ;
  assign n28944 = n28941 & n28943 ;
  assign n28945 = n16855 ^ n9416 ^ n3839 ;
  assign n28946 = n28945 ^ n20876 ^ n3678 ;
  assign n28947 = ( n10448 & ~n12709 ) | ( n10448 & n27436 ) | ( ~n12709 & n27436 ) ;
  assign n28948 = ( ~n4597 & n6525 ) | ( ~n4597 & n28947 ) | ( n6525 & n28947 ) ;
  assign n28949 = n28948 ^ n26228 ^ n1911 ;
  assign n28950 = n26540 ^ n22675 ^ n17217 ;
  assign n28951 = ( n1194 & n3542 ) | ( n1194 & ~n5580 ) | ( n3542 & ~n5580 ) ;
  assign n28952 = n28951 ^ n28498 ^ n20069 ;
  assign n28953 = n22141 ^ n13233 ^ n594 ;
  assign n28954 = n28953 ^ n28523 ^ 1'b0 ;
  assign n28955 = n21518 ^ n11957 ^ 1'b0 ;
  assign n28956 = n28954 | n28955 ;
  assign n28958 = ~n5006 & n6244 ;
  assign n28959 = ~n11636 & n28958 ;
  assign n28957 = n15268 ^ n11498 ^ 1'b0 ;
  assign n28960 = n28959 ^ n28957 ^ n10059 ;
  assign n28961 = ( n11690 & n16874 ) | ( n11690 & n28960 ) | ( n16874 & n28960 ) ;
  assign n28962 = ( ~n462 & n2907 ) | ( ~n462 & n6362 ) | ( n2907 & n6362 ) ;
  assign n28963 = n28962 ^ n27296 ^ n14022 ;
  assign n28964 = ( ~n4895 & n27771 ) | ( ~n4895 & n28963 ) | ( n27771 & n28963 ) ;
  assign n28968 = ( ~n10716 & n22132 ) | ( ~n10716 & n22465 ) | ( n22132 & n22465 ) ;
  assign n28967 = ( n10617 & n19098 ) | ( n10617 & n20673 ) | ( n19098 & n20673 ) ;
  assign n28969 = n28968 ^ n28967 ^ n8189 ;
  assign n28965 = n22740 ^ n6794 ^ 1'b0 ;
  assign n28966 = n2695 & n28965 ;
  assign n28970 = n28969 ^ n28966 ^ n15974 ;
  assign n28972 = ( ~n11011 & n13125 ) | ( ~n11011 & n26605 ) | ( n13125 & n26605 ) ;
  assign n28971 = n13510 & ~n15513 ;
  assign n28973 = n28972 ^ n28971 ^ 1'b0 ;
  assign n28974 = n28973 ^ n15172 ^ n13890 ;
  assign n28975 = n6864 ^ n5053 ^ n2835 ;
  assign n28976 = n27179 | n28975 ;
  assign n28977 = ( ~n9295 & n28974 ) | ( ~n9295 & n28976 ) | ( n28974 & n28976 ) ;
  assign n28978 = ~n5115 & n11433 ;
  assign n28979 = ~n4247 & n28978 ;
  assign n28980 = n28979 ^ n19662 ^ 1'b0 ;
  assign n28981 = ~n3804 & n28980 ;
  assign n28982 = n18209 ^ n283 ^ 1'b0 ;
  assign n28983 = n16345 ^ n15896 ^ n8871 ;
  assign n28984 = n28983 ^ n15494 ^ n8739 ;
  assign n28985 = n21530 & n26848 ;
  assign n28986 = n28985 ^ n16423 ^ 1'b0 ;
  assign n28987 = ( ~n6150 & n9976 ) | ( ~n6150 & n22727 ) | ( n9976 & n22727 ) ;
  assign n28988 = n28987 ^ n23516 ^ n8562 ;
  assign n28989 = ( n4202 & n20216 ) | ( n4202 & ~n28988 ) | ( n20216 & ~n28988 ) ;
  assign n28990 = ( n6598 & n13051 ) | ( n6598 & ~n23807 ) | ( n13051 & ~n23807 ) ;
  assign n28991 = n26782 ^ n3178 ^ 1'b0 ;
  assign n28992 = n19607 & ~n21216 ;
  assign n28993 = n16402 & n28992 ;
  assign n28994 = n5038 | n5390 ;
  assign n28995 = ( ~x91 & n3301 ) | ( ~x91 & n14268 ) | ( n3301 & n14268 ) ;
  assign n28996 = n28995 ^ n27700 ^ n17492 ;
  assign n28997 = n28994 & n28996 ;
  assign n28998 = ( n2956 & n4931 ) | ( n2956 & ~n28997 ) | ( n4931 & ~n28997 ) ;
  assign n28999 = n8186 ^ n6286 ^ n2035 ;
  assign n29000 = ( ~n3925 & n7390 ) | ( ~n3925 & n28999 ) | ( n7390 & n28999 ) ;
  assign n29001 = n5190 ^ n3725 ^ 1'b0 ;
  assign n29002 = n3969 & n29001 ;
  assign n29003 = ~n3939 & n5680 ;
  assign n29004 = ~n13948 & n29003 ;
  assign n29005 = n29004 ^ n947 ^ 1'b0 ;
  assign n29006 = n12050 & ~n29005 ;
  assign n29007 = n7740 & n29006 ;
  assign n29008 = n27791 & n29007 ;
  assign n29009 = ( ~n29000 & n29002 ) | ( ~n29000 & n29008 ) | ( n29002 & n29008 ) ;
  assign n29010 = n18972 ^ n9896 ^ 1'b0 ;
  assign n29011 = n12442 | n20958 ;
  assign n29012 = n22563 & n29011 ;
  assign n29013 = n29012 ^ x222 ^ 1'b0 ;
  assign n29014 = ( n2146 & n10345 ) | ( n2146 & ~n22585 ) | ( n10345 & ~n22585 ) ;
  assign n29015 = n14495 & n28141 ;
  assign n29016 = ~n8644 & n15370 ;
  assign n29017 = n29016 ^ n1910 ^ 1'b0 ;
  assign n29018 = n4401 & ~n20659 ;
  assign n29022 = n6918 | n18760 ;
  assign n29021 = ( n719 & ~n14606 ) | ( n719 & n25374 ) | ( ~n14606 & n25374 ) ;
  assign n29019 = n27988 ^ n24257 ^ n13008 ;
  assign n29020 = n29019 ^ n20207 ^ n18789 ;
  assign n29023 = n29022 ^ n29021 ^ n29020 ;
  assign n29024 = n11869 ^ n11392 ^ 1'b0 ;
  assign n29025 = ( n1252 & n5089 ) | ( n1252 & n29024 ) | ( n5089 & n29024 ) ;
  assign n29026 = n15813 ^ n7854 ^ n3542 ;
  assign n29031 = ( n15278 & n16951 ) | ( n15278 & ~n21423 ) | ( n16951 & ~n21423 ) ;
  assign n29032 = ( n977 & n10374 ) | ( n977 & ~n29031 ) | ( n10374 & ~n29031 ) ;
  assign n29033 = n29032 ^ n6279 ^ n1233 ;
  assign n29027 = ~n3279 & n23343 ;
  assign n29028 = n14727 & n29027 ;
  assign n29029 = ( n2858 & n27889 ) | ( n2858 & n29028 ) | ( n27889 & n29028 ) ;
  assign n29030 = n29029 ^ n19379 ^ n17006 ;
  assign n29034 = n29033 ^ n29030 ^ n28061 ;
  assign n29035 = n20054 | n27867 ;
  assign n29036 = n29035 ^ n1071 ^ 1'b0 ;
  assign n29037 = n2722 ^ n1928 ^ 1'b0 ;
  assign n29038 = n2280 & n7329 ;
  assign n29039 = ( n27759 & n29037 ) | ( n27759 & ~n29038 ) | ( n29037 & ~n29038 ) ;
  assign n29040 = n17795 ^ n4846 ^ n1381 ;
  assign n29041 = n6242 & ~n21866 ;
  assign n29042 = ~n3275 & n29041 ;
  assign n29043 = ( ~n6878 & n16926 ) | ( ~n6878 & n29042 ) | ( n16926 & n29042 ) ;
  assign n29044 = ( n10154 & ~n29040 ) | ( n10154 & n29043 ) | ( ~n29040 & n29043 ) ;
  assign n29045 = ( n3628 & n14369 ) | ( n3628 & n25522 ) | ( n14369 & n25522 ) ;
  assign n29046 = n7250 | n10543 ;
  assign n29047 = n29046 ^ n489 ^ 1'b0 ;
  assign n29048 = n5829 & ~n17801 ;
  assign n29049 = n12444 & n29048 ;
  assign n29050 = n870 & ~n29049 ;
  assign n29051 = n29050 ^ n3038 ^ 1'b0 ;
  assign n29052 = n17289 & ~n19929 ;
  assign n29053 = n29052 ^ n13809 ^ 1'b0 ;
  assign n29054 = n13375 | n29053 ;
  assign n29055 = ( n17254 & n20498 ) | ( n17254 & ~n29054 ) | ( n20498 & ~n29054 ) ;
  assign n29056 = n23304 ^ n8306 ^ n6694 ;
  assign n29061 = ~n3940 & n5206 ;
  assign n29062 = n29061 ^ n9390 ^ 1'b0 ;
  assign n29057 = n6064 & n9399 ;
  assign n29058 = n18725 & n29057 ;
  assign n29059 = n29058 ^ n20706 ^ n19315 ;
  assign n29060 = ( n13279 & ~n14221 ) | ( n13279 & n29059 ) | ( ~n14221 & n29059 ) ;
  assign n29063 = n29062 ^ n29060 ^ 1'b0 ;
  assign n29064 = n3520 | n29063 ;
  assign n29065 = n3455 ^ n1546 ^ 1'b0 ;
  assign n29066 = n14263 & n29065 ;
  assign n29068 = n28486 ^ n11891 ^ 1'b0 ;
  assign n29069 = n11851 | n29068 ;
  assign n29067 = n15086 ^ n13489 ^ n5751 ;
  assign n29070 = n29069 ^ n29067 ^ n6186 ;
  assign n29071 = ( n2116 & ~n3154 ) | ( n2116 & n29070 ) | ( ~n3154 & n29070 ) ;
  assign n29072 = n17919 ^ n9480 ^ x253 ;
  assign n29073 = n29072 ^ n9019 ^ n1730 ;
  assign n29074 = n19439 ^ n12825 ^ 1'b0 ;
  assign n29075 = n14932 ^ n4856 ^ 1'b0 ;
  assign n29076 = n28522 ^ n19045 ^ n4792 ;
  assign n29077 = ( x9 & ~n18306 ) | ( x9 & n29076 ) | ( ~n18306 & n29076 ) ;
  assign n29078 = ( n5944 & ~n8558 ) | ( n5944 & n19411 ) | ( ~n8558 & n19411 ) ;
  assign n29079 = n29078 ^ n19143 ^ n12831 ;
  assign n29080 = n29077 & ~n29079 ;
  assign n29081 = ~n9210 & n29080 ;
  assign n29082 = n10455 & n22872 ;
  assign n29083 = ~n6257 & n29082 ;
  assign n29086 = n2265 ^ n1573 ^ 1'b0 ;
  assign n29087 = ( ~n2632 & n19473 ) | ( ~n2632 & n29086 ) | ( n19473 & n29086 ) ;
  assign n29084 = n9838 ^ n9081 ^ n8327 ;
  assign n29085 = ( ~n1791 & n5219 ) | ( ~n1791 & n29084 ) | ( n5219 & n29084 ) ;
  assign n29088 = n29087 ^ n29085 ^ 1'b0 ;
  assign n29089 = ( ~n19051 & n19299 ) | ( ~n19051 & n29088 ) | ( n19299 & n29088 ) ;
  assign n29090 = n18565 ^ n10140 ^ 1'b0 ;
  assign n29091 = n8308 & n12642 ;
  assign n29092 = n29091 ^ n3535 ^ 1'b0 ;
  assign n29093 = ( n8209 & ~n23036 ) | ( n8209 & n29092 ) | ( ~n23036 & n29092 ) ;
  assign n29095 = n16945 ^ n5372 ^ 1'b0 ;
  assign n29096 = n7829 & ~n29095 ;
  assign n29097 = ( x78 & n10235 ) | ( x78 & ~n29096 ) | ( n10235 & ~n29096 ) ;
  assign n29094 = n24271 ^ n14625 ^ n8338 ;
  assign n29098 = n29097 ^ n29094 ^ n23465 ;
  assign n29099 = ( n6460 & n13396 ) | ( n6460 & ~n24827 ) | ( n13396 & ~n24827 ) ;
  assign n29100 = n29099 ^ n1946 ^ 1'b0 ;
  assign n29101 = n14487 ^ n6187 ^ n5936 ;
  assign n29102 = n4599 | n29101 ;
  assign n29103 = ~n948 & n17364 ;
  assign n29104 = n23853 ^ n10758 ^ n5038 ;
  assign n29105 = n29104 ^ n17691 ^ n6824 ;
  assign n29106 = n6161 & n22450 ;
  assign n29107 = n29105 & n29106 ;
  assign n29108 = ( n19790 & n29103 ) | ( n19790 & ~n29107 ) | ( n29103 & ~n29107 ) ;
  assign n29109 = ( n4613 & ~n5469 ) | ( n4613 & n6253 ) | ( ~n5469 & n6253 ) ;
  assign n29110 = n29109 ^ n14399 ^ x75 ;
  assign n29111 = n7743 ^ n7615 ^ 1'b0 ;
  assign n29112 = n14139 & ~n29111 ;
  assign n29113 = n29112 ^ n19711 ^ 1'b0 ;
  assign n29114 = n17332 ^ n2385 ^ 1'b0 ;
  assign n29115 = ( ~n503 & n1856 ) | ( ~n503 & n3146 ) | ( n1856 & n3146 ) ;
  assign n29116 = ( ~x66 & n15802 ) | ( ~x66 & n29115 ) | ( n15802 & n29115 ) ;
  assign n29117 = ( ~n1961 & n6979 ) | ( ~n1961 & n11124 ) | ( n6979 & n11124 ) ;
  assign n29118 = n29116 & n29117 ;
  assign n29119 = n29118 ^ n1244 ^ 1'b0 ;
  assign n29120 = n19813 ^ n18158 ^ n2729 ;
  assign n29125 = n1231 & ~n3230 ;
  assign n29126 = n29125 ^ n7450 ^ n4585 ;
  assign n29122 = n18868 ^ n17864 ^ 1'b0 ;
  assign n29123 = ~n26999 & n29122 ;
  assign n29121 = n3566 & ~n28161 ;
  assign n29124 = n29123 ^ n29121 ^ 1'b0 ;
  assign n29127 = n29126 ^ n29124 ^ n19609 ;
  assign n29128 = n29127 ^ n5201 ^ 1'b0 ;
  assign n29129 = ( n12198 & n29120 ) | ( n12198 & ~n29128 ) | ( n29120 & ~n29128 ) ;
  assign n29131 = n28405 ^ n4272 ^ 1'b0 ;
  assign n29132 = ( ~n19532 & n19554 ) | ( ~n19532 & n29131 ) | ( n19554 & n29131 ) ;
  assign n29130 = ( n13111 & n20588 ) | ( n13111 & n23387 ) | ( n20588 & n23387 ) ;
  assign n29133 = n29132 ^ n29130 ^ 1'b0 ;
  assign n29134 = n29133 ^ n14979 ^ n10532 ;
  assign n29135 = n27714 ^ n19255 ^ 1'b0 ;
  assign n29136 = n9011 ^ n645 ^ 1'b0 ;
  assign n29139 = n26512 ^ n16633 ^ n4867 ;
  assign n29140 = n29139 ^ n4848 ^ 1'b0 ;
  assign n29137 = ( n1453 & n5051 ) | ( n1453 & ~n14931 ) | ( n5051 & ~n14931 ) ;
  assign n29138 = n29137 ^ n13183 ^ 1'b0 ;
  assign n29141 = n29140 ^ n29138 ^ n12048 ;
  assign n29142 = n29141 ^ n10270 ^ n491 ;
  assign n29143 = ( n14047 & n29136 ) | ( n14047 & ~n29142 ) | ( n29136 & ~n29142 ) ;
  assign n29144 = n5600 | n29143 ;
  assign n29145 = n16669 & ~n29144 ;
  assign n29146 = ( ~n4000 & n29135 ) | ( ~n4000 & n29145 ) | ( n29135 & n29145 ) ;
  assign n29147 = ( n7521 & ~n18962 ) | ( n7521 & n25055 ) | ( ~n18962 & n25055 ) ;
  assign n29148 = n12043 ^ n565 ^ 1'b0 ;
  assign n29149 = n13357 & ~n29148 ;
  assign n29150 = n16252 ^ n1822 ^ 1'b0 ;
  assign n29151 = n2549 & n29150 ;
  assign n29152 = ~n8758 & n29151 ;
  assign n29153 = ~n26743 & n29152 ;
  assign n29155 = ~n8242 & n21976 ;
  assign n29154 = n2670 & ~n22273 ;
  assign n29156 = n29155 ^ n29154 ^ 1'b0 ;
  assign n29157 = n12189 ^ n5696 ^ n4517 ;
  assign n29158 = ( n304 & n16181 ) | ( n304 & n29157 ) | ( n16181 & n29157 ) ;
  assign n29161 = n26817 ^ n19842 ^ 1'b0 ;
  assign n29162 = n8208 & ~n29161 ;
  assign n29159 = ( n3050 & n4860 ) | ( n3050 & n5010 ) | ( n4860 & n5010 ) ;
  assign n29160 = ( n2608 & n9911 ) | ( n2608 & n29159 ) | ( n9911 & n29159 ) ;
  assign n29163 = n29162 ^ n29160 ^ n14123 ;
  assign n29164 = ( n4834 & n14425 ) | ( n4834 & n29163 ) | ( n14425 & n29163 ) ;
  assign n29165 = n13030 & n19670 ;
  assign n29166 = n29165 ^ n19886 ^ 1'b0 ;
  assign n29167 = n18029 ^ n17133 ^ 1'b0 ;
  assign n29168 = n3182 & n6875 ;
  assign n29169 = ~n6926 & n29168 ;
  assign n29170 = n21552 ^ n8000 ^ n7359 ;
  assign n29171 = ( n22344 & n29169 ) | ( n22344 & ~n29170 ) | ( n29169 & ~n29170 ) ;
  assign n29172 = n29171 ^ n20365 ^ n8728 ;
  assign n29173 = n25699 ^ n6657 ^ n573 ;
  assign n29176 = n5727 ^ n5667 ^ 1'b0 ;
  assign n29174 = n3927 & n14960 ;
  assign n29175 = ~n1006 & n29174 ;
  assign n29177 = n29176 ^ n29175 ^ n21406 ;
  assign n29179 = n11553 ^ n4588 ^ 1'b0 ;
  assign n29178 = n17500 ^ n16208 ^ n9206 ;
  assign n29180 = n29179 ^ n29178 ^ n7388 ;
  assign n29181 = n10308 ^ n3450 ^ n2670 ;
  assign n29183 = n27599 ^ n1360 ^ n321 ;
  assign n29182 = n6273 ^ n5580 ^ 1'b0 ;
  assign n29184 = n29183 ^ n29182 ^ n22809 ;
  assign n29185 = n1724 | n29184 ;
  assign n29186 = n29185 ^ n5727 ^ 1'b0 ;
  assign n29187 = n9610 ^ n1111 ^ x134 ;
  assign n29188 = n2009 | n29187 ;
  assign n29189 = n29186 & ~n29188 ;
  assign n29190 = ( ~n16999 & n19965 ) | ( ~n16999 & n29189 ) | ( n19965 & n29189 ) ;
  assign n29191 = n11000 & ~n15402 ;
  assign n29192 = n29191 ^ n1548 ^ 1'b0 ;
  assign n29193 = n29192 ^ n18184 ^ n8356 ;
  assign n29194 = n29193 ^ n16193 ^ n6644 ;
  assign n29195 = n3496 & ~n14112 ;
  assign n29196 = n22259 & n29195 ;
  assign n29197 = n29196 ^ n24337 ^ n12539 ;
  assign n29198 = n4571 & ~n15030 ;
  assign n29199 = n633 | n1345 ;
  assign n29200 = n2110 | n29199 ;
  assign n29201 = ( n909 & n4128 ) | ( n909 & ~n29200 ) | ( n4128 & ~n29200 ) ;
  assign n29202 = n11304 ^ n3049 ^ 1'b0 ;
  assign n29203 = n29201 | n29202 ;
  assign n29204 = n16638 ^ n1952 ^ 1'b0 ;
  assign n29205 = n29203 & n29204 ;
  assign n29206 = ( n11024 & n19436 ) | ( n11024 & ~n29205 ) | ( n19436 & ~n29205 ) ;
  assign n29207 = n29206 ^ n24348 ^ 1'b0 ;
  assign n29211 = n4359 ^ n1822 ^ 1'b0 ;
  assign n29212 = n5622 & ~n29211 ;
  assign n29209 = ( n7276 & n10322 ) | ( n7276 & ~n15317 ) | ( n10322 & ~n15317 ) ;
  assign n29210 = n29209 ^ n22230 ^ n9634 ;
  assign n29208 = x213 & ~n11855 ;
  assign n29213 = n29212 ^ n29210 ^ n29208 ;
  assign n29215 = n3340 & ~n8954 ;
  assign n29214 = n21394 ^ n21265 ^ 1'b0 ;
  assign n29216 = n29215 ^ n29214 ^ n12535 ;
  assign n29217 = n7056 & n21697 ;
  assign n29218 = n18533 & n29217 ;
  assign n29219 = n21506 ^ n15678 ^ n8638 ;
  assign n29220 = n7010 & ~n29219 ;
  assign n29221 = n19266 ^ n15955 ^ n4631 ;
  assign n29222 = n29221 ^ n24507 ^ n2907 ;
  assign n29223 = ( n2308 & ~n26947 ) | ( n2308 & n29222 ) | ( ~n26947 & n29222 ) ;
  assign n29224 = ~n4351 & n5941 ;
  assign n29225 = n29224 ^ n11299 ^ 1'b0 ;
  assign n29228 = n14602 ^ n14187 ^ 1'b0 ;
  assign n29226 = ( n991 & n8264 ) | ( n991 & ~n20534 ) | ( n8264 & ~n20534 ) ;
  assign n29227 = n29226 ^ n3846 ^ n1319 ;
  assign n29229 = n29228 ^ n29227 ^ n22756 ;
  assign n29230 = n29225 | n29229 ;
  assign n29231 = n29062 & ~n29230 ;
  assign n29232 = n13731 ^ n9831 ^ n7000 ;
  assign n29233 = n24627 ^ n14792 ^ n3497 ;
  assign n29234 = n13592 ^ n2989 ^ 1'b0 ;
  assign n29235 = n24307 ^ n5066 ^ 1'b0 ;
  assign n29236 = n29234 | n29235 ;
  assign n29237 = n12432 ^ n4151 ^ 1'b0 ;
  assign n29238 = n15291 & n29237 ;
  assign n29239 = n29200 ^ n2828 ^ 1'b0 ;
  assign n29240 = n3811 | n29239 ;
  assign n29241 = n29240 ^ n19326 ^ n1140 ;
  assign n29242 = ~n17863 & n29241 ;
  assign n29243 = ~n24857 & n29242 ;
  assign n29244 = ( ~n2489 & n5800 ) | ( ~n2489 & n12300 ) | ( n5800 & n12300 ) ;
  assign n29256 = ( n785 & ~n3143 ) | ( n785 & n9992 ) | ( ~n3143 & n9992 ) ;
  assign n29257 = ~n1405 & n24178 ;
  assign n29258 = n29257 ^ n11578 ^ 1'b0 ;
  assign n29259 = n29258 ^ n6892 ^ 1'b0 ;
  assign n29260 = n29256 | n29259 ;
  assign n29261 = ( n7861 & n14189 ) | ( n7861 & n29260 ) | ( n14189 & n29260 ) ;
  assign n29245 = n20180 ^ n1520 ^ n266 ;
  assign n29246 = ( ~n4337 & n12894 ) | ( ~n4337 & n29245 ) | ( n12894 & n29245 ) ;
  assign n29251 = n12043 ^ n2459 ^ 1'b0 ;
  assign n29250 = n8424 | n22997 ;
  assign n29252 = n29251 ^ n29250 ^ n2377 ;
  assign n29247 = ( n5248 & ~n7068 ) | ( n5248 & n12071 ) | ( ~n7068 & n12071 ) ;
  assign n29248 = ~n6843 & n15829 ;
  assign n29249 = n29247 & ~n29248 ;
  assign n29253 = n29252 ^ n29249 ^ 1'b0 ;
  assign n29254 = ( n2266 & ~n24987 ) | ( n2266 & n29253 ) | ( ~n24987 & n29253 ) ;
  assign n29255 = n29246 & n29254 ;
  assign n29262 = n29261 ^ n29255 ^ 1'b0 ;
  assign n29263 = n16661 & n29262 ;
  assign n29264 = ~n6901 & n7684 ;
  assign n29265 = n7385 & ~n18924 ;
  assign n29266 = n29265 ^ n13666 ^ 1'b0 ;
  assign n29267 = ( n19549 & n29264 ) | ( n19549 & n29266 ) | ( n29264 & n29266 ) ;
  assign n29268 = n16193 ^ n8692 ^ n7242 ;
  assign n29269 = n23464 & ~n29268 ;
  assign n29270 = n22841 & n29269 ;
  assign n29271 = n25755 ^ n19266 ^ n11016 ;
  assign n29272 = n29270 | n29271 ;
  assign n29273 = n29272 ^ n7486 ^ 1'b0 ;
  assign n29274 = n27199 ^ n20025 ^ 1'b0 ;
  assign n29275 = n4134 & n29274 ;
  assign n29276 = ( n25699 & ~n29273 ) | ( n25699 & n29275 ) | ( ~n29273 & n29275 ) ;
  assign n29277 = n16263 & ~n29276 ;
  assign n29281 = n1833 | n2775 ;
  assign n29278 = x189 & n12907 ;
  assign n29279 = ~n10832 & n29278 ;
  assign n29280 = n21494 | n29279 ;
  assign n29282 = n29281 ^ n29280 ^ 1'b0 ;
  assign n29283 = n4126 | n19693 ;
  assign n29284 = n29283 ^ n16297 ^ n4353 ;
  assign n29285 = ( n2480 & ~n6149 ) | ( n2480 & n12562 ) | ( ~n6149 & n12562 ) ;
  assign n29286 = n13865 & ~n29285 ;
  assign n29287 = n26613 ^ n15886 ^ 1'b0 ;
  assign n29288 = ( n2875 & n4697 ) | ( n2875 & ~n5246 ) | ( n4697 & ~n5246 ) ;
  assign n29289 = ( n1140 & n17563 ) | ( n1140 & n29288 ) | ( n17563 & n29288 ) ;
  assign n29290 = ( ~n2137 & n10334 ) | ( ~n2137 & n29289 ) | ( n10334 & n29289 ) ;
  assign n29291 = n6166 | n8020 ;
  assign n29292 = n29291 ^ n4291 ^ 1'b0 ;
  assign n29293 = ( ~n263 & n5417 ) | ( ~n263 & n9350 ) | ( n5417 & n9350 ) ;
  assign n29294 = n29293 ^ n21862 ^ 1'b0 ;
  assign n29295 = n20062 | n29294 ;
  assign n29296 = ( n11088 & n18277 ) | ( n11088 & ~n29295 ) | ( n18277 & ~n29295 ) ;
  assign n29305 = n12072 ^ n11709 ^ n11591 ;
  assign n29306 = n11831 | n29305 ;
  assign n29307 = n23363 & ~n29306 ;
  assign n29303 = n18021 & n26959 ;
  assign n29304 = ~n6575 & n29303 ;
  assign n29297 = ( n1870 & n6859 ) | ( n1870 & ~n28297 ) | ( n6859 & ~n28297 ) ;
  assign n29298 = n2984 ^ n2067 ^ n1084 ;
  assign n29299 = n29298 ^ n1599 ^ 1'b0 ;
  assign n29300 = n7152 | n27059 ;
  assign n29301 = n21360 | n29300 ;
  assign n29302 = ( n29297 & n29299 ) | ( n29297 & n29301 ) | ( n29299 & n29301 ) ;
  assign n29308 = n29307 ^ n29304 ^ n29302 ;
  assign n29309 = n682 & n28109 ;
  assign n29310 = ( n1515 & ~n10698 ) | ( n1515 & n16811 ) | ( ~n10698 & n16811 ) ;
  assign n29311 = n29310 ^ n8839 ^ n8670 ;
  assign n29312 = n19522 | n29311 ;
  assign n29313 = n27731 & ~n29312 ;
  assign n29314 = n15196 & ~n16883 ;
  assign n29315 = n29314 ^ n11819 ^ 1'b0 ;
  assign n29316 = n28457 ^ n21685 ^ n18492 ;
  assign n29317 = n29316 ^ n418 ^ 1'b0 ;
  assign n29318 = n29315 | n29317 ;
  assign n29319 = ~n2485 & n18357 ;
  assign n29320 = n28846 ^ n10389 ^ n9660 ;
  assign n29321 = x167 & n25163 ;
  assign n29322 = n1371 & n29321 ;
  assign n29323 = ( n15718 & ~n29320 ) | ( n15718 & n29322 ) | ( ~n29320 & n29322 ) ;
  assign n29324 = ( n17925 & n29319 ) | ( n17925 & ~n29323 ) | ( n29319 & ~n29323 ) ;
  assign n29325 = ( n5024 & ~n8080 ) | ( n5024 & n15961 ) | ( ~n8080 & n15961 ) ;
  assign n29326 = n3758 & ~n4619 ;
  assign n29327 = n17232 | n29326 ;
  assign n29328 = ( n23561 & n29325 ) | ( n23561 & n29327 ) | ( n29325 & n29327 ) ;
  assign n29329 = n19590 ^ n13725 ^ n3282 ;
  assign n29330 = ( n3522 & ~n3595 ) | ( n3522 & n29329 ) | ( ~n3595 & n29329 ) ;
  assign n29331 = n29330 ^ n5996 ^ n5090 ;
  assign n29332 = n3632 ^ n3504 ^ 1'b0 ;
  assign n29333 = n9104 | n29332 ;
  assign n29334 = n29333 ^ n11497 ^ n6119 ;
  assign n29335 = ~n20273 & n24524 ;
  assign n29336 = n28170 | n29335 ;
  assign n29337 = n16297 & ~n29336 ;
  assign n29338 = n3437 | n9162 ;
  assign n29339 = n10448 & ~n20391 ;
  assign n29344 = n17845 ^ n6732 ^ 1'b0 ;
  assign n29345 = x86 & n29344 ;
  assign n29340 = n17489 ^ n13535 ^ n1720 ;
  assign n29341 = ~n4803 & n7983 ;
  assign n29342 = n29340 & n29341 ;
  assign n29343 = n29342 ^ n11412 ^ 1'b0 ;
  assign n29346 = n29345 ^ n29343 ^ n4965 ;
  assign n29347 = n27089 ^ n9254 ^ n3410 ;
  assign n29349 = n9744 ^ n8374 ^ n1791 ;
  assign n29348 = n10530 ^ n6170 ^ n4176 ;
  assign n29350 = n29349 ^ n29348 ^ 1'b0 ;
  assign n29351 = n29347 & ~n29350 ;
  assign n29352 = n7224 & ~n22791 ;
  assign n29353 = n29352 ^ n755 ^ 1'b0 ;
  assign n29354 = n10371 ^ n6745 ^ n326 ;
  assign n29355 = n29354 ^ n1936 ^ 1'b0 ;
  assign n29358 = n6581 & ~n12122 ;
  assign n29359 = n7556 & n29358 ;
  assign n29356 = n15222 ^ n12323 ^ x62 ;
  assign n29357 = ~n27631 & n29356 ;
  assign n29360 = n29359 ^ n29357 ^ 1'b0 ;
  assign n29361 = ~n29355 & n29360 ;
  assign n29362 = ( n4856 & n21264 ) | ( n4856 & ~n23822 ) | ( n21264 & ~n23822 ) ;
  assign n29363 = n29362 ^ n16335 ^ n4921 ;
  assign n29364 = n3525 & n5693 ;
  assign n29365 = n14589 ^ n7574 ^ n1482 ;
  assign n29366 = ( n26933 & n29196 ) | ( n26933 & n29365 ) | ( n29196 & n29365 ) ;
  assign n29367 = ( n19256 & ~n29364 ) | ( n19256 & n29366 ) | ( ~n29364 & n29366 ) ;
  assign n29368 = n14465 ^ n4109 ^ 1'b0 ;
  assign n29369 = n29368 ^ n22680 ^ 1'b0 ;
  assign n29370 = ~n20656 & n29369 ;
  assign n29385 = ( n906 & n2137 ) | ( n906 & n5679 ) | ( n2137 & n5679 ) ;
  assign n29386 = ~n9343 & n18431 ;
  assign n29387 = ~n29385 & n29386 ;
  assign n29388 = n6118 & ~n29387 ;
  assign n29389 = n29388 ^ n23486 ^ 1'b0 ;
  assign n29390 = n29389 ^ n4168 ^ 1'b0 ;
  assign n29381 = n27676 ^ n25026 ^ n1663 ;
  assign n29375 = n9311 ^ n5484 ^ n4038 ;
  assign n29378 = ( n10022 & ~n14759 ) | ( n10022 & n20800 ) | ( ~n14759 & n20800 ) ;
  assign n29376 = x142 & ~n19002 ;
  assign n29377 = n29376 ^ n16988 ^ n2981 ;
  assign n29379 = n29378 ^ n29377 ^ 1'b0 ;
  assign n29380 = n29375 & n29379 ;
  assign n29372 = n27634 ^ n11766 ^ n961 ;
  assign n29373 = n29372 ^ n22869 ^ n7290 ;
  assign n29371 = n2949 | n16961 ;
  assign n29374 = n29373 ^ n29371 ^ 1'b0 ;
  assign n29382 = n29381 ^ n29380 ^ n29374 ;
  assign n29383 = ( ~n6190 & n27269 ) | ( ~n6190 & n29382 ) | ( n27269 & n29382 ) ;
  assign n29384 = n6663 & n29383 ;
  assign n29391 = n29390 ^ n29384 ^ 1'b0 ;
  assign n29392 = ~n1826 & n13693 ;
  assign n29393 = n21217 ^ n18922 ^ n9426 ;
  assign n29394 = n12690 & n26160 ;
  assign n29395 = ( n14206 & n23123 ) | ( n14206 & ~n29394 ) | ( n23123 & ~n29394 ) ;
  assign n29396 = n19133 | n29395 ;
  assign n29397 = n29396 ^ n26171 ^ 1'b0 ;
  assign n29398 = ( ~n10807 & n29393 ) | ( ~n10807 & n29397 ) | ( n29393 & n29397 ) ;
  assign n29399 = n29398 ^ n17120 ^ n8626 ;
  assign n29400 = n19472 ^ n6452 ^ 1'b0 ;
  assign n29401 = n20065 | n29400 ;
  assign n29402 = n5130 | n29401 ;
  assign n29403 = ( n2824 & n10953 ) | ( n2824 & n16522 ) | ( n10953 & n16522 ) ;
  assign n29404 = n5267 & ~n29403 ;
  assign n29407 = n14212 ^ n5821 ^ 1'b0 ;
  assign n29408 = n29407 ^ n25173 ^ n475 ;
  assign n29409 = n29408 ^ n20241 ^ n2678 ;
  assign n29405 = ( n9185 & ~n21200 ) | ( n9185 & n22530 ) | ( ~n21200 & n22530 ) ;
  assign n29406 = ~n23281 & n29405 ;
  assign n29410 = n29409 ^ n29406 ^ 1'b0 ;
  assign n29413 = ( n1475 & n6682 ) | ( n1475 & n6792 ) | ( n6682 & n6792 ) ;
  assign n29411 = ( n358 & n9314 ) | ( n358 & n12842 ) | ( n9314 & n12842 ) ;
  assign n29412 = n29411 ^ n4554 ^ n710 ;
  assign n29414 = n29413 ^ n29412 ^ 1'b0 ;
  assign n29415 = n27706 ^ n22005 ^ n4196 ;
  assign n29416 = ~n6692 & n19358 ;
  assign n29417 = ~n28264 & n29416 ;
  assign n29418 = n29417 ^ n16390 ^ n10813 ;
  assign n29419 = ( n1836 & ~n17078 ) | ( n1836 & n29418 ) | ( ~n17078 & n29418 ) ;
  assign n29420 = n17657 ^ n11031 ^ n5638 ;
  assign n29422 = ( n2979 & n4765 ) | ( n2979 & n11354 ) | ( n4765 & n11354 ) ;
  assign n29421 = n22101 | n24155 ;
  assign n29423 = n29422 ^ n29421 ^ 1'b0 ;
  assign n29431 = ( n12703 & n15962 ) | ( n12703 & ~n18156 ) | ( n15962 & ~n18156 ) ;
  assign n29424 = n4591 ^ n3303 ^ n1034 ;
  assign n29425 = n23395 ^ n8966 ^ 1'b0 ;
  assign n29426 = ~n3691 & n29425 ;
  assign n29427 = ( n22243 & n29424 ) | ( n22243 & ~n29426 ) | ( n29424 & ~n29426 ) ;
  assign n29428 = ( ~n9641 & n23828 ) | ( ~n9641 & n29427 ) | ( n23828 & n29427 ) ;
  assign n29429 = n25301 ^ n8339 ^ 1'b0 ;
  assign n29430 = n29428 | n29429 ;
  assign n29432 = n29431 ^ n29430 ^ 1'b0 ;
  assign n29433 = n20566 ^ n17520 ^ 1'b0 ;
  assign n29434 = n8621 | n11262 ;
  assign n29435 = n9228 | n29434 ;
  assign n29436 = n29435 ^ n23768 ^ n18273 ;
  assign n29437 = n29436 ^ n3841 ^ 1'b0 ;
  assign n29438 = ( n13043 & ~n17778 ) | ( n13043 & n21675 ) | ( ~n17778 & n21675 ) ;
  assign n29439 = n29438 ^ n18243 ^ 1'b0 ;
  assign n29440 = ~n29437 & n29439 ;
  assign n29441 = ( n7905 & n29433 ) | ( n7905 & ~n29440 ) | ( n29433 & ~n29440 ) ;
  assign n29442 = n22399 ^ n6417 ^ n4856 ;
  assign n29443 = n20058 ^ n6190 ^ 1'b0 ;
  assign n29444 = n6766 & ~n29443 ;
  assign n29445 = n29444 ^ n24685 ^ 1'b0 ;
  assign n29446 = ( n14078 & ~n18124 ) | ( n14078 & n18972 ) | ( ~n18124 & n18972 ) ;
  assign n29447 = n13345 ^ n3454 ^ 1'b0 ;
  assign n29448 = n29446 & ~n29447 ;
  assign n29450 = n18061 ^ n3103 ^ 1'b0 ;
  assign n29451 = n3007 & n29450 ;
  assign n29449 = ( ~n1527 & n9471 ) | ( ~n1527 & n9783 ) | ( n9471 & n9783 ) ;
  assign n29452 = n29451 ^ n29449 ^ 1'b0 ;
  assign n29453 = ( n9023 & n22506 ) | ( n9023 & ~n29452 ) | ( n22506 & ~n29452 ) ;
  assign n29454 = ~n3018 & n17150 ;
  assign n29455 = n13922 ^ n5570 ^ 1'b0 ;
  assign n29456 = n14252 | n29455 ;
  assign n29457 = ( n10835 & n16951 ) | ( n10835 & n29456 ) | ( n16951 & n29456 ) ;
  assign n29458 = ( n9346 & ~n22752 ) | ( n9346 & n29457 ) | ( ~n22752 & n29457 ) ;
  assign n29459 = n5637 | n9501 ;
  assign n29460 = n1456 & ~n29459 ;
  assign n29461 = n29460 ^ n26871 ^ n14782 ;
  assign n29462 = ( n4782 & n10722 ) | ( n4782 & ~n15386 ) | ( n10722 & ~n15386 ) ;
  assign n29463 = ~n591 & n9751 ;
  assign n29464 = n22523 ^ n3721 ^ 1'b0 ;
  assign n29465 = ~n19858 & n29464 ;
  assign n29466 = n12784 ^ n12640 ^ 1'b0 ;
  assign n29467 = n11076 & n29466 ;
  assign n29468 = n29040 ^ n21506 ^ n13205 ;
  assign n29469 = ~n25925 & n29468 ;
  assign n29470 = n11979 ^ n9891 ^ 1'b0 ;
  assign n29471 = ~n15509 & n29470 ;
  assign n29474 = n9601 & n22677 ;
  assign n29472 = n11479 ^ n6564 ^ 1'b0 ;
  assign n29473 = n29472 ^ n16360 ^ n12304 ;
  assign n29475 = n29474 ^ n29473 ^ 1'b0 ;
  assign n29476 = n25287 ^ n17635 ^ n3771 ;
  assign n29477 = n29476 ^ n15271 ^ n9583 ;
  assign n29478 = n15100 & ~n16064 ;
  assign n29479 = ~n5319 & n29478 ;
  assign n29480 = n29479 ^ n23465 ^ 1'b0 ;
  assign n29481 = ( ~n10939 & n12985 ) | ( ~n10939 & n29480 ) | ( n12985 & n29480 ) ;
  assign n29482 = n10344 ^ n7022 ^ n542 ;
  assign n29483 = n29482 ^ n25552 ^ 1'b0 ;
  assign n29484 = n29481 & n29483 ;
  assign n29485 = ~n10395 & n15276 ;
  assign n29486 = n26404 ^ n8860 ^ 1'b0 ;
  assign n29487 = n29486 ^ n18135 ^ n13772 ;
  assign n29488 = n4462 | n29487 ;
  assign n29489 = n18971 ^ n4808 ^ 1'b0 ;
  assign n29493 = n1821 & n4902 ;
  assign n29494 = ( n3372 & n9666 ) | ( n3372 & n29493 ) | ( n9666 & n29493 ) ;
  assign n29490 = n14048 ^ n3816 ^ 1'b0 ;
  assign n29491 = n4000 & n29490 ;
  assign n29492 = n29491 ^ n18316 ^ n4171 ;
  assign n29495 = n29494 ^ n29492 ^ n16381 ;
  assign n29498 = ( n6479 & n7452 ) | ( n6479 & n7653 ) | ( n7452 & n7653 ) ;
  assign n29499 = ( n24025 & n24546 ) | ( n24025 & ~n29498 ) | ( n24546 & ~n29498 ) ;
  assign n29496 = ~n1683 & n7309 ;
  assign n29497 = n29496 ^ n24586 ^ 1'b0 ;
  assign n29500 = n29499 ^ n29497 ^ n8039 ;
  assign n29501 = n29500 ^ n17172 ^ 1'b0 ;
  assign n29502 = n4670 & n26020 ;
  assign n29503 = n11695 & n29502 ;
  assign n29504 = n23289 ^ n6938 ^ n4438 ;
  assign n29505 = n1114 & n29504 ;
  assign n29506 = ( n4678 & n29503 ) | ( n4678 & n29505 ) | ( n29503 & n29505 ) ;
  assign n29507 = n29506 ^ n24175 ^ n866 ;
  assign n29511 = n12719 ^ n3682 ^ n1433 ;
  assign n29512 = ( n6170 & n12195 ) | ( n6170 & ~n29511 ) | ( n12195 & ~n29511 ) ;
  assign n29513 = ( n22465 & n26473 ) | ( n22465 & ~n29512 ) | ( n26473 & ~n29512 ) ;
  assign n29508 = ( ~x156 & n11780 ) | ( ~x156 & n12285 ) | ( n11780 & n12285 ) ;
  assign n29509 = ( n15816 & ~n16255 ) | ( n15816 & n29508 ) | ( ~n16255 & n29508 ) ;
  assign n29510 = n29509 ^ n7819 ^ n7189 ;
  assign n29514 = n29513 ^ n29510 ^ n23904 ;
  assign n29515 = ( ~n1725 & n4749 ) | ( ~n1725 & n17302 ) | ( n4749 & n17302 ) ;
  assign n29516 = n9157 & n11414 ;
  assign n29518 = n10082 ^ n9199 ^ n5371 ;
  assign n29517 = ~n14653 & n23469 ;
  assign n29519 = n29518 ^ n29517 ^ 1'b0 ;
  assign n29520 = ( n4889 & n15876 ) | ( n4889 & n29519 ) | ( n15876 & n29519 ) ;
  assign n29521 = n21731 ^ n13502 ^ n282 ;
  assign n29522 = n5246 & n23810 ;
  assign n29523 = n4725 & ~n13528 ;
  assign n29524 = n29523 ^ n25744 ^ 1'b0 ;
  assign n29525 = n26482 ^ n5415 ^ 1'b0 ;
  assign n29526 = ~n6724 & n29525 ;
  assign n29527 = ( n5852 & ~n27242 ) | ( n5852 & n29526 ) | ( ~n27242 & n29526 ) ;
  assign n29528 = n19216 ^ n6605 ^ 1'b0 ;
  assign n29529 = ~n13618 & n29528 ;
  assign n29530 = ( ~n7332 & n16368 ) | ( ~n7332 & n29529 ) | ( n16368 & n29529 ) ;
  assign n29531 = n29530 ^ n8339 ^ n2129 ;
  assign n29532 = n10719 | n29531 ;
  assign n29533 = n9873 ^ n6211 ^ 1'b0 ;
  assign n29534 = ( n13016 & n22557 ) | ( n13016 & n29533 ) | ( n22557 & n29533 ) ;
  assign n29535 = n8749 | n9927 ;
  assign n29536 = n18689 ^ n12280 ^ n582 ;
  assign n29537 = n29536 ^ n14934 ^ n7310 ;
  assign n29538 = n5926 ^ n4702 ^ 1'b0 ;
  assign n29539 = n9571 & n29538 ;
  assign n29540 = n29539 ^ n2714 ^ 1'b0 ;
  assign n29541 = n29537 & n29540 ;
  assign n29542 = n29541 ^ n2046 ^ 1'b0 ;
  assign n29543 = n29535 & n29542 ;
  assign n29544 = n26518 ^ n1634 ^ 1'b0 ;
  assign n29545 = n26122 & ~n29544 ;
  assign n29547 = n5950 & n28424 ;
  assign n29548 = n29547 ^ n16666 ^ 1'b0 ;
  assign n29546 = n18477 ^ n8092 ^ 1'b0 ;
  assign n29549 = n29548 ^ n29546 ^ n27165 ;
  assign n29550 = ( x34 & n15284 ) | ( x34 & ~n27434 ) | ( n15284 & ~n27434 ) ;
  assign n29551 = n29550 ^ n21130 ^ 1'b0 ;
  assign n29552 = n14373 ^ n7447 ^ 1'b0 ;
  assign n29553 = n17231 & ~n29552 ;
  assign n29554 = n29553 ^ n1719 ^ 1'b0 ;
  assign n29555 = ( ~n7142 & n29078 ) | ( ~n7142 & n29554 ) | ( n29078 & n29554 ) ;
  assign n29556 = n23449 ^ n14235 ^ n1651 ;
  assign n29557 = n29556 ^ n6959 ^ 1'b0 ;
  assign n29558 = n5076 ^ x83 ^ 1'b0 ;
  assign n29559 = ( n14016 & n14345 ) | ( n14016 & ~n16976 ) | ( n14345 & ~n16976 ) ;
  assign n29560 = n15134 ^ n4758 ^ n495 ;
  assign n29561 = n29560 ^ n21070 ^ 1'b0 ;
  assign n29562 = n29559 & ~n29561 ;
  assign n29563 = n16249 ^ n8673 ^ n5190 ;
  assign n29564 = n29563 ^ n27962 ^ n7314 ;
  assign n29565 = x33 | n29564 ;
  assign n29566 = n29565 ^ n12134 ^ 1'b0 ;
  assign n29567 = ( n1960 & ~n7768 ) | ( n1960 & n28652 ) | ( ~n7768 & n28652 ) ;
  assign n29568 = ( ~n762 & n16470 ) | ( ~n762 & n29567 ) | ( n16470 & n29567 ) ;
  assign n29569 = n26273 ^ n4115 ^ n1005 ;
  assign n29570 = n29569 ^ n24493 ^ n5574 ;
  assign n29571 = n19226 ^ n10366 ^ n909 ;
  assign n29572 = ( n7814 & n14148 ) | ( n7814 & n21835 ) | ( n14148 & n21835 ) ;
  assign n29573 = ( n15368 & n21160 ) | ( n15368 & n29572 ) | ( n21160 & n29572 ) ;
  assign n29574 = ( ~n21085 & n29571 ) | ( ~n21085 & n29573 ) | ( n29571 & n29573 ) ;
  assign n29575 = n29574 ^ n20511 ^ n3761 ;
  assign n29576 = n1897 & n29575 ;
  assign n29577 = n29576 ^ n1998 ^ 1'b0 ;
  assign n29578 = ~n462 & n14048 ;
  assign n29579 = n956 & n29578 ;
  assign n29580 = n8290 ^ n7029 ^ n6270 ;
  assign n29581 = n29580 ^ n13908 ^ n10957 ;
  assign n29584 = n11927 ^ n11216 ^ n344 ;
  assign n29582 = n1682 & n14286 ;
  assign n29583 = n29582 ^ n12790 ^ 1'b0 ;
  assign n29585 = n29584 ^ n29583 ^ n7968 ;
  assign n29586 = ( n27685 & ~n29581 ) | ( n27685 & n29585 ) | ( ~n29581 & n29585 ) ;
  assign n29587 = x163 & ~n6632 ;
  assign n29588 = ~n29586 & n29587 ;
  assign n29589 = ~n11563 & n29588 ;
  assign n29590 = ( ~n10101 & n15104 ) | ( ~n10101 & n28544 ) | ( n15104 & n28544 ) ;
  assign n29591 = n6875 & n23708 ;
  assign n29592 = n21550 & n29591 ;
  assign n29595 = n10072 ^ n4036 ^ n1242 ;
  assign n29596 = ( n12863 & n20428 ) | ( n12863 & ~n29595 ) | ( n20428 & ~n29595 ) ;
  assign n29597 = n9136 & ~n21750 ;
  assign n29598 = n29596 & n29597 ;
  assign n29593 = ~n10495 & n14377 ;
  assign n29594 = n10976 | n29593 ;
  assign n29599 = n29598 ^ n29594 ^ 1'b0 ;
  assign n29600 = n23944 ^ n14742 ^ n334 ;
  assign n29601 = n22257 ^ n1121 ^ 1'b0 ;
  assign n29602 = n23447 | n29601 ;
  assign n29603 = n29602 ^ n9999 ^ 1'b0 ;
  assign n29607 = n2266 | n16692 ;
  assign n29608 = n7709 & ~n29607 ;
  assign n29604 = ~n5714 & n13703 ;
  assign n29605 = n19901 ^ n14282 ^ n5582 ;
  assign n29606 = ( n17775 & n29604 ) | ( n17775 & n29605 ) | ( n29604 & n29605 ) ;
  assign n29609 = n29608 ^ n29606 ^ 1'b0 ;
  assign n29610 = n17846 ^ n3343 ^ 1'b0 ;
  assign n29611 = ( n3638 & n12360 ) | ( n3638 & ~n28693 ) | ( n12360 & ~n28693 ) ;
  assign n29612 = n10112 ^ n1202 ^ n1156 ;
  assign n29613 = n20314 ^ n17317 ^ n7390 ;
  assign n29614 = n15252 ^ n13961 ^ 1'b0 ;
  assign n29615 = ~n21842 & n29614 ;
  assign n29616 = ~n10755 & n16161 ;
  assign n29617 = ~n29615 & n29616 ;
  assign n29618 = n13137 & ~n29617 ;
  assign n29619 = ~n29613 & n29618 ;
  assign n29620 = ( n25198 & n29612 ) | ( n25198 & n29619 ) | ( n29612 & n29619 ) ;
  assign n29621 = n27988 ^ n21087 ^ x113 ;
  assign n29622 = n29621 ^ n19184 ^ 1'b0 ;
  assign n29623 = n5991 ^ n5953 ^ 1'b0 ;
  assign n29624 = n678 & ~n29623 ;
  assign n29625 = ( n14284 & n22635 ) | ( n14284 & ~n23308 ) | ( n22635 & ~n23308 ) ;
  assign n29626 = ~n29624 & n29625 ;
  assign n29633 = n15660 ^ n7900 ^ n2296 ;
  assign n29627 = ~n11599 & n22461 ;
  assign n29628 = n29627 ^ n10253 ^ 1'b0 ;
  assign n29629 = n17386 ^ x202 ^ 1'b0 ;
  assign n29630 = n535 & ~n29629 ;
  assign n29631 = n29630 ^ n15278 ^ 1'b0 ;
  assign n29632 = n29628 | n29631 ;
  assign n29634 = n29633 ^ n29632 ^ 1'b0 ;
  assign n29638 = ( n4697 & n6292 ) | ( n4697 & ~n14109 ) | ( n6292 & ~n14109 ) ;
  assign n29636 = n3680 | n19630 ;
  assign n29635 = n18273 ^ n5360 ^ n4581 ;
  assign n29637 = n29636 ^ n29635 ^ 1'b0 ;
  assign n29639 = n29638 ^ n29637 ^ n27849 ;
  assign n29640 = n29634 & n29639 ;
  assign n29641 = n29640 ^ n21780 ^ 1'b0 ;
  assign n29642 = n1619 | n5655 ;
  assign n29643 = ~n8030 & n10777 ;
  assign n29644 = n29643 ^ n16400 ^ 1'b0 ;
  assign n29645 = ( n5878 & n14278 ) | ( n5878 & ~n29644 ) | ( n14278 & ~n29644 ) ;
  assign n29646 = ~n25290 & n29645 ;
  assign n29647 = n29646 ^ n17713 ^ 1'b0 ;
  assign n29648 = ( n1161 & n10824 ) | ( n1161 & ~n14897 ) | ( n10824 & ~n14897 ) ;
  assign n29649 = n19038 ^ n12638 ^ n6263 ;
  assign n29650 = ~n12063 & n29649 ;
  assign n29651 = ( ~n2704 & n14733 ) | ( ~n2704 & n23904 ) | ( n14733 & n23904 ) ;
  assign n29652 = n29651 ^ n27224 ^ 1'b0 ;
  assign n29653 = n14862 ^ n9771 ^ 1'b0 ;
  assign n29654 = ~n20420 & n29653 ;
  assign n29655 = ~n4093 & n8779 ;
  assign n29656 = n28324 ^ n19671 ^ n14235 ;
  assign n29657 = n29656 ^ n14420 ^ 1'b0 ;
  assign n29658 = n9869 ^ n6774 ^ 1'b0 ;
  assign n29659 = n9855 & ~n29658 ;
  assign n29660 = n29659 ^ n5435 ^ 1'b0 ;
  assign n29661 = n5643 & n13298 ;
  assign n29662 = n8237 & n29661 ;
  assign n29663 = ( ~n14909 & n22410 ) | ( ~n14909 & n29662 ) | ( n22410 & n29662 ) ;
  assign n29664 = ( ~n17154 & n23466 ) | ( ~n17154 & n29663 ) | ( n23466 & n29663 ) ;
  assign n29665 = n29664 ^ n17915 ^ n8828 ;
  assign n29666 = n10344 ^ n3310 ^ 1'b0 ;
  assign n29669 = n2641 | n5456 ;
  assign n29667 = n17982 ^ n9921 ^ 1'b0 ;
  assign n29668 = n15364 & n29667 ;
  assign n29670 = n29669 ^ n29668 ^ 1'b0 ;
  assign n29671 = n18784 ^ n2020 ^ 1'b0 ;
  assign n29672 = ~n9742 & n26139 ;
  assign n29673 = n10115 & n29672 ;
  assign n29674 = n21249 & n28311 ;
  assign n29675 = n29674 ^ n27431 ^ n10778 ;
  assign n29676 = n10111 | n12498 ;
  assign n29677 = ( x195 & n7277 ) | ( x195 & ~n29676 ) | ( n7277 & ~n29676 ) ;
  assign n29678 = n29677 ^ n6636 ^ n4856 ;
  assign n29686 = n15844 ^ n882 ^ 1'b0 ;
  assign n29687 = n16894 | n29686 ;
  assign n29679 = n9930 & ~n10711 ;
  assign n29680 = n29679 ^ n778 ^ 1'b0 ;
  assign n29681 = n29680 ^ n22265 ^ 1'b0 ;
  assign n29682 = n7417 ^ n6999 ^ n2514 ;
  assign n29683 = n29682 ^ n18783 ^ n16965 ;
  assign n29684 = n29681 & n29683 ;
  assign n29685 = n3249 & n29684 ;
  assign n29688 = n29687 ^ n29685 ^ n2621 ;
  assign n29689 = ( n647 & n26348 ) | ( n647 & ~n29688 ) | ( n26348 & ~n29688 ) ;
  assign n29690 = n2400 & n7256 ;
  assign n29691 = n8235 & n29690 ;
  assign n29692 = n29691 ^ n7690 ^ 1'b0 ;
  assign n29693 = n29692 ^ n24057 ^ n16711 ;
  assign n29697 = ( n1904 & ~n5945 ) | ( n1904 & n8054 ) | ( ~n5945 & n8054 ) ;
  assign n29698 = n29697 ^ n7991 ^ 1'b0 ;
  assign n29694 = ( n3311 & ~n5587 ) | ( n3311 & n5890 ) | ( ~n5587 & n5890 ) ;
  assign n29695 = ( n8640 & n11080 ) | ( n8640 & ~n16960 ) | ( n11080 & ~n16960 ) ;
  assign n29696 = ( n17560 & n29694 ) | ( n17560 & n29695 ) | ( n29694 & n29695 ) ;
  assign n29699 = n29698 ^ n29696 ^ n28934 ;
  assign n29700 = n5901 & ~n29699 ;
  assign n29701 = ~n13876 & n21209 ;
  assign n29702 = n29701 ^ n17075 ^ 1'b0 ;
  assign n29703 = n18645 ^ n8983 ^ 1'b0 ;
  assign n29704 = n19477 ^ n16422 ^ n10377 ;
  assign n29705 = n29704 ^ n20318 ^ n11081 ;
  assign n29708 = n13894 ^ n5208 ^ 1'b0 ;
  assign n29706 = n2540 & ~n12471 ;
  assign n29707 = ~n12666 & n29706 ;
  assign n29709 = n29708 ^ n29707 ^ n15392 ;
  assign n29710 = n9136 ^ n2626 ^ 1'b0 ;
  assign n29711 = ~n29709 & n29710 ;
  assign n29712 = ~n9097 & n29711 ;
  assign n29713 = n6312 & n29712 ;
  assign n29714 = n29705 & ~n29713 ;
  assign n29715 = ~n29703 & n29714 ;
  assign n29716 = n4147 | n4335 ;
  assign n29717 = n29716 ^ n24139 ^ 1'b0 ;
  assign n29718 = n1818 & ~n3154 ;
  assign n29719 = n10100 & n29718 ;
  assign n29720 = n29719 ^ n21943 ^ n12385 ;
  assign n29721 = n18859 ^ n15833 ^ n7441 ;
  assign n29722 = ( n6123 & n23497 ) | ( n6123 & ~n29721 ) | ( n23497 & ~n29721 ) ;
  assign n29723 = n29722 ^ n23138 ^ n9261 ;
  assign n29724 = n29723 ^ n7216 ^ n3111 ;
  assign n29725 = n22202 ^ n19041 ^ n6424 ;
  assign n29726 = n15732 ^ n7809 ^ x152 ;
  assign n29727 = ~n9082 & n20164 ;
  assign n29728 = n29727 ^ n21990 ^ 1'b0 ;
  assign n29729 = n12392 & n29600 ;
  assign n29730 = n13189 & n17357 ;
  assign n29731 = ( n3879 & ~n20800 ) | ( n3879 & n29730 ) | ( ~n20800 & n29730 ) ;
  assign n29732 = n29731 ^ n13006 ^ n6309 ;
  assign n29733 = n9993 ^ n8911 ^ n8591 ;
  assign n29734 = ( ~n397 & n11466 ) | ( ~n397 & n12462 ) | ( n11466 & n12462 ) ;
  assign n29735 = ( ~n1100 & n29733 ) | ( ~n1100 & n29734 ) | ( n29733 & n29734 ) ;
  assign n29736 = n4910 & ~n25396 ;
  assign n29737 = n10507 & ~n29736 ;
  assign n29738 = n27044 & n29737 ;
  assign n29739 = n23863 ^ n21696 ^ n3323 ;
  assign n29740 = ( n573 & ~n9924 ) | ( n573 & n10700 ) | ( ~n9924 & n10700 ) ;
  assign n29741 = n17326 | n29740 ;
  assign n29742 = n24619 & ~n29741 ;
  assign n29743 = ~n6316 & n27428 ;
  assign n29744 = n15694 ^ n5675 ^ 1'b0 ;
  assign n29745 = ( n15992 & ~n17838 ) | ( n15992 & n29744 ) | ( ~n17838 & n29744 ) ;
  assign n29746 = n11645 & n17582 ;
  assign n29747 = n1200 & n29746 ;
  assign n29748 = n414 & n21483 ;
  assign n29749 = n29747 & n29748 ;
  assign n29750 = ( n1172 & ~n2590 ) | ( n1172 & n9900 ) | ( ~n2590 & n9900 ) ;
  assign n29751 = n5988 & ~n8538 ;
  assign n29752 = ~n29750 & n29751 ;
  assign n29753 = n29045 ^ n28101 ^ 1'b0 ;
  assign n29754 = n29752 | n29753 ;
  assign n29755 = n10156 ^ n9670 ^ 1'b0 ;
  assign n29756 = ( n5495 & ~n10999 ) | ( n5495 & n22507 ) | ( ~n10999 & n22507 ) ;
  assign n29757 = n29756 ^ n20145 ^ n6457 ;
  assign n29758 = ( n2164 & ~n2804 ) | ( n2164 & n29757 ) | ( ~n2804 & n29757 ) ;
  assign n29759 = n16200 ^ n7468 ^ 1'b0 ;
  assign n29760 = n24530 ^ n2525 ^ n1422 ;
  assign n29761 = n29760 ^ n15886 ^ 1'b0 ;
  assign n29762 = ~n29759 & n29761 ;
  assign n29763 = n4568 & ~n7107 ;
  assign n29764 = n29763 ^ n22760 ^ 1'b0 ;
  assign n29765 = ~n8087 & n11911 ;
  assign n29766 = n1202 | n13393 ;
  assign n29767 = n13738 & ~n26988 ;
  assign n29769 = x147 & n23374 ;
  assign n29770 = n29769 ^ n8087 ^ 1'b0 ;
  assign n29768 = n1460 & ~n10124 ;
  assign n29771 = n29770 ^ n29768 ^ 1'b0 ;
  assign n29772 = n3983 ^ x46 ^ 1'b0 ;
  assign n29773 = n29771 & n29772 ;
  assign n29774 = n20554 ^ n18313 ^ n2162 ;
  assign n29775 = n29773 & n29774 ;
  assign n29776 = n5774 | n8745 ;
  assign n29777 = n29776 ^ n833 ^ 1'b0 ;
  assign n29778 = n29777 ^ n19553 ^ n9721 ;
  assign n29779 = n29778 ^ n13765 ^ 1'b0 ;
  assign n29780 = n29775 & ~n29779 ;
  assign n29781 = n1697 & n3646 ;
  assign n29783 = n14446 ^ n11136 ^ n8474 ;
  assign n29782 = ~n768 & n24615 ;
  assign n29784 = n29783 ^ n29782 ^ 1'b0 ;
  assign n29785 = n6077 ^ n4209 ^ 1'b0 ;
  assign n29786 = n2014 | n29785 ;
  assign n29787 = n29786 ^ n658 ^ 1'b0 ;
  assign n29788 = ~n23839 & n29787 ;
  assign n29789 = ~n5676 & n24197 ;
  assign n29794 = n28161 ^ n7863 ^ 1'b0 ;
  assign n29795 = n8777 & ~n29794 ;
  assign n29796 = n29795 ^ n2877 ^ n545 ;
  assign n29791 = n15309 & ~n20542 ;
  assign n29790 = n14293 ^ n5135 ^ 1'b0 ;
  assign n29792 = n29791 ^ n29790 ^ n21168 ;
  assign n29793 = ( ~n13099 & n19198 ) | ( ~n13099 & n29792 ) | ( n19198 & n29792 ) ;
  assign n29797 = n29796 ^ n29793 ^ n25287 ;
  assign n29798 = ( ~n8982 & n29789 ) | ( ~n8982 & n29797 ) | ( n29789 & n29797 ) ;
  assign n29799 = n7985 | n15932 ;
  assign n29800 = ( n5262 & ~n18181 ) | ( n5262 & n18954 ) | ( ~n18181 & n18954 ) ;
  assign n29801 = ( n6199 & ~n6659 ) | ( n6199 & n14682 ) | ( ~n6659 & n14682 ) ;
  assign n29802 = n29801 ^ n12796 ^ n673 ;
  assign n29803 = ( ~n12975 & n20534 ) | ( ~n12975 & n29802 ) | ( n20534 & n29802 ) ;
  assign n29804 = ( ~n15888 & n29800 ) | ( ~n15888 & n29803 ) | ( n29800 & n29803 ) ;
  assign n29805 = ~n1241 & n3063 ;
  assign n29806 = n29805 ^ n21485 ^ 1'b0 ;
  assign n29807 = n2382 | n29806 ;
  assign n29808 = n29807 ^ n10164 ^ 1'b0 ;
  assign n29809 = n28037 ^ n2424 ^ 1'b0 ;
  assign n29810 = n27369 | n29809 ;
  assign n29811 = n29810 ^ n7870 ^ n352 ;
  assign n29812 = ( ~n13597 & n27063 ) | ( ~n13597 & n29811 ) | ( n27063 & n29811 ) ;
  assign n29813 = n23308 ^ n22755 ^ n8109 ;
  assign n29814 = ( n1763 & ~n2626 ) | ( n1763 & n26607 ) | ( ~n2626 & n26607 ) ;
  assign n29815 = n28731 & ~n29814 ;
  assign n29816 = n14838 & n29815 ;
  assign n29817 = n26142 ^ n12878 ^ n9336 ;
  assign n29818 = n17405 | n29817 ;
  assign n29819 = n15625 ^ n12066 ^ 1'b0 ;
  assign n29820 = ( ~n16831 & n27042 ) | ( ~n16831 & n29793 ) | ( n27042 & n29793 ) ;
  assign n29821 = n22971 ^ n5048 ^ 1'b0 ;
  assign n29822 = n29683 & ~n29821 ;
  assign n29823 = ( n8662 & n10150 ) | ( n8662 & ~n29822 ) | ( n10150 & ~n29822 ) ;
  assign n29826 = n11911 ^ n1209 ^ n498 ;
  assign n29827 = ( n2865 & n19290 ) | ( n2865 & n29826 ) | ( n19290 & n29826 ) ;
  assign n29824 = n14815 & n18222 ;
  assign n29825 = ~n17606 & n29824 ;
  assign n29828 = n29827 ^ n29825 ^ n9839 ;
  assign n29829 = n1068 & ~n12806 ;
  assign n29830 = n5713 & n29829 ;
  assign n29831 = n29830 ^ n7830 ^ 1'b0 ;
  assign n29832 = ( n20829 & n29500 ) | ( n20829 & n29831 ) | ( n29500 & n29831 ) ;
  assign n29833 = ( n8675 & n20661 ) | ( n8675 & n28383 ) | ( n20661 & n28383 ) ;
  assign n29834 = n29628 ^ n9555 ^ n4908 ;
  assign n29836 = n19856 ^ n19509 ^ n6707 ;
  assign n29835 = n2143 | n15795 ;
  assign n29837 = n29836 ^ n29835 ^ n12386 ;
  assign n29838 = n25408 ^ n23686 ^ n903 ;
  assign n29839 = ( n1761 & ~n2738 ) | ( n1761 & n11751 ) | ( ~n2738 & n11751 ) ;
  assign n29840 = ( ~n5394 & n11772 ) | ( ~n5394 & n29839 ) | ( n11772 & n29839 ) ;
  assign n29841 = n4747 & n21562 ;
  assign n29842 = n19221 ^ n5466 ^ n4633 ;
  assign n29843 = ( n13261 & n28534 ) | ( n13261 & n29842 ) | ( n28534 & n29842 ) ;
  assign n29844 = n19472 ^ n10045 ^ n2961 ;
  assign n29845 = n27673 ^ n26067 ^ n3517 ;
  assign n29846 = ( x144 & ~n4373 ) | ( x144 & n15051 ) | ( ~n4373 & n15051 ) ;
  assign n29847 = n1015 & n27006 ;
  assign n29848 = n29847 ^ n23947 ^ n7079 ;
  assign n29849 = ~n17118 & n29848 ;
  assign n29850 = ~n29846 & n29849 ;
  assign n29852 = n17584 ^ n12165 ^ n1805 ;
  assign n29851 = n8539 | n12035 ;
  assign n29853 = n29852 ^ n29851 ^ 1'b0 ;
  assign n29859 = n24428 ^ n3931 ^ n358 ;
  assign n29860 = ( n3113 & ~n17332 ) | ( n3113 & n29859 ) | ( ~n17332 & n29859 ) ;
  assign n29861 = n29860 ^ n6827 ^ n2133 ;
  assign n29856 = n2283 | n7039 ;
  assign n29857 = n4035 | n29856 ;
  assign n29854 = n10813 ^ n4757 ^ 1'b0 ;
  assign n29855 = n29854 ^ n27758 ^ n16421 ;
  assign n29858 = n29857 ^ n29855 ^ n21812 ;
  assign n29862 = n29861 ^ n29858 ^ n15952 ;
  assign n29865 = ( ~n9114 & n9772 ) | ( ~n9114 & n16511 ) | ( n9772 & n16511 ) ;
  assign n29863 = ~n10380 & n10602 ;
  assign n29864 = n29863 ^ n2802 ^ 1'b0 ;
  assign n29866 = n29865 ^ n29864 ^ 1'b0 ;
  assign n29867 = ~n13031 & n29866 ;
  assign n29868 = ~n2823 & n29867 ;
  assign n29869 = n848 & n29868 ;
  assign n29870 = n29869 ^ n24429 ^ n16736 ;
  assign n29871 = n5415 & n10649 ;
  assign n29872 = n4043 & n29871 ;
  assign n29873 = n1928 | n29872 ;
  assign n29874 = n29873 ^ n14993 ^ n5690 ;
  assign n29875 = n14139 ^ n12299 ^ 1'b0 ;
  assign n29876 = ( ~n18206 & n22250 ) | ( ~n18206 & n29875 ) | ( n22250 & n29875 ) ;
  assign n29877 = ( n831 & ~n12898 ) | ( n831 & n29876 ) | ( ~n12898 & n29876 ) ;
  assign n29878 = n12419 ^ n10900 ^ 1'b0 ;
  assign n29879 = n29878 ^ n11455 ^ 1'b0 ;
  assign n29882 = n26817 ^ n17803 ^ n15506 ;
  assign n29880 = n18687 ^ n2134 ^ n1424 ;
  assign n29881 = n8132 | n29880 ;
  assign n29883 = n29882 ^ n29881 ^ 1'b0 ;
  assign n29884 = n8360 | n15204 ;
  assign n29885 = n24543 ^ n24061 ^ n15398 ;
  assign n29886 = n26474 & ~n29885 ;
  assign n29887 = n29886 ^ n5104 ^ 1'b0 ;
  assign n29888 = n10079 ^ n8591 ^ 1'b0 ;
  assign n29889 = ( n17278 & n24424 ) | ( n17278 & ~n29888 ) | ( n24424 & ~n29888 ) ;
  assign n29890 = ( n487 & ~n9733 ) | ( n487 & n29889 ) | ( ~n9733 & n29889 ) ;
  assign n29891 = n19108 | n29890 ;
  assign n29892 = n29891 ^ n16174 ^ 1'b0 ;
  assign n29893 = n20493 ^ n10731 ^ n4019 ;
  assign n29894 = ~n22115 & n29893 ;
  assign n29895 = n5508 & n29894 ;
  assign n29896 = n25242 ^ n17605 ^ 1'b0 ;
  assign n29897 = ( n4373 & n9029 ) | ( n4373 & ~n16275 ) | ( n9029 & ~n16275 ) ;
  assign n29898 = ( n3072 & n4564 ) | ( n3072 & n7075 ) | ( n4564 & n7075 ) ;
  assign n29899 = ~n3340 & n6298 ;
  assign n29900 = ( n3575 & n29898 ) | ( n3575 & n29899 ) | ( n29898 & n29899 ) ;
  assign n29901 = ~x6 & n22952 ;
  assign n29902 = n2028 ^ n1832 ^ 1'b0 ;
  assign n29903 = n29902 ^ n6645 ^ 1'b0 ;
  assign n29904 = n5872 | n29903 ;
  assign n29905 = ( ~n6905 & n29901 ) | ( ~n6905 & n29904 ) | ( n29901 & n29904 ) ;
  assign n29906 = ( ~n29897 & n29900 ) | ( ~n29897 & n29905 ) | ( n29900 & n29905 ) ;
  assign n29907 = n24560 ^ n22955 ^ n9402 ;
  assign n29908 = ~n6051 & n29907 ;
  assign n29909 = n29908 ^ n15382 ^ 1'b0 ;
  assign n29910 = ( ~n7729 & n11651 ) | ( ~n7729 & n26901 ) | ( n11651 & n26901 ) ;
  assign n29911 = n29910 ^ n11345 ^ 1'b0 ;
  assign n29912 = n29911 ^ n26231 ^ n17631 ;
  assign n29913 = n26561 ^ n3688 ^ 1'b0 ;
  assign n29914 = n4894 & n11442 ;
  assign n29915 = ( ~n1727 & n4456 ) | ( ~n1727 & n29914 ) | ( n4456 & n29914 ) ;
  assign n29921 = n4100 | n6269 ;
  assign n29919 = n22213 ^ n6634 ^ n1116 ;
  assign n29917 = n23011 ^ n15783 ^ n3478 ;
  assign n29918 = n4516 & ~n29917 ;
  assign n29920 = n29919 ^ n29918 ^ 1'b0 ;
  assign n29916 = n10574 ^ n9538 ^ 1'b0 ;
  assign n29922 = n29921 ^ n29920 ^ n29916 ;
  assign n29923 = n7523 | n10176 ;
  assign n29924 = ( ~n21105 & n21109 ) | ( ~n21105 & n22750 ) | ( n21109 & n22750 ) ;
  assign n29925 = ( ~n13599 & n15368 ) | ( ~n13599 & n29924 ) | ( n15368 & n29924 ) ;
  assign n29926 = n29925 ^ n1352 ^ 1'b0 ;
  assign n29927 = n8424 ^ n4935 ^ 1'b0 ;
  assign n29928 = n29927 ^ n23219 ^ 1'b0 ;
  assign n29929 = ( ~n1603 & n2457 ) | ( ~n1603 & n10517 ) | ( n2457 & n10517 ) ;
  assign n29930 = ( n13959 & n28157 ) | ( n13959 & n28588 ) | ( n28157 & n28588 ) ;
  assign n29931 = n29930 ^ n968 ^ 1'b0 ;
  assign n29932 = ~n20908 & n29931 ;
  assign n29933 = n7044 | n11912 ;
  assign n29934 = n14890 | n29933 ;
  assign n29935 = ( n2350 & n5208 ) | ( n2350 & ~n8230 ) | ( n5208 & ~n8230 ) ;
  assign n29936 = n2041 & ~n18882 ;
  assign n29937 = n11634 & n29936 ;
  assign n29938 = ( n8662 & ~n15744 ) | ( n8662 & n29937 ) | ( ~n15744 & n29937 ) ;
  assign n29939 = n29938 ^ n20523 ^ 1'b0 ;
  assign n29940 = ~n29935 & n29939 ;
  assign n29941 = ( ~n12716 & n29934 ) | ( ~n12716 & n29940 ) | ( n29934 & n29940 ) ;
  assign n29942 = n14044 ^ n6161 ^ 1'b0 ;
  assign n29943 = n29942 ^ n28152 ^ n25085 ;
  assign n29944 = ( ~n10086 & n22101 ) | ( ~n10086 & n26959 ) | ( n22101 & n26959 ) ;
  assign n29945 = n29674 ^ n1207 ^ 1'b0 ;
  assign n29946 = n18164 ^ n8892 ^ 1'b0 ;
  assign n29947 = n29946 ^ n23593 ^ n16325 ;
  assign n29948 = ~n24213 & n24241 ;
  assign n29949 = ~n24563 & n29948 ;
  assign n29950 = n9940 | n20415 ;
  assign n29951 = ~n26798 & n29950 ;
  assign n29952 = ~n25773 & n29951 ;
  assign n29953 = ( n766 & ~n6411 ) | ( n766 & n13084 ) | ( ~n6411 & n13084 ) ;
  assign n29954 = n8470 & ~n19155 ;
  assign n29955 = ~n10169 & n29954 ;
  assign n29956 = n29955 ^ n26789 ^ n7728 ;
  assign n29957 = ~n8635 & n13220 ;
  assign n29958 = ~n27037 & n29957 ;
  assign n29959 = n29958 ^ n8083 ^ n6816 ;
  assign n29960 = ~n636 & n8759 ;
  assign n29961 = n29960 ^ n13709 ^ 1'b0 ;
  assign n29962 = n10243 & ~n29961 ;
  assign n29963 = n29959 & n29962 ;
  assign n29964 = n4272 | n13449 ;
  assign n29965 = n29964 ^ n25641 ^ 1'b0 ;
  assign n29966 = n29965 ^ n24519 ^ n9788 ;
  assign n29967 = n16735 | n20594 ;
  assign n29968 = ( n659 & ~n23694 ) | ( n659 & n29967 ) | ( ~n23694 & n29967 ) ;
  assign n29969 = ( n5488 & ~n17787 ) | ( n5488 & n29968 ) | ( ~n17787 & n29968 ) ;
  assign n29970 = n25216 | n29969 ;
  assign n29971 = n29966 | n29970 ;
  assign n29972 = n29920 ^ n19439 ^ 1'b0 ;
  assign n29973 = ( n8377 & n16625 ) | ( n8377 & n24594 ) | ( n16625 & n24594 ) ;
  assign n29974 = n29973 ^ n13744 ^ n3454 ;
  assign n29975 = n29974 ^ n9509 ^ 1'b0 ;
  assign n29976 = ~n29972 & n29975 ;
  assign n29977 = n2566 | n22189 ;
  assign n29978 = n8321 ^ n3736 ^ 1'b0 ;
  assign n29979 = ( n13130 & n20643 ) | ( n13130 & n26388 ) | ( n20643 & n26388 ) ;
  assign n29984 = n12773 ^ n3954 ^ n2570 ;
  assign n29983 = n14523 ^ n4703 ^ x80 ;
  assign n29985 = n29984 ^ n29983 ^ 1'b0 ;
  assign n29981 = ~n2636 & n9568 ;
  assign n29982 = n29981 ^ n3448 ^ 1'b0 ;
  assign n29980 = ( n2451 & n6497 ) | ( n2451 & n16831 ) | ( n6497 & n16831 ) ;
  assign n29986 = n29985 ^ n29982 ^ n29980 ;
  assign n29987 = n28833 ^ n19350 ^ n9411 ;
  assign n29992 = n16019 ^ n13351 ^ 1'b0 ;
  assign n29993 = n29992 ^ n7493 ^ n5888 ;
  assign n29988 = ( ~n6441 & n7261 ) | ( ~n6441 & n20398 ) | ( n7261 & n20398 ) ;
  assign n29989 = n29988 ^ n18861 ^ 1'b0 ;
  assign n29990 = ( n3418 & ~n15389 ) | ( n3418 & n29989 ) | ( ~n15389 & n29989 ) ;
  assign n29991 = n29990 ^ n18629 ^ n4748 ;
  assign n29994 = n29993 ^ n29991 ^ n26542 ;
  assign n29995 = ~n7348 & n29994 ;
  assign n29996 = n25982 & n29995 ;
  assign n29997 = n29987 & n29996 ;
  assign n29998 = n21525 ^ n6544 ^ n2148 ;
  assign n29999 = n29998 ^ n4449 ^ 1'b0 ;
  assign n30000 = n29999 ^ n16314 ^ n1605 ;
  assign n30001 = n18986 ^ n13936 ^ 1'b0 ;
  assign n30002 = n18183 ^ n17509 ^ n1649 ;
  assign n30003 = ( ~n1019 & n13720 ) | ( ~n1019 & n30002 ) | ( n13720 & n30002 ) ;
  assign n30004 = n7246 | n30003 ;
  assign n30005 = n13746 & ~n30004 ;
  assign n30009 = ( n1283 & n1485 ) | ( n1283 & ~n6601 ) | ( n1485 & ~n6601 ) ;
  assign n30010 = n30009 ^ n14555 ^ n4572 ;
  assign n30011 = n30010 ^ n25220 ^ n1607 ;
  assign n30007 = n5334 | n25097 ;
  assign n30008 = n6556 & ~n30007 ;
  assign n30012 = n30011 ^ n30008 ^ n4051 ;
  assign n30006 = n17015 ^ n9898 ^ n988 ;
  assign n30013 = n30012 ^ n30006 ^ n14012 ;
  assign n30014 = n825 & n5896 ;
  assign n30015 = n19943 & ~n29875 ;
  assign n30016 = n14678 & ~n30015 ;
  assign n30024 = n4957 ^ n1709 ^ 1'b0 ;
  assign n30025 = ~n14572 & n30024 ;
  assign n30022 = ( n1324 & ~n3789 ) | ( n1324 & n10421 ) | ( ~n3789 & n10421 ) ;
  assign n30023 = n30022 ^ n17207 ^ n4793 ;
  assign n30017 = ( n2111 & n2212 ) | ( n2111 & ~n10521 ) | ( n2212 & ~n10521 ) ;
  assign n30018 = ~n14296 & n30017 ;
  assign n30019 = n30018 ^ n12588 ^ 1'b0 ;
  assign n30020 = n17748 | n30019 ;
  assign n30021 = n30020 ^ n20091 ^ 1'b0 ;
  assign n30026 = n30025 ^ n30023 ^ n30021 ;
  assign n30027 = n30026 ^ n6813 ^ n6361 ;
  assign n30028 = ~n21241 & n30027 ;
  assign n30029 = n17855 ^ n10458 ^ n807 ;
  assign n30030 = n14702 & ~n29791 ;
  assign n30031 = n7644 ^ n4038 ^ 1'b0 ;
  assign n30032 = n2329 | n30031 ;
  assign n30033 = ( n279 & n23727 ) | ( n279 & n30032 ) | ( n23727 & n30032 ) ;
  assign n30034 = n269 & ~n4329 ;
  assign n30035 = ~n8669 & n30034 ;
  assign n30036 = n4523 ^ n3240 ^ n2350 ;
  assign n30037 = ( ~n13897 & n30035 ) | ( ~n13897 & n30036 ) | ( n30035 & n30036 ) ;
  assign n30038 = ( ~n15628 & n30033 ) | ( ~n15628 & n30037 ) | ( n30033 & n30037 ) ;
  assign n30039 = n15056 ^ n6680 ^ n3819 ;
  assign n30040 = ( ~n1016 & n25432 ) | ( ~n1016 & n30039 ) | ( n25432 & n30039 ) ;
  assign n30041 = n30040 ^ n27434 ^ n25564 ;
  assign n30043 = n28764 ^ n27060 ^ n5414 ;
  assign n30044 = n13880 | n30043 ;
  assign n30045 = n3761 | n30044 ;
  assign n30042 = n12021 & n13685 ;
  assign n30046 = n30045 ^ n30042 ^ 1'b0 ;
  assign n30047 = n21510 ^ n4677 ^ 1'b0 ;
  assign n30054 = n4789 ^ n4671 ^ n1589 ;
  assign n30055 = ( n11661 & n15329 ) | ( n11661 & ~n30054 ) | ( n15329 & ~n30054 ) ;
  assign n30056 = n24589 | n30055 ;
  assign n30057 = n30056 ^ n263 ^ 1'b0 ;
  assign n30058 = n30057 ^ n11327 ^ n261 ;
  assign n30048 = n17508 ^ n6591 ^ n2097 ;
  assign n30049 = n30048 ^ n22125 ^ n18166 ;
  assign n30050 = n4143 & n8617 ;
  assign n30051 = n30050 ^ n15535 ^ 1'b0 ;
  assign n30052 = ( ~n1743 & n22097 ) | ( ~n1743 & n30051 ) | ( n22097 & n30051 ) ;
  assign n30053 = ( n26653 & n30049 ) | ( n26653 & ~n30052 ) | ( n30049 & ~n30052 ) ;
  assign n30059 = n30058 ^ n30053 ^ n29885 ;
  assign n30060 = n30059 ^ n27364 ^ n15464 ;
  assign n30061 = n2782 | n14523 ;
  assign n30062 = n19792 ^ n11552 ^ n7176 ;
  assign n30063 = ( n15480 & n30061 ) | ( n15480 & ~n30062 ) | ( n30061 & ~n30062 ) ;
  assign n30064 = n25978 ^ n19658 ^ n16364 ;
  assign n30065 = ~n7910 & n16180 ;
  assign n30066 = ( n24856 & ~n30064 ) | ( n24856 & n30065 ) | ( ~n30064 & n30065 ) ;
  assign n30067 = ~n20648 & n25173 ;
  assign n30068 = ( ~n6685 & n16047 ) | ( ~n6685 & n30067 ) | ( n16047 & n30067 ) ;
  assign n30070 = n27023 ^ n15287 ^ 1'b0 ;
  assign n30071 = n16776 & n30070 ;
  assign n30069 = n438 | n21340 ;
  assign n30072 = n30071 ^ n30069 ^ 1'b0 ;
  assign n30073 = n12241 ^ n5494 ^ 1'b0 ;
  assign n30074 = n30073 ^ n27248 ^ 1'b0 ;
  assign n30075 = n2052 & n30074 ;
  assign n30076 = n30075 ^ n29510 ^ n16345 ;
  assign n30077 = n4366 & n15173 ;
  assign n30078 = n30076 & n30077 ;
  assign n30079 = ( n817 & n5214 ) | ( n817 & n27042 ) | ( n5214 & n27042 ) ;
  assign n30080 = n2228 & ~n9717 ;
  assign n30081 = ~n11553 & n30080 ;
  assign n30082 = n8567 | n15123 ;
  assign n30083 = ( ~n12827 & n30081 ) | ( ~n12827 & n30082 ) | ( n30081 & n30082 ) ;
  assign n30084 = n30083 ^ n23567 ^ n23021 ;
  assign n30085 = n22551 ^ n4747 ^ 1'b0 ;
  assign n30086 = n6229 & ~n30085 ;
  assign n30087 = n30086 ^ n23842 ^ 1'b0 ;
  assign n30088 = n21587 ^ n17626 ^ 1'b0 ;
  assign n30089 = n22622 ^ n13065 ^ n10430 ;
  assign n30090 = n30089 ^ n19494 ^ 1'b0 ;
  assign n30091 = n12744 & n30090 ;
  assign n30092 = ( n7457 & n23748 ) | ( n7457 & n27860 ) | ( n23748 & n27860 ) ;
  assign n30093 = n12420 ^ n4658 ^ n2362 ;
  assign n30094 = n16925 ^ n5942 ^ n5651 ;
  assign n30095 = n1716 | n9183 ;
  assign n30096 = n30095 ^ n12876 ^ 1'b0 ;
  assign n30097 = n13097 & ~n30096 ;
  assign n30098 = n30097 ^ n5824 ^ 1'b0 ;
  assign n30099 = n12638 & n27076 ;
  assign n30100 = n30099 ^ n14186 ^ 1'b0 ;
  assign n30101 = n24960 ^ n12483 ^ n10087 ;
  assign n30102 = ( n9030 & n28963 ) | ( n9030 & ~n30101 ) | ( n28963 & ~n30101 ) ;
  assign n30104 = ( n8021 & n12271 ) | ( n8021 & ~n16671 ) | ( n12271 & ~n16671 ) ;
  assign n30103 = n2591 & ~n9446 ;
  assign n30105 = n30104 ^ n30103 ^ n11942 ;
  assign n30106 = ( ~n2105 & n12065 ) | ( ~n2105 & n15293 ) | ( n12065 & n15293 ) ;
  assign n30107 = n27094 ^ n8348 ^ 1'b0 ;
  assign n30108 = n30106 & n30107 ;
  assign n30109 = n6767 | n14749 ;
  assign n30110 = n30026 ^ n4855 ^ 1'b0 ;
  assign n30111 = n21889 ^ n12912 ^ 1'b0 ;
  assign n30113 = ~n1719 & n4203 ;
  assign n30112 = n22856 ^ n370 ^ 1'b0 ;
  assign n30114 = n30113 ^ n30112 ^ n18488 ;
  assign n30115 = ~n3073 & n3416 ;
  assign n30116 = n30115 ^ n21277 ^ 1'b0 ;
  assign n30117 = n30116 ^ n27211 ^ 1'b0 ;
  assign n30118 = n30114 | n30117 ;
  assign n30119 = n21842 ^ n19636 ^ n19033 ;
  assign n30122 = n6596 & n13118 ;
  assign n30123 = n30122 ^ n11600 ^ 1'b0 ;
  assign n30120 = n19471 ^ n1529 ^ 1'b0 ;
  assign n30121 = n22953 | n30120 ;
  assign n30124 = n30123 ^ n30121 ^ n1394 ;
  assign n30125 = n30124 ^ n24722 ^ n17332 ;
  assign n30126 = n30125 ^ n24703 ^ n15727 ;
  assign n30127 = n1292 | n11994 ;
  assign n30128 = n30127 ^ n1729 ^ 1'b0 ;
  assign n30129 = ~n10619 & n30128 ;
  assign n30130 = n7570 | n17572 ;
  assign n30131 = n30130 ^ n29175 ^ n15149 ;
  assign n30132 = n30131 ^ n24806 ^ n13506 ;
  assign n30133 = n11369 ^ n10152 ^ n3635 ;
  assign n30134 = ( n12451 & n20524 ) | ( n12451 & ~n26679 ) | ( n20524 & ~n26679 ) ;
  assign n30135 = ( ~n17736 & n30133 ) | ( ~n17736 & n30134 ) | ( n30133 & n30134 ) ;
  assign n30137 = ( n1601 & n6272 ) | ( n1601 & n18552 ) | ( n6272 & n18552 ) ;
  assign n30136 = n17811 ^ n11882 ^ 1'b0 ;
  assign n30138 = n30137 ^ n30136 ^ n13224 ;
  assign n30139 = n24985 ^ n12034 ^ x156 ;
  assign n30140 = ( n6296 & n18814 ) | ( n6296 & ~n30139 ) | ( n18814 & ~n30139 ) ;
  assign n30141 = n17391 ^ n17185 ^ n12025 ;
  assign n30142 = n9332 ^ n1914 ^ 1'b0 ;
  assign n30143 = n3837 & n16048 ;
  assign n30144 = ~n30142 & n30143 ;
  assign n30145 = n30141 & n30144 ;
  assign n30146 = n29359 ^ n24433 ^ n15309 ;
  assign n30147 = n4293 | n16989 ;
  assign n30148 = n20521 & ~n30147 ;
  assign n30149 = n30148 ^ n14497 ^ n10402 ;
  assign n30150 = n30149 ^ n8269 ^ n681 ;
  assign n30151 = n22942 ^ n20035 ^ n12831 ;
  assign n30156 = n5585 ^ n1921 ^ 1'b0 ;
  assign n30152 = n17254 ^ n8560 ^ 1'b0 ;
  assign n30153 = n8839 & n30152 ;
  assign n30154 = n9811 ^ n9162 ^ 1'b0 ;
  assign n30155 = ( n7948 & n30153 ) | ( n7948 & ~n30154 ) | ( n30153 & ~n30154 ) ;
  assign n30157 = n30156 ^ n30155 ^ n20407 ;
  assign n30158 = n30157 ^ n424 ^ 1'b0 ;
  assign n30159 = n30158 ^ n1593 ^ 1'b0 ;
  assign n30160 = n7070 ^ n1528 ^ 1'b0 ;
  assign n30161 = n30159 & n30160 ;
  assign n30162 = ( n10574 & n16701 ) | ( n10574 & n21518 ) | ( n16701 & n21518 ) ;
  assign n30163 = n3609 ^ n549 ^ n502 ;
  assign n30164 = ~n598 & n30163 ;
  assign n30165 = ~n274 & n4531 ;
  assign n30166 = n30165 ^ n850 ^ 1'b0 ;
  assign n30167 = n30166 ^ n10988 ^ 1'b0 ;
  assign n30168 = n15047 | n30167 ;
  assign n30169 = ( n20262 & n27612 ) | ( n20262 & ~n30168 ) | ( n27612 & ~n30168 ) ;
  assign n30173 = n13886 ^ n3758 ^ n598 ;
  assign n30174 = n30173 ^ n14299 ^ n1616 ;
  assign n30170 = n5619 | n16954 ;
  assign n30171 = n30170 ^ n29935 ^ 1'b0 ;
  assign n30172 = ( n8037 & n15841 ) | ( n8037 & n30171 ) | ( n15841 & n30171 ) ;
  assign n30175 = n30174 ^ n30172 ^ n10561 ;
  assign n30176 = n1681 | n18169 ;
  assign n30177 = ( n3915 & n28474 ) | ( n3915 & n30176 ) | ( n28474 & n30176 ) ;
  assign n30178 = n19271 & ~n26370 ;
  assign n30179 = n30178 ^ n11206 ^ 1'b0 ;
  assign n30180 = n30179 ^ n15066 ^ 1'b0 ;
  assign n30181 = n30177 | n30180 ;
  assign n30182 = n291 | n11826 ;
  assign n30183 = n30182 ^ n10328 ^ 1'b0 ;
  assign n30184 = ( n8710 & n28105 ) | ( n8710 & ~n30183 ) | ( n28105 & ~n30183 ) ;
  assign n30185 = ~n668 & n3185 ;
  assign n30186 = n30185 ^ n10175 ^ 1'b0 ;
  assign n30187 = ~n11234 & n30186 ;
  assign n30188 = ( n20536 & n25906 ) | ( n20536 & n30187 ) | ( n25906 & n30187 ) ;
  assign n30189 = n5023 & ~n20594 ;
  assign n30190 = ~n3846 & n30189 ;
  assign n30191 = ( n28590 & n29383 ) | ( n28590 & n30190 ) | ( n29383 & n30190 ) ;
  assign n30193 = n2794 & n7362 ;
  assign n30192 = n5054 & n23211 ;
  assign n30194 = n30193 ^ n30192 ^ 1'b0 ;
  assign n30195 = ~n8750 & n20328 ;
  assign n30196 = n30195 ^ n14861 ^ 1'b0 ;
  assign n30197 = ( n14775 & n15819 ) | ( n14775 & ~n29088 ) | ( n15819 & ~n29088 ) ;
  assign n30198 = ~n1789 & n8501 ;
  assign n30199 = n30198 ^ n7727 ^ 1'b0 ;
  assign n30200 = ~n5078 & n30199 ;
  assign n30201 = ~n9913 & n30200 ;
  assign n30202 = ~n12336 & n30201 ;
  assign n30203 = ( n10128 & n15041 ) | ( n10128 & n22407 ) | ( n15041 & n22407 ) ;
  assign n30204 = n14850 & ~n24271 ;
  assign n30205 = n30203 & n30204 ;
  assign n30206 = n30179 ^ n26853 ^ n2094 ;
  assign n30207 = ~n12672 & n30206 ;
  assign n30208 = n10980 ^ n8848 ^ 1'b0 ;
  assign n30209 = ( n16447 & n30092 ) | ( n16447 & ~n30208 ) | ( n30092 & ~n30208 ) ;
  assign n30210 = n28908 ^ n4752 ^ 1'b0 ;
  assign n30211 = ( ~n11710 & n14078 ) | ( ~n11710 & n30210 ) | ( n14078 & n30210 ) ;
  assign n30212 = n29209 ^ n20513 ^ n978 ;
  assign n30213 = n4579 ^ n1746 ^ 1'b0 ;
  assign n30214 = n30212 & ~n30213 ;
  assign n30217 = n19146 ^ n15084 ^ n1685 ;
  assign n30218 = n16830 ^ n2203 ^ 1'b0 ;
  assign n30219 = ~n11639 & n30218 ;
  assign n30220 = ( n8901 & ~n30217 ) | ( n8901 & n30219 ) | ( ~n30217 & n30219 ) ;
  assign n30215 = x196 & n21369 ;
  assign n30216 = n30215 ^ n12090 ^ 1'b0 ;
  assign n30221 = n30220 ^ n30216 ^ n8582 ;
  assign n30222 = n12419 ^ n9934 ^ 1'b0 ;
  assign n30223 = n10672 ^ n9202 ^ n2593 ;
  assign n30224 = ( n8766 & n23533 ) | ( n8766 & ~n30223 ) | ( n23533 & ~n30223 ) ;
  assign n30225 = ~n9219 & n25857 ;
  assign n30226 = n30225 ^ n11506 ^ 1'b0 ;
  assign n30227 = ( x163 & n4733 ) | ( x163 & ~n16548 ) | ( n4733 & ~n16548 ) ;
  assign n30228 = n6244 & n30227 ;
  assign n30229 = ~n11189 & n30228 ;
  assign n30230 = n27766 | n30229 ;
  assign n30231 = n13277 & ~n24638 ;
  assign n30232 = ~n9970 & n30231 ;
  assign n30233 = x107 & n14065 ;
  assign n30234 = ~n8548 & n30233 ;
  assign n30235 = n1588 & ~n30234 ;
  assign n30236 = ( n1297 & ~n4452 ) | ( n1297 & n7861 ) | ( ~n4452 & n7861 ) ;
  assign n30237 = n30236 ^ n23539 ^ n17686 ;
  assign n30238 = n30237 ^ n29210 ^ n9853 ;
  assign n30239 = n10332 | n11652 ;
  assign n30240 = n30238 & ~n30239 ;
  assign n30241 = ( ~n1761 & n16891 ) | ( ~n1761 & n26416 ) | ( n16891 & n26416 ) ;
  assign n30242 = x240 & n938 ;
  assign n30243 = n1108 & n30242 ;
  assign n30244 = n30243 ^ n27678 ^ n21628 ;
  assign n30245 = ( n6790 & n11439 ) | ( n6790 & ~n16695 ) | ( n11439 & ~n16695 ) ;
  assign n30250 = n13317 | n14471 ;
  assign n30251 = n19472 & ~n30250 ;
  assign n30249 = ( n16607 & n26711 ) | ( n16607 & n27242 ) | ( n26711 & n27242 ) ;
  assign n30246 = n15089 & n15742 ;
  assign n30247 = n30246 ^ n28915 ^ 1'b0 ;
  assign n30248 = n30247 ^ n8189 ^ n4459 ;
  assign n30252 = n30251 ^ n30249 ^ n30248 ;
  assign n30253 = n25682 & ~n28595 ;
  assign n30254 = n14911 ^ n3642 ^ 1'b0 ;
  assign n30255 = ( n24167 & ~n25509 ) | ( n24167 & n30254 ) | ( ~n25509 & n30254 ) ;
  assign n30256 = n21039 & ~n21500 ;
  assign n30257 = n7745 ^ n4501 ^ 1'b0 ;
  assign n30258 = n7195 | n30257 ;
  assign n30259 = n4894 & ~n27418 ;
  assign n30260 = ~n4086 & n30259 ;
  assign n30261 = n1152 | n30260 ;
  assign n30262 = n23678 | n30261 ;
  assign n30265 = n2643 | n10129 ;
  assign n30263 = ( ~n10130 & n13086 ) | ( ~n10130 & n13718 ) | ( n13086 & n13718 ) ;
  assign n30264 = n4424 & ~n30263 ;
  assign n30266 = n30265 ^ n30264 ^ 1'b0 ;
  assign n30267 = n5185 ^ n653 ^ n530 ;
  assign n30268 = ( n3438 & ~n3813 ) | ( n3438 & n30267 ) | ( ~n3813 & n30267 ) ;
  assign n30269 = n30268 ^ n27965 ^ 1'b0 ;
  assign n30270 = ( ~n5678 & n9742 ) | ( ~n5678 & n29359 ) | ( n9742 & n29359 ) ;
  assign n30271 = n22770 ^ n4168 ^ 1'b0 ;
  assign n30272 = n28754 ^ n10280 ^ 1'b0 ;
  assign n30275 = n9238 ^ n3116 ^ n987 ;
  assign n30276 = n30275 ^ n7004 ^ 1'b0 ;
  assign n30277 = ~n8134 & n30276 ;
  assign n30273 = n22498 ^ n18921 ^ n1079 ;
  assign n30274 = n30273 ^ n24751 ^ n1003 ;
  assign n30278 = n30277 ^ n30274 ^ n883 ;
  assign n30279 = n27761 ^ n22171 ^ 1'b0 ;
  assign n30281 = n11451 & ~n14680 ;
  assign n30280 = n14382 & n15656 ;
  assign n30282 = n30281 ^ n30280 ^ n2894 ;
  assign n30283 = n3725 & n20619 ;
  assign n30284 = n18403 & n30283 ;
  assign n30285 = ( n7101 & n28571 ) | ( n7101 & n30284 ) | ( n28571 & n30284 ) ;
  assign n30286 = ~n20396 & n30285 ;
  assign n30287 = n22494 ^ n7907 ^ n4470 ;
  assign n30288 = n30287 ^ n8345 ^ n3562 ;
  assign n30289 = ( n10091 & ~n20974 ) | ( n10091 & n30288 ) | ( ~n20974 & n30288 ) ;
  assign n30290 = n22790 ^ n21604 ^ n15654 ;
  assign n30291 = ( ~n1898 & n28963 ) | ( ~n1898 & n30290 ) | ( n28963 & n30290 ) ;
  assign n30292 = n13662 | n18773 ;
  assign n30293 = n30292 ^ n5866 ^ 1'b0 ;
  assign n30294 = ( n3261 & n12560 ) | ( n3261 & ~n19654 ) | ( n12560 & ~n19654 ) ;
  assign n30295 = n30294 ^ n23032 ^ n6594 ;
  assign n30296 = ( ~n8269 & n12927 ) | ( ~n8269 & n25445 ) | ( n12927 & n25445 ) ;
  assign n30297 = ( n1695 & n10163 ) | ( n1695 & ~n30296 ) | ( n10163 & ~n30296 ) ;
  assign n30298 = ( n4192 & ~n12812 ) | ( n4192 & n30297 ) | ( ~n12812 & n30297 ) ;
  assign n30299 = n14034 ^ n9467 ^ 1'b0 ;
  assign n30300 = ~n11206 & n30299 ;
  assign n30301 = ( ~n27180 & n30298 ) | ( ~n27180 & n30300 ) | ( n30298 & n30300 ) ;
  assign n30302 = n28416 ^ n13794 ^ n11106 ;
  assign n30303 = n30302 ^ x53 ^ 1'b0 ;
  assign n30304 = n30303 ^ n8187 ^ n5830 ;
  assign n30305 = ( n9206 & ~n20233 ) | ( n9206 & n29595 ) | ( ~n20233 & n29595 ) ;
  assign n30306 = ( ~n4890 & n16257 ) | ( ~n4890 & n30305 ) | ( n16257 & n30305 ) ;
  assign n30307 = n30306 ^ n10677 ^ 1'b0 ;
  assign n30308 = n22555 & n30307 ;
  assign n30309 = ~n5417 & n14892 ;
  assign n30310 = n27505 ^ n14407 ^ 1'b0 ;
  assign n30311 = n14250 & n30310 ;
  assign n30312 = ~n30309 & n30311 ;
  assign n30313 = n30312 ^ n12419 ^ 1'b0 ;
  assign n30314 = n329 | n8393 ;
  assign n30315 = n22629 & ~n30314 ;
  assign n30318 = n13875 ^ n10227 ^ n1750 ;
  assign n30319 = ( ~n3947 & n15951 ) | ( ~n3947 & n30318 ) | ( n15951 & n30318 ) ;
  assign n30320 = n30319 ^ n5462 ^ n3128 ;
  assign n30316 = n17960 ^ n17490 ^ 1'b0 ;
  assign n30317 = n20205 | n30316 ;
  assign n30321 = n30320 ^ n30317 ^ 1'b0 ;
  assign n30322 = n7039 | n7184 ;
  assign n30323 = n30128 ^ n14931 ^ n987 ;
  assign n30324 = ( n27876 & n30322 ) | ( n27876 & ~n30323 ) | ( n30322 & ~n30323 ) ;
  assign n30325 = ( n1508 & ~n10447 ) | ( n1508 & n12306 ) | ( ~n10447 & n12306 ) ;
  assign n30327 = n941 | n7522 ;
  assign n30328 = n30327 ^ n7460 ^ 1'b0 ;
  assign n30326 = n28317 ^ n16389 ^ n8087 ;
  assign n30329 = n30328 ^ n30326 ^ n8205 ;
  assign n30330 = n30329 ^ n26328 ^ n4726 ;
  assign n30331 = ( n15774 & ~n26605 ) | ( n15774 & n30330 ) | ( ~n26605 & n30330 ) ;
  assign n30332 = n26529 ^ n1009 ^ n986 ;
  assign n30333 = ( n7944 & ~n25831 ) | ( n7944 & n30332 ) | ( ~n25831 & n30332 ) ;
  assign n30334 = n25698 ^ n6985 ^ 1'b0 ;
  assign n30335 = n7961 & ~n11773 ;
  assign n30336 = n11573 | n30335 ;
  assign n30337 = ( ~n5182 & n5593 ) | ( ~n5182 & n13701 ) | ( n5593 & n13701 ) ;
  assign n30338 = n30337 ^ x139 ^ 1'b0 ;
  assign n30339 = n13296 ^ n7188 ^ 1'b0 ;
  assign n30340 = ( ~n1586 & n9154 ) | ( ~n1586 & n9438 ) | ( n9154 & n9438 ) ;
  assign n30341 = n30340 ^ n24777 ^ n15615 ;
  assign n30342 = n30341 ^ n29088 ^ n696 ;
  assign n30348 = n16964 ^ n8088 ^ n2825 ;
  assign n30345 = n1865 & ~n2194 ;
  assign n30346 = ( n6915 & n11991 ) | ( n6915 & ~n30345 ) | ( n11991 & ~n30345 ) ;
  assign n30343 = ~n13604 & n25886 ;
  assign n30344 = n30343 ^ n1685 ^ 1'b0 ;
  assign n30347 = n30346 ^ n30344 ^ n20998 ;
  assign n30349 = n30348 ^ n30347 ^ n19399 ;
  assign n30350 = ( n2706 & ~n6444 ) | ( n2706 & n27520 ) | ( ~n6444 & n27520 ) ;
  assign n30351 = ( ~n2173 & n12001 ) | ( ~n2173 & n18991 ) | ( n12001 & n18991 ) ;
  assign n30353 = n29662 ^ n12040 ^ n323 ;
  assign n30352 = n15214 ^ n13119 ^ n4294 ;
  assign n30354 = n30353 ^ n30352 ^ n18889 ;
  assign n30355 = ( ~n9775 & n30351 ) | ( ~n9775 & n30354 ) | ( n30351 & n30354 ) ;
  assign n30356 = ~n30350 & n30355 ;
  assign n30357 = ~n21075 & n30356 ;
  assign n30360 = n19445 ^ n13659 ^ 1'b0 ;
  assign n30361 = ~n768 & n30360 ;
  assign n30358 = n25929 ^ n14017 ^ n3985 ;
  assign n30359 = n11001 & n30358 ;
  assign n30362 = n30361 ^ n30359 ^ 1'b0 ;
  assign n30363 = ( ~n3799 & n6963 ) | ( ~n3799 & n20131 ) | ( n6963 & n20131 ) ;
  assign n30364 = ( n1457 & n11125 ) | ( n1457 & ~n29431 ) | ( n11125 & ~n29431 ) ;
  assign n30365 = n4189 | n10007 ;
  assign n30366 = n30365 ^ n28999 ^ 1'b0 ;
  assign n30367 = n8241 ^ n8135 ^ n485 ;
  assign n30368 = ( ~n17576 & n30366 ) | ( ~n17576 & n30367 ) | ( n30366 & n30367 ) ;
  assign n30371 = ~n6255 & n11748 ;
  assign n30369 = n11879 & ~n26637 ;
  assign n30370 = n11188 & n30369 ;
  assign n30372 = n30371 ^ n30370 ^ n17867 ;
  assign n30373 = n30372 ^ n12069 ^ n1593 ;
  assign n30376 = n1590 ^ n944 ^ 1'b0 ;
  assign n30377 = n30376 ^ n8180 ^ n3134 ;
  assign n30378 = n30377 ^ n7270 ^ n5956 ;
  assign n30374 = n21640 ^ n17499 ^ 1'b0 ;
  assign n30375 = ~n17302 & n30374 ;
  assign n30379 = n30378 ^ n30375 ^ n1570 ;
  assign n30380 = n19893 ^ n11236 ^ 1'b0 ;
  assign n30381 = n30379 | n30380 ;
  assign n30382 = n30381 ^ n7658 ^ 1'b0 ;
  assign n30383 = n22462 ^ n13962 ^ n13052 ;
  assign n30384 = n30383 ^ n7211 ^ 1'b0 ;
  assign n30385 = n7316 & n30384 ;
  assign n30386 = n27468 ^ n9949 ^ 1'b0 ;
  assign n30387 = n3226 & n30386 ;
  assign n30388 = n30387 ^ n10912 ^ 1'b0 ;
  assign n30389 = ~n30385 & n30388 ;
  assign n30390 = n14401 ^ n13784 ^ n2457 ;
  assign n30391 = n1886 & ~n3649 ;
  assign n30392 = n14042 & n30391 ;
  assign n30393 = ( ~n11554 & n21342 ) | ( ~n11554 & n30392 ) | ( n21342 & n30392 ) ;
  assign n30394 = ~n30390 & n30393 ;
  assign n30395 = ~n30389 & n30394 ;
  assign n30396 = ~n23056 & n27037 ;
  assign n30397 = ~n16182 & n30396 ;
  assign n30398 = ~n13306 & n20324 ;
  assign n30399 = n30398 ^ n12469 ^ n11075 ;
  assign n30400 = n23451 ^ n13465 ^ n4576 ;
  assign n30401 = ( n6784 & n10640 ) | ( n6784 & n16955 ) | ( n10640 & n16955 ) ;
  assign n30402 = n28077 | n30341 ;
  assign n30403 = n18870 | n30402 ;
  assign n30404 = n9986 ^ n2793 ^ n456 ;
  assign n30405 = n1208 & ~n20647 ;
  assign n30406 = n30404 & n30405 ;
  assign n30407 = n14667 & ~n30406 ;
  assign n30408 = ~n30403 & n30407 ;
  assign n30409 = ~n5984 & n12353 ;
  assign n30410 = n21018 & n30409 ;
  assign n30411 = n30410 ^ n20216 ^ n17840 ;
  assign n30412 = ( n30401 & n30408 ) | ( n30401 & ~n30411 ) | ( n30408 & ~n30411 ) ;
  assign n30413 = ( x218 & n4460 ) | ( x218 & n6253 ) | ( n4460 & n6253 ) ;
  assign n30414 = ( n9818 & ~n14628 ) | ( n9818 & n30413 ) | ( ~n14628 & n30413 ) ;
  assign n30415 = n7977 & n30414 ;
  assign n30416 = n23184 & n30415 ;
  assign n30420 = n6442 & n7169 ;
  assign n30421 = n30420 ^ n25704 ^ n2931 ;
  assign n30417 = n5326 & ~n17756 ;
  assign n30418 = n16950 ^ n6015 ^ 1'b0 ;
  assign n30419 = ~n30417 & n30418 ;
  assign n30422 = n30421 ^ n30419 ^ n22532 ;
  assign n30426 = n14870 ^ n13836 ^ n4029 ;
  assign n30424 = ( ~n6572 & n14775 ) | ( ~n6572 & n27338 ) | ( n14775 & n27338 ) ;
  assign n30423 = ~n1257 & n3374 ;
  assign n30425 = n30424 ^ n30423 ^ n17270 ;
  assign n30427 = n30426 ^ n30425 ^ n18962 ;
  assign n30428 = n5414 ^ n4866 ^ n637 ;
  assign n30429 = ~n11201 & n30428 ;
  assign n30430 = n9913 ^ n4178 ^ n3431 ;
  assign n30431 = ( n9830 & n19159 ) | ( n9830 & ~n21248 ) | ( n19159 & ~n21248 ) ;
  assign n30432 = ( n2911 & ~n30430 ) | ( n2911 & n30431 ) | ( ~n30430 & n30431 ) ;
  assign n30433 = n18391 ^ n17069 ^ n15245 ;
  assign n30434 = n12895 & n26119 ;
  assign n30436 = n404 & ~n12221 ;
  assign n30435 = ( n4609 & n10982 ) | ( n4609 & ~n28239 ) | ( n10982 & ~n28239 ) ;
  assign n30437 = n30436 ^ n30435 ^ n5362 ;
  assign n30438 = n22163 & n30437 ;
  assign n30439 = n30438 ^ n3517 ^ n2685 ;
  assign n30440 = n1071 & ~n6271 ;
  assign n30441 = n30440 ^ n19585 ^ 1'b0 ;
  assign n30442 = n7950 ^ n5185 ^ 1'b0 ;
  assign n30443 = n13826 ^ n4626 ^ 1'b0 ;
  assign n30446 = n17855 ^ n7475 ^ n6942 ;
  assign n30444 = ( ~n2650 & n15952 ) | ( ~n2650 & n25220 ) | ( n15952 & n25220 ) ;
  assign n30445 = n30444 ^ n13830 ^ n6318 ;
  assign n30447 = n30446 ^ n30445 ^ n19362 ;
  assign n30448 = n30447 ^ n12707 ^ n8780 ;
  assign n30451 = n27987 ^ n14895 ^ n14586 ;
  assign n30449 = n15543 ^ n9792 ^ n3596 ;
  assign n30450 = n30449 ^ n18644 ^ n1085 ;
  assign n30452 = n30451 ^ n30450 ^ n15455 ;
  assign n30453 = ( n5511 & n9436 ) | ( n5511 & ~n18484 ) | ( n9436 & ~n18484 ) ;
  assign n30454 = n7332 | n24787 ;
  assign n30455 = n30454 ^ n14540 ^ 1'b0 ;
  assign n30456 = ( n1110 & n1606 ) | ( n1110 & n12053 ) | ( n1606 & n12053 ) ;
  assign n30457 = ( n11611 & n12952 ) | ( n11611 & n30456 ) | ( n12952 & n30456 ) ;
  assign n30458 = ( n10703 & ~n26429 ) | ( n10703 & n30457 ) | ( ~n26429 & n30457 ) ;
  assign n30460 = n2630 & n9679 ;
  assign n30461 = n30460 ^ n24571 ^ 1'b0 ;
  assign n30459 = n23741 | n27938 ;
  assign n30462 = n30461 ^ n30459 ^ 1'b0 ;
  assign n30464 = n13613 ^ n12658 ^ n4046 ;
  assign n30463 = n12340 ^ n11382 ^ n1332 ;
  assign n30465 = n30464 ^ n30463 ^ n27585 ;
  assign n30466 = n30465 ^ n947 ^ 1'b0 ;
  assign n30467 = n7730 ^ n3934 ^ 1'b0 ;
  assign n30468 = ~n10845 & n30467 ;
  assign n30469 = n7947 & n30468 ;
  assign n30470 = n30469 ^ n17197 ^ n3668 ;
  assign n30471 = n8900 & ~n13900 ;
  assign n30472 = ~n30470 & n30471 ;
  assign n30473 = n29438 ^ n11637 ^ 1'b0 ;
  assign n30474 = n7309 & ~n30473 ;
  assign n30475 = ~n7828 & n17300 ;
  assign n30476 = n30475 ^ n28214 ^ 1'b0 ;
  assign n30477 = ( ~n526 & n7082 ) | ( ~n526 & n30476 ) | ( n7082 & n30476 ) ;
  assign n30478 = ( ~n14338 & n26351 ) | ( ~n14338 & n30477 ) | ( n26351 & n30477 ) ;
  assign n30479 = n18002 & ~n27046 ;
  assign n30480 = ~n30478 & n30479 ;
  assign n30481 = n23721 ^ n2509 ^ 1'b0 ;
  assign n30482 = n30480 | n30481 ;
  assign n30483 = n9531 ^ n5141 ^ n3338 ;
  assign n30484 = ( n21791 & ~n25795 ) | ( n21791 & n30483 ) | ( ~n25795 & n30483 ) ;
  assign n30485 = n13640 | n19477 ;
  assign n30486 = n30485 ^ n23994 ^ n14285 ;
  assign n30487 = n30486 ^ n17099 ^ n14678 ;
  assign n30488 = n23253 ^ n10931 ^ n1697 ;
  assign n30489 = n30488 ^ n27257 ^ n2240 ;
  assign n30495 = n19303 ^ x27 ^ 1'b0 ;
  assign n30496 = ~n1565 & n30495 ;
  assign n30490 = ( ~n334 & n4097 ) | ( ~n334 & n4136 ) | ( n4097 & n4136 ) ;
  assign n30491 = n30490 ^ n6747 ^ 1'b0 ;
  assign n30492 = n11838 & ~n30491 ;
  assign n30493 = ( n2244 & n22154 ) | ( n2244 & n30492 ) | ( n22154 & n30492 ) ;
  assign n30494 = n30493 ^ n23235 ^ n9289 ;
  assign n30497 = n30496 ^ n30494 ^ 1'b0 ;
  assign n30498 = n5106 | n30497 ;
  assign n30499 = n5155 & ~n7397 ;
  assign n30500 = n30499 ^ n3081 ^ 1'b0 ;
  assign n30501 = n30500 ^ n4188 ^ 1'b0 ;
  assign n30502 = n2579 | n11526 ;
  assign n30503 = n6036 & ~n30502 ;
  assign n30504 = n15764 | n30503 ;
  assign n30505 = n30504 ^ n24707 ^ 1'b0 ;
  assign n30506 = ( n13674 & n30501 ) | ( n13674 & n30505 ) | ( n30501 & n30505 ) ;
  assign n30507 = ( n9516 & n10344 ) | ( n9516 & ~n21620 ) | ( n10344 & ~n21620 ) ;
  assign n30508 = ~n9766 & n25673 ;
  assign n30509 = ~n1666 & n30508 ;
  assign n30510 = n30509 ^ n21419 ^ 1'b0 ;
  assign n30511 = ~n2758 & n30510 ;
  assign n30512 = ~n15581 & n30511 ;
  assign n30513 = ~n30507 & n30512 ;
  assign n30514 = ( ~n13294 & n29029 ) | ( ~n13294 & n30513 ) | ( n29029 & n30513 ) ;
  assign n30515 = n17531 | n19774 ;
  assign n30516 = n30515 ^ n17041 ^ 1'b0 ;
  assign n30517 = ( n16379 & n28387 ) | ( n16379 & n30516 ) | ( n28387 & n30516 ) ;
  assign n30518 = n20311 ^ n5473 ^ 1'b0 ;
  assign n30519 = n9350 | n30518 ;
  assign n30522 = ( n257 & n20784 ) | ( n257 & ~n23865 ) | ( n20784 & ~n23865 ) ;
  assign n30520 = ~n12998 & n21807 ;
  assign n30521 = n30520 ^ n7994 ^ 1'b0 ;
  assign n30523 = n30522 ^ n30521 ^ n8398 ;
  assign n30524 = n27443 ^ n8782 ^ 1'b0 ;
  assign n30535 = ~n9197 & n17813 ;
  assign n30534 = n11068 ^ n9706 ^ n9689 ;
  assign n30526 = n15034 ^ n3538 ^ 1'b0 ;
  assign n30528 = x108 | n2706 ;
  assign n30529 = n7577 | n30528 ;
  assign n30527 = ( ~n4923 & n8211 ) | ( ~n4923 & n16481 ) | ( n8211 & n16481 ) ;
  assign n30530 = n30529 ^ n30527 ^ n18397 ;
  assign n30531 = ~n30526 & n30530 ;
  assign n30525 = n3963 | n22453 ;
  assign n30532 = n30531 ^ n30525 ^ 1'b0 ;
  assign n30533 = n30532 ^ n27299 ^ n17150 ;
  assign n30536 = n30535 ^ n30534 ^ n30533 ;
  assign n30537 = n16443 ^ n12578 ^ 1'b0 ;
  assign n30538 = n12577 & ~n30537 ;
  assign n30539 = n28854 & n30538 ;
  assign n30540 = n12535 ^ n7021 ^ 1'b0 ;
  assign n30541 = ( n779 & n4663 ) | ( n779 & n11679 ) | ( n4663 & n11679 ) ;
  assign n30542 = n325 | n30541 ;
  assign n30543 = n30542 ^ n24387 ^ 1'b0 ;
  assign n30544 = ( n5947 & ~n13489 ) | ( n5947 & n23318 ) | ( ~n13489 & n23318 ) ;
  assign n30545 = ~n8576 & n18860 ;
  assign n30546 = n6704 & ~n25639 ;
  assign n30547 = n30546 ^ n10950 ^ 1'b0 ;
  assign n30548 = n9535 & n15046 ;
  assign n30549 = ~n30547 & n30548 ;
  assign n30553 = n8933 ^ n4603 ^ 1'b0 ;
  assign n30552 = n17079 ^ n6682 ^ 1'b0 ;
  assign n30550 = n8115 | n15535 ;
  assign n30551 = n30550 ^ n18617 ^ 1'b0 ;
  assign n30554 = n30553 ^ n30552 ^ n30551 ;
  assign n30555 = ( n5062 & n7603 ) | ( n5062 & n17038 ) | ( n7603 & n17038 ) ;
  assign n30556 = ~n1708 & n4039 ;
  assign n30557 = ( n4388 & ~n17045 ) | ( n4388 & n30556 ) | ( ~n17045 & n30556 ) ;
  assign n30558 = ( ~n13908 & n14513 ) | ( ~n13908 & n30557 ) | ( n14513 & n30557 ) ;
  assign n30559 = n3089 & ~n30558 ;
  assign n30560 = n12776 & n30559 ;
  assign n30561 = ~n3799 & n28768 ;
  assign n30562 = n30561 ^ n16914 ^ 1'b0 ;
  assign n30563 = n26834 ^ n14643 ^ n2583 ;
  assign n30564 = n15544 & ~n28572 ;
  assign n30565 = ( n7286 & n30563 ) | ( n7286 & ~n30564 ) | ( n30563 & ~n30564 ) ;
  assign n30566 = ( x112 & n19454 ) | ( x112 & ~n30565 ) | ( n19454 & ~n30565 ) ;
  assign n30567 = n3481 & ~n25584 ;
  assign n30574 = n10705 ^ n8167 ^ n589 ;
  assign n30568 = n2885 & ~n9230 ;
  assign n30569 = n20466 & n30568 ;
  assign n30570 = ( n2667 & n10461 ) | ( n2667 & ~n11750 ) | ( n10461 & ~n11750 ) ;
  assign n30571 = n9310 & n30570 ;
  assign n30572 = n30571 ^ n9012 ^ 1'b0 ;
  assign n30573 = ( ~n10665 & n30569 ) | ( ~n10665 & n30572 ) | ( n30569 & n30572 ) ;
  assign n30575 = n30574 ^ n30573 ^ n23178 ;
  assign n30576 = ( ~n1862 & n2097 ) | ( ~n1862 & n4544 ) | ( n2097 & n4544 ) ;
  assign n30577 = n14110 ^ n13063 ^ 1'b0 ;
  assign n30578 = n18994 & ~n30577 ;
  assign n30579 = n30578 ^ n12670 ^ 1'b0 ;
  assign n30580 = ~n30576 & n30579 ;
  assign n30581 = n11679 & ~n16531 ;
  assign n30582 = n30581 ^ n7307 ^ 1'b0 ;
  assign n30583 = ( n11328 & n16122 ) | ( n11328 & n18242 ) | ( n16122 & n18242 ) ;
  assign n30584 = ~n24365 & n24516 ;
  assign n30585 = n29659 ^ n15275 ^ n9209 ;
  assign n30586 = ( n2838 & n16150 ) | ( n2838 & n21163 ) | ( n16150 & n21163 ) ;
  assign n30587 = ( ~n14151 & n30585 ) | ( ~n14151 & n30586 ) | ( n30585 & n30586 ) ;
  assign n30588 = n30587 ^ n21042 ^ n14449 ;
  assign n30589 = ( x204 & n1761 ) | ( x204 & n11496 ) | ( n1761 & n11496 ) ;
  assign n30590 = ( n15284 & n21628 ) | ( n15284 & n30589 ) | ( n21628 & n30589 ) ;
  assign n30591 = ( n4668 & n6877 ) | ( n4668 & ~n30590 ) | ( n6877 & ~n30590 ) ;
  assign n30592 = ( n14849 & n26388 ) | ( n14849 & n30591 ) | ( n26388 & n30591 ) ;
  assign n30593 = n10642 & n13577 ;
  assign n30594 = n575 & ~n3210 ;
  assign n30595 = n30594 ^ n21954 ^ 1'b0 ;
  assign n30596 = n17088 & ~n29452 ;
  assign n30597 = n14533 ^ n11962 ^ 1'b0 ;
  assign n30598 = ~n7797 & n30597 ;
  assign n30599 = ~n30596 & n30598 ;
  assign n30600 = ( ~n552 & n4196 ) | ( ~n552 & n17372 ) | ( n4196 & n17372 ) ;
  assign n30601 = ~n4713 & n19820 ;
  assign n30602 = ( ~n7444 & n9745 ) | ( ~n7444 & n30601 ) | ( n9745 & n30601 ) ;
  assign n30603 = n30600 | n30602 ;
  assign n30604 = n30603 ^ n8585 ^ 1'b0 ;
  assign n30605 = ( n15396 & n16588 ) | ( n15396 & ~n30604 ) | ( n16588 & ~n30604 ) ;
  assign n30615 = n16543 ^ n12133 ^ n5144 ;
  assign n30610 = n441 | n15421 ;
  assign n30611 = n30610 ^ n19248 ^ 1'b0 ;
  assign n30612 = n30611 ^ n14684 ^ 1'b0 ;
  assign n30613 = n30612 ^ n25380 ^ n4470 ;
  assign n30614 = n26494 & ~n30613 ;
  assign n30616 = n30615 ^ n30614 ^ 1'b0 ;
  assign n30606 = n8009 & ~n10858 ;
  assign n30607 = n3054 & n30606 ;
  assign n30608 = ( n7629 & ~n21757 ) | ( n7629 & n30607 ) | ( ~n21757 & n30607 ) ;
  assign n30609 = n30608 ^ n18304 ^ 1'b0 ;
  assign n30617 = n30616 ^ n30609 ^ n7415 ;
  assign n30618 = n4997 | n17057 ;
  assign n30619 = ( n3061 & n3432 ) | ( n3061 & ~n30618 ) | ( n3432 & ~n30618 ) ;
  assign n30620 = n2765 & n4507 ;
  assign n30621 = n30463 & n30620 ;
  assign n30622 = n21174 | n30621 ;
  assign n30623 = n9370 & ~n30622 ;
  assign n30624 = n27913 ^ n4670 ^ n2947 ;
  assign n30625 = n16721 ^ n7034 ^ 1'b0 ;
  assign n30626 = ~n30624 & n30625 ;
  assign n30627 = n8804 & ~n30626 ;
  assign n30628 = n5616 & n13119 ;
  assign n30629 = n30627 & n30628 ;
  assign n30630 = n24971 ^ n5352 ^ n622 ;
  assign n30631 = n13996 & n22406 ;
  assign n30632 = ~n30630 & n30631 ;
  assign n30633 = n24389 | n30632 ;
  assign n30634 = n1308 | n30633 ;
  assign n30635 = n4563 ^ n298 ^ 1'b0 ;
  assign n30636 = ~n6221 & n11428 ;
  assign n30637 = ( n16521 & n17125 ) | ( n16521 & n30636 ) | ( n17125 & n30636 ) ;
  assign n30638 = n18485 ^ n12571 ^ n8153 ;
  assign n30639 = n17370 & ~n18264 ;
  assign n30640 = n30639 ^ n23835 ^ n7954 ;
  assign n30644 = n19155 ^ n9040 ^ n6732 ;
  assign n30642 = ( ~n9223 & n22100 ) | ( ~n9223 & n23676 ) | ( n22100 & n23676 ) ;
  assign n30641 = n27926 ^ n12043 ^ n4993 ;
  assign n30643 = n30642 ^ n30641 ^ n2442 ;
  assign n30645 = n30644 ^ n30643 ^ n27485 ;
  assign n30646 = n8564 ^ n8376 ^ 1'b0 ;
  assign n30647 = ( n6088 & ~n7494 ) | ( n6088 & n10569 ) | ( ~n7494 & n10569 ) ;
  assign n30648 = ( n571 & ~n5638 ) | ( n571 & n30647 ) | ( ~n5638 & n30647 ) ;
  assign n30649 = n9034 ^ n7111 ^ n4935 ;
  assign n30650 = n10695 | n30649 ;
  assign n30651 = n8310 | n30650 ;
  assign n30652 = n30651 ^ n6717 ^ 1'b0 ;
  assign n30653 = n8305 | n11305 ;
  assign n30654 = n5519 ^ n2837 ^ 1'b0 ;
  assign n30655 = ( n1019 & n15566 ) | ( n1019 & ~n30654 ) | ( n15566 & ~n30654 ) ;
  assign n30656 = n8063 ^ n6495 ^ 1'b0 ;
  assign n30657 = n4238 | n30656 ;
  assign n30658 = n30657 ^ n4792 ^ 1'b0 ;
  assign n30659 = ~n956 & n1946 ;
  assign n30660 = n3450 & n30659 ;
  assign n30661 = n23538 & ~n30660 ;
  assign n30662 = n16720 & n30661 ;
  assign n30663 = n30662 ^ n17038 ^ n1060 ;
  assign n30664 = n30663 ^ n24063 ^ n8427 ;
  assign n30665 = ( n12073 & n14453 ) | ( n12073 & n14702 ) | ( n14453 & n14702 ) ;
  assign n30666 = n30665 ^ n13462 ^ n11282 ;
  assign n30667 = n30666 ^ n11165 ^ n7828 ;
  assign n30670 = ( n8481 & n9721 ) | ( n8481 & ~n12133 ) | ( n9721 & ~n12133 ) ;
  assign n30668 = ( n1457 & n3265 ) | ( n1457 & ~n14436 ) | ( n3265 & ~n14436 ) ;
  assign n30669 = ( n4137 & n26267 ) | ( n4137 & ~n30668 ) | ( n26267 & ~n30668 ) ;
  assign n30671 = n30670 ^ n30669 ^ 1'b0 ;
  assign n30672 = n8554 | n30671 ;
  assign n30673 = ( n2009 & n30667 ) | ( n2009 & ~n30672 ) | ( n30667 & ~n30672 ) ;
  assign n30674 = ( n1971 & ~n4886 ) | ( n1971 & n7218 ) | ( ~n4886 & n7218 ) ;
  assign n30675 = n8351 ^ n3165 ^ 1'b0 ;
  assign n30676 = n21332 ^ n1517 ^ 1'b0 ;
  assign n30677 = n30675 & ~n30676 ;
  assign n30678 = n30677 ^ n16093 ^ n8370 ;
  assign n30679 = ( n19290 & n30674 ) | ( n19290 & n30678 ) | ( n30674 & n30678 ) ;
  assign n30680 = ( n1194 & ~n1251 ) | ( n1194 & n9988 ) | ( ~n1251 & n9988 ) ;
  assign n30681 = n4896 & ~n6052 ;
  assign n30682 = n30680 & n30681 ;
  assign n30683 = n30682 ^ n6005 ^ 1'b0 ;
  assign n30684 = ( ~n1573 & n11316 ) | ( ~n1573 & n30683 ) | ( n11316 & n30683 ) ;
  assign n30685 = n28678 ^ n2971 ^ 1'b0 ;
  assign n30686 = ( n3151 & n5367 ) | ( n3151 & n7635 ) | ( n5367 & n7635 ) ;
  assign n30687 = n30686 ^ n30163 ^ n11176 ;
  assign n30688 = n27394 ^ n16552 ^ 1'b0 ;
  assign n30689 = n30688 ^ n19739 ^ n14625 ;
  assign n30690 = n30689 ^ n7654 ^ 1'b0 ;
  assign n30691 = n26999 ^ n6883 ^ 1'b0 ;
  assign n30692 = ~n20501 & n30691 ;
  assign n30693 = ~n5374 & n30692 ;
  assign n30694 = n2627 & n2629 ;
  assign n30695 = n30694 ^ n4012 ^ 1'b0 ;
  assign n30696 = ( n4672 & ~n9272 ) | ( n4672 & n27023 ) | ( ~n9272 & n27023 ) ;
  assign n30697 = ( n6890 & n30695 ) | ( n6890 & ~n30696 ) | ( n30695 & ~n30696 ) ;
  assign n30698 = n3519 & n16886 ;
  assign n30699 = ( n7805 & ~n11437 ) | ( n7805 & n30698 ) | ( ~n11437 & n30698 ) ;
  assign n30700 = ( ~n5482 & n7876 ) | ( ~n5482 & n17174 ) | ( n7876 & n17174 ) ;
  assign n30701 = n15124 & ~n30700 ;
  assign n30702 = n16289 & n30701 ;
  assign n30703 = n30702 ^ n29986 ^ 1'b0 ;
  assign n30704 = n23428 ^ n4143 ^ n3041 ;
  assign n30705 = ~n14775 & n30704 ;
  assign n30706 = n19109 & n30705 ;
  assign n30707 = n23842 & ~n30706 ;
  assign n30708 = n30707 ^ n21511 ^ 1'b0 ;
  assign n30709 = ~n3347 & n10929 ;
  assign n30712 = ~n3334 & n6383 ;
  assign n30713 = n30712 ^ n405 ^ 1'b0 ;
  assign n30711 = ( n473 & n1587 ) | ( n473 & n5882 ) | ( n1587 & n5882 ) ;
  assign n30710 = n15654 ^ n7166 ^ 1'b0 ;
  assign n30714 = n30713 ^ n30711 ^ n30710 ;
  assign n30715 = ~n30709 & n30714 ;
  assign n30716 = ~n23231 & n30715 ;
  assign n30717 = n4543 ^ n3928 ^ n2947 ;
  assign n30718 = n30717 ^ n5546 ^ 1'b0 ;
  assign n30719 = n21836 & ~n30718 ;
  assign n30720 = n7937 ^ n7723 ^ n306 ;
  assign n30721 = n30720 ^ n23319 ^ n530 ;
  assign n30722 = n15915 ^ n9524 ^ n2886 ;
  assign n30723 = n25694 ^ n20808 ^ 1'b0 ;
  assign n30724 = n2028 & n27590 ;
  assign n30725 = ~n1856 & n30724 ;
  assign n30726 = ~n16759 & n20317 ;
  assign n30727 = n11955 ^ n3601 ^ 1'b0 ;
  assign n30728 = n30720 | n30727 ;
  assign n30729 = n15542 & n24691 ;
  assign n30730 = n23601 & n30729 ;
  assign n30731 = ( n5400 & n30728 ) | ( n5400 & ~n30730 ) | ( n30728 & ~n30730 ) ;
  assign n30733 = n13589 ^ n1373 ^ 1'b0 ;
  assign n30734 = ~n7428 & n30733 ;
  assign n30732 = n5380 & n18159 ;
  assign n30735 = n30734 ^ n30732 ^ 1'b0 ;
  assign n30736 = n2069 | n30735 ;
  assign n30737 = n15724 | n30736 ;
  assign n30738 = ~n16771 & n30737 ;
  assign n30739 = n14712 ^ n7443 ^ 1'b0 ;
  assign n30740 = ~n5050 & n30739 ;
  assign n30741 = ~n28581 & n30740 ;
  assign n30742 = n19238 ^ n13583 ^ n8551 ;
  assign n30743 = n30742 ^ n15902 ^ 1'b0 ;
  assign n30744 = n30743 ^ n13817 ^ x146 ;
  assign n30745 = n2009 | n2164 ;
  assign n30746 = n30744 | n30745 ;
  assign n30747 = n22355 ^ n13782 ^ 1'b0 ;
  assign n30749 = n30366 ^ n27755 ^ n2547 ;
  assign n30748 = n15270 ^ n11556 ^ 1'b0 ;
  assign n30750 = n30749 ^ n30748 ^ n7137 ;
  assign n30751 = n5230 ^ n1664 ^ 1'b0 ;
  assign n30752 = n30750 & ~n30751 ;
  assign n30753 = n8923 | n14510 ;
  assign n30754 = n30752 | n30753 ;
  assign n30755 = n21490 & ~n27198 ;
  assign n30757 = ( n11491 & n13471 ) | ( n11491 & ~n26638 ) | ( n13471 & ~n26638 ) ;
  assign n30756 = ( ~n19878 & n23544 ) | ( ~n19878 & n29183 ) | ( n23544 & n29183 ) ;
  assign n30758 = n30757 ^ n30756 ^ x227 ;
  assign n30759 = n20237 ^ n18080 ^ n2326 ;
  assign n30761 = ~n4987 & n20226 ;
  assign n30762 = ~n1433 & n30761 ;
  assign n30763 = ( n8435 & n12375 ) | ( n8435 & ~n30762 ) | ( n12375 & ~n30762 ) ;
  assign n30760 = ( n7617 & ~n22631 ) | ( n7617 & n24657 ) | ( ~n22631 & n24657 ) ;
  assign n30764 = n30763 ^ n30760 ^ n27198 ;
  assign n30766 = ~n5184 & n15945 ;
  assign n30765 = n21525 ^ n11114 ^ 1'b0 ;
  assign n30767 = n30766 ^ n30765 ^ n27617 ;
  assign n30769 = ~n12274 & n20752 ;
  assign n30770 = n30769 ^ n9113 ^ 1'b0 ;
  assign n30768 = n22053 | n30722 ;
  assign n30771 = n30770 ^ n30768 ^ 1'b0 ;
  assign n30774 = ~n366 & n18896 ;
  assign n30775 = n30774 ^ n8464 ^ 1'b0 ;
  assign n30772 = n1737 | n2728 ;
  assign n30773 = n30772 ^ n20446 ^ 1'b0 ;
  assign n30776 = n30775 ^ n30773 ^ n18710 ;
  assign n30777 = ( ~n2173 & n22202 ) | ( ~n2173 & n24562 ) | ( n22202 & n24562 ) ;
  assign n30778 = n6851 ^ n6812 ^ n2154 ;
  assign n30779 = ( n4277 & n4459 ) | ( n4277 & ~n30778 ) | ( n4459 & ~n30778 ) ;
  assign n30780 = n24338 ^ n20478 ^ 1'b0 ;
  assign n30781 = ~n17302 & n30780 ;
  assign n30782 = n19578 ^ n19036 ^ n4859 ;
  assign n30783 = n29656 ^ n6301 ^ 1'b0 ;
  assign n30784 = n13267 ^ n7670 ^ n6952 ;
  assign n30785 = ( n7262 & n28051 ) | ( n7262 & ~n30784 ) | ( n28051 & ~n30784 ) ;
  assign n30786 = n16883 ^ n13202 ^ 1'b0 ;
  assign n30787 = n16187 | n30786 ;
  assign n30788 = n993 | n30787 ;
  assign n30789 = n30788 ^ n2382 ^ n1808 ;
  assign n30790 = ( n5738 & n16950 ) | ( n5738 & ~n23452 ) | ( n16950 & ~n23452 ) ;
  assign n30791 = n30790 ^ n12622 ^ n6041 ;
  assign n30792 = ( ~n8515 & n11102 ) | ( ~n8515 & n16471 ) | ( n11102 & n16471 ) ;
  assign n30793 = n30792 ^ n5214 ^ n470 ;
  assign n30794 = n30793 ^ n23216 ^ n10169 ;
  assign n30795 = ( n3667 & ~n8100 ) | ( n3667 & n17772 ) | ( ~n8100 & n17772 ) ;
  assign n30799 = n23080 ^ n7489 ^ n2941 ;
  assign n30796 = n15172 ^ n14010 ^ 1'b0 ;
  assign n30797 = n6708 & n30796 ;
  assign n30798 = n22413 & n30797 ;
  assign n30800 = n30799 ^ n30798 ^ 1'b0 ;
  assign n30801 = n3156 & ~n3686 ;
  assign n30802 = ~n4190 & n30801 ;
  assign n30804 = n13386 ^ n7035 ^ n2332 ;
  assign n30803 = n21140 ^ n2800 ^ 1'b0 ;
  assign n30805 = n30804 ^ n30803 ^ n6582 ;
  assign n30806 = n30805 ^ n16352 ^ n4831 ;
  assign n30807 = n14398 ^ n1853 ^ 1'b0 ;
  assign n30808 = n7798 ^ n7475 ^ 1'b0 ;
  assign n30809 = ( n578 & ~n30807 ) | ( n578 & n30808 ) | ( ~n30807 & n30808 ) ;
  assign n30810 = n30809 ^ n7514 ^ n1014 ;
  assign n30811 = ( n2762 & ~n17748 ) | ( n2762 & n30810 ) | ( ~n17748 & n30810 ) ;
  assign n30812 = n30811 ^ n29600 ^ x248 ;
  assign n30814 = n916 | n16657 ;
  assign n30815 = n8111 & ~n30814 ;
  assign n30813 = n22356 ^ n14116 ^ n8915 ;
  assign n30816 = n30815 ^ n30813 ^ n1394 ;
  assign n30817 = n25422 ^ n11001 ^ 1'b0 ;
  assign n30818 = n2561 | n3313 ;
  assign n30819 = n30817 | n30818 ;
  assign n30820 = ~n7197 & n8620 ;
  assign n30821 = n19671 & n30820 ;
  assign n30822 = n3889 & ~n30821 ;
  assign n30823 = n30822 ^ n20884 ^ 1'b0 ;
  assign n30824 = n30823 ^ n17107 ^ n894 ;
  assign n30825 = ( n843 & n17140 ) | ( n843 & ~n25867 ) | ( n17140 & ~n25867 ) ;
  assign n30826 = n16905 & ~n26266 ;
  assign n30827 = ~n6743 & n30826 ;
  assign n30828 = ( n4009 & n11163 ) | ( n4009 & ~n27848 ) | ( n11163 & ~n27848 ) ;
  assign n30829 = ( ~n13852 & n30827 ) | ( ~n13852 & n30828 ) | ( n30827 & n30828 ) ;
  assign n30830 = ( ~n2321 & n10562 ) | ( ~n2321 & n13031 ) | ( n10562 & n13031 ) ;
  assign n30831 = n30830 ^ n29373 ^ n17829 ;
  assign n30832 = ( ~n5572 & n24705 ) | ( ~n5572 & n30831 ) | ( n24705 & n30831 ) ;
  assign n30833 = n28039 ^ n9069 ^ n5948 ;
  assign n30834 = n23067 | n27157 ;
  assign n30835 = n817 | n30834 ;
  assign n30836 = n2987 ^ n2392 ^ 1'b0 ;
  assign n30837 = ~n27574 & n30836 ;
  assign n30839 = ~n2736 & n17319 ;
  assign n30838 = n27866 ^ n24149 ^ n10054 ;
  assign n30840 = n30839 ^ n30838 ^ n13505 ;
  assign n30841 = n2573 & ~n7456 ;
  assign n30842 = n3130 & n30841 ;
  assign n30843 = ( ~n12557 & n14333 ) | ( ~n12557 & n30842 ) | ( n14333 & n30842 ) ;
  assign n30844 = n2116 ^ n1998 ^ 1'b0 ;
  assign n30845 = n3002 & ~n6599 ;
  assign n30846 = n30845 ^ n10650 ^ 1'b0 ;
  assign n30847 = ( n4330 & n30844 ) | ( n4330 & ~n30846 ) | ( n30844 & ~n30846 ) ;
  assign n30848 = ~n932 & n13664 ;
  assign n30849 = ( n2141 & ~n30847 ) | ( n2141 & n30848 ) | ( ~n30847 & n30848 ) ;
  assign n30850 = ( ~n21780 & n30843 ) | ( ~n21780 & n30849 ) | ( n30843 & n30849 ) ;
  assign n30851 = n19982 ^ n9586 ^ 1'b0 ;
  assign n30852 = n21319 | n30851 ;
  assign n30853 = n24060 & n30128 ;
  assign n30854 = n30853 ^ n17857 ^ 1'b0 ;
  assign n30855 = n14227 ^ n11719 ^ n10132 ;
  assign n30856 = n21216 ^ n10191 ^ 1'b0 ;
  assign n30857 = n30855 | n30856 ;
  assign n30858 = n3393 & n10892 ;
  assign n30859 = ~n2437 & n30858 ;
  assign n30860 = ( n3462 & n4707 ) | ( n3462 & ~n5392 ) | ( n4707 & ~n5392 ) ;
  assign n30861 = n30860 ^ n5121 ^ 1'b0 ;
  assign n30862 = ~n30859 & n30861 ;
  assign n30863 = n30862 ^ n9829 ^ 1'b0 ;
  assign n30864 = ( n7589 & ~n16556 ) | ( n7589 & n30863 ) | ( ~n16556 & n30863 ) ;
  assign n30865 = n30864 ^ n19742 ^ n19653 ;
  assign n30866 = n3052 & ~n8947 ;
  assign n30867 = n30866 ^ n16321 ^ 1'b0 ;
  assign n30868 = n3766 ^ n2447 ^ 1'b0 ;
  assign n30869 = n30868 ^ n7240 ^ n1770 ;
  assign n30870 = ( n19911 & ~n30867 ) | ( n19911 & n30869 ) | ( ~n30867 & n30869 ) ;
  assign n30871 = n17841 ^ n11188 ^ n2271 ;
  assign n30872 = n30871 ^ n17345 ^ n677 ;
  assign n30873 = n30872 ^ n15987 ^ n3552 ;
  assign n30876 = n1088 | n6781 ;
  assign n30877 = n30876 ^ n2617 ^ 1'b0 ;
  assign n30874 = n1473 | n12361 ;
  assign n30875 = ( n15072 & n15560 ) | ( n15072 & n30874 ) | ( n15560 & n30874 ) ;
  assign n30878 = n30877 ^ n30875 ^ 1'b0 ;
  assign n30879 = ~n30873 & n30878 ;
  assign n30880 = n1611 | n3356 ;
  assign n30881 = n30880 ^ n14026 ^ n12696 ;
  assign n30882 = n16989 ^ n13381 ^ 1'b0 ;
  assign n30883 = ~n4097 & n8933 ;
  assign n30884 = ( n1252 & n4651 ) | ( n1252 & n14381 ) | ( n4651 & n14381 ) ;
  assign n30885 = ( ~x221 & n30883 ) | ( ~x221 & n30884 ) | ( n30883 & n30884 ) ;
  assign n30886 = ( n11071 & n20748 ) | ( n11071 & n30885 ) | ( n20748 & n30885 ) ;
  assign n30887 = n10207 & ~n10730 ;
  assign n30888 = n30886 & n30887 ;
  assign n30889 = n20071 ^ n2433 ^ 1'b0 ;
  assign n30890 = ( n19512 & ~n21054 ) | ( n19512 & n30889 ) | ( ~n21054 & n30889 ) ;
  assign n30898 = ( n3813 & ~n10784 ) | ( n3813 & n19930 ) | ( ~n10784 & n19930 ) ;
  assign n30899 = n30898 ^ n13226 ^ n10356 ;
  assign n30900 = n30899 ^ n18969 ^ 1'b0 ;
  assign n30891 = n19130 ^ n8897 ^ n5952 ;
  assign n30892 = n30891 ^ n8896 ^ 1'b0 ;
  assign n30893 = n13035 | n30892 ;
  assign n30894 = n22487 ^ n21804 ^ n2964 ;
  assign n30895 = n30894 ^ n30660 ^ n17940 ;
  assign n30896 = n30895 ^ n21745 ^ n2510 ;
  assign n30897 = ( n2021 & n30893 ) | ( n2021 & n30896 ) | ( n30893 & n30896 ) ;
  assign n30901 = n30900 ^ n30897 ^ n13849 ;
  assign n30904 = ( n12025 & n13949 ) | ( n12025 & ~n15298 ) | ( n13949 & ~n15298 ) ;
  assign n30903 = n28405 ^ n23850 ^ n4954 ;
  assign n30902 = n14513 ^ n7186 ^ n4006 ;
  assign n30905 = n30904 ^ n30903 ^ n30902 ;
  assign n30906 = n27255 ^ n20370 ^ n2742 ;
  assign n30907 = ( n14305 & n18060 ) | ( n14305 & n30906 ) | ( n18060 & n30906 ) ;
  assign n30908 = ( n825 & ~n4446 ) | ( n825 & n13657 ) | ( ~n4446 & n13657 ) ;
  assign n30909 = n30908 ^ n449 ^ 1'b0 ;
  assign n30910 = n15959 ^ n11139 ^ 1'b0 ;
  assign n30911 = n17312 ^ n10447 ^ n7732 ;
  assign n30912 = ( n20344 & n22701 ) | ( n20344 & n30911 ) | ( n22701 & n30911 ) ;
  assign n30921 = n28777 ^ n4736 ^ n507 ;
  assign n30918 = n27244 ^ n15284 ^ 1'b0 ;
  assign n30919 = n15232 | n30918 ;
  assign n30913 = n30869 ^ n3247 ^ 1'b0 ;
  assign n30914 = n7830 & ~n30913 ;
  assign n30915 = n7705 & ~n30914 ;
  assign n30916 = n13275 | n26389 ;
  assign n30917 = n30915 & ~n30916 ;
  assign n30920 = n30919 ^ n30917 ^ n13554 ;
  assign n30922 = n30921 ^ n30920 ^ n16336 ;
  assign n30923 = n18284 ^ n17592 ^ 1'b0 ;
  assign n30924 = n7062 & ~n30923 ;
  assign n30925 = ~n30922 & n30924 ;
  assign n30926 = n20777 ^ n15691 ^ 1'b0 ;
  assign n30927 = ( n1524 & n30925 ) | ( n1524 & n30926 ) | ( n30925 & n30926 ) ;
  assign n30928 = n26377 ^ n9883 ^ n2680 ;
  assign n30929 = ( ~x168 & n9951 ) | ( ~x168 & n25833 ) | ( n9951 & n25833 ) ;
  assign n30930 = ( ~n5307 & n30928 ) | ( ~n5307 & n30929 ) | ( n30928 & n30929 ) ;
  assign n30931 = ( n1226 & n7130 ) | ( n1226 & n30590 ) | ( n7130 & n30590 ) ;
  assign n30932 = n10986 | n27577 ;
  assign n30933 = n30932 ^ n5547 ^ 1'b0 ;
  assign n30934 = ( ~n25008 & n30931 ) | ( ~n25008 & n30933 ) | ( n30931 & n30933 ) ;
  assign n30935 = ( ~n15642 & n18848 ) | ( ~n15642 & n30934 ) | ( n18848 & n30934 ) ;
  assign n30936 = ~n2643 & n4285 ;
  assign n30937 = ~n5593 & n30936 ;
  assign n30938 = n30937 ^ n16911 ^ 1'b0 ;
  assign n30939 = ( n18889 & n26710 ) | ( n18889 & ~n30938 ) | ( n26710 & ~n30938 ) ;
  assign n30942 = n20685 ^ n19617 ^ 1'b0 ;
  assign n30943 = n20576 & n30942 ;
  assign n30944 = n7572 & n30943 ;
  assign n30940 = n21782 ^ n17230 ^ 1'b0 ;
  assign n30941 = n7002 | n30940 ;
  assign n30945 = n30944 ^ n30941 ^ n11093 ;
  assign n30946 = n4751 & n6977 ;
  assign n30947 = ( n3952 & n26634 ) | ( n3952 & n30946 ) | ( n26634 & n30946 ) ;
  assign n30948 = ( ~n9535 & n9655 ) | ( ~n9535 & n19364 ) | ( n9655 & n19364 ) ;
  assign n30949 = n7845 ^ n2224 ^ 1'b0 ;
  assign n30950 = n12108 & n30949 ;
  assign n30956 = n4723 ^ n1614 ^ 1'b0 ;
  assign n30957 = n30956 ^ n23507 ^ n15533 ;
  assign n30951 = n408 & n14934 ;
  assign n30952 = ~n12687 & n30951 ;
  assign n30953 = ( n4620 & ~n21056 ) | ( n4620 & n30952 ) | ( ~n21056 & n30952 ) ;
  assign n30954 = n26921 & ~n30953 ;
  assign n30955 = ~n24815 & n30954 ;
  assign n30958 = n30957 ^ n30955 ^ n4268 ;
  assign n30962 = ~n6864 & n27732 ;
  assign n30963 = n30962 ^ n14904 ^ 1'b0 ;
  assign n30959 = n8099 ^ n7436 ^ 1'b0 ;
  assign n30960 = n18450 ^ n11284 ^ 1'b0 ;
  assign n30961 = n30959 & ~n30960 ;
  assign n30964 = n30963 ^ n30961 ^ n27916 ;
  assign n30965 = n4112 & ~n5056 ;
  assign n30966 = ~n3096 & n30965 ;
  assign n30967 = ( n3710 & n13331 ) | ( n3710 & ~n30966 ) | ( n13331 & ~n30966 ) ;
  assign n30968 = ( ~n14847 & n20215 ) | ( ~n14847 & n29131 ) | ( n20215 & n29131 ) ;
  assign n30969 = n28227 ^ n15959 ^ n8707 ;
  assign n30975 = n27836 ^ n12210 ^ n5687 ;
  assign n30970 = ( ~n1748 & n5894 ) | ( ~n1748 & n9540 ) | ( n5894 & n9540 ) ;
  assign n30971 = n30970 ^ n2411 ^ 1'b0 ;
  assign n30972 = n30971 ^ n6444 ^ 1'b0 ;
  assign n30973 = ~n1838 & n30972 ;
  assign n30974 = ~n24775 & n30973 ;
  assign n30976 = n30975 ^ n30974 ^ 1'b0 ;
  assign n30977 = n400 | n23516 ;
  assign n30978 = n10660 & ~n30977 ;
  assign n30979 = ( n6124 & ~n20571 ) | ( n6124 & n30978 ) | ( ~n20571 & n30978 ) ;
  assign n30980 = n29136 ^ n25308 ^ n12586 ;
  assign n30981 = ( ~n12310 & n15158 ) | ( ~n12310 & n30980 ) | ( n15158 & n30980 ) ;
  assign n30982 = n21603 ^ n14007 ^ n2581 ;
  assign n30983 = n21351 & n30982 ;
  assign n30984 = n19337 ^ n458 ^ x104 ;
  assign n30985 = ( n14366 & ~n21725 ) | ( n14366 & n30984 ) | ( ~n21725 & n30984 ) ;
  assign n30986 = n17626 & n30985 ;
  assign n30987 = n30986 ^ n2893 ^ 1'b0 ;
  assign n30988 = n30987 ^ n29681 ^ n26779 ;
  assign n30989 = n18996 ^ n8289 ^ n4338 ;
  assign n30990 = n13597 | n16538 ;
  assign n30991 = ( n7632 & n11507 ) | ( n7632 & ~n18436 ) | ( n11507 & ~n18436 ) ;
  assign n30992 = ~n13886 & n30991 ;
  assign n30993 = ( n16812 & n19781 ) | ( n16812 & ~n30992 ) | ( n19781 & ~n30992 ) ;
  assign n30994 = n22433 ^ n19774 ^ n14090 ;
  assign n30995 = n28029 ^ n16072 ^ n9398 ;
  assign n30996 = n20336 ^ n6996 ^ n4100 ;
  assign n30997 = n30996 ^ n14197 ^ n13510 ;
  assign n30998 = ~n474 & n30997 ;
  assign n30999 = n1299 & n30998 ;
  assign n31000 = ~n3948 & n17612 ;
  assign n31001 = n31000 ^ n29345 ^ n24026 ;
  assign n31002 = ( n10804 & n17317 ) | ( n10804 & ~n17363 ) | ( n17317 & ~n17363 ) ;
  assign n31003 = n16094 | n31002 ;
  assign n31004 = ( n6329 & n6585 ) | ( n6329 & n15291 ) | ( n6585 & n15291 ) ;
  assign n31005 = n31004 ^ n12810 ^ n10939 ;
  assign n31006 = x99 | n7757 ;
  assign n31007 = n31006 ^ n18374 ^ 1'b0 ;
  assign n31008 = n10353 ^ n2849 ^ 1'b0 ;
  assign n31009 = ( n3963 & ~n31007 ) | ( n3963 & n31008 ) | ( ~n31007 & n31008 ) ;
  assign n31010 = n24818 ^ n14865 ^ n12107 ;
  assign n31011 = n21632 & n23397 ;
  assign n31012 = n31010 & n31011 ;
  assign n31013 = n6071 & ~n22337 ;
  assign n31014 = n30678 & n31013 ;
  assign n31016 = ~n6272 & n24827 ;
  assign n31015 = n9780 & n15148 ;
  assign n31017 = n31016 ^ n31015 ^ n12438 ;
  assign n31018 = n3219 & n5611 ;
  assign n31019 = n29440 & ~n31018 ;
  assign n31020 = n31019 ^ n29752 ^ 1'b0 ;
  assign n31021 = ( n8298 & n31017 ) | ( n8298 & n31020 ) | ( n31017 & n31020 ) ;
  assign n31022 = n29486 ^ n22091 ^ 1'b0 ;
  assign n31023 = n2535 ^ n635 ^ 1'b0 ;
  assign n31024 = n10915 & ~n31023 ;
  assign n31025 = ( n6774 & n8270 ) | ( n6774 & ~n31024 ) | ( n8270 & ~n31024 ) ;
  assign n31026 = n25787 ^ n11972 ^ n1863 ;
  assign n31027 = n31026 ^ n11131 ^ n5115 ;
  assign n31028 = n11131 ^ n10886 ^ n9150 ;
  assign n31029 = n31028 ^ n11855 ^ 1'b0 ;
  assign n31030 = n1007 & n30924 ;
  assign n31031 = n31029 & ~n31030 ;
  assign n31032 = n14388 | n28355 ;
  assign n31033 = n31032 ^ n15329 ^ 1'b0 ;
  assign n31034 = n31033 ^ n18733 ^ 1'b0 ;
  assign n31035 = n31034 ^ n19296 ^ n3053 ;
  assign n31036 = ( n1001 & n1599 ) | ( n1001 & n11406 ) | ( n1599 & n11406 ) ;
  assign n31037 = n19424 & n31036 ;
  assign n31038 = n6722 ^ n4764 ^ 1'b0 ;
  assign n31039 = ~n3331 & n29204 ;
  assign n31040 = n19304 ^ n17663 ^ n12151 ;
  assign n31041 = ( n8371 & n17762 ) | ( n8371 & ~n23053 ) | ( n17762 & ~n23053 ) ;
  assign n31046 = n13596 & ~n15300 ;
  assign n31047 = ~n21336 & n31046 ;
  assign n31048 = ( ~n7051 & n23678 ) | ( ~n7051 & n31047 ) | ( n23678 & n31047 ) ;
  assign n31042 = ( n2432 & n12739 ) | ( n2432 & n13854 ) | ( n12739 & n13854 ) ;
  assign n31043 = ( x215 & ~n9202 ) | ( x215 & n21377 ) | ( ~n9202 & n21377 ) ;
  assign n31044 = n31042 & ~n31043 ;
  assign n31045 = n2825 & n31044 ;
  assign n31049 = n31048 ^ n31045 ^ n7046 ;
  assign n31050 = n31049 ^ n13823 ^ 1'b0 ;
  assign n31051 = n24737 ^ n14397 ^ n11021 ;
  assign n31052 = n7372 ^ n5951 ^ n705 ;
  assign n31053 = ( n885 & ~n16640 ) | ( n885 & n31052 ) | ( ~n16640 & n31052 ) ;
  assign n31054 = ( n7770 & n28168 ) | ( n7770 & ~n31053 ) | ( n28168 & ~n31053 ) ;
  assign n31055 = n15714 ^ n13776 ^ n991 ;
  assign n31056 = n31055 ^ n19007 ^ n271 ;
  assign n31057 = n6866 & ~n31056 ;
  assign n31058 = n7774 | n16283 ;
  assign n31059 = n31058 ^ n12705 ^ 1'b0 ;
  assign n31060 = ( n15741 & n19041 ) | ( n15741 & ~n24578 ) | ( n19041 & ~n24578 ) ;
  assign n31063 = n16527 ^ n13811 ^ n11160 ;
  assign n31061 = x212 & ~n21981 ;
  assign n31062 = ~n14308 & n31061 ;
  assign n31064 = n31063 ^ n31062 ^ n7676 ;
  assign n31065 = n14795 ^ n12367 ^ n2352 ;
  assign n31066 = n31065 ^ n16459 ^ n6099 ;
  assign n31067 = n4344 ^ n2580 ^ 1'b0 ;
  assign n31068 = n26748 ^ n4257 ^ 1'b0 ;
  assign n31069 = n4616 & n31068 ;
  assign n31070 = n12847 & ~n26505 ;
  assign n31071 = n5562 & ~n20996 ;
  assign n31072 = ( n6921 & ~n11724 ) | ( n6921 & n22132 ) | ( ~n11724 & n22132 ) ;
  assign n31074 = n30340 ^ n26741 ^ x39 ;
  assign n31073 = n12703 ^ n8968 ^ n8611 ;
  assign n31075 = n31074 ^ n31073 ^ 1'b0 ;
  assign n31076 = n31072 & ~n31075 ;
  assign n31081 = n3073 ^ n2157 ^ 1'b0 ;
  assign n31078 = n25942 ^ n6654 ^ 1'b0 ;
  assign n31079 = n1887 | n31078 ;
  assign n31080 = ( ~n2343 & n17106 ) | ( ~n2343 & n31079 ) | ( n17106 & n31079 ) ;
  assign n31077 = ( n6930 & ~n8067 ) | ( n6930 & n25535 ) | ( ~n8067 & n25535 ) ;
  assign n31082 = n31081 ^ n31080 ^ n31077 ;
  assign n31083 = n18010 ^ n1734 ^ 1'b0 ;
  assign n31084 = ( n31076 & n31082 ) | ( n31076 & ~n31083 ) | ( n31082 & ~n31083 ) ;
  assign n31085 = n19429 & n19890 ;
  assign n31086 = n3587 & n12416 ;
  assign n31087 = ~n31085 & n31086 ;
  assign n31088 = n31087 ^ n26835 ^ n5201 ;
  assign n31089 = n23272 ^ n23123 ^ n2363 ;
  assign n31090 = n20105 & n31089 ;
  assign n31091 = n31090 ^ n5711 ^ 1'b0 ;
  assign n31092 = n31091 ^ n24315 ^ n18418 ;
  assign n31093 = n7114 & n26942 ;
  assign n31094 = ~n15565 & n28821 ;
  assign n31095 = ~n1327 & n31094 ;
  assign n31096 = n30709 ^ n25714 ^ n25579 ;
  assign n31097 = n22726 ^ n13100 ^ 1'b0 ;
  assign n31099 = n16249 ^ n5842 ^ n2888 ;
  assign n31100 = n31099 ^ n5918 ^ 1'b0 ;
  assign n31101 = ~n5917 & n31100 ;
  assign n31098 = ( n5802 & ~n13798 ) | ( n5802 & n20193 ) | ( ~n13798 & n20193 ) ;
  assign n31102 = n31101 ^ n31098 ^ n19823 ;
  assign n31103 = n25693 ^ n9218 ^ n2383 ;
  assign n31104 = ( n31097 & ~n31102 ) | ( n31097 & n31103 ) | ( ~n31102 & n31103 ) ;
  assign n31105 = ( n1820 & ~n4212 ) | ( n1820 & n30754 ) | ( ~n4212 & n30754 ) ;
  assign n31106 = n19836 ^ n15247 ^ 1'b0 ;
  assign n31107 = n6241 & ~n14859 ;
  assign n31108 = n31107 ^ n13838 ^ n2883 ;
  assign n31109 = n27632 ^ n20856 ^ n20673 ;
  assign n31111 = n10188 & n25635 ;
  assign n31112 = ( n7700 & ~n19888 ) | ( n7700 & n31111 ) | ( ~n19888 & n31111 ) ;
  assign n31113 = ( n12007 & ~n15145 ) | ( n12007 & n31112 ) | ( ~n15145 & n31112 ) ;
  assign n31110 = n28787 ^ n27890 ^ n15667 ;
  assign n31114 = n31113 ^ n31110 ^ n11242 ;
  assign n31115 = ( n16739 & n31109 ) | ( n16739 & ~n31114 ) | ( n31109 & ~n31114 ) ;
  assign n31116 = n20130 ^ n8492 ^ 1'b0 ;
  assign n31117 = ( n1933 & n11365 ) | ( n1933 & n29446 ) | ( n11365 & n29446 ) ;
  assign n31118 = n13592 ^ n10943 ^ 1'b0 ;
  assign n31119 = n12704 & n31118 ;
  assign n31120 = n22859 & ~n30054 ;
  assign n31121 = ~n20450 & n31120 ;
  assign n31122 = n28734 ^ n15483 ^ n11139 ;
  assign n31123 = ~n2008 & n16905 ;
  assign n31124 = n31123 ^ n20286 ^ 1'b0 ;
  assign n31125 = ( n7849 & n24366 ) | ( n7849 & n31124 ) | ( n24366 & n31124 ) ;
  assign n31126 = ~n13689 & n14719 ;
  assign n31127 = n31126 ^ n10330 ^ 1'b0 ;
  assign n31128 = n31127 ^ n18583 ^ n4470 ;
  assign n31129 = n19639 ^ n4709 ^ 1'b0 ;
  assign n31130 = n490 & n5561 ;
  assign n31131 = n31130 ^ n5823 ^ 1'b0 ;
  assign n31132 = n1691 & n2417 ;
  assign n31133 = n31132 ^ n22003 ^ n12576 ;
  assign n31134 = n31133 ^ n9366 ^ 1'b0 ;
  assign n31136 = ( n1173 & ~n9756 ) | ( n1173 & n19455 ) | ( ~n9756 & n19455 ) ;
  assign n31135 = ( n7306 & n14064 ) | ( n7306 & n28558 ) | ( n14064 & n28558 ) ;
  assign n31137 = n31136 ^ n31135 ^ n20934 ;
  assign n31138 = n9914 | n31137 ;
  assign n31139 = n14771 ^ n1017 ^ 1'b0 ;
  assign n31140 = ( n1516 & n2447 ) | ( n1516 & ~n31139 ) | ( n2447 & ~n31139 ) ;
  assign n31141 = ( n8602 & n9369 ) | ( n8602 & ~n26844 ) | ( n9369 & ~n26844 ) ;
  assign n31142 = n31141 ^ n10846 ^ n2841 ;
  assign n31143 = ~n10154 & n22310 ;
  assign n31144 = n3353 & n22370 ;
  assign n31145 = n7609 & n31144 ;
  assign n31146 = n24148 & ~n31145 ;
  assign n31147 = n12806 ^ n6417 ^ n2105 ;
  assign n31148 = n27547 | n29572 ;
  assign n31149 = ( n2516 & n31147 ) | ( n2516 & n31148 ) | ( n31147 & n31148 ) ;
  assign n31150 = n11587 ^ n7558 ^ n4330 ;
  assign n31151 = ( n5149 & ~n27562 ) | ( n5149 & n31150 ) | ( ~n27562 & n31150 ) ;
  assign n31152 = n847 | n6894 ;
  assign n31153 = n31152 ^ n7050 ^ 1'b0 ;
  assign n31154 = n22349 ^ n9422 ^ 1'b0 ;
  assign n31155 = n31153 & ~n31154 ;
  assign n31156 = n5163 & ~n27404 ;
  assign n31157 = n21989 ^ n20596 ^ n18538 ;
  assign n31158 = n31157 ^ n6428 ^ 1'b0 ;
  assign n31159 = n9186 & n31158 ;
  assign n31160 = n31156 & n31159 ;
  assign n31161 = n31160 ^ n15822 ^ 1'b0 ;
  assign n31162 = n9613 ^ n7928 ^ n3010 ;
  assign n31163 = n705 & ~n3733 ;
  assign n31164 = ~n31162 & n31163 ;
  assign n31165 = ( n10433 & n14790 ) | ( n10433 & ~n15324 ) | ( n14790 & ~n15324 ) ;
  assign n31166 = ( n1141 & n10381 ) | ( n1141 & n31165 ) | ( n10381 & n31165 ) ;
  assign n31167 = n13754 ^ n1006 ^ 1'b0 ;
  assign n31168 = n3704 | n31167 ;
  assign n31169 = n27645 ^ n24179 ^ 1'b0 ;
  assign n31170 = n15926 ^ n15470 ^ n9118 ;
  assign n31171 = n31170 ^ n26550 ^ n20581 ;
  assign n31172 = ~n2767 & n28453 ;
  assign n31173 = n3929 & n31172 ;
  assign n31174 = ( n7672 & ~n9371 ) | ( n7672 & n31173 ) | ( ~n9371 & n31173 ) ;
  assign n31175 = n31174 ^ n30319 ^ n2670 ;
  assign n31176 = ( n31169 & n31171 ) | ( n31169 & ~n31175 ) | ( n31171 & ~n31175 ) ;
  assign n31178 = ( n6160 & n14533 ) | ( n6160 & ~n23914 ) | ( n14533 & ~n23914 ) ;
  assign n31177 = n17713 ^ n3620 ^ 1'b0 ;
  assign n31179 = n31178 ^ n31177 ^ 1'b0 ;
  assign n31180 = n18285 ^ n14152 ^ 1'b0 ;
  assign n31181 = n19850 | n20329 ;
  assign n31182 = n21055 & ~n31181 ;
  assign n31183 = n18996 & n19853 ;
  assign n31184 = n19679 ^ n16242 ^ n11139 ;
  assign n31185 = n31184 ^ n24444 ^ n4924 ;
  assign n31186 = n27207 ^ n23413 ^ 1'b0 ;
  assign n31187 = n13441 & n31186 ;
  assign n31188 = n31187 ^ n12841 ^ 1'b0 ;
  assign n31189 = n473 | n3502 ;
  assign n31190 = ~n5883 & n31189 ;
  assign n31191 = n15164 ^ n13274 ^ 1'b0 ;
  assign n31192 = n17093 ^ n2151 ^ 1'b0 ;
  assign n31193 = ( n1510 & n31191 ) | ( n1510 & n31192 ) | ( n31191 & n31192 ) ;
  assign n31194 = ( n19477 & n19815 ) | ( n19477 & n31193 ) | ( n19815 & n31193 ) ;
  assign n31195 = n24687 & ~n31194 ;
  assign n31196 = n31195 ^ n18185 ^ 1'b0 ;
  assign n31197 = n6394 & ~n9804 ;
  assign n31198 = n8540 & n31197 ;
  assign n31199 = n31198 ^ n5503 ^ 1'b0 ;
  assign n31200 = n18159 ^ n9324 ^ 1'b0 ;
  assign n31201 = ~n18767 & n31200 ;
  assign n31202 = ( n333 & n18397 ) | ( n333 & ~n31201 ) | ( n18397 & ~n31201 ) ;
  assign n31203 = ( ~n13738 & n26624 ) | ( ~n13738 & n31202 ) | ( n26624 & n31202 ) ;
  assign n31204 = n28395 ^ n7113 ^ 1'b0 ;
  assign n31205 = n15659 ^ n3771 ^ 1'b0 ;
  assign n31206 = ( ~n18549 & n31150 ) | ( ~n18549 & n31205 ) | ( n31150 & n31205 ) ;
  assign n31207 = ( n5924 & n12345 ) | ( n5924 & ~n20596 ) | ( n12345 & ~n20596 ) ;
  assign n31208 = ~n16304 & n31207 ;
  assign n31209 = n23807 ^ n13321 ^ 1'b0 ;
  assign n31210 = n11208 | n31209 ;
  assign n31211 = n12103 ^ x214 ^ x177 ;
  assign n31212 = n31211 ^ n14057 ^ n13875 ;
  assign n31213 = n2836 & n9308 ;
  assign n31214 = n31213 ^ n30436 ^ n16931 ;
  assign n31215 = n27135 ^ n8752 ^ 1'b0 ;
  assign n31216 = ( n18198 & n31214 ) | ( n18198 & n31215 ) | ( n31214 & n31215 ) ;
  assign n31217 = ( n4525 & n11149 ) | ( n4525 & ~n16378 ) | ( n11149 & ~n16378 ) ;
  assign n31218 = ( n4216 & ~n23440 ) | ( n4216 & n31217 ) | ( ~n23440 & n31217 ) ;
  assign n31219 = ( n10020 & n16300 ) | ( n10020 & n31218 ) | ( n16300 & n31218 ) ;
  assign n31220 = n11529 ^ n622 ^ 1'b0 ;
  assign n31221 = n18672 ^ n5753 ^ 1'b0 ;
  assign n31222 = ( n29288 & n31220 ) | ( n29288 & ~n31221 ) | ( n31220 & ~n31221 ) ;
  assign n31223 = n31222 ^ n3045 ^ 1'b0 ;
  assign n31224 = n31223 ^ n19626 ^ 1'b0 ;
  assign n31225 = n22974 & ~n31224 ;
  assign n31226 = ~n12535 & n31225 ;
  assign n31227 = n17437 ^ n12470 ^ 1'b0 ;
  assign n31228 = n14286 & n31227 ;
  assign n31229 = ( n3431 & ~n15835 ) | ( n3431 & n28410 ) | ( ~n15835 & n28410 ) ;
  assign n31230 = n31229 ^ n8327 ^ n1026 ;
  assign n31231 = n5534 ^ n1196 ^ 1'b0 ;
  assign n31232 = ~n27046 & n31231 ;
  assign n31233 = n29241 & n31232 ;
  assign n31234 = n21451 & n31233 ;
  assign n31241 = ( n2068 & n10352 ) | ( n2068 & ~n26188 ) | ( n10352 & ~n26188 ) ;
  assign n31237 = n3966 | n6179 ;
  assign n31238 = n18819 ^ n17101 ^ 1'b0 ;
  assign n31239 = n31237 | n31238 ;
  assign n31236 = n28239 ^ n6621 ^ 1'b0 ;
  assign n31240 = n31239 ^ n31236 ^ n28915 ;
  assign n31242 = n31241 ^ n31240 ^ n1146 ;
  assign n31235 = n22892 | n25008 ;
  assign n31243 = n31242 ^ n31235 ^ 1'b0 ;
  assign n31244 = n1476 & ~n21496 ;
  assign n31245 = n31244 ^ n28027 ^ 1'b0 ;
  assign n31246 = ~n21264 & n31245 ;
  assign n31247 = n31246 ^ n27142 ^ 1'b0 ;
  assign n31248 = ( n3651 & n7808 ) | ( n3651 & ~n22017 ) | ( n7808 & ~n22017 ) ;
  assign n31249 = n31248 ^ n22182 ^ n3271 ;
  assign n31250 = n6557 ^ n4306 ^ n2710 ;
  assign n31251 = ( n17600 & n28760 ) | ( n17600 & n31250 ) | ( n28760 & n31250 ) ;
  assign n31252 = n345 | n12282 ;
  assign n31253 = x126 ^ x108 ^ 1'b0 ;
  assign n31254 = ~n3483 & n31253 ;
  assign n31255 = n31254 ^ n10745 ^ n8632 ;
  assign n31257 = n2510 ^ n1064 ^ 1'b0 ;
  assign n31258 = n2849 & n31257 ;
  assign n31259 = n31258 ^ n5904 ^ 1'b0 ;
  assign n31256 = ( n6951 & ~n7207 ) | ( n6951 & n9911 ) | ( ~n7207 & n9911 ) ;
  assign n31260 = n31259 ^ n31256 ^ n21306 ;
  assign n31261 = ( ~n3244 & n31255 ) | ( ~n3244 & n31260 ) | ( n31255 & n31260 ) ;
  assign n31262 = ( ~n2019 & n3221 ) | ( ~n2019 & n25752 ) | ( n3221 & n25752 ) ;
  assign n31263 = ~n7842 & n31262 ;
  assign n31264 = n31263 ^ n17427 ^ 1'b0 ;
  assign n31265 = n10272 ^ n8930 ^ 1'b0 ;
  assign n31266 = n18400 & n31265 ;
  assign n31267 = n3150 ^ n1663 ^ 1'b0 ;
  assign n31268 = n30148 | n31267 ;
  assign n31275 = ( ~n2057 & n7332 ) | ( ~n2057 & n15299 ) | ( n7332 & n15299 ) ;
  assign n31276 = n17513 & ~n31275 ;
  assign n31277 = n31276 ^ n7643 ^ 1'b0 ;
  assign n31278 = n31277 ^ n9949 ^ n1408 ;
  assign n31272 = n3460 ^ n2807 ^ 1'b0 ;
  assign n31269 = n13824 ^ n10725 ^ 1'b0 ;
  assign n31270 = n11252 & n12577 ;
  assign n31271 = n31269 & n31270 ;
  assign n31273 = n31272 ^ n31271 ^ n6029 ;
  assign n31274 = n31273 ^ n24202 ^ n7659 ;
  assign n31279 = n31278 ^ n31274 ^ n12644 ;
  assign n31280 = ( ~n4834 & n15146 ) | ( ~n4834 & n18289 ) | ( n15146 & n18289 ) ;
  assign n31281 = ( n12481 & n20444 ) | ( n12481 & ~n31280 ) | ( n20444 & ~n31280 ) ;
  assign n31282 = n31281 ^ n9709 ^ n4404 ;
  assign n31283 = ( n6240 & n12563 ) | ( n6240 & ~n24492 ) | ( n12563 & ~n24492 ) ;
  assign n31284 = n18729 ^ n15959 ^ 1'b0 ;
  assign n31285 = n31283 & n31284 ;
  assign n31286 = n29842 ^ n5831 ^ n3355 ;
  assign n31287 = n1610 | n28161 ;
  assign n31288 = n31287 ^ n17364 ^ 1'b0 ;
  assign n31289 = n31288 ^ n7860 ^ 1'b0 ;
  assign n31290 = n28580 ^ n15825 ^ n7550 ;
  assign n31291 = n31290 ^ n17062 ^ n7739 ;
  assign n31292 = n16266 & n31291 ;
  assign n31293 = n17170 ^ n12048 ^ n4899 ;
  assign n31294 = n31293 ^ n23871 ^ n18563 ;
  assign n31295 = ( n4221 & n11553 ) | ( n4221 & n19119 ) | ( n11553 & n19119 ) ;
  assign n31296 = ~n13554 & n14621 ;
  assign n31297 = n8578 & n31296 ;
  assign n31298 = ( ~n2499 & n9074 ) | ( ~n2499 & n10415 ) | ( n9074 & n10415 ) ;
  assign n31299 = ( n376 & ~n31297 ) | ( n376 & n31298 ) | ( ~n31297 & n31298 ) ;
  assign n31301 = ( ~n842 & n3528 ) | ( ~n842 & n9294 ) | ( n3528 & n9294 ) ;
  assign n31302 = ( n11180 & n21110 ) | ( n11180 & ~n24252 ) | ( n21110 & ~n24252 ) ;
  assign n31303 = n31301 & n31302 ;
  assign n31300 = ~n12987 & n15128 ;
  assign n31304 = n31303 ^ n31300 ^ n18663 ;
  assign n31305 = n13456 & n25690 ;
  assign n31306 = n914 & n31305 ;
  assign n31307 = n25215 ^ n3141 ^ 1'b0 ;
  assign n31308 = n17398 | n31307 ;
  assign n31309 = n8881 & n24203 ;
  assign n31311 = n13982 ^ n8117 ^ n2251 ;
  assign n31310 = ( n12850 & n12887 ) | ( n12850 & ~n13273 ) | ( n12887 & ~n13273 ) ;
  assign n31312 = n31311 ^ n31310 ^ n19479 ;
  assign n31313 = n20226 & ~n20899 ;
  assign n31314 = ( ~n3393 & n21209 ) | ( ~n3393 & n31313 ) | ( n21209 & n31313 ) ;
  assign n31315 = n23664 ^ n13759 ^ n13027 ;
  assign n31316 = ( n5221 & ~n7693 ) | ( n5221 & n31315 ) | ( ~n7693 & n31315 ) ;
  assign n31317 = ( n12107 & n31097 ) | ( n12107 & n31316 ) | ( n31097 & n31316 ) ;
  assign n31319 = ~n7789 & n11081 ;
  assign n31320 = n31319 ^ n20540 ^ 1'b0 ;
  assign n31318 = ( n7946 & ~n15581 ) | ( n7946 & n20588 ) | ( ~n15581 & n20588 ) ;
  assign n31321 = n31320 ^ n31318 ^ n26911 ;
  assign n31322 = n15502 | n27593 ;
  assign n31323 = n31322 ^ n5490 ^ 1'b0 ;
  assign n31324 = n27437 & n31323 ;
  assign n31325 = ~n27255 & n31324 ;
  assign n31326 = n25780 ^ n1596 ^ 1'b0 ;
  assign n31327 = n17200 ^ n11151 ^ 1'b0 ;
  assign n31328 = n1711 & ~n31327 ;
  assign n31329 = n29636 | n31328 ;
  assign n31330 = n6918 & ~n31329 ;
  assign n31331 = ~n31326 & n31330 ;
  assign n31332 = n579 & ~n12390 ;
  assign n31333 = ( n4971 & n14976 ) | ( n4971 & ~n31332 ) | ( n14976 & ~n31332 ) ;
  assign n31334 = ( n2051 & n10800 ) | ( n2051 & n31202 ) | ( n10800 & n31202 ) ;
  assign n31335 = ( n7829 & ~n8428 ) | ( n7829 & n31334 ) | ( ~n8428 & n31334 ) ;
  assign n31336 = n10486 ^ n9594 ^ 1'b0 ;
  assign n31337 = n5323 & n31336 ;
  assign n31338 = ( n5415 & ~n27618 ) | ( n5415 & n31337 ) | ( ~n27618 & n31337 ) ;
  assign n31339 = n7635 ^ n2550 ^ 1'b0 ;
  assign n31340 = ~n961 & n31339 ;
  assign n31341 = n31340 ^ n6919 ^ x67 ;
  assign n31342 = n27352 & ~n31341 ;
  assign n31343 = ~n31338 & n31342 ;
  assign n31344 = n346 & ~n21053 ;
  assign n31345 = n13945 & n31344 ;
  assign n31346 = n11870 ^ n1130 ^ 1'b0 ;
  assign n31347 = n11053 ^ n7471 ^ n5318 ;
  assign n31348 = ( n7628 & n31346 ) | ( n7628 & n31347 ) | ( n31346 & n31347 ) ;
  assign n31349 = n31348 ^ n12930 ^ n9385 ;
  assign n31350 = ( x211 & ~n31345 ) | ( x211 & n31349 ) | ( ~n31345 & n31349 ) ;
  assign n31351 = ( n2835 & n31343 ) | ( n2835 & n31350 ) | ( n31343 & n31350 ) ;
  assign n31352 = n31137 ^ n30516 ^ n15956 ;
  assign n31353 = ( ~n3097 & n16825 ) | ( ~n3097 & n20486 ) | ( n16825 & n20486 ) ;
  assign n31354 = ( n2904 & n4314 ) | ( n2904 & ~n26047 ) | ( n4314 & ~n26047 ) ;
  assign n31355 = n16918 ^ n15517 ^ n8777 ;
  assign n31356 = ( n11312 & n15187 ) | ( n11312 & n16332 ) | ( n15187 & n16332 ) ;
  assign n31357 = ( ~n31354 & n31355 ) | ( ~n31354 & n31356 ) | ( n31355 & n31356 ) ;
  assign n31358 = ( n5389 & n28808 ) | ( n5389 & ~n31357 ) | ( n28808 & ~n31357 ) ;
  assign n31359 = n7566 ^ n1090 ^ 1'b0 ;
  assign n31360 = n31359 ^ n28580 ^ n15113 ;
  assign n31361 = n31360 ^ n28974 ^ n8008 ;
  assign n31362 = ( n6642 & n11479 ) | ( n6642 & n23085 ) | ( n11479 & n23085 ) ;
  assign n31363 = ( n11804 & n22086 ) | ( n11804 & ~n31362 ) | ( n22086 & ~n31362 ) ;
  assign n31364 = n5575 | n31363 ;
  assign n31368 = n24697 ^ n7573 ^ n3327 ;
  assign n31366 = n6475 ^ n5592 ^ n902 ;
  assign n31365 = ( n341 & ~n865 ) | ( n341 & n2400 ) | ( ~n865 & n2400 ) ;
  assign n31367 = n31366 ^ n31365 ^ 1'b0 ;
  assign n31369 = n31368 ^ n31367 ^ n20005 ;
  assign n31370 = ( n8488 & n16381 ) | ( n8488 & ~n23744 ) | ( n16381 & ~n23744 ) ;
  assign n31371 = n2877 & n16569 ;
  assign n31372 = ( n8327 & n16083 ) | ( n8327 & n28375 ) | ( n16083 & n28375 ) ;
  assign n31373 = n31372 ^ n7633 ^ x138 ;
  assign n31374 = ( n7885 & n9123 ) | ( n7885 & ~n28963 ) | ( n9123 & ~n28963 ) ;
  assign n31375 = n31374 ^ n15277 ^ n11800 ;
  assign n31376 = n7640 & n15725 ;
  assign n31377 = ~n17157 & n31376 ;
  assign n31378 = n2955 ^ n1752 ^ 1'b0 ;
  assign n31379 = n29493 | n31378 ;
  assign n31380 = ( n2199 & n23095 ) | ( n2199 & ~n26109 ) | ( n23095 & ~n26109 ) ;
  assign n31381 = ( n6040 & ~n16170 ) | ( n6040 & n22106 ) | ( ~n16170 & n22106 ) ;
  assign n31382 = n14544 ^ n11603 ^ 1'b0 ;
  assign n31383 = ( ~n2997 & n21456 ) | ( ~n2997 & n31382 ) | ( n21456 & n31382 ) ;
  assign n31388 = n9704 ^ n8528 ^ n3750 ;
  assign n31389 = n31388 ^ n12790 ^ n9964 ;
  assign n31384 = n18395 ^ n10644 ^ n6912 ;
  assign n31385 = n18258 | n31384 ;
  assign n31386 = n8895 | n31385 ;
  assign n31387 = ~n7480 & n31386 ;
  assign n31390 = n31389 ^ n31387 ^ 1'b0 ;
  assign n31391 = ( n30302 & n31383 ) | ( n30302 & ~n31390 ) | ( n31383 & ~n31390 ) ;
  assign n31392 = n28729 ^ n25079 ^ 1'b0 ;
  assign n31394 = n12037 ^ n5958 ^ n1672 ;
  assign n31393 = ( ~x22 & n4442 ) | ( ~x22 & n25244 ) | ( n4442 & n25244 ) ;
  assign n31395 = n31394 ^ n31393 ^ n28524 ;
  assign n31396 = ( n4296 & n5965 ) | ( n4296 & ~n8085 ) | ( n5965 & ~n8085 ) ;
  assign n31397 = n31396 ^ n11477 ^ n10112 ;
  assign n31398 = n7919 | n31397 ;
  assign n31399 = n983 | n14727 ;
  assign n31400 = n4984 & ~n30880 ;
  assign n31401 = ( n3981 & n24957 ) | ( n3981 & n31400 ) | ( n24957 & n31400 ) ;
  assign n31402 = n17966 & n31401 ;
  assign n31403 = n31399 & n31402 ;
  assign n31404 = n24521 | n26327 ;
  assign n31405 = ( n6699 & ~n9763 ) | ( n6699 & n14439 ) | ( ~n9763 & n14439 ) ;
  assign n31406 = n31405 ^ n22345 ^ n17822 ;
  assign n31407 = ( n3784 & ~n7297 ) | ( n3784 & n27924 ) | ( ~n7297 & n27924 ) ;
  assign n31408 = ( ~n31404 & n31406 ) | ( ~n31404 & n31407 ) | ( n31406 & n31407 ) ;
  assign n31409 = n5367 | n12031 ;
  assign n31410 = n4732 | n31409 ;
  assign n31411 = ( ~n18844 & n27167 ) | ( ~n18844 & n31410 ) | ( n27167 & n31410 ) ;
  assign n31412 = n26335 ^ n15858 ^ 1'b0 ;
  assign n31415 = n1200 | n12119 ;
  assign n31413 = n9706 & n17798 ;
  assign n31414 = ~n7914 & n31413 ;
  assign n31416 = n31415 ^ n31414 ^ n7944 ;
  assign n31417 = n4509 & n31416 ;
  assign n31418 = n6441 & n31417 ;
  assign n31419 = n27577 ^ n14482 ^ 1'b0 ;
  assign n31420 = ~n9003 & n31419 ;
  assign n31421 = n7088 ^ n3050 ^ 1'b0 ;
  assign n31422 = n24581 ^ n6164 ^ n2558 ;
  assign n31423 = ( n8874 & ~n18239 ) | ( n8874 & n24628 ) | ( ~n18239 & n24628 ) ;
  assign n31424 = n4204 & ~n31423 ;
  assign n31425 = ~n31422 & n31424 ;
  assign n31427 = n18834 ^ n5179 ^ 1'b0 ;
  assign n31428 = n3525 & ~n31427 ;
  assign n31429 = n30275 & n31428 ;
  assign n31430 = n31429 ^ n5847 ^ 1'b0 ;
  assign n31426 = n24083 ^ n19082 ^ n1500 ;
  assign n31431 = n31430 ^ n31426 ^ 1'b0 ;
  assign n31432 = n26571 ^ n3776 ^ 1'b0 ;
  assign n31433 = n15288 & n31432 ;
  assign n31434 = n21262 & n31433 ;
  assign n31435 = n12777 & n31434 ;
  assign n31436 = n9642 ^ n3125 ^ n3099 ;
  assign n31437 = ( n6670 & n31435 ) | ( n6670 & ~n31436 ) | ( n31435 & ~n31436 ) ;
  assign n31438 = n6280 & ~n22765 ;
  assign n31439 = x33 & ~n12281 ;
  assign n31440 = n31439 ^ n25738 ^ 1'b0 ;
  assign n31441 = n31440 ^ n12020 ^ 1'b0 ;
  assign n31442 = n31441 ^ n30026 ^ n17839 ;
  assign n31443 = ( n4152 & ~n13092 ) | ( n4152 & n31442 ) | ( ~n13092 & n31442 ) ;
  assign n31444 = n4919 | n15049 ;
  assign n31445 = n4830 & n7862 ;
  assign n31446 = ~n31444 & n31445 ;
  assign n31447 = n31446 ^ n18978 ^ 1'b0 ;
  assign n31448 = n5613 & ~n26361 ;
  assign n31449 = n31448 ^ n20542 ^ n12815 ;
  assign n31450 = n26965 ^ n24476 ^ n14888 ;
  assign n31451 = n15076 ^ n10899 ^ n10560 ;
  assign n31452 = n31451 ^ n9778 ^ 1'b0 ;
  assign n31453 = n12940 & ~n31452 ;
  assign n31454 = n29097 & n31453 ;
  assign n31455 = n5712 & n12477 ;
  assign n31456 = n13796 | n31455 ;
  assign n31457 = n23660 & ~n31456 ;
  assign n31458 = n2175 & ~n13916 ;
  assign n31459 = ~n23637 & n31458 ;
  assign n31460 = n8401 & ~n27652 ;
  assign n31461 = n31460 ^ n15442 ^ n12724 ;
  assign n31462 = ( n4506 & n15852 ) | ( n4506 & n23225 ) | ( n15852 & n23225 ) ;
  assign n31463 = n31462 ^ n19300 ^ n8239 ;
  assign n31464 = n17437 & n21668 ;
  assign n31465 = n7444 & n31464 ;
  assign n31466 = ( ~n16121 & n30173 ) | ( ~n16121 & n31465 ) | ( n30173 & n31465 ) ;
  assign n31467 = n7288 & n16457 ;
  assign n31468 = n15382 | n31467 ;
  assign n31469 = n31468 ^ n11905 ^ 1'b0 ;
  assign n31470 = ( n6887 & n9104 ) | ( n6887 & n12241 ) | ( n9104 & n12241 ) ;
  assign n31471 = n16637 | n19637 ;
  assign n31472 = n26322 & ~n31471 ;
  assign n31473 = ( ~n14384 & n31470 ) | ( ~n14384 & n31472 ) | ( n31470 & n31472 ) ;
  assign n31474 = n30106 ^ n28243 ^ n18990 ;
  assign n31475 = n18141 ^ n16726 ^ 1'b0 ;
  assign n31476 = n11503 ^ n9705 ^ 1'b0 ;
  assign n31477 = n12708 & ~n31476 ;
  assign n31478 = n31477 ^ n20745 ^ n13976 ;
  assign n31480 = n21957 ^ n15491 ^ n3786 ;
  assign n31479 = ~n29974 & n31131 ;
  assign n31481 = n31480 ^ n31479 ^ 1'b0 ;
  assign n31485 = n11679 & ~n15990 ;
  assign n31482 = n14823 ^ n4731 ^ n4463 ;
  assign n31483 = ( ~n19884 & n26525 ) | ( ~n19884 & n31482 ) | ( n26525 & n31482 ) ;
  assign n31484 = n10553 & n31483 ;
  assign n31486 = n31485 ^ n31484 ^ n5006 ;
  assign n31487 = n31486 ^ n20027 ^ 1'b0 ;
  assign n31488 = n11092 & ~n31487 ;
  assign n31489 = n10508 ^ n1903 ^ 1'b0 ;
  assign n31490 = n31489 ^ n13418 ^ 1'b0 ;
  assign n31491 = ( ~n10605 & n22675 ) | ( ~n10605 & n26093 ) | ( n22675 & n26093 ) ;
  assign n31492 = n3389 & ~n25344 ;
  assign n31493 = ~n18029 & n31492 ;
  assign n31494 = ( x112 & ~n1162 ) | ( x112 & n2417 ) | ( ~n1162 & n2417 ) ;
  assign n31495 = ( x249 & n19390 ) | ( x249 & ~n29182 ) | ( n19390 & ~n29182 ) ;
  assign n31496 = ( n22290 & n29682 ) | ( n22290 & n31495 ) | ( n29682 & n31495 ) ;
  assign n31497 = ( ~n23135 & n31494 ) | ( ~n23135 & n31496 ) | ( n31494 & n31496 ) ;
  assign n31498 = ( n1555 & n2107 ) | ( n1555 & ~n2264 ) | ( n2107 & ~n2264 ) ;
  assign n31499 = n22142 | n31498 ;
  assign n31500 = n31499 ^ n7687 ^ 1'b0 ;
  assign n31510 = n16382 ^ n8946 ^ n4257 ;
  assign n31511 = n30570 & n31510 ;
  assign n31512 = ~n21191 & n31511 ;
  assign n31508 = n30959 ^ n16378 ^ n5750 ;
  assign n31506 = n19579 ^ n12880 ^ 1'b0 ;
  assign n31507 = ~n20870 & n31506 ;
  assign n31501 = n22330 ^ n13603 ^ 1'b0 ;
  assign n31502 = n7546 & n31501 ;
  assign n31503 = ( n3799 & n5037 ) | ( n3799 & n15365 ) | ( n5037 & n15365 ) ;
  assign n31504 = n31503 ^ n25420 ^ n5189 ;
  assign n31505 = ( n8384 & ~n31502 ) | ( n8384 & n31504 ) | ( ~n31502 & n31504 ) ;
  assign n31509 = n31508 ^ n31507 ^ n31505 ;
  assign n31513 = n31512 ^ n31509 ^ n6120 ;
  assign n31514 = ( n8318 & n21497 ) | ( n8318 & n31150 ) | ( n21497 & n31150 ) ;
  assign n31515 = n1513 | n22418 ;
  assign n31516 = n13452 | n17617 ;
  assign n31517 = n31516 ^ n1883 ^ 1'b0 ;
  assign n31518 = n3097 & n15362 ;
  assign n31519 = n31518 ^ n11622 ^ 1'b0 ;
  assign n31522 = n24202 ^ n9168 ^ n7423 ;
  assign n31523 = n2768 & n31522 ;
  assign n31524 = ~n29518 & n31523 ;
  assign n31520 = n7589 & n16664 ;
  assign n31521 = ~n11793 & n31520 ;
  assign n31525 = n31524 ^ n31521 ^ n7315 ;
  assign n31526 = ( n14986 & n18087 ) | ( n14986 & n31290 ) | ( n18087 & n31290 ) ;
  assign n31527 = ( n6046 & ~n8903 ) | ( n6046 & n10700 ) | ( ~n8903 & n10700 ) ;
  assign n31529 = ( ~n17325 & n21870 ) | ( ~n17325 & n22653 ) | ( n21870 & n22653 ) ;
  assign n31528 = n2843 & n4566 ;
  assign n31530 = n31529 ^ n31528 ^ 1'b0 ;
  assign n31531 = ( n29925 & n31527 ) | ( n29925 & ~n31530 ) | ( n31527 & ~n31530 ) ;
  assign n31532 = n5976 & ~n18583 ;
  assign n31533 = n31532 ^ n1391 ^ 1'b0 ;
  assign n31539 = ( n3005 & n6725 ) | ( n3005 & n11938 ) | ( n6725 & n11938 ) ;
  assign n31540 = n19853 | n31539 ;
  assign n31541 = n2050 & ~n13270 ;
  assign n31542 = n31541 ^ n22154 ^ 1'b0 ;
  assign n31543 = ( ~n953 & n31540 ) | ( ~n953 & n31542 ) | ( n31540 & n31542 ) ;
  assign n31534 = n10152 ^ n7729 ^ n5104 ;
  assign n31535 = ( ~n1047 & n1907 ) | ( ~n1047 & n12843 ) | ( n1907 & n12843 ) ;
  assign n31536 = n7169 & n10296 ;
  assign n31537 = ( n31534 & ~n31535 ) | ( n31534 & n31536 ) | ( ~n31535 & n31536 ) ;
  assign n31538 = n25252 & n31537 ;
  assign n31544 = n31543 ^ n31538 ^ 1'b0 ;
  assign n31553 = ( n3688 & n6543 ) | ( n3688 & n17462 ) | ( n6543 & n17462 ) ;
  assign n31549 = n2751 ^ n2559 ^ 1'b0 ;
  assign n31550 = n31549 ^ n16133 ^ n10818 ;
  assign n31551 = n10513 | n31550 ;
  assign n31552 = ( n16731 & n21788 ) | ( n16731 & ~n31551 ) | ( n21788 & ~n31551 ) ;
  assign n31554 = n31553 ^ n31552 ^ n19231 ;
  assign n31545 = ( n14236 & n22737 ) | ( n14236 & n28032 ) | ( n22737 & n28032 ) ;
  assign n31546 = n31545 ^ n17211 ^ 1'b0 ;
  assign n31547 = n6110 | n31546 ;
  assign n31548 = n7706 & ~n31547 ;
  assign n31555 = n31554 ^ n31548 ^ 1'b0 ;
  assign n31556 = n13321 ^ n3291 ^ n2199 ;
  assign n31557 = n31556 ^ n19854 ^ n13370 ;
  assign n31558 = n31394 & ~n31557 ;
  assign n31559 = n30563 ^ n27940 ^ n21291 ;
  assign n31560 = n31559 ^ n17812 ^ n13948 ;
  assign n31561 = n18397 ^ n14693 ^ n8122 ;
  assign n31562 = n31561 ^ n7592 ^ n3858 ;
  assign n31563 = n14094 | n31562 ;
  assign n31564 = n30684 ^ n19706 ^ 1'b0 ;
  assign n31565 = n3308 & ~n31564 ;
  assign n31568 = n11563 ^ n7540 ^ 1'b0 ;
  assign n31566 = n8639 ^ n8347 ^ 1'b0 ;
  assign n31567 = n31566 ^ n7743 ^ n5407 ;
  assign n31569 = n31568 ^ n31567 ^ n9312 ;
  assign n31570 = n12329 ^ n10761 ^ 1'b0 ;
  assign n31571 = ~n15108 & n31570 ;
  assign n31572 = ( ~n22824 & n31569 ) | ( ~n22824 & n31571 ) | ( n31569 & n31571 ) ;
  assign n31573 = n4924 & n6645 ;
  assign n31574 = n31573 ^ n3912 ^ 1'b0 ;
  assign n31575 = n31574 ^ n18658 ^ 1'b0 ;
  assign n31576 = ~n31572 & n31575 ;
  assign n31577 = ( ~n9918 & n10448 ) | ( ~n9918 & n19546 ) | ( n10448 & n19546 ) ;
  assign n31578 = n18491 ^ n7378 ^ 1'b0 ;
  assign n31579 = ~n24768 & n31578 ;
  assign n31580 = n31579 ^ n9602 ^ n3926 ;
  assign n31581 = ( n7029 & n15444 ) | ( n7029 & n17690 ) | ( n15444 & n17690 ) ;
  assign n31582 = ( ~n31577 & n31580 ) | ( ~n31577 & n31581 ) | ( n31580 & n31581 ) ;
  assign n31583 = ( n15566 & n20597 ) | ( n15566 & ~n29539 ) | ( n20597 & ~n29539 ) ;
  assign n31584 = ( ~n10801 & n20504 ) | ( ~n10801 & n30862 ) | ( n20504 & n30862 ) ;
  assign n31585 = ( ~n13169 & n28239 ) | ( ~n13169 & n30384 ) | ( n28239 & n30384 ) ;
  assign n31586 = n17265 ^ n1448 ^ 1'b0 ;
  assign n31587 = n25809 & ~n31586 ;
  assign n31588 = ( n5394 & n7103 ) | ( n5394 & ~n31587 ) | ( n7103 & ~n31587 ) ;
  assign n31589 = n5495 ^ n4130 ^ 1'b0 ;
  assign n31592 = n3853 & ~n7283 ;
  assign n31593 = ~n10716 & n31592 ;
  assign n31590 = n553 | n3895 ;
  assign n31591 = n31590 ^ n30446 ^ n13197 ;
  assign n31594 = n31593 ^ n31591 ^ n27740 ;
  assign n31595 = n31589 & n31594 ;
  assign n31596 = n31588 & n31595 ;
  assign n31597 = ~n18821 & n20645 ;
  assign n31598 = n31597 ^ n16896 ^ 1'b0 ;
  assign n31599 = n31598 ^ n8146 ^ 1'b0 ;
  assign n31600 = n7013 & ~n31599 ;
  assign n31601 = n21271 ^ n649 ^ 1'b0 ;
  assign n31602 = ( n9246 & n15327 ) | ( n9246 & n16573 ) | ( n15327 & n16573 ) ;
  assign n31603 = ( ~n2357 & n10473 ) | ( ~n2357 & n14837 ) | ( n10473 & n14837 ) ;
  assign n31604 = ( ~n20946 & n31602 ) | ( ~n20946 & n31603 ) | ( n31602 & n31603 ) ;
  assign n31605 = ( n8196 & ~n14232 ) | ( n8196 & n15187 ) | ( ~n14232 & n15187 ) ;
  assign n31606 = n12491 | n20616 ;
  assign n31607 = n31605 & ~n31606 ;
  assign n31608 = ( ~n9138 & n31604 ) | ( ~n9138 & n31607 ) | ( n31604 & n31607 ) ;
  assign n31609 = ( n9589 & ~n16130 ) | ( n9589 & n17421 ) | ( ~n16130 & n17421 ) ;
  assign n31615 = ~n2593 & n7843 ;
  assign n31616 = n31615 ^ n7542 ^ 1'b0 ;
  assign n31610 = n3717 ^ n575 ^ 1'b0 ;
  assign n31611 = n7759 | n31610 ;
  assign n31612 = n31611 ^ n17393 ^ n3530 ;
  assign n31613 = n8342 & n31612 ;
  assign n31614 = ~n4454 & n31613 ;
  assign n31617 = n31616 ^ n31614 ^ n12716 ;
  assign n31618 = n23106 ^ n20902 ^ 1'b0 ;
  assign n31619 = n5833 & n31618 ;
  assign n31620 = n10133 ^ n9123 ^ n1848 ;
  assign n31621 = ~n30503 & n31620 ;
  assign n31622 = n18732 & ~n31621 ;
  assign n31623 = n15911 & n31622 ;
  assign n31624 = ( n12562 & n13689 ) | ( n12562 & ~n20288 ) | ( n13689 & ~n20288 ) ;
  assign n31625 = ~n11594 & n16267 ;
  assign n31626 = ~n23274 & n31625 ;
  assign n31627 = n11603 & ~n20787 ;
  assign n31628 = n28665 & n31627 ;
  assign n31629 = n9458 | n11032 ;
  assign n31630 = n12675 | n31629 ;
  assign n31631 = ~n31628 & n31630 ;
  assign n31633 = n26956 ^ n19200 ^ n4562 ;
  assign n31632 = ~n16615 & n16901 ;
  assign n31634 = n31633 ^ n31632 ^ 1'b0 ;
  assign n31635 = ( n10033 & ~n10663 ) | ( n10033 & n30942 ) | ( ~n10663 & n30942 ) ;
  assign n31638 = n924 & ~n6681 ;
  assign n31637 = ( ~n3117 & n10697 ) | ( ~n3117 & n23500 ) | ( n10697 & n23500 ) ;
  assign n31636 = n3931 & n26572 ;
  assign n31639 = n31638 ^ n31637 ^ n31636 ;
  assign n31640 = n31635 | n31639 ;
  assign n31641 = n31640 ^ n13386 ^ 1'b0 ;
  assign n31642 = ( n18359 & n19725 ) | ( n18359 & ~n25494 ) | ( n19725 & ~n25494 ) ;
  assign n31643 = ( ~n12992 & n14860 ) | ( ~n12992 & n22603 ) | ( n14860 & n22603 ) ;
  assign n31644 = n31643 ^ n7043 ^ n5548 ;
  assign n31647 = n10739 ^ n7503 ^ n2438 ;
  assign n31648 = ( ~n15109 & n24301 ) | ( ~n15109 & n31647 ) | ( n24301 & n31647 ) ;
  assign n31645 = ( n11429 & n13002 ) | ( n11429 & ~n22080 ) | ( n13002 & ~n22080 ) ;
  assign n31646 = n31645 ^ n14271 ^ 1'b0 ;
  assign n31649 = n31648 ^ n31646 ^ n12640 ;
  assign n31650 = n8046 & n9897 ;
  assign n31651 = n31650 ^ n27926 ^ 1'b0 ;
  assign n31652 = ( n16504 & ~n31649 ) | ( n16504 & n31651 ) | ( ~n31649 & n31651 ) ;
  assign n31653 = n24178 ^ n20992 ^ n9674 ;
  assign n31654 = n19131 ^ n17574 ^ 1'b0 ;
  assign n31655 = n25235 & ~n31654 ;
  assign n31656 = n8145 | n18010 ;
  assign n31657 = n31656 ^ n13688 ^ 1'b0 ;
  assign n31658 = n31655 & ~n31657 ;
  assign n31659 = n31658 ^ n12561 ^ n9655 ;
  assign n31660 = n29031 ^ n12484 ^ n12102 ;
  assign n31661 = ( n330 & n11670 ) | ( n330 & n31660 ) | ( n11670 & n31660 ) ;
  assign n31662 = n24541 ^ n11308 ^ n3325 ;
  assign n31663 = n31662 ^ n10447 ^ n10310 ;
  assign n31665 = n10322 ^ n6891 ^ n2633 ;
  assign n31664 = ( n834 & n4341 ) | ( n834 & n21440 ) | ( n4341 & n21440 ) ;
  assign n31666 = n31665 ^ n31664 ^ 1'b0 ;
  assign n31667 = ( n1448 & ~n18295 ) | ( n1448 & n19711 ) | ( ~n18295 & n19711 ) ;
  assign n31668 = n31568 ^ n20042 ^ n16443 ;
  assign n31669 = n22192 ^ n19903 ^ 1'b0 ;
  assign n31670 = n31668 & n31669 ;
  assign n31671 = n7753 & n14565 ;
  assign n31672 = n31671 ^ n5757 ^ 1'b0 ;
  assign n31673 = ( n3963 & ~n6317 ) | ( n3963 & n31672 ) | ( ~n6317 & n31672 ) ;
  assign n31674 = n1218 | n4484 ;
  assign n31675 = n12551 | n31674 ;
  assign n31676 = ~n14638 & n18173 ;
  assign n31677 = ~n31675 & n31676 ;
  assign n31678 = n4801 & ~n17730 ;
  assign n31679 = n5429 & n31678 ;
  assign n31680 = n5918 | n31679 ;
  assign n31681 = n31677 & ~n31680 ;
  assign n31682 = n31681 ^ n20157 ^ n6468 ;
  assign n31683 = ( n3775 & ~n21172 ) | ( n3775 & n25232 ) | ( ~n21172 & n25232 ) ;
  assign n31684 = n13452 & ~n22987 ;
  assign n31685 = ( n5237 & ~n7562 ) | ( n5237 & n15633 ) | ( ~n7562 & n15633 ) ;
  assign n31686 = n31685 ^ n29990 ^ n11199 ;
  assign n31687 = n22311 ^ n1753 ^ 1'b0 ;
  assign n31688 = n31604 & n31687 ;
  assign n31689 = x220 & ~n18825 ;
  assign n31690 = n14017 | n31689 ;
  assign n31691 = ( n4498 & n13419 ) | ( n4498 & ~n14856 ) | ( n13419 & ~n14856 ) ;
  assign n31692 = n13844 ^ n3282 ^ n3124 ;
  assign n31693 = ( n7185 & n25516 ) | ( n7185 & ~n31692 ) | ( n25516 & ~n31692 ) ;
  assign n31694 = n2608 | n3596 ;
  assign n31695 = n31694 ^ n4141 ^ 1'b0 ;
  assign n31696 = ( ~n1164 & n5338 ) | ( ~n1164 & n27216 ) | ( n5338 & n27216 ) ;
  assign n31697 = ~n2283 & n10764 ;
  assign n31698 = n31697 ^ n25773 ^ n5856 ;
  assign n31699 = n31698 ^ n12782 ^ n1594 ;
  assign n31700 = n22599 ^ n11923 ^ 1'b0 ;
  assign n31701 = n14490 & ~n31700 ;
  assign n31702 = n2659 & n31701 ;
  assign n31703 = n31702 ^ n17988 ^ 1'b0 ;
  assign n31704 = n13817 ^ n11941 ^ 1'b0 ;
  assign n31705 = n8494 | n31704 ;
  assign n31706 = n5593 & ~n7523 ;
  assign n31707 = n31705 & n31706 ;
  assign n31708 = n31707 ^ n16515 ^ n8676 ;
  assign n31709 = n31703 | n31708 ;
  assign n31710 = n2619 ^ n2583 ^ n1929 ;
  assign n31711 = ( n28684 & n30263 ) | ( n28684 & ~n31710 ) | ( n30263 & ~n31710 ) ;
  assign n31712 = n7859 & ~n28176 ;
  assign n31713 = ~n31711 & n31712 ;
  assign n31714 = n27736 ^ n15392 ^ n12818 ;
  assign n31715 = n31714 ^ n19483 ^ 1'b0 ;
  assign n31716 = n8806 | n10155 ;
  assign n31717 = n31716 ^ n8985 ^ 1'b0 ;
  assign n31718 = n26963 ^ n16477 ^ 1'b0 ;
  assign n31719 = n1664 | n31718 ;
  assign n31722 = n2927 & n4772 ;
  assign n31720 = n7108 | n10072 ;
  assign n31721 = n31720 ^ n16515 ^ 1'b0 ;
  assign n31723 = n31722 ^ n31721 ^ n6801 ;
  assign n31724 = ( n4305 & n14746 ) | ( n4305 & n31723 ) | ( n14746 & n31723 ) ;
  assign n31725 = n31724 ^ n21204 ^ n8099 ;
  assign n31726 = ~n3276 & n31725 ;
  assign n31727 = ( n914 & n5794 ) | ( n914 & ~n12037 ) | ( n5794 & ~n12037 ) ;
  assign n31728 = n13130 & n31727 ;
  assign n31729 = n6031 | n31728 ;
  assign n31730 = ( ~n5463 & n12198 ) | ( ~n5463 & n18938 ) | ( n12198 & n18938 ) ;
  assign n31731 = n31730 ^ n18868 ^ n5941 ;
  assign n31732 = n30680 ^ n6159 ^ n4245 ;
  assign n31733 = n14943 ^ n14556 ^ n2378 ;
  assign n31734 = n31733 ^ n9465 ^ n4798 ;
  assign n31740 = n25168 ^ n7156 ^ 1'b0 ;
  assign n31735 = n12673 ^ n8566 ^ n2264 ;
  assign n31736 = n31735 ^ n7914 ^ n1959 ;
  assign n31737 = n31736 ^ n24237 ^ 1'b0 ;
  assign n31738 = n20798 & n31737 ;
  assign n31739 = n4502 & n31738 ;
  assign n31741 = n31740 ^ n31739 ^ 1'b0 ;
  assign n31742 = n27839 ^ n5656 ^ n5209 ;
  assign n31743 = n5231 & ~n31742 ;
  assign n31744 = n28754 ^ n6460 ^ n5467 ;
  assign n31745 = n9915 & ~n16692 ;
  assign n31746 = n2342 & n31745 ;
  assign n31747 = n31746 ^ n4701 ^ 1'b0 ;
  assign n31748 = n31747 ^ n2240 ^ n672 ;
  assign n31749 = ( n2958 & n31744 ) | ( n2958 & n31748 ) | ( n31744 & n31748 ) ;
  assign n31750 = n2609 & n20759 ;
  assign n31751 = ( x135 & ~n4582 ) | ( x135 & n31750 ) | ( ~n4582 & n31750 ) ;
  assign n31752 = ( n3416 & n28517 ) | ( n3416 & ~n31751 ) | ( n28517 & ~n31751 ) ;
  assign n31753 = n12117 | n25563 ;
  assign n31754 = n31753 ^ n21804 ^ 1'b0 ;
  assign n31755 = n18127 ^ n17247 ^ n17197 ;
  assign n31756 = ( n8424 & n22218 ) | ( n8424 & ~n31755 ) | ( n22218 & ~n31755 ) ;
  assign n31757 = n10329 ^ n7925 ^ n4261 ;
  assign n31758 = ( n7092 & ~n26279 ) | ( n7092 & n31757 ) | ( ~n26279 & n31757 ) ;
  assign n31759 = ( n2187 & n2476 ) | ( n2187 & ~n3944 ) | ( n2476 & ~n3944 ) ;
  assign n31760 = n31759 ^ n22762 ^ 1'b0 ;
  assign n31761 = n14653 & n31760 ;
  assign n31762 = n17357 ^ n1490 ^ 1'b0 ;
  assign n31763 = n31762 ^ n21804 ^ n2275 ;
  assign n31764 = n4175 ^ n3387 ^ 1'b0 ;
  assign n31765 = n30589 & ~n31764 ;
  assign n31766 = ( ~n1491 & n2697 ) | ( ~n1491 & n31765 ) | ( n2697 & n31765 ) ;
  assign n31767 = n16268 ^ n10549 ^ 1'b0 ;
  assign n31768 = ~n4468 & n5482 ;
  assign n31769 = n4087 & n31768 ;
  assign n31770 = n20661 & ~n31769 ;
  assign n31772 = n13844 ^ n3944 ^ n3542 ;
  assign n31771 = ~n13538 & n19089 ;
  assign n31773 = n31772 ^ n31771 ^ 1'b0 ;
  assign n31774 = n31773 ^ n5641 ^ 1'b0 ;
  assign n31775 = ~n11601 & n31774 ;
  assign n31777 = n2961 ^ n657 ^ 1'b0 ;
  assign n31776 = ~n8953 & n18470 ;
  assign n31778 = n31777 ^ n31776 ^ 1'b0 ;
  assign n31779 = ~n2552 & n31778 ;
  assign n31780 = n585 & n1023 ;
  assign n31781 = ~x185 & n31780 ;
  assign n31782 = ( n4846 & ~n5513 ) | ( n4846 & n31781 ) | ( ~n5513 & n31781 ) ;
  assign n31783 = ( n3288 & n9892 ) | ( n3288 & ~n12062 ) | ( n9892 & ~n12062 ) ;
  assign n31784 = ( n4342 & ~n22713 ) | ( n4342 & n31783 ) | ( ~n22713 & n31783 ) ;
  assign n31785 = ( ~n29752 & n31782 ) | ( ~n29752 & n31784 ) | ( n31782 & n31784 ) ;
  assign n31786 = n29847 ^ n2885 ^ 1'b0 ;
  assign n31787 = n25805 | n31786 ;
  assign n31788 = ~n31785 & n31787 ;
  assign n31789 = n25558 ^ n5623 ^ n578 ;
  assign n31790 = ( n3578 & n18538 ) | ( n3578 & ~n31789 ) | ( n18538 & ~n31789 ) ;
  assign n31791 = n2556 & n24985 ;
  assign n31792 = n31791 ^ n19981 ^ 1'b0 ;
  assign n31793 = ( ~n22567 & n31790 ) | ( ~n22567 & n31792 ) | ( n31790 & n31792 ) ;
  assign n31794 = n10456 ^ n6206 ^ n759 ;
  assign n31795 = ( n1078 & ~n10910 ) | ( n1078 & n31794 ) | ( ~n10910 & n31794 ) ;
  assign n31796 = ( ~n3638 & n9910 ) | ( ~n3638 & n15770 ) | ( n9910 & n15770 ) ;
  assign n31797 = ( n8907 & n14192 ) | ( n8907 & ~n18551 ) | ( n14192 & ~n18551 ) ;
  assign n31798 = n14050 ^ n7385 ^ n4705 ;
  assign n31799 = n12900 ^ n11652 ^ n2909 ;
  assign n31800 = ( n3673 & n9553 ) | ( n3673 & n12894 ) | ( n9553 & n12894 ) ;
  assign n31801 = n301 & n21582 ;
  assign n31802 = n31801 ^ n4985 ^ 1'b0 ;
  assign n31803 = n2689 & n31802 ;
  assign n31804 = n31803 ^ n21739 ^ n9608 ;
  assign n31805 = n31800 | n31804 ;
  assign n31806 = ~n6802 & n13048 ;
  assign n31807 = n28295 & n31806 ;
  assign n31808 = n4169 & n19236 ;
  assign n31809 = n31808 ^ n2899 ^ 1'b0 ;
  assign n31810 = ~n3151 & n31809 ;
  assign n31811 = n5437 & ~n31810 ;
  assign n31812 = n565 | n2824 ;
  assign n31813 = n31812 ^ n9477 ^ 1'b0 ;
  assign n31814 = n31813 ^ n25108 ^ n4286 ;
  assign n31815 = ( n9393 & n22273 ) | ( n9393 & n27547 ) | ( n22273 & n27547 ) ;
  assign n31816 = ( ~n982 & n7761 ) | ( ~n982 & n9282 ) | ( n7761 & n9282 ) ;
  assign n31817 = n6045 & n22682 ;
  assign n31818 = ( n7237 & n12939 ) | ( n7237 & n31817 ) | ( n12939 & n31817 ) ;
  assign n31819 = n25489 ^ n18604 ^ 1'b0 ;
  assign n31821 = n10985 ^ n4859 ^ 1'b0 ;
  assign n31822 = n2750 & ~n31821 ;
  assign n31820 = n6236 & ~n8543 ;
  assign n31823 = n31822 ^ n31820 ^ 1'b0 ;
  assign n31824 = ( n5548 & n5744 ) | ( n5548 & n15571 ) | ( n5744 & n15571 ) ;
  assign n31825 = n1508 & ~n31824 ;
  assign n31826 = ~n27858 & n31825 ;
  assign n31827 = n25582 ^ n15868 ^ n14644 ;
  assign n31828 = n31827 ^ n31426 ^ n17975 ;
  assign n31829 = ( ~n3223 & n8444 ) | ( ~n3223 & n9530 ) | ( n8444 & n9530 ) ;
  assign n31830 = n19029 ^ n3052 ^ 1'b0 ;
  assign n31831 = n31830 ^ n14407 ^ 1'b0 ;
  assign n31832 = n23933 | n31831 ;
  assign n31833 = ( ~n24455 & n31829 ) | ( ~n24455 & n31832 ) | ( n31829 & n31832 ) ;
  assign n31834 = n22777 ^ n7327 ^ 1'b0 ;
  assign n31835 = n10899 & n31834 ;
  assign n31836 = ( n847 & n19960 ) | ( n847 & ~n31835 ) | ( n19960 & ~n31835 ) ;
  assign n31837 = n31836 ^ n28250 ^ n23997 ;
  assign n31838 = n23308 ^ n19299 ^ x184 ;
  assign n31839 = ~n1931 & n23501 ;
  assign n31840 = n31839 ^ n4930 ^ 1'b0 ;
  assign n31841 = ~n20353 & n31840 ;
  assign n31842 = ( n6990 & n22174 ) | ( n6990 & n31841 ) | ( n22174 & n31841 ) ;
  assign n31843 = x70 & n8875 ;
  assign n31844 = ~n4514 & n31843 ;
  assign n31845 = n21342 & n31844 ;
  assign n31847 = n19531 ^ n11130 ^ n6547 ;
  assign n31846 = ( ~n4998 & n18773 ) | ( ~n4998 & n25888 ) | ( n18773 & n25888 ) ;
  assign n31848 = n31847 ^ n31846 ^ n1487 ;
  assign n31849 = n20399 ^ n7111 ^ 1'b0 ;
  assign n31850 = n12427 | n31849 ;
  assign n31851 = ( ~x39 & n476 ) | ( ~x39 & n21309 ) | ( n476 & n21309 ) ;
  assign n31852 = ( n5260 & n31850 ) | ( n5260 & n31851 ) | ( n31850 & n31851 ) ;
  assign n31853 = n9874 | n25116 ;
  assign n31854 = ( ~n15238 & n21907 ) | ( ~n15238 & n27220 ) | ( n21907 & n27220 ) ;
  assign n31855 = ( n9674 & n18552 ) | ( n9674 & n20261 ) | ( n18552 & n20261 ) ;
  assign n31856 = n10581 & n31855 ;
  assign n31857 = ~n552 & n31856 ;
  assign n31858 = n1753 & ~n31857 ;
  assign n31859 = n31858 ^ n16156 ^ 1'b0 ;
  assign n31860 = n8680 & ~n19806 ;
  assign n31861 = n3764 & ~n20366 ;
  assign n31862 = ~n31860 & n31861 ;
  assign n31863 = ( n7328 & n10525 ) | ( n7328 & ~n24266 ) | ( n10525 & ~n24266 ) ;
  assign n31864 = ( ~x121 & n5575 ) | ( ~x121 & n21075 ) | ( n5575 & n21075 ) ;
  assign n31865 = n31864 ^ n3002 ^ 1'b0 ;
  assign n31866 = ( ~n27290 & n31863 ) | ( ~n27290 & n31865 ) | ( n31863 & n31865 ) ;
  assign n31867 = n6894 & n27011 ;
  assign n31868 = n9309 ^ n9166 ^ 1'b0 ;
  assign n31869 = n9512 & ~n31868 ;
  assign n31870 = n31869 ^ n6816 ^ 1'b0 ;
  assign n31871 = n1194 | n20880 ;
  assign n31872 = n31871 ^ n16110 ^ n14047 ;
  assign n31873 = ( n8364 & ~n28310 ) | ( n8364 & n31872 ) | ( ~n28310 & n31872 ) ;
  assign n31874 = ( n1585 & n15672 ) | ( n1585 & n24477 ) | ( n15672 & n24477 ) ;
  assign n31875 = ( n754 & n8279 ) | ( n754 & ~n31874 ) | ( n8279 & ~n31874 ) ;
  assign n31876 = n12363 | n13187 ;
  assign n31877 = n31876 ^ n1870 ^ 1'b0 ;
  assign n31878 = n12079 & ~n20909 ;
  assign n31879 = ~n31877 & n31878 ;
  assign n31880 = n26646 ^ n4939 ^ 1'b0 ;
  assign n31881 = n2104 & n28198 ;
  assign n31882 = n31881 ^ n10780 ^ 1'b0 ;
  assign n31883 = n7155 | n31882 ;
  assign n31884 = n6368 | n10959 ;
  assign n31885 = n31884 ^ n30009 ^ 1'b0 ;
  assign n31886 = n14507 & ~n28970 ;
  assign n31887 = n3401 & n31886 ;
  assign n31888 = n31887 ^ n26430 ^ 1'b0 ;
  assign n31889 = n7832 & ~n31888 ;
  assign n31890 = n15144 & n15468 ;
  assign n31891 = n23975 & n31890 ;
  assign n31892 = ( n1759 & ~n15846 ) | ( n1759 & n31891 ) | ( ~n15846 & n31891 ) ;
  assign n31893 = n31892 ^ n30275 ^ n6109 ;
  assign n31894 = ~n8161 & n31893 ;
  assign n31895 = n31894 ^ n3678 ^ 1'b0 ;
  assign n31896 = n3720 | n20292 ;
  assign n31897 = n2827 & ~n31896 ;
  assign n31898 = n28384 & ~n31897 ;
  assign n31899 = n29569 ^ n13094 ^ n2334 ;
  assign n31900 = ( n6882 & n22860 ) | ( n6882 & ~n31899 ) | ( n22860 & ~n31899 ) ;
  assign n31901 = n10197 | n19834 ;
  assign n31902 = n31901 ^ n1305 ^ 1'b0 ;
  assign n31903 = n31902 ^ n13677 ^ n3260 ;
  assign n31904 = ( n10623 & n31900 ) | ( n10623 & n31903 ) | ( n31900 & n31903 ) ;
  assign n31905 = ~n11226 & n22863 ;
  assign n31906 = n20420 ^ n8465 ^ 1'b0 ;
  assign n31907 = n12891 ^ n10868 ^ 1'b0 ;
  assign n31908 = n1210 | n31907 ;
  assign n31909 = ( ~n882 & n6603 ) | ( ~n882 & n7986 ) | ( n6603 & n7986 ) ;
  assign n31910 = n25303 ^ n19422 ^ 1'b0 ;
  assign n31911 = ~n31909 & n31910 ;
  assign n31912 = n20856 ^ n14890 ^ 1'b0 ;
  assign n31913 = ( ~n634 & n11364 ) | ( ~n634 & n31912 ) | ( n11364 & n31912 ) ;
  assign n31914 = n31913 ^ n10922 ^ 1'b0 ;
  assign n31915 = n975 ^ n791 ^ 1'b0 ;
  assign n31916 = n31915 ^ n28419 ^ n20503 ;
  assign n31917 = n31855 ^ n27405 ^ n8095 ;
  assign n31918 = n12873 ^ n10206 ^ n8887 ;
  assign n31919 = ( ~n16984 & n24363 ) | ( ~n16984 & n26742 ) | ( n24363 & n26742 ) ;
  assign n31920 = n31919 ^ n13798 ^ n6733 ;
  assign n31924 = n4937 & ~n20150 ;
  assign n31925 = n31924 ^ n23829 ^ 1'b0 ;
  assign n31926 = ( n15129 & n23730 ) | ( n15129 & n31925 ) | ( n23730 & n31925 ) ;
  assign n31921 = ( ~n2081 & n4196 ) | ( ~n2081 & n20033 ) | ( n4196 & n20033 ) ;
  assign n31922 = n31921 ^ n24084 ^ 1'b0 ;
  assign n31923 = ~n31866 & n31922 ;
  assign n31927 = n31926 ^ n31923 ^ 1'b0 ;
  assign n31928 = ( n1629 & n6543 ) | ( n1629 & n13674 ) | ( n6543 & n13674 ) ;
  assign n31929 = ( x155 & n25445 ) | ( x155 & ~n31928 ) | ( n25445 & ~n31928 ) ;
  assign n31930 = ( n5823 & n7703 ) | ( n5823 & n31929 ) | ( n7703 & n31929 ) ;
  assign n31931 = ( ~n4705 & n12956 ) | ( ~n4705 & n31930 ) | ( n12956 & n31930 ) ;
  assign n31932 = ~n18865 & n31931 ;
  assign n31937 = n1098 & n7991 ;
  assign n31938 = n31937 ^ n10418 ^ 1'b0 ;
  assign n31933 = ( ~n4480 & n8611 ) | ( ~n4480 & n11920 ) | ( n8611 & n11920 ) ;
  assign n31934 = ~n3336 & n31933 ;
  assign n31935 = n4048 & n31934 ;
  assign n31936 = ( n3813 & ~n6915 ) | ( n3813 & n31935 ) | ( ~n6915 & n31935 ) ;
  assign n31939 = n31938 ^ n31936 ^ n11696 ;
  assign n31940 = n24196 ^ n10267 ^ 1'b0 ;
  assign n31941 = n31940 ^ n28144 ^ n26000 ;
  assign n31942 = n24960 ^ n21924 ^ n4050 ;
  assign n31943 = n31942 ^ n30414 ^ n23035 ;
  assign n31944 = n27542 ^ n16076 ^ n11915 ;
  assign n31945 = ( ~n6738 & n7310 ) | ( ~n6738 & n23149 ) | ( n7310 & n23149 ) ;
  assign n31946 = x170 & ~n31945 ;
  assign n31947 = n31946 ^ n22628 ^ 1'b0 ;
  assign n31948 = n8522 | n10526 ;
  assign n31949 = ( n5503 & n17764 ) | ( n5503 & n31948 ) | ( n17764 & n31948 ) ;
  assign n31950 = n17977 ^ n4925 ^ n4340 ;
  assign n31951 = n31950 ^ n26847 ^ n26121 ;
  assign n31952 = ( ~n7977 & n8930 ) | ( ~n7977 & n13315 ) | ( n8930 & n13315 ) ;
  assign n31953 = n7658 & n11747 ;
  assign n31954 = n31953 ^ n17205 ^ 1'b0 ;
  assign n31955 = n4819 ^ n933 ^ 1'b0 ;
  assign n31956 = ( ~x5 & n10583 ) | ( ~x5 & n31955 ) | ( n10583 & n31955 ) ;
  assign n31957 = n20502 ^ n17466 ^ n13854 ;
  assign n31958 = n23303 | n31957 ;
  assign n31959 = n31956 & ~n31958 ;
  assign n31960 = n18775 ^ n14805 ^ n12859 ;
  assign n31961 = n15283 ^ n1956 ^ 1'b0 ;
  assign n31962 = x21 & ~n1762 ;
  assign n31963 = ~n4888 & n31962 ;
  assign n31964 = n31961 & ~n31963 ;
  assign n31965 = ( n2523 & n11664 ) | ( n2523 & n14793 ) | ( n11664 & n14793 ) ;
  assign n31966 = n31965 ^ n23053 ^ 1'b0 ;
  assign n31967 = n30128 ^ n9102 ^ n6851 ;
  assign n31968 = n11608 & ~n28895 ;
  assign n31969 = n23415 ^ n12274 ^ 1'b0 ;
  assign n31970 = n9313 & n31969 ;
  assign n31971 = n7654 & ~n31970 ;
  assign n31972 = ( n13425 & n28157 ) | ( n13425 & ~n31971 ) | ( n28157 & ~n31971 ) ;
  assign n31973 = ( n2332 & n15875 ) | ( n2332 & ~n31972 ) | ( n15875 & ~n31972 ) ;
  assign n31974 = n16274 ^ n11203 ^ 1'b0 ;
  assign n31975 = ~n31973 & n31974 ;
  assign n31976 = n29236 ^ n26503 ^ n17861 ;
  assign n31977 = ( n2381 & n5800 ) | ( n2381 & ~n10431 ) | ( n5800 & ~n10431 ) ;
  assign n31978 = n16288 ^ n8166 ^ 1'b0 ;
  assign n31979 = ( ~n16714 & n28496 ) | ( ~n16714 & n30348 ) | ( n28496 & n30348 ) ;
  assign n31980 = ( n31977 & n31978 ) | ( n31977 & n31979 ) | ( n31978 & n31979 ) ;
  assign n31981 = ( n19856 & n26298 ) | ( n19856 & n31980 ) | ( n26298 & n31980 ) ;
  assign n31982 = n17270 ^ n15634 ^ n2697 ;
  assign n31983 = n15990 ^ n5790 ^ n2057 ;
  assign n31984 = ( n19061 & n25055 ) | ( n19061 & ~n31983 ) | ( n25055 & ~n31983 ) ;
  assign n31985 = ( n17257 & ~n28235 ) | ( n17257 & n31984 ) | ( ~n28235 & n31984 ) ;
  assign n31986 = ( n15530 & ~n24252 ) | ( n15530 & n31755 ) | ( ~n24252 & n31755 ) ;
  assign n31987 = n31986 ^ n25578 ^ n3858 ;
  assign n31988 = ( n1251 & n15364 ) | ( n1251 & ~n28097 ) | ( n15364 & ~n28097 ) ;
  assign n31989 = n20388 & n31988 ;
  assign n31990 = n31989 ^ n8262 ^ 1'b0 ;
  assign n31991 = n4437 & n10328 ;
  assign n31992 = n13782 ^ n8895 ^ n1293 ;
  assign n31994 = ( n3619 & n3953 ) | ( n3619 & n16559 ) | ( n3953 & n16559 ) ;
  assign n31993 = ( n16124 & ~n25727 ) | ( n16124 & n29750 ) | ( ~n25727 & n29750 ) ;
  assign n31995 = n31994 ^ n31993 ^ n17695 ;
  assign n31996 = n31995 ^ n26359 ^ 1'b0 ;
  assign n31997 = n18324 & ~n31996 ;
  assign n31998 = n31997 ^ n29107 ^ n2145 ;
  assign n31999 = n30432 ^ n21717 ^ n16652 ;
  assign n32005 = n4247 ^ n3322 ^ n1586 ;
  assign n32000 = n7742 ^ n6512 ^ 1'b0 ;
  assign n32001 = n13466 | n32000 ;
  assign n32002 = ( n6538 & n16441 ) | ( n6538 & ~n32001 ) | ( n16441 & ~n32001 ) ;
  assign n32003 = n32002 ^ n8173 ^ 1'b0 ;
  assign n32004 = ~n18898 & n32003 ;
  assign n32006 = n32005 ^ n32004 ^ n3365 ;
  assign n32007 = n14509 ^ n7294 ^ n656 ;
  assign n32008 = ( n8977 & ~n14995 ) | ( n8977 & n19394 ) | ( ~n14995 & n19394 ) ;
  assign n32009 = n11317 ^ n5014 ^ 1'b0 ;
  assign n32010 = ( ~n735 & n15039 ) | ( ~n735 & n32009 ) | ( n15039 & n32009 ) ;
  assign n32011 = n32010 ^ n15178 ^ n10398 ;
  assign n32012 = n30991 ^ n20091 ^ 1'b0 ;
  assign n32013 = ~n32011 & n32012 ;
  assign n32014 = ~n5055 & n32013 ;
  assign n32015 = n32008 & n32014 ;
  assign n32016 = n28523 ^ n11295 ^ 1'b0 ;
  assign n32017 = n6638 | n32016 ;
  assign n32018 = n6946 | n18115 ;
  assign n32019 = n32018 ^ n3630 ^ 1'b0 ;
  assign n32020 = n28817 ^ n7260 ^ n3119 ;
  assign n32021 = ( ~n17552 & n32019 ) | ( ~n17552 & n32020 ) | ( n32019 & n32020 ) ;
  assign n32022 = ( n2235 & ~n3638 ) | ( n2235 & n31979 ) | ( ~n3638 & n31979 ) ;
  assign n32023 = ( ~n2324 & n3919 ) | ( ~n2324 & n12362 ) | ( n3919 & n12362 ) ;
  assign n32024 = n25297 ^ n9045 ^ n673 ;
  assign n32025 = ( ~n6246 & n13334 ) | ( ~n6246 & n32024 ) | ( n13334 & n32024 ) ;
  assign n32026 = n7118 ^ n2933 ^ 1'b0 ;
  assign n32027 = n9771 & n32026 ;
  assign n32028 = n32027 ^ n19923 ^ 1'b0 ;
  assign n32029 = n5126 | n28840 ;
  assign n32030 = n310 & ~n32029 ;
  assign n32031 = n13888 ^ n4457 ^ n2910 ;
  assign n32032 = n32031 ^ n23413 ^ n21450 ;
  assign n32033 = n32032 ^ n5235 ^ n1256 ;
  assign n32034 = n32033 ^ n31626 ^ n8254 ;
  assign n32035 = n20553 ^ n11895 ^ n6245 ;
  assign n32036 = n31275 ^ n26624 ^ n9516 ;
  assign n32037 = n32036 ^ n17792 ^ n9839 ;
  assign n32038 = n1055 | n32037 ;
  assign n32039 = n32035 | n32038 ;
  assign n32040 = n8384 | n22204 ;
  assign n32041 = n3613 & ~n32040 ;
  assign n32042 = n26501 ^ n24864 ^ n9884 ;
  assign n32043 = ( ~n4533 & n22159 ) | ( ~n4533 & n32042 ) | ( n22159 & n32042 ) ;
  assign n32046 = ( n4164 & ~n11965 ) | ( n4164 & n16081 ) | ( ~n11965 & n16081 ) ;
  assign n32044 = n24830 ^ n4318 ^ n2760 ;
  assign n32045 = ( ~n13264 & n19257 ) | ( ~n13264 & n32044 ) | ( n19257 & n32044 ) ;
  assign n32047 = n32046 ^ n32045 ^ n2299 ;
  assign n32048 = ( ~n7415 & n8253 ) | ( ~n7415 & n32047 ) | ( n8253 & n32047 ) ;
  assign n32049 = ( n4570 & n5824 ) | ( n4570 & ~n11564 ) | ( n5824 & ~n11564 ) ;
  assign n32050 = ( n6784 & ~n13787 ) | ( n6784 & n28014 ) | ( ~n13787 & n28014 ) ;
  assign n32051 = ( n13944 & n16182 ) | ( n13944 & ~n32050 ) | ( n16182 & ~n32050 ) ;
  assign n32052 = n32051 ^ n28501 ^ n1487 ;
  assign n32053 = n4311 & n24361 ;
  assign n32054 = n1495 ^ n1284 ^ n1046 ;
  assign n32055 = ( n8733 & ~n13016 ) | ( n8733 & n32054 ) | ( ~n13016 & n32054 ) ;
  assign n32056 = ( ~n1382 & n1796 ) | ( ~n1382 & n32055 ) | ( n1796 & n32055 ) ;
  assign n32057 = n16405 ^ n10163 ^ 1'b0 ;
  assign n32058 = n32057 ^ n20678 ^ n9949 ;
  assign n32059 = ( n4003 & ~n8448 ) | ( n4003 & n10673 ) | ( ~n8448 & n10673 ) ;
  assign n32060 = n32059 ^ n19979 ^ 1'b0 ;
  assign n32061 = n9353 & n32060 ;
  assign n32062 = n32058 | n32061 ;
  assign n32063 = n21530 ^ n20588 ^ n17517 ;
  assign n32064 = n25475 ^ n8777 ^ n4501 ;
  assign n32065 = ( n10187 & ~n20239 ) | ( n10187 & n25481 ) | ( ~n20239 & n25481 ) ;
  assign n32066 = ~n16880 & n32065 ;
  assign n32067 = ( n10743 & n14525 ) | ( n10743 & n17484 ) | ( n14525 & n17484 ) ;
  assign n32068 = n32067 ^ n4594 ^ 1'b0 ;
  assign n32069 = n32066 & n32068 ;
  assign n32070 = ~n10211 & n20525 ;
  assign n32071 = n13482 | n32070 ;
  assign n32072 = n32071 ^ n1997 ^ 1'b0 ;
  assign n32073 = ( ~n22913 & n30874 ) | ( ~n22913 & n32072 ) | ( n30874 & n32072 ) ;
  assign n32074 = n32073 ^ n9356 ^ 1'b0 ;
  assign n32075 = n1998 & n23510 ;
  assign n32076 = ~n32074 & n32075 ;
  assign n32077 = n2309 | n15004 ;
  assign n32078 = n12944 | n32077 ;
  assign n32079 = n32078 ^ n26412 ^ n7445 ;
  assign n32080 = n24908 | n32079 ;
  assign n32085 = ( ~n5739 & n16732 ) | ( ~n5739 & n31556 ) | ( n16732 & n31556 ) ;
  assign n32086 = ( n7327 & n10525 ) | ( n7327 & n15943 ) | ( n10525 & n15943 ) ;
  assign n32087 = n2226 | n32086 ;
  assign n32088 = ~n3523 & n32087 ;
  assign n32089 = n32085 & n32088 ;
  assign n32083 = n3447 | n8122 ;
  assign n32084 = n2545 & ~n32083 ;
  assign n32081 = n7774 ^ n7442 ^ n1746 ;
  assign n32082 = ( ~n15717 & n23201 ) | ( ~n15717 & n32081 ) | ( n23201 & n32081 ) ;
  assign n32090 = n32089 ^ n32084 ^ n32082 ;
  assign n32091 = n19776 | n26541 ;
  assign n32092 = n7221 & n22502 ;
  assign n32093 = ~n17764 & n32092 ;
  assign n32094 = ( n11349 & n16453 ) | ( n11349 & ~n26751 ) | ( n16453 & ~n26751 ) ;
  assign n32095 = n2872 | n11773 ;
  assign n32096 = n32095 ^ n13921 ^ 1'b0 ;
  assign n32097 = n25109 ^ n5956 ^ n4263 ;
  assign n32098 = n32097 ^ n16638 ^ n3374 ;
  assign n32099 = n5037 & n32098 ;
  assign n32100 = n2449 & n32099 ;
  assign n32101 = n32096 & n32100 ;
  assign n32102 = n32101 ^ n27094 ^ n12580 ;
  assign n32103 = n5878 ^ n5065 ^ 1'b0 ;
  assign n32104 = ( n3723 & n4169 ) | ( n3723 & ~n32103 ) | ( n4169 & ~n32103 ) ;
  assign n32105 = n16649 ^ n15306 ^ n13950 ;
  assign n32106 = n32105 ^ n19210 ^ n14611 ;
  assign n32107 = n20369 ^ n11459 ^ 1'b0 ;
  assign n32108 = n26825 | n32107 ;
  assign n32109 = n32106 | n32108 ;
  assign n32110 = n31157 ^ n30611 ^ 1'b0 ;
  assign n32111 = ( n798 & n21025 ) | ( n798 & n32110 ) | ( n21025 & n32110 ) ;
  assign n32112 = n15401 & n32111 ;
  assign n32113 = n32112 ^ n19271 ^ 1'b0 ;
  assign n32114 = n10896 & ~n27750 ;
  assign n32115 = n5806 & n32114 ;
  assign n32116 = n1433 & ~n28297 ;
  assign n32117 = n6015 | n32116 ;
  assign n32118 = n3125 & ~n32117 ;
  assign n32119 = ( ~x245 & n1457 ) | ( ~x245 & n8374 ) | ( n1457 & n8374 ) ;
  assign n32120 = ( n9128 & n32118 ) | ( n9128 & n32119 ) | ( n32118 & n32119 ) ;
  assign n32121 = n18661 ^ n11716 ^ n525 ;
  assign n32123 = ( n2861 & n5080 ) | ( n2861 & n6596 ) | ( n5080 & n6596 ) ;
  assign n32122 = n9487 ^ n5883 ^ 1'b0 ;
  assign n32124 = n32123 ^ n32122 ^ x28 ;
  assign n32125 = ( n26998 & n32121 ) | ( n26998 & ~n32124 ) | ( n32121 & ~n32124 ) ;
  assign n32126 = ( x187 & n32120 ) | ( x187 & ~n32125 ) | ( n32120 & ~n32125 ) ;
  assign n32127 = n1449 & ~n12339 ;
  assign n32128 = n32127 ^ n17824 ^ n4248 ;
  assign n32129 = ( n14950 & n24991 ) | ( n14950 & n32128 ) | ( n24991 & n32128 ) ;
  assign n32131 = n31197 ^ n12090 ^ n644 ;
  assign n32130 = n18797 & ~n30055 ;
  assign n32132 = n32131 ^ n32130 ^ n21217 ;
  assign n32133 = n32132 ^ n17758 ^ n467 ;
  assign n32134 = n9096 | n32133 ;
  assign n32135 = n12186 ^ n7864 ^ 1'b0 ;
  assign n32136 = n3496 | n32135 ;
  assign n32137 = n30987 ^ n23416 ^ 1'b0 ;
  assign n32138 = ~n5755 & n32137 ;
  assign n32139 = n24908 | n32138 ;
  assign n32140 = ( ~n3385 & n8749 ) | ( ~n3385 & n10602 ) | ( n8749 & n10602 ) ;
  assign n32141 = n13153 & ~n29196 ;
  assign n32142 = ~n14383 & n32141 ;
  assign n32143 = n32142 ^ n19429 ^ n13828 ;
  assign n32144 = ( n11327 & n27109 ) | ( n11327 & ~n32143 ) | ( n27109 & ~n32143 ) ;
  assign n32145 = ( ~n3568 & n7565 ) | ( ~n3568 & n16297 ) | ( n7565 & n16297 ) ;
  assign n32146 = n351 & n23818 ;
  assign n32147 = ~n22853 & n32146 ;
  assign n32148 = n32147 ^ n19656 ^ n12086 ;
  assign n32149 = n21866 ^ x70 ^ 1'b0 ;
  assign n32150 = n17045 | n32149 ;
  assign n32151 = n32150 ^ n18904 ^ n7853 ;
  assign n32152 = n32151 ^ n26699 ^ n284 ;
  assign n32153 = n2233 & n2722 ;
  assign n32154 = n32153 ^ n825 ^ 1'b0 ;
  assign n32155 = ( n22884 & ~n29279 ) | ( n22884 & n31103 ) | ( ~n29279 & n31103 ) ;
  assign n32156 = n20190 ^ n17514 ^ n5999 ;
  assign n32157 = n9142 ^ n2509 ^ 1'b0 ;
  assign n32158 = n32157 ^ n13708 ^ n1524 ;
  assign n32159 = n16011 & n32158 ;
  assign n32160 = ( n23595 & ~n32156 ) | ( n23595 & n32159 ) | ( ~n32156 & n32159 ) ;
  assign n32161 = n5411 ^ n3757 ^ n3515 ;
  assign n32162 = n32161 ^ n22728 ^ n5789 ;
  assign n32163 = n32162 ^ n10206 ^ 1'b0 ;
  assign n32164 = n32163 ^ n30574 ^ n5169 ;
  assign n32165 = n30234 ^ n12476 ^ n8862 ;
  assign n32166 = n31202 ^ n8955 ^ n1710 ;
  assign n32168 = n22442 ^ n21637 ^ n17326 ;
  assign n32167 = n6029 | n13949 ;
  assign n32169 = n32168 ^ n32167 ^ n14305 ;
  assign n32170 = n30675 ^ n24292 ^ n2390 ;
  assign n32171 = ( n15640 & n26875 ) | ( n15640 & ~n27028 ) | ( n26875 & ~n27028 ) ;
  assign n32172 = n26942 ^ n19754 ^ n3111 ;
  assign n32173 = n27857 ^ n24618 ^ n271 ;
  assign n32174 = n32173 ^ n27520 ^ n8547 ;
  assign n32175 = n19813 ^ n11244 ^ n3864 ;
  assign n32176 = n15178 & ~n19453 ;
  assign n32177 = n32175 & n32176 ;
  assign n32178 = n32177 ^ n4141 ^ n3282 ;
  assign n32179 = n1268 ^ n331 ^ 1'b0 ;
  assign n32180 = n12914 | n32179 ;
  assign n32181 = n31191 ^ n2527 ^ 1'b0 ;
  assign n32182 = n8075 & n9189 ;
  assign n32183 = ~n24932 & n32182 ;
  assign n32189 = n24170 ^ n14936 ^ n7282 ;
  assign n32187 = n10721 ^ n10316 ^ n9670 ;
  assign n32184 = n1787 & n24447 ;
  assign n32185 = n5657 & n32184 ;
  assign n32186 = n7594 | n32185 ;
  assign n32188 = n32187 ^ n32186 ^ 1'b0 ;
  assign n32190 = n32189 ^ n32188 ^ 1'b0 ;
  assign n32191 = n24466 ^ n15343 ^ n9557 ;
  assign n32200 = n30488 ^ n9222 ^ 1'b0 ;
  assign n32192 = ~n1369 & n28457 ;
  assign n32193 = n26766 & n32192 ;
  assign n32194 = n32193 ^ n25472 ^ 1'b0 ;
  assign n32196 = n6983 ^ n1555 ^ 1'b0 ;
  assign n32197 = n1797 & ~n32196 ;
  assign n32195 = n21313 ^ n18167 ^ n4518 ;
  assign n32198 = n32197 ^ n32195 ^ n1823 ;
  assign n32199 = n32194 | n32198 ;
  assign n32201 = n32200 ^ n32199 ^ 1'b0 ;
  assign n32202 = ( n10022 & n15124 ) | ( n10022 & ~n29077 ) | ( n15124 & ~n29077 ) ;
  assign n32203 = ( n1305 & ~n16020 ) | ( n1305 & n32202 ) | ( ~n16020 & n32202 ) ;
  assign n32205 = n3949 & n8503 ;
  assign n32204 = n25914 | n30915 ;
  assign n32206 = n32205 ^ n32204 ^ 1'b0 ;
  assign n32208 = n17448 ^ n10023 ^ n4289 ;
  assign n32207 = n25596 ^ n15372 ^ n6060 ;
  assign n32209 = n32208 ^ n32207 ^ 1'b0 ;
  assign n32210 = ( n766 & n2800 ) | ( n766 & ~n2837 ) | ( n2800 & ~n2837 ) ;
  assign n32211 = ( ~n6265 & n8861 ) | ( ~n6265 & n10037 ) | ( n8861 & n10037 ) ;
  assign n32212 = ( n4733 & n10851 ) | ( n4733 & ~n18530 ) | ( n10851 & ~n18530 ) ;
  assign n32213 = ( n5724 & n32211 ) | ( n5724 & ~n32212 ) | ( n32211 & ~n32212 ) ;
  assign n32214 = n7044 ^ x172 ^ 1'b0 ;
  assign n32215 = n32214 ^ n11330 ^ n8707 ;
  assign n32216 = n32215 ^ n25512 ^ 1'b0 ;
  assign n32218 = n10051 & ~n11481 ;
  assign n32217 = ~n1106 & n9774 ;
  assign n32219 = n32218 ^ n32217 ^ 1'b0 ;
  assign n32220 = n32219 ^ n29858 ^ n18715 ;
  assign n32221 = n9972 ^ n5858 ^ 1'b0 ;
  assign n32222 = n5092 | n32221 ;
  assign n32223 = ( n3072 & n23011 ) | ( n3072 & n28661 ) | ( n23011 & n28661 ) ;
  assign n32224 = n32223 ^ n20005 ^ 1'b0 ;
  assign n32225 = ~n32222 & n32224 ;
  assign n32226 = ( n2638 & ~n9315 ) | ( n2638 & n22737 ) | ( ~n9315 & n22737 ) ;
  assign n32227 = n30915 ^ n9441 ^ 1'b0 ;
  assign n32228 = n8643 | n32227 ;
  assign n32229 = n25323 ^ n23653 ^ 1'b0 ;
  assign n32231 = n24026 ^ n12237 ^ n10333 ;
  assign n32232 = n32231 ^ n24802 ^ n22078 ;
  assign n32230 = ( ~n1783 & n11984 ) | ( ~n1783 & n30319 ) | ( n11984 & n30319 ) ;
  assign n32233 = n32232 ^ n32230 ^ n29826 ;
  assign n32234 = ( n10161 & ~n19240 ) | ( n10161 & n31675 ) | ( ~n19240 & n31675 ) ;
  assign n32235 = n32234 ^ n6151 ^ 1'b0 ;
  assign n32236 = n32235 ^ n19095 ^ n14696 ;
  assign n32237 = n2041 & n12464 ;
  assign n32238 = ~n16793 & n32237 ;
  assign n32239 = n32238 ^ n13458 ^ n3868 ;
  assign n32245 = n28901 ^ n7120 ^ n4952 ;
  assign n32241 = n5324 & ~n6865 ;
  assign n32242 = n32241 ^ n9789 ^ n5878 ;
  assign n32243 = ( n1310 & n18006 ) | ( n1310 & n32242 ) | ( n18006 & n32242 ) ;
  assign n32240 = ( n2766 & ~n23069 ) | ( n2766 & n28643 ) | ( ~n23069 & n28643 ) ;
  assign n32244 = n32243 ^ n32240 ^ n8188 ;
  assign n32246 = n32245 ^ n32244 ^ n27834 ;
  assign n32247 = n24383 ^ n7322 ^ 1'b0 ;
  assign n32248 = ~n5956 & n24125 ;
  assign n32249 = ( ~n26178 & n26273 ) | ( ~n26178 & n32248 ) | ( n26273 & n32248 ) ;
  assign n32250 = ~n1144 & n3271 ;
  assign n32251 = ~n7832 & n32250 ;
  assign n32252 = ( n25160 & ~n28838 ) | ( n25160 & n32251 ) | ( ~n28838 & n32251 ) ;
  assign n32253 = n4408 | n13796 ;
  assign n32254 = n10920 | n32253 ;
  assign n32255 = n12398 & ~n18836 ;
  assign n32256 = ~n32254 & n32255 ;
  assign n32257 = n32256 ^ n25408 ^ 1'b0 ;
  assign n32258 = n3157 & ~n32257 ;
  assign n32259 = n25857 ^ n20643 ^ 1'b0 ;
  assign n32260 = n16436 & n32259 ;
  assign n32265 = ( n13100 & n13150 ) | ( n13100 & n17649 ) | ( n13150 & n17649 ) ;
  assign n32266 = n32265 ^ n23409 ^ n9911 ;
  assign n32261 = ( n3200 & n3410 ) | ( n3200 & ~n14523 ) | ( n3410 & ~n14523 ) ;
  assign n32262 = ( ~n5214 & n12450 ) | ( ~n5214 & n22765 ) | ( n12450 & n22765 ) ;
  assign n32263 = n15962 ^ n12910 ^ n2903 ;
  assign n32264 = ( n32261 & n32262 ) | ( n32261 & ~n32263 ) | ( n32262 & ~n32263 ) ;
  assign n32267 = n32266 ^ n32264 ^ n16971 ;
  assign n32268 = n32267 ^ n15589 ^ 1'b0 ;
  assign n32269 = n11794 ^ n5466 ^ 1'b0 ;
  assign n32270 = ( n1582 & n1588 ) | ( n1582 & ~n4826 ) | ( n1588 & ~n4826 ) ;
  assign n32271 = ( n23798 & n28752 ) | ( n23798 & n32270 ) | ( n28752 & n32270 ) ;
  assign n32272 = ( ~n21526 & n32269 ) | ( ~n21526 & n32271 ) | ( n32269 & n32271 ) ;
  assign n32273 = ( n1256 & n6210 ) | ( n1256 & ~n9344 ) | ( n6210 & ~n9344 ) ;
  assign n32274 = n32273 ^ n20105 ^ n348 ;
  assign n32275 = n9436 | n27686 ;
  assign n32276 = n23653 & ~n32275 ;
  assign n32277 = n21245 ^ n14431 ^ n11789 ;
  assign n32278 = n20462 ^ n641 ^ 1'b0 ;
  assign n32279 = ~n32277 & n32278 ;
  assign n32280 = n4538 | n16446 ;
  assign n32281 = n32280 ^ n17775 ^ 1'b0 ;
  assign n32282 = n32281 ^ n26998 ^ n17299 ;
  assign n32283 = n32282 ^ n22233 ^ n6682 ;
  assign n32284 = n5496 & n9945 ;
  assign n32285 = n28760 & n32284 ;
  assign n32292 = n2343 & ~n17773 ;
  assign n32293 = n8947 & n32292 ;
  assign n32289 = ~n3734 & n11397 ;
  assign n32290 = n32289 ^ n21920 ^ 1'b0 ;
  assign n32291 = n7469 & ~n32290 ;
  assign n32294 = n32293 ^ n32291 ^ n7411 ;
  assign n32286 = n13396 ^ n8294 ^ n7971 ;
  assign n32287 = n32286 ^ n20515 ^ n7522 ;
  assign n32288 = ( n9614 & n25582 ) | ( n9614 & ~n32287 ) | ( n25582 & ~n32287 ) ;
  assign n32295 = n32294 ^ n32288 ^ n21040 ;
  assign n32296 = n32295 ^ n26856 ^ 1'b0 ;
  assign n32297 = n3865 | n32296 ;
  assign n32298 = n12559 ^ n3597 ^ n622 ;
  assign n32299 = n26067 ^ n1068 ^ 1'b0 ;
  assign n32300 = ( n15255 & ~n18203 ) | ( n15255 & n22861 ) | ( ~n18203 & n22861 ) ;
  assign n32304 = n19626 ^ n4384 ^ n1748 ;
  assign n32305 = n32304 ^ n20329 ^ n4431 ;
  assign n32301 = n8430 & ~n22174 ;
  assign n32302 = n20320 & n32301 ;
  assign n32303 = n32302 ^ n6166 ^ 1'b0 ;
  assign n32306 = n32305 ^ n32303 ^ n10058 ;
  assign n32307 = n17029 & ~n30424 ;
  assign n32308 = n5506 ^ n2477 ^ 1'b0 ;
  assign n32309 = ~n27573 & n32308 ;
  assign n32310 = n6359 ^ n2548 ^ n2205 ;
  assign n32311 = ( n12855 & n28911 ) | ( n12855 & ~n32310 ) | ( n28911 & ~n32310 ) ;
  assign n32312 = ( x4 & n11476 ) | ( x4 & ~n13220 ) | ( n11476 & ~n13220 ) ;
  assign n32313 = ( n1750 & n17056 ) | ( n1750 & n32312 ) | ( n17056 & n32312 ) ;
  assign n32314 = n26324 ^ n20748 ^ 1'b0 ;
  assign n32315 = n19730 | n32314 ;
  assign n32316 = n16771 ^ n7539 ^ 1'b0 ;
  assign n32317 = n27617 & ~n32316 ;
  assign n32318 = n23950 & n32317 ;
  assign n32319 = n32318 ^ n24839 ^ 1'b0 ;
  assign n32320 = n18733 ^ n13034 ^ n278 ;
  assign n32321 = n32320 ^ n7505 ^ 1'b0 ;
  assign n32322 = ~n32319 & n32321 ;
  assign n32323 = n13615 ^ n9393 ^ 1'b0 ;
  assign n32324 = ~n10251 & n30565 ;
  assign n32325 = n32323 & n32324 ;
  assign n32326 = n28259 ^ n13466 ^ n2674 ;
  assign n32327 = n5877 ^ n2997 ^ 1'b0 ;
  assign n32328 = n13799 ^ n3128 ^ n515 ;
  assign n32329 = n32328 ^ n6571 ^ 1'b0 ;
  assign n32330 = n14148 & ~n25025 ;
  assign n32332 = n12368 ^ n2341 ^ 1'b0 ;
  assign n32331 = n3423 & ~n13610 ;
  assign n32333 = n32332 ^ n32331 ^ 1'b0 ;
  assign n32334 = n14926 & ~n32333 ;
  assign n32335 = n32334 ^ n4735 ^ 1'b0 ;
  assign n32336 = n8569 | n18828 ;
  assign n32337 = n32336 ^ n25004 ^ 1'b0 ;
  assign n32338 = ( n1528 & ~n5352 ) | ( n1528 & n14017 ) | ( ~n5352 & n14017 ) ;
  assign n32343 = n21010 ^ n17100 ^ 1'b0 ;
  assign n32339 = n3182 & ~n23865 ;
  assign n32340 = n32339 ^ n21348 ^ 1'b0 ;
  assign n32341 = n32340 ^ n22907 ^ n3235 ;
  assign n32342 = ( n11065 & n20603 ) | ( n11065 & ~n32341 ) | ( n20603 & ~n32341 ) ;
  assign n32344 = n32343 ^ n32342 ^ n8557 ;
  assign n32345 = n28665 ^ n10037 ^ 1'b0 ;
  assign n32346 = n23133 & n32345 ;
  assign n32347 = ( ~n10943 & n20816 ) | ( ~n10943 & n24086 ) | ( n20816 & n24086 ) ;
  assign n32348 = ~n3785 & n10778 ;
  assign n32349 = ( ~n3408 & n10309 ) | ( ~n3408 & n26335 ) | ( n10309 & n26335 ) ;
  assign n32350 = ~n7778 & n21661 ;
  assign n32351 = ( n8901 & n18182 ) | ( n8901 & n32350 ) | ( n18182 & n32350 ) ;
  assign n32352 = n14069 & ~n32351 ;
  assign n32353 = n16595 ^ n8233 ^ 1'b0 ;
  assign n32354 = n3990 | n32353 ;
  assign n32355 = n32354 ^ n20619 ^ n9086 ;
  assign n32356 = ~n17730 & n25395 ;
  assign n32357 = n32356 ^ n15955 ^ 1'b0 ;
  assign n32358 = ( n12691 & n32355 ) | ( n12691 & ~n32357 ) | ( n32355 & ~n32357 ) ;
  assign n32359 = ~n6965 & n26937 ;
  assign n32360 = n32359 ^ n27065 ^ 1'b0 ;
  assign n32361 = ( n4180 & n9780 ) | ( n4180 & ~n12409 ) | ( n9780 & ~n12409 ) ;
  assign n32362 = n32361 ^ n11312 ^ n7256 ;
  assign n32363 = n14794 ^ n9065 ^ 1'b0 ;
  assign n32364 = ( ~n7907 & n32362 ) | ( ~n7907 & n32363 ) | ( n32362 & n32363 ) ;
  assign n32365 = n21226 ^ n10862 ^ 1'b0 ;
  assign n32366 = n6809 & n32365 ;
  assign n32367 = ( x222 & n16697 ) | ( x222 & ~n31645 ) | ( n16697 & ~n31645 ) ;
  assign n32368 = n1070 & n10958 ;
  assign n32369 = n32368 ^ n8644 ^ 1'b0 ;
  assign n32370 = n32367 & ~n32369 ;
  assign n32371 = ( n27914 & n32366 ) | ( n27914 & n32370 ) | ( n32366 & n32370 ) ;
  assign n32380 = n10662 & n25296 ;
  assign n32381 = ~n11682 & n32380 ;
  assign n32372 = n882 & ~n7622 ;
  assign n32373 = n310 & n32372 ;
  assign n32374 = ~n325 & n7803 ;
  assign n32375 = n32374 ^ n4106 ^ 1'b0 ;
  assign n32376 = n32375 ^ x49 ^ 1'b0 ;
  assign n32377 = ( n9370 & n30306 ) | ( n9370 & ~n32376 ) | ( n30306 & ~n32376 ) ;
  assign n32378 = ~n32373 & n32377 ;
  assign n32379 = ~n20071 & n32378 ;
  assign n32382 = n32381 ^ n32379 ^ n27399 ;
  assign n32383 = n32185 ^ n28547 ^ n4040 ;
  assign n32384 = ~n2083 & n5482 ;
  assign n32385 = n32384 ^ n18980 ^ 1'b0 ;
  assign n32386 = ( n1421 & ~n7349 ) | ( n1421 & n12193 ) | ( ~n7349 & n12193 ) ;
  assign n32387 = ~n31839 & n32386 ;
  assign n32388 = ~n21259 & n32387 ;
  assign n32389 = n10414 ^ n6593 ^ n5828 ;
  assign n32390 = n32389 ^ n31942 ^ n18172 ;
  assign n32391 = n23644 ^ n681 ^ 1'b0 ;
  assign n32392 = n7341 | n32391 ;
  assign n32393 = ( n1700 & n32230 ) | ( n1700 & ~n32392 ) | ( n32230 & ~n32392 ) ;
  assign n32394 = n32393 ^ n13143 ^ n12603 ;
  assign n32395 = n8537 & ~n19233 ;
  assign n32396 = n32395 ^ n21494 ^ n4925 ;
  assign n32397 = n27220 ^ n11553 ^ 1'b0 ;
  assign n32398 = ~n9701 & n32397 ;
  assign n32399 = n6027 & n32398 ;
  assign n32400 = n3305 | n11183 ;
  assign n32401 = n1757 & n30179 ;
  assign n32402 = n18120 | n32401 ;
  assign n32403 = n13586 & n15253 ;
  assign n32404 = ~n32402 & n32403 ;
  assign n32405 = n14931 ^ n11536 ^ 1'b0 ;
  assign n32406 = n32405 ^ n27111 ^ 1'b0 ;
  assign n32407 = n32404 | n32406 ;
  assign n32408 = n14058 ^ n3333 ^ n1877 ;
  assign n32409 = n12367 ^ n12143 ^ n7788 ;
  assign n32410 = n32409 ^ n21115 ^ n8092 ;
  assign n32411 = n14515 ^ n5511 ^ n1808 ;
  assign n32412 = n32411 ^ n20351 ^ 1'b0 ;
  assign n32416 = n24088 ^ n20221 ^ n16591 ;
  assign n32413 = ~n3249 & n21908 ;
  assign n32414 = n32413 ^ x164 ^ 1'b0 ;
  assign n32415 = n32414 ^ n18689 ^ n15274 ;
  assign n32417 = n32416 ^ n32415 ^ n3287 ;
  assign n32418 = ( n22188 & n27207 ) | ( n22188 & ~n28007 ) | ( n27207 & ~n28007 ) ;
  assign n32420 = ( n1198 & n5055 ) | ( n1198 & n10139 ) | ( n5055 & n10139 ) ;
  assign n32419 = n723 & ~n6878 ;
  assign n32421 = n32420 ^ n32419 ^ 1'b0 ;
  assign n32422 = n4593 ^ n4419 ^ 1'b0 ;
  assign n32423 = n32421 | n32422 ;
  assign n32424 = n738 | n32423 ;
  assign n32425 = ( ~n12516 & n20254 ) | ( ~n12516 & n31986 ) | ( n20254 & n31986 ) ;
  assign n32426 = n32425 ^ n3904 ^ 1'b0 ;
  assign n32427 = ( x73 & n14281 ) | ( x73 & n32426 ) | ( n14281 & n32426 ) ;
  assign n32428 = n18946 ^ n7882 ^ n5727 ;
  assign n32429 = ( ~n1032 & n2222 ) | ( ~n1032 & n5072 ) | ( n2222 & n5072 ) ;
  assign n32430 = n3437 & ~n8147 ;
  assign n32431 = ( n32428 & ~n32429 ) | ( n32428 & n32430 ) | ( ~n32429 & n32430 ) ;
  assign n32432 = ( n6399 & ~n16047 ) | ( n6399 & n32431 ) | ( ~n16047 & n32431 ) ;
  assign n32433 = ~n2183 & n6144 ;
  assign n32434 = n24103 & n32433 ;
  assign n32435 = n18713 & n30141 ;
  assign n32436 = n32354 & n32435 ;
  assign n32437 = ( n31751 & ~n32434 ) | ( n31751 & n32436 ) | ( ~n32434 & n32436 ) ;
  assign n32438 = ( n7492 & n8089 ) | ( n7492 & ~n24230 ) | ( n8089 & ~n24230 ) ;
  assign n32439 = ( n6141 & ~n20536 ) | ( n6141 & n32438 ) | ( ~n20536 & n32438 ) ;
  assign n32440 = n32439 ^ n26464 ^ n2224 ;
  assign n32441 = n11032 ^ n921 ^ 1'b0 ;
  assign n32442 = n5284 & ~n32441 ;
  assign n32443 = n5599 ^ n5002 ^ 1'b0 ;
  assign n32444 = ~n7097 & n32443 ;
  assign n32445 = ( n27242 & n27861 ) | ( n27242 & ~n32444 ) | ( n27861 & ~n32444 ) ;
  assign n32446 = ( n8918 & ~n26642 ) | ( n8918 & n32445 ) | ( ~n26642 & n32445 ) ;
  assign n32447 = ( n29847 & n32442 ) | ( n29847 & ~n32446 ) | ( n32442 & ~n32446 ) ;
  assign n32448 = ~n19110 & n24955 ;
  assign n32449 = n12886 & n17743 ;
  assign n32450 = n2468 & ~n19409 ;
  assign n32451 = n15962 | n23453 ;
  assign n32452 = n7487 & ~n32451 ;
  assign n32453 = x155 & n4487 ;
  assign n32454 = n9058 & ~n32453 ;
  assign n32455 = n11554 & n32454 ;
  assign n32456 = n17215 ^ n4093 ^ 1'b0 ;
  assign n32457 = n24142 ^ n8447 ^ 1'b0 ;
  assign n32458 = n14246 ^ n977 ^ 1'b0 ;
  assign n32459 = n17999 | n32458 ;
  assign n32460 = n32459 ^ n797 ^ 1'b0 ;
  assign n32461 = n12239 ^ n9594 ^ n6888 ;
  assign n32462 = ( n6469 & n6494 ) | ( n6469 & ~n32461 ) | ( n6494 & ~n32461 ) ;
  assign n32463 = n11938 & ~n28925 ;
  assign n32464 = n32463 ^ n10822 ^ 1'b0 ;
  assign n32468 = n10152 ^ n9454 ^ n2163 ;
  assign n32465 = ( ~n2926 & n10952 ) | ( ~n2926 & n11110 ) | ( n10952 & n11110 ) ;
  assign n32466 = n3284 & n32465 ;
  assign n32467 = n32466 ^ n2070 ^ 1'b0 ;
  assign n32469 = n32468 ^ n32467 ^ n24859 ;
  assign n32470 = n24175 ^ n18642 ^ n5176 ;
  assign n32471 = n32470 ^ n31832 ^ n15121 ;
  assign n32472 = n32471 ^ n7516 ^ 1'b0 ;
  assign n32473 = ( ~n32464 & n32469 ) | ( ~n32464 & n32472 ) | ( n32469 & n32472 ) ;
  assign n32477 = n29141 ^ n25674 ^ n18361 ;
  assign n32478 = n32477 ^ n30887 ^ 1'b0 ;
  assign n32479 = n449 | n32478 ;
  assign n32474 = n20339 ^ n18527 ^ n11889 ;
  assign n32475 = n32474 ^ n14446 ^ n1695 ;
  assign n32476 = n32475 ^ n13196 ^ n1629 ;
  assign n32480 = n32479 ^ n32476 ^ n13982 ;
  assign n32481 = x21 & n1976 ;
  assign n32482 = n32481 ^ n17378 ^ 1'b0 ;
  assign n32483 = n9267 ^ n2417 ^ 1'b0 ;
  assign n32484 = n32483 ^ n15945 ^ n4147 ;
  assign n32485 = ( n9785 & n21617 ) | ( n9785 & n32484 ) | ( n21617 & n32484 ) ;
  assign n32486 = n32485 ^ n14443 ^ x18 ;
  assign n32487 = n6951 | n17964 ;
  assign n32488 = ( n15925 & n31832 ) | ( n15925 & ~n32487 ) | ( n31832 & ~n32487 ) ;
  assign n32489 = n32488 ^ n15132 ^ n4866 ;
  assign n32490 = n15442 ^ n9883 ^ n6286 ;
  assign n32491 = ( n4217 & ~n15093 ) | ( n4217 & n32490 ) | ( ~n15093 & n32490 ) ;
  assign n32492 = ( ~n1062 & n3496 ) | ( ~n1062 & n32491 ) | ( n3496 & n32491 ) ;
  assign n32493 = ( n505 & ~n4636 ) | ( n505 & n27631 ) | ( ~n4636 & n27631 ) ;
  assign n32494 = ( n3999 & ~n24123 ) | ( n3999 & n32493 ) | ( ~n24123 & n32493 ) ;
  assign n32495 = ( ~n6975 & n17526 ) | ( ~n6975 & n18432 ) | ( n17526 & n18432 ) ;
  assign n32496 = ( n6663 & ~n31017 ) | ( n6663 & n32495 ) | ( ~n31017 & n32495 ) ;
  assign n32497 = n18188 ^ n2661 ^ 1'b0 ;
  assign n32498 = n1359 & ~n32497 ;
  assign n32499 = n5611 & n32498 ;
  assign n32500 = n12056 ^ n5795 ^ n3276 ;
  assign n32501 = n32500 ^ n1087 ^ 1'b0 ;
  assign n32502 = ( n1500 & n21816 ) | ( n1500 & n23010 ) | ( n21816 & n23010 ) ;
  assign n32503 = ~n8911 & n32502 ;
  assign n32504 = n21452 | n32503 ;
  assign n32505 = n32472 & ~n32504 ;
  assign n32506 = n32501 & n32505 ;
  assign n32507 = n5185 & ~n13938 ;
  assign n32508 = ( n23446 & n31462 ) | ( n23446 & n32507 ) | ( n31462 & n32507 ) ;
  assign n32509 = n7153 & ~n29225 ;
  assign n32510 = n13813 ^ n4640 ^ 1'b0 ;
  assign n32511 = n32510 ^ n30149 ^ n8456 ;
  assign n32512 = n20642 ^ n9596 ^ 1'b0 ;
  assign n32513 = ( n2356 & n15795 ) | ( n2356 & n17486 ) | ( n15795 & n17486 ) ;
  assign n32514 = n19219 | n32513 ;
  assign n32515 = n19591 & ~n32514 ;
  assign n32516 = n32515 ^ n14463 ^ 1'b0 ;
  assign n32517 = n27689 ^ n13675 ^ n12510 ;
  assign n32518 = n18980 ^ n17880 ^ 1'b0 ;
  assign n32519 = n32517 | n32518 ;
  assign n32520 = n5669 & n6577 ;
  assign n32521 = n32520 ^ n8790 ^ 1'b0 ;
  assign n32522 = ( x81 & n21332 ) | ( x81 & n28653 ) | ( n21332 & n28653 ) ;
  assign n32523 = n4697 ^ n2589 ^ 1'b0 ;
  assign n32525 = n22325 ^ n17319 ^ n2971 ;
  assign n32524 = n13284 | n18571 ;
  assign n32526 = n32525 ^ n32524 ^ 1'b0 ;
  assign n32527 = ( n4507 & n6552 ) | ( n4507 & ~n17900 ) | ( n6552 & ~n17900 ) ;
  assign n32528 = ( n2099 & ~n8383 ) | ( n2099 & n32527 ) | ( ~n8383 & n32527 ) ;
  assign n32529 = n32528 ^ n2801 ^ 1'b0 ;
  assign n32530 = n10617 ^ n2475 ^ 1'b0 ;
  assign n32531 = n32530 ^ n6669 ^ n6474 ;
  assign n32532 = n17040 ^ n8956 ^ n2597 ;
  assign n32533 = n25160 ^ n8530 ^ n5475 ;
  assign n32534 = n27841 & ~n32533 ;
  assign n32535 = n32532 & ~n32534 ;
  assign n32536 = ~n8045 & n32535 ;
  assign n32537 = ( n5480 & n21609 ) | ( n5480 & ~n32536 ) | ( n21609 & ~n32536 ) ;
  assign n32541 = ( x240 & n2083 ) | ( x240 & ~n11526 ) | ( n2083 & ~n11526 ) ;
  assign n32538 = n4494 ^ n1675 ^ 1'b0 ;
  assign n32539 = n3452 & n32538 ;
  assign n32540 = n32539 ^ n7313 ^ n3885 ;
  assign n32542 = n32541 ^ n32540 ^ 1'b0 ;
  assign n32543 = n6547 | n6840 ;
  assign n32544 = n1143 & ~n32543 ;
  assign n32545 = n32544 ^ n23003 ^ n1945 ;
  assign n32546 = n1399 & n26613 ;
  assign n32547 = n32546 ^ n17536 ^ 1'b0 ;
  assign n32548 = ( n16731 & ~n30860 ) | ( n16731 & n32547 ) | ( ~n30860 & n32547 ) ;
  assign n32549 = n12016 ^ n906 ^ 1'b0 ;
  assign n32550 = ( n5293 & n16187 ) | ( n5293 & n17027 ) | ( n16187 & n17027 ) ;
  assign n32551 = ( n22456 & n32420 ) | ( n22456 & ~n32550 ) | ( n32420 & ~n32550 ) ;
  assign n32552 = n6301 | n24024 ;
  assign n32553 = n32551 | n32552 ;
  assign n32554 = n23856 ^ n9040 ^ n1580 ;
  assign n32555 = n21255 ^ n19669 ^ n5924 ;
  assign n32556 = n10332 ^ n5854 ^ n1496 ;
  assign n32557 = ( n15988 & ~n32555 ) | ( n15988 & n32556 ) | ( ~n32555 & n32556 ) ;
  assign n32558 = n32557 ^ n8992 ^ n2205 ;
  assign n32559 = ( n2708 & n10951 ) | ( n2708 & n12658 ) | ( n10951 & n12658 ) ;
  assign n32560 = n29910 & ~n32559 ;
  assign n32561 = ~n330 & n32560 ;
  assign n32562 = ( n11766 & n28355 ) | ( n11766 & ~n32561 ) | ( n28355 & ~n32561 ) ;
  assign n32563 = ( n17519 & n18395 ) | ( n17519 & n26586 ) | ( n18395 & n26586 ) ;
  assign n32564 = ( ~n3204 & n10317 ) | ( ~n3204 & n11631 ) | ( n10317 & n11631 ) ;
  assign n32565 = n32564 ^ n11424 ^ 1'b0 ;
  assign n32566 = n19606 ^ n6889 ^ 1'b0 ;
  assign n32567 = n32565 & n32566 ;
  assign n32568 = n10548 & ~n32567 ;
  assign n32569 = ( n1040 & n19017 ) | ( n1040 & n32568 ) | ( n19017 & n32568 ) ;
  assign n32572 = n3872 & ~n7132 ;
  assign n32571 = n18971 | n19255 ;
  assign n32573 = n32572 ^ n32571 ^ 1'b0 ;
  assign n32570 = n28859 ^ n15155 ^ n2315 ;
  assign n32574 = n32573 ^ n32570 ^ n2021 ;
  assign n32575 = n27686 ^ n21915 ^ 1'b0 ;
  assign n32576 = n32574 | n32575 ;
  assign n32577 = n16513 ^ n15047 ^ n4048 ;
  assign n32578 = ( n1500 & ~n16701 ) | ( n1500 & n32577 ) | ( ~n16701 & n32577 ) ;
  assign n32580 = n26452 ^ n5387 ^ 1'b0 ;
  assign n32581 = n18117 & ~n32580 ;
  assign n32579 = n30644 ^ n14204 ^ n8481 ;
  assign n32582 = n32581 ^ n32579 ^ n5640 ;
  assign n32583 = ( n5679 & n20449 ) | ( n5679 & ~n32582 ) | ( n20449 & ~n32582 ) ;
  assign n32584 = n11889 ^ n10664 ^ 1'b0 ;
  assign n32585 = n6006 & ~n14291 ;
  assign n32586 = n32585 ^ n10834 ^ 1'b0 ;
  assign n32587 = n11238 ^ n9650 ^ n573 ;
  assign n32588 = ~n23943 & n32587 ;
  assign n32589 = ~n32586 & n32588 ;
  assign n32590 = n25397 ^ n13226 ^ n9313 ;
  assign n32591 = n18642 ^ n7632 ^ n6728 ;
  assign n32592 = n5998 | n18150 ;
  assign n32593 = n21359 & ~n32592 ;
  assign n32594 = n32593 ^ n23537 ^ 1'b0 ;
  assign n32595 = ( n21172 & n32591 ) | ( n21172 & ~n32594 ) | ( n32591 & ~n32594 ) ;
  assign n32596 = ( n14421 & n29019 ) | ( n14421 & n32595 ) | ( n29019 & n32595 ) ;
  assign n32597 = ( n355 & n16348 ) | ( n355 & n25039 ) | ( n16348 & n25039 ) ;
  assign n32598 = ( ~n12439 & n15354 ) | ( ~n12439 & n18108 ) | ( n15354 & n18108 ) ;
  assign n32599 = ( n1995 & n32597 ) | ( n1995 & ~n32598 ) | ( n32597 & ~n32598 ) ;
  assign n32600 = n22557 & n32599 ;
  assign n32601 = n17983 ^ n17697 ^ n5138 ;
  assign n32604 = n2859 ^ n2488 ^ 1'b0 ;
  assign n32605 = ~n29935 & n32604 ;
  assign n32606 = n32605 ^ n5370 ^ n2621 ;
  assign n32607 = ( n591 & ~n1446 ) | ( n591 & n32606 ) | ( ~n1446 & n32606 ) ;
  assign n32602 = n20324 ^ n7937 ^ 1'b0 ;
  assign n32603 = ~n6496 & n32602 ;
  assign n32608 = n32607 ^ n32603 ^ 1'b0 ;
  assign n32609 = n7139 | n17869 ;
  assign n32610 = ( ~n5660 & n5757 ) | ( ~n5660 & n7903 ) | ( n5757 & n7903 ) ;
  assign n32611 = n32610 ^ n5026 ^ 1'b0 ;
  assign n32612 = n5945 & n32611 ;
  assign n32613 = n12045 | n14917 ;
  assign n32614 = n32613 ^ n26531 ^ 1'b0 ;
  assign n32615 = n856 | n32614 ;
  assign n32616 = ( n4502 & ~n32612 ) | ( n4502 & n32615 ) | ( ~n32612 & n32615 ) ;
  assign n32617 = n26566 ^ n10298 ^ n7827 ;
  assign n32618 = ( ~n21747 & n26444 ) | ( ~n21747 & n32617 ) | ( n26444 & n32617 ) ;
  assign n32619 = n32618 ^ n30193 ^ n2794 ;
  assign n32620 = n29802 ^ n24305 ^ n15370 ;
  assign n32621 = ( n7478 & n28218 ) | ( n7478 & ~n32620 ) | ( n28218 & ~n32620 ) ;
  assign n32623 = ( n4702 & n7745 ) | ( n4702 & ~n11483 ) | ( n7745 & ~n11483 ) ;
  assign n32622 = n26912 ^ n15531 ^ n8696 ;
  assign n32624 = n32623 ^ n32622 ^ n10540 ;
  assign n32625 = ( n9433 & n28161 ) | ( n9433 & n32624 ) | ( n28161 & n32624 ) ;
  assign n32626 = ( n4024 & ~n7163 ) | ( n4024 & n8686 ) | ( ~n7163 & n8686 ) ;
  assign n32627 = x17 & ~n32626 ;
  assign n32628 = n1532 | n28022 ;
  assign n32629 = n6508 & ~n16773 ;
  assign n32630 = n32629 ^ n25833 ^ n16509 ;
  assign n32631 = ( n13090 & ~n25056 ) | ( n13090 & n32630 ) | ( ~n25056 & n32630 ) ;
  assign n32633 = n11596 ^ n9350 ^ n6234 ;
  assign n32634 = ( n5330 & n23990 ) | ( n5330 & ~n32633 ) | ( n23990 & ~n32633 ) ;
  assign n32632 = n15498 | n18753 ;
  assign n32635 = n32634 ^ n32632 ^ 1'b0 ;
  assign n32636 = n32635 ^ n26959 ^ n5090 ;
  assign n32637 = n14187 & n26514 ;
  assign n32638 = n16196 | n32637 ;
  assign n32639 = n32638 ^ n21848 ^ 1'b0 ;
  assign n32640 = n22568 ^ n20494 ^ 1'b0 ;
  assign n32641 = n32639 & n32640 ;
  assign n32642 = n18071 ^ n15628 ^ n2203 ;
  assign n32643 = n32642 ^ n27030 ^ n2089 ;
  assign n32644 = ( ~n32636 & n32641 ) | ( ~n32636 & n32643 ) | ( n32641 & n32643 ) ;
  assign n32645 = n26952 ^ n25772 ^ n25193 ;
  assign n32646 = n9903 ^ n6204 ^ 1'b0 ;
  assign n32647 = n11255 & n18537 ;
  assign n32648 = n32647 ^ n10660 ^ 1'b0 ;
  assign n32649 = ( ~n7382 & n23535 ) | ( ~n7382 & n24044 ) | ( n23535 & n24044 ) ;
  assign n32650 = n32649 ^ n1339 ^ 1'b0 ;
  assign n32651 = n9008 & n32650 ;
  assign n32652 = n32651 ^ n6010 ^ 1'b0 ;
  assign n32653 = n3555 & n13901 ;
  assign n32654 = ( ~n1221 & n22982 ) | ( ~n1221 & n32653 ) | ( n22982 & n32653 ) ;
  assign n32655 = ( n8446 & ~n9639 ) | ( n8446 & n32654 ) | ( ~n9639 & n32654 ) ;
  assign n32656 = n24197 ^ n16391 ^ 1'b0 ;
  assign n32657 = ( n25599 & n26309 ) | ( n25599 & ~n32656 ) | ( n26309 & ~n32656 ) ;
  assign n32658 = n2664 & ~n15858 ;
  assign n32659 = n32658 ^ n21003 ^ 1'b0 ;
  assign n32660 = ( n9679 & n17730 ) | ( n9679 & ~n32659 ) | ( n17730 & ~n32659 ) ;
  assign n32661 = ( n22490 & n24078 ) | ( n22490 & ~n32660 ) | ( n24078 & ~n32660 ) ;
  assign n32662 = n16493 ^ n4644 ^ x161 ;
  assign n32663 = n27171 ^ n12808 ^ n3577 ;
  assign n32664 = ~n23151 & n32663 ;
  assign n32665 = ( ~n17289 & n32662 ) | ( ~n17289 & n32664 ) | ( n32662 & n32664 ) ;
  assign n32666 = n13631 ^ n11529 ^ n7072 ;
  assign n32667 = n6762 | n32666 ;
  assign n32669 = ~n958 & n9125 ;
  assign n32670 = n22087 & n32669 ;
  assign n32668 = ( n6760 & ~n11657 ) | ( n6760 & n23074 ) | ( ~n11657 & n23074 ) ;
  assign n32671 = n32670 ^ n32668 ^ n1860 ;
  assign n32672 = ( n1165 & ~n11847 ) | ( n1165 & n32671 ) | ( ~n11847 & n32671 ) ;
  assign n32673 = ~n9018 & n12988 ;
  assign n32674 = n28554 ^ n6776 ^ 1'b0 ;
  assign n32675 = n32674 ^ n17966 ^ 1'b0 ;
  assign n32678 = n11884 & n15247 ;
  assign n32676 = n26335 ^ n14652 ^ n6558 ;
  assign n32677 = ( x63 & n23341 ) | ( x63 & ~n32676 ) | ( n23341 & ~n32676 ) ;
  assign n32679 = n32678 ^ n32677 ^ n5331 ;
  assign n32680 = n29492 ^ n22413 ^ n12787 ;
  assign n32681 = n772 & n11356 ;
  assign n32682 = n5478 & n32681 ;
  assign n32683 = n18979 ^ n7488 ^ 1'b0 ;
  assign n32684 = n6850 & n32683 ;
  assign n32685 = n18778 ^ n16927 ^ n7136 ;
  assign n32686 = n32685 ^ n27577 ^ n17583 ;
  assign n32689 = ~n3865 & n20576 ;
  assign n32690 = n32689 ^ n13384 ^ 1'b0 ;
  assign n32687 = n30361 ^ n10186 ^ 1'b0 ;
  assign n32688 = ( n26969 & ~n27739 ) | ( n26969 & n32687 ) | ( ~n27739 & n32687 ) ;
  assign n32691 = n32690 ^ n32688 ^ n25228 ;
  assign n32692 = ( n341 & n1452 ) | ( n341 & n9083 ) | ( n1452 & n9083 ) ;
  assign n32693 = n18242 & ~n32692 ;
  assign n32694 = n26438 ^ n5994 ^ 1'b0 ;
  assign n32695 = n5024 & ~n6307 ;
  assign n32696 = n7085 ^ n4498 ^ 1'b0 ;
  assign n32697 = n1856 & n32696 ;
  assign n32699 = n9914 & n17265 ;
  assign n32700 = n1127 & n32699 ;
  assign n32698 = ( ~n3025 & n8193 ) | ( ~n3025 & n23904 ) | ( n8193 & n23904 ) ;
  assign n32701 = n32700 ^ n32698 ^ n25972 ;
  assign n32702 = x10 & ~n20395 ;
  assign n32703 = n32702 ^ n24203 ^ n20015 ;
  assign n32704 = ( ~n2627 & n2939 ) | ( ~n2627 & n32703 ) | ( n2939 & n32703 ) ;
  assign n32706 = n14495 | n27046 ;
  assign n32707 = n32706 ^ n19960 ^ n10939 ;
  assign n32705 = n31495 ^ n13008 ^ n7554 ;
  assign n32708 = n32707 ^ n32705 ^ 1'b0 ;
  assign n32709 = n15898 & n32708 ;
  assign n32710 = n11183 ^ n9458 ^ n1243 ;
  assign n32711 = ( n6745 & n26034 ) | ( n6745 & n32710 ) | ( n26034 & n32710 ) ;
  assign n32712 = n16139 ^ n13823 ^ n11999 ;
  assign n32713 = n32712 ^ n2363 ^ 1'b0 ;
  assign n32714 = ( ~n2907 & n14857 ) | ( ~n2907 & n32713 ) | ( n14857 & n32713 ) ;
  assign n32715 = n32714 ^ n21181 ^ n16766 ;
  assign n32716 = n14681 ^ n13338 ^ n10998 ;
  assign n32717 = ( n331 & n26062 ) | ( n331 & n32716 ) | ( n26062 & n32716 ) ;
  assign n32718 = ( ~n22787 & n24643 ) | ( ~n22787 & n25896 ) | ( n24643 & n25896 ) ;
  assign n32719 = ( n6457 & n8012 ) | ( n6457 & ~n22397 ) | ( n8012 & ~n22397 ) ;
  assign n32720 = n32719 ^ n20301 ^ n5829 ;
  assign n32721 = n32720 ^ n20208 ^ 1'b0 ;
  assign n32722 = n24573 & ~n32721 ;
  assign n32723 = n18601 ^ n13110 ^ n3529 ;
  assign n32724 = n24727 & ~n32723 ;
  assign n32725 = n32724 ^ n27202 ^ 1'b0 ;
  assign n32726 = n32720 ^ n12777 ^ n8374 ;
  assign n32727 = n3644 ^ n3529 ^ 1'b0 ;
  assign n32728 = n5524 & ~n32727 ;
  assign n32729 = n32728 ^ n18149 ^ n11896 ;
  assign n32730 = n32729 ^ n27881 ^ n25314 ;
  assign n32731 = n32730 ^ n2894 ^ 1'b0 ;
  assign n32732 = ~n32726 & n32731 ;
  assign n32733 = n18967 & ~n22180 ;
  assign n32734 = n29827 ^ n16660 ^ n5802 ;
  assign n32735 = n26571 ^ x134 ^ 1'b0 ;
  assign n32736 = n12373 ^ n5576 ^ 1'b0 ;
  assign n32737 = ~n8136 & n32736 ;
  assign n32738 = n28228 ^ n4570 ^ 1'b0 ;
  assign n32739 = n24317 ^ n16998 ^ n4375 ;
  assign n32740 = n13045 ^ n9605 ^ n708 ;
  assign n32741 = n16184 | n32740 ;
  assign n32742 = n32741 ^ n4792 ^ n3288 ;
  assign n32747 = ~n9997 & n19226 ;
  assign n32744 = n8067 ^ n5828 ^ 1'b0 ;
  assign n32745 = n4661 & ~n32744 ;
  assign n32743 = n26701 ^ n25198 ^ n7843 ;
  assign n32746 = n32745 ^ n32743 ^ n18909 ;
  assign n32748 = n32747 ^ n32746 ^ n26693 ;
  assign n32749 = n10519 | n32748 ;
  assign n32750 = n2573 | n32749 ;
  assign n32751 = n29955 ^ n13928 ^ n11496 ;
  assign n32754 = n1480 & ~n20340 ;
  assign n32755 = n2880 & n32754 ;
  assign n32752 = n20380 ^ n17760 ^ 1'b0 ;
  assign n32753 = ( n11115 & n15450 ) | ( n11115 & ~n32752 ) | ( n15450 & ~n32752 ) ;
  assign n32756 = n32755 ^ n32753 ^ 1'b0 ;
  assign n32757 = n32751 & n32756 ;
  assign n32758 = n3962 & ~n12322 ;
  assign n32759 = n32758 ^ n29002 ^ 1'b0 ;
  assign n32760 = ( n5880 & ~n6052 ) | ( n5880 & n28755 ) | ( ~n6052 & n28755 ) ;
  assign n32761 = n24815 ^ n9851 ^ n3782 ;
  assign n32762 = n32761 ^ n12019 ^ n7460 ;
  assign n32763 = n3701 ^ n1611 ^ 1'b0 ;
  assign n32764 = n16358 ^ n14097 ^ n9528 ;
  assign n32765 = n9106 & ~n22372 ;
  assign n32766 = ~n10264 & n32765 ;
  assign n32767 = n32766 ^ x64 ^ 1'b0 ;
  assign n32768 = n32764 | n32767 ;
  assign n32769 = ( n1826 & n2041 ) | ( n1826 & ~n9484 ) | ( n2041 & ~n9484 ) ;
  assign n32770 = n11384 ^ n1132 ^ x236 ;
  assign n32771 = ( n8864 & ~n12284 ) | ( n8864 & n32770 ) | ( ~n12284 & n32770 ) ;
  assign n32772 = n32771 ^ n4501 ^ x215 ;
  assign n32773 = n32772 ^ n15229 ^ 1'b0 ;
  assign n32774 = n32769 & ~n32773 ;
  assign n32775 = n6675 & ~n12066 ;
  assign n32776 = ~n13245 & n32775 ;
  assign n32777 = x128 & ~n29935 ;
  assign n32778 = n32777 ^ n802 ^ 1'b0 ;
  assign n32779 = n9238 ^ n6541 ^ n4971 ;
  assign n32780 = n25483 & ~n32779 ;
  assign n32781 = ~n13443 & n31604 ;
  assign n32782 = n32781 ^ n26720 ^ 1'b0 ;
  assign n32783 = n32533 & n32782 ;
  assign n32784 = ~n17426 & n30112 ;
  assign n32785 = n28067 ^ n27336 ^ 1'b0 ;
  assign n32786 = n22242 & n32785 ;
  assign n32787 = n549 | n11226 ;
  assign n32788 = n9144 | n32787 ;
  assign n32789 = ( n19575 & ~n28597 ) | ( n19575 & n32788 ) | ( ~n28597 & n32788 ) ;
  assign n32790 = ( n740 & ~n4529 ) | ( n740 & n25876 ) | ( ~n4529 & n25876 ) ;
  assign n32791 = n32790 ^ n25468 ^ 1'b0 ;
  assign n32792 = n23840 ^ n21165 ^ n7910 ;
  assign n32793 = n16237 ^ n4897 ^ 1'b0 ;
  assign n32794 = ( n2334 & n3217 ) | ( n2334 & ~n25120 ) | ( n3217 & ~n25120 ) ;
  assign n32795 = ( n4933 & n29991 ) | ( n4933 & n32794 ) | ( n29991 & n32794 ) ;
  assign n32796 = n14144 ^ n12566 ^ n2816 ;
  assign n32797 = n32796 ^ n22859 ^ 1'b0 ;
  assign n32798 = n26665 ^ n17150 ^ n3092 ;
  assign n32799 = ~n21958 & n32798 ;
  assign n32800 = n15873 ^ n2336 ^ 1'b0 ;
  assign n32801 = n9701 | n32800 ;
  assign n32802 = ( ~x104 & n6737 ) | ( ~x104 & n32801 ) | ( n6737 & n32801 ) ;
  assign n32803 = ~n18552 & n32802 ;
  assign n32806 = n7832 & n13066 ;
  assign n32807 = n32806 ^ n29529 ^ 1'b0 ;
  assign n32808 = n1570 | n15147 ;
  assign n32809 = n32807 & ~n32808 ;
  assign n32804 = n16993 ^ n13034 ^ 1'b0 ;
  assign n32805 = ~n22710 & n32804 ;
  assign n32810 = n32809 ^ n32805 ^ n12236 ;
  assign n32811 = n32595 ^ n20438 ^ n9597 ;
  assign n32812 = n32811 ^ n17751 ^ 1'b0 ;
  assign n32813 = n27637 ^ n1042 ^ n895 ;
  assign n32814 = n14516 ^ n12627 ^ n8537 ;
  assign n32815 = n5464 & n8598 ;
  assign n32816 = n5053 & n19845 ;
  assign n32817 = n13583 & n32816 ;
  assign n32818 = n5660 & n22573 ;
  assign n32819 = ~n15090 & n32818 ;
  assign n32820 = ( n2804 & ~n17276 ) | ( n2804 & n32819 ) | ( ~n17276 & n32819 ) ;
  assign n32821 = n6459 | n32820 ;
  assign n32822 = n23940 | n32821 ;
  assign n32823 = n14006 ^ n9067 ^ n3945 ;
  assign n32824 = n15608 ^ n10611 ^ 1'b0 ;
  assign n32825 = n32823 | n32824 ;
  assign n32826 = ( n4384 & ~n4456 ) | ( n4384 & n11374 ) | ( ~n4456 & n11374 ) ;
  assign n32827 = n32826 ^ n3383 ^ x21 ;
  assign n32828 = n27653 ^ n6922 ^ n2648 ;
  assign n32829 = ( n28422 & n32827 ) | ( n28422 & n32828 ) | ( n32827 & n32828 ) ;
  assign n32830 = ( ~n1500 & n32825 ) | ( ~n1500 & n32829 ) | ( n32825 & n32829 ) ;
  assign n32831 = n4844 & n32493 ;
  assign n32835 = ( ~n23272 & n25813 ) | ( ~n23272 & n31646 ) | ( n25813 & n31646 ) ;
  assign n32833 = ( ~n6062 & n6295 ) | ( ~n6062 & n24381 ) | ( n6295 & n24381 ) ;
  assign n32832 = n18872 ^ n12208 ^ n10334 ;
  assign n32834 = n32833 ^ n32832 ^ 1'b0 ;
  assign n32836 = n32835 ^ n32834 ^ n6077 ;
  assign n32837 = n14445 ^ n10531 ^ 1'b0 ;
  assign n32838 = n32837 ^ n11584 ^ 1'b0 ;
  assign n32839 = n24019 & n32838 ;
  assign n32840 = ( n3309 & n7322 ) | ( n3309 & n21304 ) | ( n7322 & n21304 ) ;
  assign n32841 = n12221 ^ n11920 ^ n8472 ;
  assign n32842 = n32415 ^ n24878 ^ n14620 ;
  assign n32843 = n16186 ^ n7828 ^ n2388 ;
  assign n32844 = ( ~n7382 & n27976 ) | ( ~n7382 & n32843 ) | ( n27976 & n32843 ) ;
  assign n32845 = n5464 | n20647 ;
  assign n32846 = n25998 & ~n32845 ;
  assign n32847 = ( n12153 & n22790 ) | ( n12153 & ~n32846 ) | ( n22790 & ~n32846 ) ;
  assign n32848 = ~n1681 & n32847 ;
  assign n32849 = n2422 & n32848 ;
  assign n32850 = ~n12817 & n18512 ;
  assign n32851 = ( ~n2910 & n11591 ) | ( ~n2910 & n25596 ) | ( n11591 & n25596 ) ;
  assign n32852 = n32851 ^ n12476 ^ n11158 ;
  assign n32853 = n32852 ^ n6771 ^ 1'b0 ;
  assign n32854 = n32853 ^ n24099 ^ n1884 ;
  assign n32855 = ~n7990 & n9070 ;
  assign n32856 = n32855 ^ n1087 ^ 1'b0 ;
  assign n32857 = n21018 ^ n10017 ^ 1'b0 ;
  assign n32858 = n32857 ^ n27669 ^ n20827 ;
  assign n32859 = ( n14016 & n32856 ) | ( n14016 & ~n32858 ) | ( n32856 & ~n32858 ) ;
  assign n32860 = n2350 & ~n5274 ;
  assign n32861 = n32860 ^ n23018 ^ n17487 ;
  assign n32862 = n32861 ^ n21469 ^ 1'b0 ;
  assign n32863 = n8253 & ~n32862 ;
  assign n32864 = n14043 & n21457 ;
  assign n32865 = n32864 ^ n2694 ^ 1'b0 ;
  assign n32866 = ( n7389 & n9064 ) | ( n7389 & n32865 ) | ( n9064 & n32865 ) ;
  assign n32867 = n13852 ^ n7272 ^ 1'b0 ;
  assign n32868 = n2599 | n32867 ;
  assign n32869 = n16047 ^ n14175 ^ n9028 ;
  assign n32870 = ( n19412 & n32868 ) | ( n19412 & ~n32869 ) | ( n32868 & ~n32869 ) ;
  assign n32871 = n24407 ^ n14280 ^ 1'b0 ;
  assign n32872 = n32871 ^ n25273 ^ n11005 ;
  assign n32873 = ( n15010 & n25641 ) | ( n15010 & n32872 ) | ( n25641 & n32872 ) ;
  assign n32875 = n31255 ^ n5789 ^ n1578 ;
  assign n32874 = n31291 ^ n18141 ^ n13031 ;
  assign n32876 = n32875 ^ n32874 ^ n24136 ;
  assign n32877 = n12999 ^ n9137 ^ n5630 ;
  assign n32878 = n27396 ^ n14668 ^ 1'b0 ;
  assign n32879 = n32877 & ~n32878 ;
  assign n32880 = ( n11170 & n22831 ) | ( n11170 & ~n32879 ) | ( n22831 & ~n32879 ) ;
  assign n32881 = n6755 ^ n995 ^ n350 ;
  assign n32882 = n32881 ^ n21050 ^ n9892 ;
  assign n32883 = n32882 ^ n32151 ^ n3895 ;
  assign n32884 = n32883 ^ n20369 ^ n13532 ;
  assign n32886 = n24624 ^ n5595 ^ 1'b0 ;
  assign n32885 = n13505 & ~n30247 ;
  assign n32887 = n32886 ^ n32885 ^ 1'b0 ;
  assign n32888 = n1636 | n8367 ;
  assign n32889 = n22450 | n32888 ;
  assign n32890 = n32889 ^ n29132 ^ n3050 ;
  assign n32891 = ( n12392 & n18701 ) | ( n12392 & ~n32890 ) | ( n18701 & ~n32890 ) ;
  assign n32892 = n8621 ^ n8085 ^ 1'b0 ;
  assign n32893 = n1990 & ~n32892 ;
  assign n32894 = n32893 ^ n28026 ^ n4170 ;
  assign n32895 = ( n975 & n3592 ) | ( n975 & ~n21681 ) | ( n3592 & ~n21681 ) ;
  assign n32896 = n32895 ^ n27302 ^ n5124 ;
  assign n32897 = n667 | n32896 ;
  assign n32898 = n15289 | n32897 ;
  assign n32899 = ( n5080 & n8547 ) | ( n5080 & n25693 ) | ( n8547 & n25693 ) ;
  assign n32900 = ( n8697 & n26231 ) | ( n8697 & n32899 ) | ( n26231 & n32899 ) ;
  assign n32901 = n32900 ^ n30666 ^ n3415 ;
  assign n32902 = ~n9829 & n32901 ;
  assign n32903 = ( n10895 & ~n29671 ) | ( n10895 & n32902 ) | ( ~n29671 & n32902 ) ;
  assign n32904 = ( n7764 & n11280 ) | ( n7764 & n13478 ) | ( n11280 & n13478 ) ;
  assign n32905 = ~n1508 & n19491 ;
  assign n32906 = n32905 ^ n20371 ^ 1'b0 ;
  assign n32907 = n7124 | n32906 ;
  assign n32908 = ( ~n4539 & n12677 ) | ( ~n4539 & n32907 ) | ( n12677 & n32907 ) ;
  assign n32909 = ( n13073 & n23671 ) | ( n13073 & n24816 ) | ( n23671 & n24816 ) ;
  assign n32910 = ( n7711 & n24246 ) | ( n7711 & ~n32909 ) | ( n24246 & ~n32909 ) ;
  assign n32912 = n19606 ^ n10114 ^ n4126 ;
  assign n32911 = ( n3619 & ~n8569 ) | ( n3619 & n32263 ) | ( ~n8569 & n32263 ) ;
  assign n32913 = n32912 ^ n32911 ^ n18453 ;
  assign n32914 = n4010 ^ n3335 ^ 1'b0 ;
  assign n32915 = n30139 & ~n32914 ;
  assign n32916 = ~n32913 & n32915 ;
  assign n32917 = n32916 ^ n27117 ^ 1'b0 ;
  assign n32919 = ( n2059 & ~n4300 ) | ( n2059 & n14745 ) | ( ~n4300 & n14745 ) ;
  assign n32918 = n438 & n14773 ;
  assign n32920 = n32919 ^ n32918 ^ 1'b0 ;
  assign n32922 = n26729 ^ n13803 ^ n7942 ;
  assign n32921 = n32317 ^ n26103 ^ n8248 ;
  assign n32923 = n32922 ^ n32921 ^ n3016 ;
  assign n32924 = ( n13607 & n26373 ) | ( n13607 & ~n32923 ) | ( n26373 & ~n32923 ) ;
  assign n32925 = n20744 ^ n2369 ^ n566 ;
  assign n32927 = n9063 ^ n534 ^ n526 ;
  assign n32928 = ( n17583 & ~n19902 ) | ( n17583 & n32927 ) | ( ~n19902 & n32927 ) ;
  assign n32926 = n30903 ^ n30877 ^ n29629 ;
  assign n32929 = n32928 ^ n32926 ^ n15411 ;
  assign n32930 = n3775 ^ n1713 ^ x203 ;
  assign n32931 = ( n5172 & n21274 ) | ( n5172 & ~n32930 ) | ( n21274 & ~n32930 ) ;
  assign n32935 = n12334 ^ n5184 ^ n959 ;
  assign n32937 = n23253 ^ n18733 ^ n3901 ;
  assign n32938 = ( ~n4771 & n19869 ) | ( ~n4771 & n32937 ) | ( n19869 & n32937 ) ;
  assign n32936 = ~n7869 & n9180 ;
  assign n32939 = n32938 ^ n32936 ^ 1'b0 ;
  assign n32940 = ( ~n11271 & n15100 ) | ( ~n11271 & n32939 ) | ( n15100 & n32939 ) ;
  assign n32941 = n25810 & ~n32940 ;
  assign n32942 = n32941 ^ n30348 ^ 1'b0 ;
  assign n32943 = n32935 & ~n32942 ;
  assign n32932 = n13100 ^ n5044 ^ 1'b0 ;
  assign n32933 = n10998 ^ n2328 ^ 1'b0 ;
  assign n32934 = ( ~n23975 & n32932 ) | ( ~n23975 & n32933 ) | ( n32932 & n32933 ) ;
  assign n32944 = n32943 ^ n32934 ^ 1'b0 ;
  assign n32945 = ~n18585 & n32944 ;
  assign n32946 = ( n5668 & n7193 ) | ( n5668 & ~n15776 ) | ( n7193 & ~n15776 ) ;
  assign n32947 = ( n15425 & n20635 ) | ( n15425 & n32946 ) | ( n20635 & n32946 ) ;
  assign n32948 = ( n511 & n1999 ) | ( n511 & ~n13533 ) | ( n1999 & ~n13533 ) ;
  assign n32949 = n32948 ^ n17683 ^ n2777 ;
  assign n32950 = n8646 & ~n9813 ;
  assign n32951 = n22401 ^ n17183 ^ n3213 ;
  assign n32952 = n8009 & n24608 ;
  assign n32953 = ~n32951 & n32952 ;
  assign n32954 = ~n1629 & n9416 ;
  assign n32955 = n27363 ^ n19175 ^ 1'b0 ;
  assign n32956 = ~n32954 & n32955 ;
  assign n32957 = ( ~n18615 & n32953 ) | ( ~n18615 & n32956 ) | ( n32953 & n32956 ) ;
  assign n32958 = n32809 ^ n27263 ^ x225 ;
  assign n32959 = ( n349 & ~n27577 ) | ( n349 & n32958 ) | ( ~n27577 & n32958 ) ;
  assign n32960 = n10287 ^ n6663 ^ 1'b0 ;
  assign n32961 = n26697 | n32960 ;
  assign n32962 = n32961 ^ n5585 ^ 1'b0 ;
  assign n32963 = n10635 & ~n17477 ;
  assign n32964 = ( n20788 & ~n24048 ) | ( n20788 & n31291 ) | ( ~n24048 & n31291 ) ;
  assign n32965 = n7188 & n13006 ;
  assign n32966 = n32965 ^ n7108 ^ 1'b0 ;
  assign n32967 = ~n32232 & n32966 ;
  assign n32968 = n2598 & n32967 ;
  assign n32969 = ( ~n15727 & n22015 ) | ( ~n15727 & n22030 ) | ( n22015 & n22030 ) ;
  assign n32970 = n28584 ^ n25087 ^ n14127 ;
  assign n32971 = n8430 | n16273 ;
  assign n32972 = ( n26562 & n28020 ) | ( n26562 & ~n32971 ) | ( n28020 & ~n32971 ) ;
  assign n32973 = n25173 ^ n20623 ^ n19792 ;
  assign n32974 = n6478 ^ n3909 ^ 1'b0 ;
  assign n32975 = n32973 & ~n32974 ;
  assign n32978 = ( n6582 & n9941 ) | ( n6582 & ~n17732 ) | ( n9941 & ~n17732 ) ;
  assign n32976 = n19404 ^ n4373 ^ n336 ;
  assign n32977 = n11694 & n32976 ;
  assign n32979 = n32978 ^ n32977 ^ 1'b0 ;
  assign n32980 = x126 & ~n6103 ;
  assign n32981 = n32980 ^ n2859 ^ 1'b0 ;
  assign n32982 = ( n1392 & n4352 ) | ( n1392 & ~n20330 ) | ( n4352 & ~n20330 ) ;
  assign n32983 = ( n11756 & n32981 ) | ( n11756 & n32982 ) | ( n32981 & n32982 ) ;
  assign n32984 = n28451 ^ n21338 ^ n1710 ;
  assign n32986 = n13603 ^ n1973 ^ 1'b0 ;
  assign n32985 = ( n18566 & ~n24744 ) | ( n18566 & n31077 ) | ( ~n24744 & n31077 ) ;
  assign n32987 = n32986 ^ n32985 ^ 1'b0 ;
  assign n32988 = ( n3317 & ~n7167 ) | ( n3317 & n18873 ) | ( ~n7167 & n18873 ) ;
  assign n32989 = ( n5939 & n13686 ) | ( n5939 & ~n16758 ) | ( n13686 & ~n16758 ) ;
  assign n32990 = n19684 | n32989 ;
  assign n32991 = n32990 ^ n12045 ^ 1'b0 ;
  assign n32992 = n32991 ^ n15965 ^ n7299 ;
  assign n32993 = ( n4507 & n14084 ) | ( n4507 & ~n23983 ) | ( n14084 & ~n23983 ) ;
  assign n32994 = ~n6872 & n32993 ;
  assign n32995 = ~n6933 & n32994 ;
  assign n32996 = ( ~n20707 & n27926 ) | ( ~n20707 & n32995 ) | ( n27926 & n32995 ) ;
  assign n32997 = n17682 ^ n4192 ^ n3642 ;
  assign n32998 = n981 & n5964 ;
  assign n32999 = n1433 & n32998 ;
  assign n33000 = ( n1625 & ~n7742 ) | ( n1625 & n32999 ) | ( ~n7742 & n32999 ) ;
  assign n33001 = ( n11128 & n13960 ) | ( n11128 & n20853 ) | ( n13960 & n20853 ) ;
  assign n33002 = n33000 & ~n33001 ;
  assign n33003 = ~n18904 & n24863 ;
  assign n33004 = n9431 | n33003 ;
  assign n33005 = n31438 & ~n33004 ;
  assign n33006 = n9746 & ~n33005 ;
  assign n33007 = n28039 ^ n20669 ^ 1'b0 ;
  assign n33008 = n7473 ^ n846 ^ 1'b0 ;
  assign n33009 = n33008 ^ n14170 ^ n6292 ;
  assign n33010 = n33009 ^ n17686 ^ n14135 ;
  assign n33011 = n11608 & n16370 ;
  assign n33012 = n33011 ^ n12412 ^ n2392 ;
  assign n33013 = n7442 ^ n5787 ^ 1'b0 ;
  assign n33014 = n33013 ^ n8606 ^ n1741 ;
  assign n33015 = ( n12878 & n33012 ) | ( n12878 & n33014 ) | ( n33012 & n33014 ) ;
  assign n33016 = n16949 | n30842 ;
  assign n33017 = n33016 ^ n7149 ^ 1'b0 ;
  assign n33018 = n33017 ^ n13236 ^ n3193 ;
  assign n33019 = n26274 ^ n15850 ^ n1728 ;
  assign n33020 = ( n4042 & n4476 ) | ( n4042 & n33019 ) | ( n4476 & n33019 ) ;
  assign n33021 = n33018 & n33020 ;
  assign n33022 = n5640 & ~n33002 ;
  assign n33023 = ( n1902 & n29097 ) | ( n1902 & ~n33022 ) | ( n29097 & ~n33022 ) ;
  assign n33024 = ( n3508 & ~n6043 ) | ( n3508 & n11244 ) | ( ~n6043 & n11244 ) ;
  assign n33025 = n33024 ^ n2892 ^ 1'b0 ;
  assign n33026 = n7405 & ~n20441 ;
  assign n33027 = n33026 ^ n1205 ^ 1'b0 ;
  assign n33028 = n12151 ^ n12121 ^ 1'b0 ;
  assign n33029 = n5209 & n25023 ;
  assign n33030 = n33028 & n33029 ;
  assign n33031 = n12188 ^ x68 ^ 1'b0 ;
  assign n33032 = n33031 ^ n14344 ^ n5976 ;
  assign n33033 = n9869 ^ n8335 ^ n6437 ;
  assign n33034 = n33033 ^ n15368 ^ n12277 ;
  assign n33035 = n9009 | n17303 ;
  assign n33036 = n10384 & ~n33035 ;
  assign n33038 = ( ~n4150 & n8371 ) | ( ~n4150 & n13674 ) | ( n8371 & n13674 ) ;
  assign n33037 = ~n9580 & n24335 ;
  assign n33039 = n33038 ^ n33037 ^ n29569 ;
  assign n33040 = ~n1022 & n10780 ;
  assign n33041 = n33040 ^ n8772 ^ 1'b0 ;
  assign n33042 = n33041 ^ n6769 ^ 1'b0 ;
  assign n33043 = ~n1597 & n33042 ;
  assign n33044 = n33043 ^ n13757 ^ n7317 ;
  assign n33045 = n1958 & ~n33044 ;
  assign n33046 = ~n1529 & n33045 ;
  assign n33047 = n33046 ^ n19994 ^ 1'b0 ;
  assign n33048 = ~n33039 & n33047 ;
  assign n33049 = ( n4256 & ~n9991 ) | ( n4256 & n21177 ) | ( ~n9991 & n21177 ) ;
  assign n33050 = n18011 ^ n12281 ^ n11384 ;
  assign n33051 = ( n12574 & n33049 ) | ( n12574 & ~n33050 ) | ( n33049 & ~n33050 ) ;
  assign n33052 = n25091 & ~n26530 ;
  assign n33053 = n23056 ^ n20337 ^ 1'b0 ;
  assign n33054 = n2610 ^ x80 ^ 1'b0 ;
  assign n33055 = n9418 & ~n33054 ;
  assign n33056 = n13303 ^ n12630 ^ n11673 ;
  assign n33057 = n33056 ^ n23439 ^ 1'b0 ;
  assign n33058 = ( n6318 & ~n15352 ) | ( n6318 & n29499 ) | ( ~n15352 & n29499 ) ;
  assign n33059 = n8508 ^ n6938 ^ n825 ;
  assign n33060 = ( n7601 & ~n11942 ) | ( n7601 & n25395 ) | ( ~n11942 & n25395 ) ;
  assign n33061 = ( n12809 & n33059 ) | ( n12809 & n33060 ) | ( n33059 & n33060 ) ;
  assign n33062 = n33061 ^ n12699 ^ n10180 ;
  assign n33063 = ( ~n775 & n3390 ) | ( ~n775 & n11455 ) | ( n3390 & n11455 ) ;
  assign n33064 = n28226 ^ n20899 ^ n14712 ;
  assign n33065 = ( n8254 & n33063 ) | ( n8254 & n33064 ) | ( n33063 & n33064 ) ;
  assign n33066 = n12557 ^ n4126 ^ 1'b0 ;
  assign n33067 = ( ~n11501 & n16013 ) | ( ~n11501 & n33066 ) | ( n16013 & n33066 ) ;
  assign n33068 = n33067 ^ n23720 ^ 1'b0 ;
  assign n33069 = n27984 & ~n33068 ;
  assign n33070 = n9670 & ~n23593 ;
  assign n33071 = ( n9278 & ~n9877 ) | ( n9278 & n33070 ) | ( ~n9877 & n33070 ) ;
  assign n33072 = n13350 & n17324 ;
  assign n33073 = n14231 ^ n6373 ^ n2171 ;
  assign n33074 = n33073 ^ n27839 ^ n15626 ;
  assign n33075 = n33074 ^ n32127 ^ n11165 ;
  assign n33076 = n23115 ^ n20434 ^ 1'b0 ;
  assign n33077 = n33076 ^ n22198 ^ n11120 ;
  assign n33078 = ( n6164 & n32179 ) | ( n6164 & n33077 ) | ( n32179 & n33077 ) ;
  assign n33080 = n20538 ^ n802 ^ 1'b0 ;
  assign n33079 = n31328 ^ n17753 ^ n17516 ;
  assign n33081 = n33080 ^ n33079 ^ n19043 ;
  assign n33082 = n18994 ^ n2473 ^ 1'b0 ;
  assign n33084 = ( n6834 & n7546 ) | ( n6834 & n19621 ) | ( n7546 & n19621 ) ;
  assign n33085 = n10442 & ~n29731 ;
  assign n33086 = ~n33084 & n33085 ;
  assign n33083 = n23357 ^ n5145 ^ 1'b0 ;
  assign n33087 = n33086 ^ n33083 ^ n3553 ;
  assign n33088 = n739 & ~n10328 ;
  assign n33089 = n10670 & n33088 ;
  assign n33090 = n33089 ^ n5243 ^ 1'b0 ;
  assign n33091 = ( n10701 & n23641 ) | ( n10701 & ~n30381 ) | ( n23641 & ~n30381 ) ;
  assign n33092 = n8352 ^ n7681 ^ n6628 ;
  assign n33093 = n33092 ^ n30887 ^ n22833 ;
  assign n33094 = ( ~n15751 & n31288 ) | ( ~n15751 & n33093 ) | ( n31288 & n33093 ) ;
  assign n33095 = ( n12450 & n14990 ) | ( n12450 & n20853 ) | ( n14990 & n20853 ) ;
  assign n33096 = n33095 ^ n4883 ^ n1273 ;
  assign n33097 = ~n3919 & n8401 ;
  assign n33098 = n13205 | n33097 ;
  assign n33099 = n33098 ^ n29556 ^ 1'b0 ;
  assign n33104 = n2570 | n16081 ;
  assign n33100 = n1992 & n20867 ;
  assign n33101 = n33100 ^ n11820 ^ 1'b0 ;
  assign n33102 = ~n16525 & n33101 ;
  assign n33103 = n33102 ^ n10446 ^ 1'b0 ;
  assign n33105 = n33104 ^ n33103 ^ n28136 ;
  assign n33109 = n13906 ^ n4226 ^ 1'b0 ;
  assign n33110 = n7113 & n33109 ;
  assign n33111 = ~n3874 & n33110 ;
  assign n33112 = ( n5017 & n11703 ) | ( n5017 & ~n33111 ) | ( n11703 & ~n33111 ) ;
  assign n33106 = n16940 ^ n16657 ^ n11389 ;
  assign n33107 = ~n2599 & n33106 ;
  assign n33108 = n33107 ^ n24597 ^ 1'b0 ;
  assign n33113 = n33112 ^ n33108 ^ n8205 ;
  assign n33114 = ~n4558 & n7112 ;
  assign n33115 = ~n5399 & n33114 ;
  assign n33116 = n14299 ^ n11806 ^ 1'b0 ;
  assign n33117 = ~n9306 & n13266 ;
  assign n33118 = n6654 | n33117 ;
  assign n33119 = ( n8705 & n12108 ) | ( n8705 & n13482 ) | ( n12108 & n13482 ) ;
  assign n33120 = ( n24703 & ~n33118 ) | ( n24703 & n33119 ) | ( ~n33118 & n33119 ) ;
  assign n33121 = ( n33115 & ~n33116 ) | ( n33115 & n33120 ) | ( ~n33116 & n33120 ) ;
  assign n33122 = n3358 ^ n1019 ^ 1'b0 ;
  assign n33123 = n2768 & ~n33122 ;
  assign n33126 = n2383 | n8099 ;
  assign n33127 = n12035 & ~n33126 ;
  assign n33128 = n33127 ^ n28664 ^ n5951 ;
  assign n33124 = n25274 ^ n15738 ^ n355 ;
  assign n33125 = n33124 ^ n10918 ^ 1'b0 ;
  assign n33129 = n33128 ^ n33125 ^ n26079 ;
  assign n33130 = n14895 & n31521 ;
  assign n33131 = ( n12759 & ~n27720 ) | ( n12759 & n33130 ) | ( ~n27720 & n33130 ) ;
  assign n33132 = n13558 ^ n3450 ^ 1'b0 ;
  assign n33133 = ( n372 & ~n984 ) | ( n372 & n33132 ) | ( ~n984 & n33132 ) ;
  assign n33134 = n9358 & n27406 ;
  assign n33135 = ( n19619 & ~n33133 ) | ( n19619 & n33134 ) | ( ~n33133 & n33134 ) ;
  assign n33136 = n17526 ^ n12064 ^ 1'b0 ;
  assign n33137 = n28531 ^ n17697 ^ n8043 ;
  assign n33138 = n33137 ^ n11108 ^ n3433 ;
  assign n33139 = ( n4316 & ~n33136 ) | ( n4316 & n33138 ) | ( ~n33136 & n33138 ) ;
  assign n33140 = ~n9660 & n33139 ;
  assign n33141 = ( n28058 & n30666 ) | ( n28058 & n33140 ) | ( n30666 & n33140 ) ;
  assign n33145 = n5847 & n7345 ;
  assign n33146 = n5957 | n33145 ;
  assign n33142 = n25996 ^ n3754 ^ 1'b0 ;
  assign n33143 = ( n9536 & n19518 ) | ( n9536 & n33142 ) | ( n19518 & n33142 ) ;
  assign n33144 = ( n5470 & ~n7525 ) | ( n5470 & n33143 ) | ( ~n7525 & n33143 ) ;
  assign n33147 = n33146 ^ n33144 ^ n15633 ;
  assign n33148 = n24202 ^ n20466 ^ x70 ;
  assign n33149 = n26329 ^ n9100 ^ n3777 ;
  assign n33150 = ( x198 & n2555 ) | ( x198 & ~n12098 ) | ( n2555 & ~n12098 ) ;
  assign n33151 = n16539 ^ n4651 ^ 1'b0 ;
  assign n33152 = n27830 ^ n404 ^ 1'b0 ;
  assign n33153 = n29115 & ~n33152 ;
  assign n33154 = n1957 | n12332 ;
  assign n33155 = n33153 | n33154 ;
  assign n33156 = n5810 ^ x40 ^ 1'b0 ;
  assign n33157 = n33156 ^ n23067 ^ n10362 ;
  assign n33158 = n18538 ^ n15703 ^ n5890 ;
  assign n33159 = n28322 | n28549 ;
  assign n33160 = n24054 & ~n33159 ;
  assign n33161 = n16900 | n31028 ;
  assign n33162 = ( n10593 & n16615 ) | ( n10593 & ~n23134 ) | ( n16615 & ~n23134 ) ;
  assign n33163 = n13596 & n16728 ;
  assign n33164 = n33163 ^ n13016 ^ n6783 ;
  assign n33165 = ~n2777 & n21074 ;
  assign n33166 = n33165 ^ n20438 ^ 1'b0 ;
  assign n33167 = ~n3318 & n33166 ;
  assign n33168 = n22623 ^ n15602 ^ n631 ;
  assign n33169 = x52 | n33168 ;
  assign n33170 = n14649 & n23773 ;
  assign n33171 = ( n6823 & ~n7667 ) | ( n6823 & n27482 ) | ( ~n7667 & n27482 ) ;
  assign n33172 = n20604 & ~n27114 ;
  assign n33173 = n33172 ^ n24186 ^ 1'b0 ;
  assign n33174 = n13823 ^ n9411 ^ n497 ;
  assign n33175 = n33174 ^ n1756 ^ 1'b0 ;
  assign n33176 = x186 & n33175 ;
  assign n33177 = n22443 ^ n11336 ^ 1'b0 ;
  assign n33178 = n33176 & n33177 ;
  assign n33179 = n16973 ^ n4710 ^ 1'b0 ;
  assign n33180 = n33178 & ~n33179 ;
  assign n33181 = n33180 ^ n4188 ^ 1'b0 ;
  assign n33182 = n33173 | n33181 ;
  assign n33183 = ( ~n3164 & n6119 ) | ( ~n3164 & n25818 ) | ( n6119 & n25818 ) ;
  assign n33184 = n6523 & n10373 ;
  assign n33185 = n33184 ^ n9003 ^ 1'b0 ;
  assign n33186 = n33185 ^ n23069 ^ n12535 ;
  assign n33187 = n15519 ^ n7451 ^ n406 ;
  assign n33188 = ( n404 & n13787 ) | ( n404 & ~n17267 ) | ( n13787 & ~n17267 ) ;
  assign n33189 = n33188 ^ n29176 ^ n10233 ;
  assign n33191 = n22218 ^ n10101 ^ n1950 ;
  assign n33190 = ~n30584 & n31298 ;
  assign n33192 = n33191 ^ n33190 ^ 1'b0 ;
  assign n33193 = ( n27526 & n33189 ) | ( n27526 & ~n33192 ) | ( n33189 & ~n33192 ) ;
  assign n33194 = n28722 & n33193 ;
  assign n33195 = n27231 & n33194 ;
  assign n33196 = ~n20131 & n26100 ;
  assign n33197 = n11208 | n25961 ;
  assign n33198 = n15886 & ~n33197 ;
  assign n33199 = ~n14606 & n33198 ;
  assign n33200 = ( n8862 & n12883 ) | ( n8862 & ~n32633 ) | ( n12883 & ~n32633 ) ;
  assign n33201 = n3288 & n33200 ;
  assign n33202 = ( n6687 & n28330 ) | ( n6687 & ~n33201 ) | ( n28330 & ~n33201 ) ;
  assign n33203 = ( ~n3352 & n12800 ) | ( ~n3352 & n33202 ) | ( n12800 & n33202 ) ;
  assign n33204 = ( n7128 & ~n12578 ) | ( n7128 & n33203 ) | ( ~n12578 & n33203 ) ;
  assign n33205 = n15846 & n23571 ;
  assign n33206 = ( ~n15858 & n28521 ) | ( ~n15858 & n33205 ) | ( n28521 & n33205 ) ;
  assign n33207 = n14180 | n20491 ;
  assign n33208 = ~n1487 & n33207 ;
  assign n33209 = n33208 ^ n10973 ^ 1'b0 ;
  assign n33210 = ( ~x6 & n2633 ) | ( ~x6 & n13909 ) | ( n2633 & n13909 ) ;
  assign n33211 = n33210 ^ n4673 ^ 1'b0 ;
  assign n33212 = ( ~n1958 & n10241 ) | ( ~n1958 & n33211 ) | ( n10241 & n33211 ) ;
  assign n33213 = n20216 ^ n12245 ^ n5038 ;
  assign n33214 = n11119 ^ n7293 ^ 1'b0 ;
  assign n33215 = n33214 ^ n14127 ^ 1'b0 ;
  assign n33216 = ( n12853 & ~n14163 ) | ( n12853 & n14308 ) | ( ~n14163 & n14308 ) ;
  assign n33217 = ( n11220 & n12330 ) | ( n11220 & n33216 ) | ( n12330 & n33216 ) ;
  assign n33218 = n33217 ^ n8071 ^ 1'b0 ;
  assign n33219 = ( n10087 & n13457 ) | ( n10087 & ~n15300 ) | ( n13457 & ~n15300 ) ;
  assign n33220 = n2644 & ~n13724 ;
  assign n33221 = ~n33219 & n33220 ;
  assign n33222 = n3482 | n16597 ;
  assign n33223 = ( n24386 & ~n27338 ) | ( n24386 & n33222 ) | ( ~n27338 & n33222 ) ;
  assign n33224 = n25417 | n33223 ;
  assign n33225 = ~n9463 & n25410 ;
  assign n33226 = n33225 ^ n24391 ^ 1'b0 ;
  assign n33227 = n19231 ^ n2410 ^ n754 ;
  assign n33228 = n17215 | n33227 ;
  assign n33229 = ( ~n15309 & n23272 ) | ( ~n15309 & n32926 ) | ( n23272 & n32926 ) ;
  assign n33230 = n9086 & n14434 ;
  assign n33231 = ( n14159 & ~n24444 ) | ( n14159 & n33230 ) | ( ~n24444 & n33230 ) ;
  assign n33232 = n28351 ^ n5618 ^ 1'b0 ;
  assign n33233 = n22812 & ~n33232 ;
  assign n33234 = n21719 & n32465 ;
  assign n33235 = ~n33233 & n33234 ;
  assign n33236 = ( ~n4128 & n5878 ) | ( ~n4128 & n21148 ) | ( n5878 & n21148 ) ;
  assign n33237 = n33236 ^ n17819 ^ n2652 ;
  assign n33238 = n3991 | n22843 ;
  assign n33239 = n33237 & ~n33238 ;
  assign n33240 = ~n16434 & n25432 ;
  assign n33241 = n24600 ^ n22842 ^ n8492 ;
  assign n33244 = ( ~n9900 & n9911 ) | ( ~n9900 & n15941 ) | ( n9911 & n15941 ) ;
  assign n33245 = n33244 ^ n3899 ^ 1'b0 ;
  assign n33242 = n11851 ^ n4427 ^ 1'b0 ;
  assign n33243 = ~n9947 & n33242 ;
  assign n33246 = n33245 ^ n33243 ^ 1'b0 ;
  assign n33247 = n28101 & n33246 ;
  assign n33248 = n33241 & n33247 ;
  assign n33249 = ( ~n18184 & n21005 ) | ( ~n18184 & n33248 ) | ( n21005 & n33248 ) ;
  assign n33251 = n9836 ^ n5259 ^ n4417 ;
  assign n33252 = n33251 ^ n6977 ^ n802 ;
  assign n33253 = n33252 ^ n31127 ^ n5002 ;
  assign n33250 = n7713 ^ n768 ^ 1'b0 ;
  assign n33254 = n33253 ^ n33250 ^ n23806 ;
  assign n33255 = x10 & n17154 ;
  assign n33256 = n18946 & n33255 ;
  assign n33257 = n33256 ^ n27974 ^ 1'b0 ;
  assign n33258 = n27092 & ~n33257 ;
  assign n33259 = n31872 ^ n16517 ^ n10144 ;
  assign n33260 = ( ~n3639 & n8071 ) | ( ~n3639 & n28566 ) | ( n8071 & n28566 ) ;
  assign n33261 = n14292 ^ n3088 ^ 1'b0 ;
  assign n33262 = ~n1324 & n33261 ;
  assign n33263 = n33262 ^ n25787 ^ n13945 ;
  assign n33264 = ( n31250 & ~n33260 ) | ( n31250 & n33263 ) | ( ~n33260 & n33263 ) ;
  assign n33265 = ( n25954 & ~n33259 ) | ( n25954 & n33264 ) | ( ~n33259 & n33264 ) ;
  assign n33266 = n14310 ^ n13675 ^ n12774 ;
  assign n33267 = n15322 ^ n14382 ^ 1'b0 ;
  assign n33268 = n19660 ^ n18251 ^ n16940 ;
  assign n33269 = n33268 ^ n4372 ^ 1'b0 ;
  assign n33270 = n21692 & n33269 ;
  assign n33271 = ( n3365 & n13635 ) | ( n3365 & n21798 ) | ( n13635 & n21798 ) ;
  assign n33272 = n13249 | n19531 ;
  assign n33273 = n33272 ^ n24126 ^ 1'b0 ;
  assign n33274 = ( n16925 & n21945 ) | ( n16925 & ~n33273 ) | ( n21945 & ~n33273 ) ;
  assign n33275 = ( ~n11852 & n33271 ) | ( ~n11852 & n33274 ) | ( n33271 & n33274 ) ;
  assign n33276 = ( ~n25529 & n25629 ) | ( ~n25529 & n27677 ) | ( n25629 & n27677 ) ;
  assign n33277 = n33276 ^ n17550 ^ n308 ;
  assign n33278 = n668 | n3034 ;
  assign n33279 = n3936 ^ n1916 ^ 1'b0 ;
  assign n33280 = ( n1082 & n7726 ) | ( n1082 & ~n33279 ) | ( n7726 & ~n33279 ) ;
  assign n33281 = ( n431 & ~n20738 ) | ( n431 & n28540 ) | ( ~n20738 & n28540 ) ;
  assign n33284 = n23037 ^ n19637 ^ 1'b0 ;
  assign n33283 = n3265 & n14968 ;
  assign n33282 = ( n4139 & n7367 ) | ( n4139 & ~n15330 ) | ( n7367 & ~n15330 ) ;
  assign n33285 = n33284 ^ n33283 ^ n33282 ;
  assign n33286 = ( n3856 & ~n22527 ) | ( n3856 & n33285 ) | ( ~n22527 & n33285 ) ;
  assign n33287 = n860 & ~n9611 ;
  assign n33288 = ~n3309 & n14926 ;
  assign n33289 = n33287 & n33288 ;
  assign n33290 = n1709 | n10274 ;
  assign n33291 = n5443 & ~n33290 ;
  assign n33292 = n33291 ^ n6213 ^ n3999 ;
  assign n33293 = n19566 & n33292 ;
  assign n33294 = n8819 & n18024 ;
  assign n33295 = n33294 ^ n33127 ^ n4477 ;
  assign n33300 = x83 | n3706 ;
  assign n33296 = ( n3556 & ~n7347 ) | ( n3556 & n16692 ) | ( ~n7347 & n16692 ) ;
  assign n33297 = n33296 ^ n15693 ^ n4798 ;
  assign n33298 = n33297 ^ n5852 ^ n558 ;
  assign n33299 = ( n3775 & n23998 ) | ( n3775 & ~n33298 ) | ( n23998 & ~n33298 ) ;
  assign n33301 = n33300 ^ n33299 ^ n6263 ;
  assign n33302 = n15064 ^ n820 ^ 1'b0 ;
  assign n33303 = n5482 & n26627 ;
  assign n33304 = n6979 ^ n6544 ^ 1'b0 ;
  assign n33305 = n3362 & ~n33304 ;
  assign n33306 = n33303 & n33305 ;
  assign n33307 = n33306 ^ n1842 ^ 1'b0 ;
  assign n33308 = n29085 ^ n2076 ^ 1'b0 ;
  assign n33309 = n4830 & n32678 ;
  assign n33310 = ( ~n12479 & n33308 ) | ( ~n12479 & n33309 ) | ( n33308 & n33309 ) ;
  assign n33311 = n12036 & ~n14083 ;
  assign n33312 = n33311 ^ n27286 ^ 1'b0 ;
  assign n33313 = n20025 & n33312 ;
  assign n33314 = ~n7988 & n25575 ;
  assign n33315 = ( n5513 & n13045 ) | ( n5513 & n33314 ) | ( n13045 & n33314 ) ;
  assign n33316 = n24207 ^ n16707 ^ n3998 ;
  assign n33317 = n19348 & ~n33316 ;
  assign n33318 = n27867 & n33317 ;
  assign n33319 = n2696 | n4272 ;
  assign n33320 = n29636 ^ n24444 ^ 1'b0 ;
  assign n33321 = n28936 ^ n16632 ^ n3429 ;
  assign n33322 = n33321 ^ n24500 ^ n912 ;
  assign n33323 = n10892 ^ n2073 ^ 1'b0 ;
  assign n33324 = n33323 ^ n28654 ^ n17473 ;
  assign n33326 = ~n13530 & n15061 ;
  assign n33327 = ( n7480 & n15204 ) | ( n7480 & n33326 ) | ( n15204 & n33326 ) ;
  assign n33328 = n7917 | n33327 ;
  assign n33325 = n8506 ^ n7371 ^ n6484 ;
  assign n33329 = n33328 ^ n33325 ^ n27431 ;
  assign n33330 = n17271 ^ n17247 ^ 1'b0 ;
  assign n33331 = n5860 & n33330 ;
  assign n33332 = n30438 ^ n5064 ^ 1'b0 ;
  assign n33333 = n866 & ~n33332 ;
  assign n33334 = n7393 & ~n17758 ;
  assign n33335 = n8386 ^ n2922 ^ 1'b0 ;
  assign n33336 = n17175 & n33335 ;
  assign n33337 = n33336 ^ n23521 ^ n10867 ;
  assign n33338 = ~n8720 & n33337 ;
  assign n33339 = ~n33334 & n33338 ;
  assign n33340 = n33339 ^ n27774 ^ n15931 ;
  assign n33341 = n30896 ^ n4670 ^ 1'b0 ;
  assign n33342 = n26122 ^ n6357 ^ 1'b0 ;
  assign n33343 = n13834 & n33342 ;
  assign n33344 = n33343 ^ n20285 ^ n18174 ;
  assign n33345 = n16154 ^ n12806 ^ 1'b0 ;
  assign n33346 = ~n30670 & n33345 ;
  assign n33347 = ( n7254 & n24100 ) | ( n7254 & n33346 ) | ( n24100 & n33346 ) ;
  assign n33348 = n10762 ^ n8156 ^ 1'b0 ;
  assign n33349 = n752 | n33348 ;
  assign n33350 = n8668 & ~n33349 ;
  assign n33351 = n13460 & n14063 ;
  assign n33352 = n12442 & n17278 ;
  assign n33353 = ~n13001 & n33352 ;
  assign n33354 = n28416 | n33353 ;
  assign n33355 = n33351 & ~n33354 ;
  assign n33356 = n22052 ^ n8905 ^ 1'b0 ;
  assign n33357 = ~n23486 & n33356 ;
  assign n33358 = ( n2031 & n24843 ) | ( n2031 & ~n33357 ) | ( n24843 & ~n33357 ) ;
  assign n33361 = n32001 ^ n18251 ^ 1'b0 ;
  assign n33362 = n5482 & n33361 ;
  assign n33360 = n11428 & n13327 ;
  assign n33359 = n6052 | n11211 ;
  assign n33363 = n33362 ^ n33360 ^ n33359 ;
  assign n33369 = n12066 ^ n3826 ^ 1'b0 ;
  assign n33368 = n28684 ^ n8976 ^ n6899 ;
  assign n33364 = n26070 ^ n15535 ^ 1'b0 ;
  assign n33365 = n15786 | n33364 ;
  assign n33366 = n15597 ^ n1587 ^ 1'b0 ;
  assign n33367 = n33365 | n33366 ;
  assign n33370 = n33369 ^ n33368 ^ n33367 ;
  assign n33371 = n25076 ^ n1107 ^ 1'b0 ;
  assign n33372 = n22653 ^ n21111 ^ 1'b0 ;
  assign n33373 = n33371 & n33372 ;
  assign n33374 = ( n28573 & n28628 ) | ( n28573 & ~n33373 ) | ( n28628 & ~n33373 ) ;
  assign n33375 = n1722 ^ n723 ^ n488 ;
  assign n33376 = n33375 ^ n28917 ^ n15207 ;
  assign n33377 = n33376 ^ n11005 ^ 1'b0 ;
  assign n33378 = ~n1403 & n33377 ;
  assign n33379 = n33378 ^ n24130 ^ 1'b0 ;
  assign n33380 = ~n5142 & n33379 ;
  assign n33381 = ( ~n4757 & n5952 ) | ( ~n4757 & n12922 ) | ( n5952 & n12922 ) ;
  assign n33382 = n33381 ^ n13382 ^ n12719 ;
  assign n33383 = n33382 ^ n32886 ^ 1'b0 ;
  assign n33384 = n7986 & ~n33383 ;
  assign n33385 = n22016 ^ n14590 ^ 1'b0 ;
  assign n33386 = n2073 | n33385 ;
  assign n33387 = n14571 ^ n11198 ^ n3130 ;
  assign n33388 = n18000 ^ n8694 ^ 1'b0 ;
  assign n33389 = ~n33387 & n33388 ;
  assign n33390 = n8363 & n33389 ;
  assign n33391 = n33390 ^ n4738 ^ 1'b0 ;
  assign n33392 = n30010 & ~n33391 ;
  assign n33393 = ( n8551 & ~n13989 ) | ( n8551 & n15022 ) | ( ~n13989 & n15022 ) ;
  assign n33394 = n29487 ^ n9283 ^ n1833 ;
  assign n33395 = n7367 & ~n28722 ;
  assign n33396 = n28913 ^ n9835 ^ n2060 ;
  assign n33397 = n18275 & n33396 ;
  assign n33398 = n33397 ^ n23524 ^ n14823 ;
  assign n33399 = n33398 ^ n11107 ^ 1'b0 ;
  assign n33400 = n14945 ^ n3034 ^ 1'b0 ;
  assign n33401 = n23660 | n33400 ;
  assign n33402 = n33401 ^ n28784 ^ n18066 ;
  assign n33403 = n16198 ^ n13474 ^ n2974 ;
  assign n33404 = ( n20691 & n27270 ) | ( n20691 & n33403 ) | ( n27270 & n33403 ) ;
  assign n33405 = n11194 ^ n1783 ^ 1'b0 ;
  assign n33406 = ( n21104 & ~n23810 ) | ( n21104 & n33405 ) | ( ~n23810 & n33405 ) ;
  assign n33407 = ( n2231 & n8012 ) | ( n2231 & n29225 ) | ( n8012 & n29225 ) ;
  assign n33408 = n31984 ^ n1967 ^ 1'b0 ;
  assign n33409 = ~n10434 & n33408 ;
  assign n33414 = ( n3158 & n5188 ) | ( n3158 & n28770 ) | ( n5188 & n28770 ) ;
  assign n33410 = n13883 ^ n11858 ^ n7774 ;
  assign n33411 = n4638 ^ n1476 ^ 1'b0 ;
  assign n33412 = n33410 | n33411 ;
  assign n33413 = n27076 & ~n33412 ;
  assign n33415 = n33414 ^ n33413 ^ 1'b0 ;
  assign n33416 = n25714 ^ n9127 ^ n2663 ;
  assign n33417 = ( n620 & n17833 ) | ( n620 & n22809 ) | ( n17833 & n22809 ) ;
  assign n33418 = ( n7305 & n10033 ) | ( n7305 & ~n20216 ) | ( n10033 & ~n20216 ) ;
  assign n33419 = n4721 | n4869 ;
  assign n33420 = n18330 | n33419 ;
  assign n33421 = n18399 ^ n2948 ^ 1'b0 ;
  assign n33422 = ~n27042 & n33421 ;
  assign n33423 = n19259 ^ n12361 ^ n4182 ;
  assign n33424 = n31223 ^ n22371 ^ n3058 ;
  assign n33425 = n10639 & n12843 ;
  assign n33426 = ( n13921 & n25500 ) | ( n13921 & ~n33425 ) | ( n25500 & ~n33425 ) ;
  assign n33427 = n33426 ^ n11719 ^ n6271 ;
  assign n33428 = n22096 ^ n11547 ^ n5978 ;
  assign n33429 = ( n7167 & ~n10217 ) | ( n7167 & n33428 ) | ( ~n10217 & n33428 ) ;
  assign n33430 = n4156 ^ n4036 ^ 1'b0 ;
  assign n33431 = ( ~n9589 & n15715 ) | ( ~n9589 & n33430 ) | ( n15715 & n33430 ) ;
  assign n33432 = x72 & ~n5746 ;
  assign n33433 = n33432 ^ n9515 ^ 1'b0 ;
  assign n33434 = n5145 & n33433 ;
  assign n33435 = n13384 & n33434 ;
  assign n33436 = ( ~n2988 & n23069 ) | ( ~n2988 & n33435 ) | ( n23069 & n33435 ) ;
  assign n33439 = n4970 ^ n592 ^ 1'b0 ;
  assign n33440 = x72 & n33439 ;
  assign n33441 = ( ~n12015 & n31494 ) | ( ~n12015 & n33440 ) | ( n31494 & n33440 ) ;
  assign n33437 = ( n14575 & n22247 ) | ( n14575 & ~n23995 ) | ( n22247 & ~n23995 ) ;
  assign n33438 = n33437 ^ n29791 ^ n2036 ;
  assign n33442 = n33441 ^ n33438 ^ n4869 ;
  assign n33443 = ( n20844 & n33436 ) | ( n20844 & n33442 ) | ( n33436 & n33442 ) ;
  assign n33444 = n16378 ^ n6490 ^ 1'b0 ;
  assign n33445 = n33444 ^ n25087 ^ n24960 ;
  assign n33446 = n20509 & n24493 ;
  assign n33447 = n6651 & n33446 ;
  assign n33448 = ( ~n1254 & n9927 ) | ( ~n1254 & n14870 ) | ( n9927 & n14870 ) ;
  assign n33449 = ( n5478 & n15881 ) | ( n5478 & n33448 ) | ( n15881 & n33448 ) ;
  assign n33450 = ~n33447 & n33449 ;
  assign n33451 = n10161 & n13284 ;
  assign n33452 = n29062 ^ n20407 ^ n5434 ;
  assign n33453 = ~n453 & n33452 ;
  assign n33454 = ~n33451 & n33453 ;
  assign n33455 = n10973 & n28243 ;
  assign n33459 = n23129 ^ n21220 ^ n8820 ;
  assign n33456 = n28848 ^ n20221 ^ n12376 ;
  assign n33457 = n28554 & n33456 ;
  assign n33458 = n33457 ^ n30680 ^ 1'b0 ;
  assign n33460 = n33459 ^ n33458 ^ n813 ;
  assign n33464 = n12398 ^ n5883 ^ 1'b0 ;
  assign n33461 = n18295 ^ n14062 ^ n405 ;
  assign n33462 = n910 ^ n764 ^ 1'b0 ;
  assign n33463 = n33461 & n33462 ;
  assign n33465 = n33464 ^ n33463 ^ n3230 ;
  assign n33466 = ( n3592 & ~n8328 ) | ( n3592 & n12121 ) | ( ~n8328 & n12121 ) ;
  assign n33467 = n33466 ^ n11082 ^ 1'b0 ;
  assign n33468 = n14921 & ~n28792 ;
  assign n33469 = n33468 ^ n11774 ^ 1'b0 ;
  assign n33470 = ( n8389 & n9839 ) | ( n8389 & ~n20104 ) | ( n9839 & ~n20104 ) ;
  assign n33471 = ( n343 & n8896 ) | ( n343 & ~n14911 ) | ( n8896 & ~n14911 ) ;
  assign n33472 = n19084 | n33471 ;
  assign n33473 = n33470 | n33472 ;
  assign n33474 = n1339 & ~n13935 ;
  assign n33475 = n33474 ^ n17861 ^ 1'b0 ;
  assign n33476 = ~n2043 & n19323 ;
  assign n33477 = n6632 | n33476 ;
  assign n33478 = n33475 | n33477 ;
  assign n33479 = n33478 ^ n16509 ^ n5385 ;
  assign n33480 = n14239 & n33479 ;
  assign n33481 = n33480 ^ n3918 ^ 1'b0 ;
  assign n33482 = n33481 ^ n27610 ^ n25888 ;
  assign n33483 = n12801 ^ n2488 ^ 1'b0 ;
  assign n33484 = ~n16661 & n33483 ;
  assign n33485 = ~n4281 & n33484 ;
  assign n33486 = ~n12151 & n33485 ;
  assign n33487 = ( n19642 & n24108 ) | ( n19642 & ~n33486 ) | ( n24108 & ~n33486 ) ;
  assign n33488 = n30793 ^ n26474 ^ n2377 ;
  assign n33489 = ( ~n890 & n21600 ) | ( ~n890 & n31579 ) | ( n21600 & n31579 ) ;
  assign n33490 = n33489 ^ n15311 ^ n2086 ;
  assign n33491 = n33490 ^ n6337 ^ 1'b0 ;
  assign n33492 = n4752 & n7142 ;
  assign n33493 = ~n27481 & n33492 ;
  assign n33494 = ~n28149 & n33493 ;
  assign n33495 = n20512 ^ n6970 ^ n4205 ;
  assign n33496 = ( n2770 & n11475 ) | ( n2770 & n33495 ) | ( n11475 & n33495 ) ;
  assign n33497 = n33496 ^ n11827 ^ n5462 ;
  assign n33498 = n25109 ^ n24764 ^ n19156 ;
  assign n33499 = n33498 ^ n32629 ^ 1'b0 ;
  assign n33500 = n33499 ^ n33282 ^ n12126 ;
  assign n33501 = n28324 ^ n28274 ^ n15693 ;
  assign n33502 = n33501 ^ n1373 ^ 1'b0 ;
  assign n33503 = ~n11489 & n18030 ;
  assign n33504 = n2052 & ~n11947 ;
  assign n33505 = n33504 ^ n6781 ^ 1'b0 ;
  assign n33506 = n4159 ^ n4120 ^ 1'b0 ;
  assign n33507 = n32528 ^ n3849 ^ n3725 ;
  assign n33508 = ~n27025 & n31932 ;
  assign n33509 = n33508 ^ n6445 ^ 1'b0 ;
  assign n33510 = n18215 & n19387 ;
  assign n33511 = n8236 & n33510 ;
  assign n33514 = ( ~n3557 & n7732 ) | ( ~n3557 & n10137 ) | ( n7732 & n10137 ) ;
  assign n33512 = n1682 & n24392 ;
  assign n33513 = n33512 ^ n8164 ^ 1'b0 ;
  assign n33515 = n33514 ^ n33513 ^ n3579 ;
  assign n33516 = ( n2400 & n14413 ) | ( n2400 & n25532 ) | ( n14413 & n25532 ) ;
  assign n33517 = ~n25328 & n33516 ;
  assign n33518 = ( n5549 & ~n11955 ) | ( n5549 & n33056 ) | ( ~n11955 & n33056 ) ;
  assign n33519 = n10370 ^ n8107 ^ n2720 ;
  assign n33520 = ( n14579 & ~n29354 ) | ( n14579 & n33519 ) | ( ~n29354 & n33519 ) ;
  assign n33521 = ~n19962 & n20373 ;
  assign n33522 = n33521 ^ n27406 ^ 1'b0 ;
  assign n33523 = ( n6619 & n14926 ) | ( n6619 & n30251 ) | ( n14926 & n30251 ) ;
  assign n33524 = n4169 & ~n16782 ;
  assign n33525 = n33524 ^ n28719 ^ 1'b0 ;
  assign n33526 = n33523 & n33525 ;
  assign n33527 = n12617 & n33526 ;
  assign n33528 = n4853 & ~n18771 ;
  assign n33529 = n11962 | n20942 ;
  assign n33530 = ( n9785 & ~n22140 ) | ( n9785 & n33529 ) | ( ~n22140 & n33529 ) ;
  assign n33531 = n11920 & ~n30562 ;
  assign n33532 = n7118 & ~n32008 ;
  assign n33533 = n12899 & ~n33532 ;
  assign n33534 = n8543 ^ n8111 ^ 1'b0 ;
  assign n33535 = ( n1346 & n2828 ) | ( n1346 & n8754 ) | ( n2828 & n8754 ) ;
  assign n33536 = n15583 | n33535 ;
  assign n33537 = n33536 ^ n4467 ^ 1'b0 ;
  assign n33538 = n33537 ^ n23762 ^ 1'b0 ;
  assign n33539 = n23691 & ~n33538 ;
  assign n33540 = n2832 ^ n2474 ^ n1769 ;
  assign n33541 = n2681 | n33540 ;
  assign n33542 = n33539 & ~n33541 ;
  assign n33543 = ( n1695 & n4250 ) | ( n1695 & n6544 ) | ( n4250 & n6544 ) ;
  assign n33544 = ( n14567 & ~n28210 ) | ( n14567 & n33543 ) | ( ~n28210 & n33543 ) ;
  assign n33547 = n3054 | n10364 ;
  assign n33545 = n526 & n3597 ;
  assign n33546 = ( n7574 & n8904 ) | ( n7574 & ~n33545 ) | ( n8904 & ~n33545 ) ;
  assign n33548 = n33547 ^ n33546 ^ n26688 ;
  assign n33549 = ( n5992 & n6861 ) | ( n5992 & n21722 ) | ( n6861 & n21722 ) ;
  assign n33550 = n33549 ^ n17378 ^ n14571 ;
  assign n33552 = n10282 ^ n7002 ^ 1'b0 ;
  assign n33553 = ~n21570 & n33552 ;
  assign n33551 = ~n19822 & n21494 ;
  assign n33554 = n33553 ^ n33551 ^ 1'b0 ;
  assign n33555 = n23106 ^ n16741 ^ n1945 ;
  assign n33556 = ( n15354 & ~n17332 ) | ( n15354 & n19210 ) | ( ~n17332 & n19210 ) ;
  assign n33557 = n33556 ^ n17109 ^ n7809 ;
  assign n33558 = n29169 ^ n8891 ^ 1'b0 ;
  assign n33559 = n20890 ^ n3404 ^ x161 ;
  assign n33560 = ( n33557 & ~n33558 ) | ( n33557 & n33559 ) | ( ~n33558 & n33559 ) ;
  assign n33561 = n14250 ^ n9287 ^ 1'b0 ;
  assign n33568 = n23152 ^ n15155 ^ 1'b0 ;
  assign n33569 = n9972 & ~n33568 ;
  assign n33570 = ( ~n6657 & n13663 ) | ( ~n6657 & n33569 ) | ( n13663 & n33569 ) ;
  assign n33564 = n18397 ^ n8819 ^ n8432 ;
  assign n33562 = n10547 & n14711 ;
  assign n33563 = ~n12058 & n33562 ;
  assign n33565 = n33564 ^ n33563 ^ n3050 ;
  assign n33566 = ( n22556 & n27391 ) | ( n22556 & n33565 ) | ( n27391 & n33565 ) ;
  assign n33567 = n3209 & ~n33566 ;
  assign n33571 = n33570 ^ n33567 ^ 1'b0 ;
  assign n33572 = n33571 ^ n21875 ^ 1'b0 ;
  assign n33573 = n14652 ^ n7495 ^ n4075 ;
  assign n33574 = n33573 ^ n15964 ^ 1'b0 ;
  assign n33575 = n14851 ^ x237 ^ 1'b0 ;
  assign n33576 = n33575 ^ n19239 ^ 1'b0 ;
  assign n33577 = n33576 ^ n13779 ^ n7830 ;
  assign n33578 = n4109 ^ n3483 ^ 1'b0 ;
  assign n33579 = ~n2678 & n33578 ;
  assign n33580 = x221 & n33579 ;
  assign n33581 = n33580 ^ n25662 ^ 1'b0 ;
  assign n33582 = ( n927 & ~n1365 ) | ( n927 & n16207 ) | ( ~n1365 & n16207 ) ;
  assign n33584 = n18644 ^ n17690 ^ 1'b0 ;
  assign n33585 = ( n8603 & ~n23501 ) | ( n8603 & n33584 ) | ( ~n23501 & n33584 ) ;
  assign n33586 = n23726 & n33585 ;
  assign n33587 = n33586 ^ n10612 ^ 1'b0 ;
  assign n33583 = n13100 & n27737 ;
  assign n33588 = n33587 ^ n33583 ^ 1'b0 ;
  assign n33589 = n27072 | n33588 ;
  assign n33592 = n11428 ^ n6833 ^ n3218 ;
  assign n33593 = ( ~n8390 & n11442 ) | ( ~n8390 & n33592 ) | ( n11442 & n33592 ) ;
  assign n33591 = n15822 ^ n14257 ^ n8166 ;
  assign n33590 = n2912 ^ x173 ^ 1'b0 ;
  assign n33594 = n33593 ^ n33591 ^ n33590 ;
  assign n33595 = n4973 ^ n2529 ^ 1'b0 ;
  assign n33596 = ~n17827 & n33595 ;
  assign n33597 = n4570 ^ n2729 ^ 1'b0 ;
  assign n33598 = n33597 ^ n24356 ^ 1'b0 ;
  assign n33599 = ~n2390 & n33598 ;
  assign n33600 = n6401 ^ n4591 ^ n3043 ;
  assign n33601 = n33600 ^ n30553 ^ n4492 ;
  assign n33602 = n7671 & ~n33601 ;
  assign n33603 = n33602 ^ n4303 ^ 1'b0 ;
  assign n33604 = n4566 & n10464 ;
  assign n33605 = n13863 & n33604 ;
  assign n33606 = ( n2089 & ~n33603 ) | ( n2089 & n33605 ) | ( ~n33603 & n33605 ) ;
  assign n33607 = n10514 & n10589 ;
  assign n33608 = n17824 ^ n4487 ^ 1'b0 ;
  assign n33609 = n33608 ^ n31240 ^ n11997 ;
  assign n33610 = ( n2036 & ~n9358 ) | ( n2036 & n10471 ) | ( ~n9358 & n10471 ) ;
  assign n33611 = ( n24084 & n28501 ) | ( n24084 & ~n33610 ) | ( n28501 & ~n33610 ) ;
  assign n33612 = n33611 ^ n27818 ^ 1'b0 ;
  assign n33613 = ~n32861 & n33612 ;
  assign n33614 = n10200 ^ n5421 ^ n5405 ;
  assign n33615 = n33614 ^ n29955 ^ n17342 ;
  assign n33616 = n33615 ^ n29109 ^ n15916 ;
  assign n33617 = ~n8577 & n33616 ;
  assign n33618 = n27232 ^ n22631 ^ n5969 ;
  assign n33620 = ( n8913 & n8916 ) | ( n8913 & n24827 ) | ( n8916 & n24827 ) ;
  assign n33621 = n33620 ^ n13703 ^ 1'b0 ;
  assign n33622 = n13536 & ~n33621 ;
  assign n33619 = ( n1561 & ~n3775 ) | ( n1561 & n5771 ) | ( ~n3775 & n5771 ) ;
  assign n33623 = n33622 ^ n33619 ^ 1'b0 ;
  assign n33624 = ~n2527 & n33101 ;
  assign n33625 = n13086 & n33624 ;
  assign n33626 = n26959 ^ n20821 ^ n19969 ;
  assign n33627 = n10345 | n25488 ;
  assign n33628 = n33627 ^ n12569 ^ 1'b0 ;
  assign n33629 = n14964 ^ n3979 ^ 1'b0 ;
  assign n33630 = ( n3367 & n33139 ) | ( n3367 & ~n33629 ) | ( n33139 & ~n33629 ) ;
  assign n33631 = ( n26907 & n33628 ) | ( n26907 & n33630 ) | ( n33628 & n33630 ) ;
  assign n33634 = n21329 ^ n11409 ^ 1'b0 ;
  assign n33632 = n7703 ^ n849 ^ 1'b0 ;
  assign n33633 = n33632 ^ n24779 ^ n1218 ;
  assign n33635 = n33634 ^ n33633 ^ 1'b0 ;
  assign n33636 = ( n13636 & ~n32846 ) | ( n13636 & n33635 ) | ( ~n32846 & n33635 ) ;
  assign n33637 = n19828 ^ n15582 ^ n6799 ;
  assign n33638 = n4934 & n26373 ;
  assign n33639 = ( n9380 & n33637 ) | ( n9380 & n33638 ) | ( n33637 & n33638 ) ;
  assign n33640 = n8699 | n21993 ;
  assign n33641 = n33640 ^ n27277 ^ 1'b0 ;
  assign n33642 = ~n2083 & n33641 ;
  assign n33643 = n33642 ^ n3274 ^ n619 ;
  assign n33646 = n17299 ^ n15175 ^ n6106 ;
  assign n33644 = n13964 & n14540 ;
  assign n33645 = n16749 & n33644 ;
  assign n33647 = n33646 ^ n33645 ^ n8156 ;
  assign n33648 = n17759 ^ n5965 ^ n3525 ;
  assign n33649 = n11211 ^ n9656 ^ n8169 ;
  assign n33650 = ( ~n13567 & n27108 ) | ( ~n13567 & n33649 ) | ( n27108 & n33649 ) ;
  assign n33651 = ( n10354 & ~n24483 ) | ( n10354 & n29305 ) | ( ~n24483 & n29305 ) ;
  assign n33652 = n32671 ^ n3538 ^ x246 ;
  assign n33653 = ( n33650 & ~n33651 ) | ( n33650 & n33652 ) | ( ~n33651 & n33652 ) ;
  assign n33654 = ( ~x163 & n2208 ) | ( ~x163 & n9030 ) | ( n2208 & n9030 ) ;
  assign n33655 = n14568 & ~n33654 ;
  assign n33656 = n33655 ^ n30686 ^ 1'b0 ;
  assign n33657 = n33656 ^ n9210 ^ 1'b0 ;
  assign n33658 = ( n657 & n19143 ) | ( n657 & ~n21108 ) | ( n19143 & ~n21108 ) ;
  assign n33659 = ( ~n6372 & n30569 ) | ( ~n6372 & n31297 ) | ( n30569 & n31297 ) ;
  assign n33660 = n29588 ^ n25844 ^ n9991 ;
  assign n33661 = ( n18990 & ~n21059 ) | ( n18990 & n24915 ) | ( ~n21059 & n24915 ) ;
  assign n33663 = n8124 | n13114 ;
  assign n33664 = n33663 ^ n8481 ^ 1'b0 ;
  assign n33665 = ( n3430 & n9382 ) | ( n3430 & ~n33664 ) | ( n9382 & ~n33664 ) ;
  assign n33662 = ~n8367 & n9945 ;
  assign n33666 = n33665 ^ n33662 ^ 1'b0 ;
  assign n33667 = ~n16158 & n21812 ;
  assign n33668 = n12282 & n33667 ;
  assign n33669 = n25831 ^ n25827 ^ n6461 ;
  assign n33670 = ( n20773 & n27083 ) | ( n20773 & n33669 ) | ( n27083 & n33669 ) ;
  assign n33671 = n14518 ^ n9670 ^ n3781 ;
  assign n33672 = n33671 ^ n26455 ^ n444 ;
  assign n33673 = ~n11859 & n27417 ;
  assign n33674 = n33673 ^ n14912 ^ 1'b0 ;
  assign n33676 = n7819 ^ n7699 ^ 1'b0 ;
  assign n33675 = n6321 & n8054 ;
  assign n33677 = n33676 ^ n33675 ^ 1'b0 ;
  assign n33678 = ( n2838 & ~n10960 ) | ( n2838 & n20568 ) | ( ~n10960 & n20568 ) ;
  assign n33682 = n21259 ^ n20933 ^ n5688 ;
  assign n33681 = ( n7884 & n9208 ) | ( n7884 & n11967 ) | ( n9208 & n11967 ) ;
  assign n33679 = n11799 ^ n2055 ^ 1'b0 ;
  assign n33680 = n23208 & n33679 ;
  assign n33683 = n33682 ^ n33681 ^ n33680 ;
  assign n33684 = n6996 | n27481 ;
  assign n33685 = n2877 & ~n33684 ;
  assign n33686 = n18992 ^ n17476 ^ n12932 ;
  assign n33687 = n30828 & ~n33686 ;
  assign n33688 = n7995 & n33687 ;
  assign n33689 = n19157 ^ n18209 ^ 1'b0 ;
  assign n33690 = ~n3296 & n33689 ;
  assign n33691 = n1465 & ~n12298 ;
  assign n33692 = n33691 ^ n15397 ^ 1'b0 ;
  assign n33693 = ( n6343 & ~n22982 ) | ( n6343 & n33692 ) | ( ~n22982 & n33692 ) ;
  assign n33694 = ( n31313 & ~n33690 ) | ( n31313 & n33693 ) | ( ~n33690 & n33693 ) ;
  assign n33696 = n26052 ^ n19089 ^ 1'b0 ;
  assign n33697 = n13173 | n33696 ;
  assign n33698 = n33697 ^ n19991 ^ n1729 ;
  assign n33695 = ( ~n10655 & n14350 ) | ( ~n10655 & n22172 ) | ( n14350 & n22172 ) ;
  assign n33699 = n33698 ^ n33695 ^ n19858 ;
  assign n33700 = ( n2170 & n33694 ) | ( n2170 & n33699 ) | ( n33694 & n33699 ) ;
  assign n33701 = ( ~n21388 & n23271 ) | ( ~n21388 & n28292 ) | ( n23271 & n28292 ) ;
  assign n33702 = ( n1890 & n16014 ) | ( n1890 & ~n25241 ) | ( n16014 & ~n25241 ) ;
  assign n33703 = ~n932 & n30468 ;
  assign n33704 = n7468 & n33703 ;
  assign n33707 = n20462 ^ n16652 ^ 1'b0 ;
  assign n33705 = n2819 & n8886 ;
  assign n33706 = ( ~n593 & n12991 ) | ( ~n593 & n33705 ) | ( n12991 & n33705 ) ;
  assign n33708 = n33707 ^ n33706 ^ n23229 ;
  assign n33709 = ( n17822 & n33704 ) | ( n17822 & n33708 ) | ( n33704 & n33708 ) ;
  assign n33710 = ( n2462 & n5405 ) | ( n2462 & ~n16487 ) | ( n5405 & ~n16487 ) ;
  assign n33711 = n33710 ^ n28916 ^ x78 ;
  assign n33712 = n14303 ^ n6842 ^ 1'b0 ;
  assign n33713 = ( n1031 & n26766 ) | ( n1031 & ~n33712 ) | ( n26766 & ~n33712 ) ;
  assign n33714 = n18656 ^ n11330 ^ 1'b0 ;
  assign n33715 = ( n5529 & ~n8621 ) | ( n5529 & n33714 ) | ( ~n8621 & n33714 ) ;
  assign n33716 = n6186 & ~n8729 ;
  assign n33717 = n6809 & ~n16818 ;
  assign n33718 = n31062 & n33717 ;
  assign n33719 = n9085 ^ n5878 ^ 1'b0 ;
  assign n33720 = n33719 ^ n27496 ^ n25785 ;
  assign n33721 = n26020 ^ n24458 ^ 1'b0 ;
  assign n33722 = ~n366 & n27654 ;
  assign n33723 = n15301 ^ n655 ^ x169 ;
  assign n33724 = ( ~n17022 & n30437 ) | ( ~n17022 & n33723 ) | ( n30437 & n33723 ) ;
  assign n33725 = ( n869 & n7277 ) | ( n869 & n10356 ) | ( n7277 & n10356 ) ;
  assign n33726 = ( n10167 & ~n33724 ) | ( n10167 & n33725 ) | ( ~n33724 & n33725 ) ;
  assign n33727 = n24307 ^ n12491 ^ 1'b0 ;
  assign n33728 = n10469 ^ n10226 ^ n1359 ;
  assign n33729 = ( n8212 & n9565 ) | ( n8212 & n33728 ) | ( n9565 & n33728 ) ;
  assign n33730 = ( n429 & ~n8013 ) | ( n429 & n8710 ) | ( ~n8013 & n8710 ) ;
  assign n33731 = ( n27366 & ~n33729 ) | ( n27366 & n33730 ) | ( ~n33729 & n33730 ) ;
  assign n33732 = n16209 ^ n431 ^ 1'b0 ;
  assign n33733 = n33731 | n33732 ;
  assign n33734 = n6712 & ~n32660 ;
  assign n33736 = n3338 ^ n3152 ^ 1'b0 ;
  assign n33735 = n31451 ^ n6475 ^ 1'b0 ;
  assign n33737 = n33736 ^ n33735 ^ n915 ;
  assign n33739 = n7240 & ~n18838 ;
  assign n33738 = n6810 | n22589 ;
  assign n33740 = n33739 ^ n33738 ^ n16609 ;
  assign n33742 = n4014 ^ n3694 ^ 1'b0 ;
  assign n33741 = n18835 | n26013 ;
  assign n33743 = n33742 ^ n33741 ^ 1'b0 ;
  assign n33744 = n33743 ^ n12016 ^ 1'b0 ;
  assign n33745 = n7545 | n33744 ;
  assign n33746 = n15879 & ~n33745 ;
  assign n33747 = n33746 ^ n5881 ^ 1'b0 ;
  assign n33748 = n4534 | n33747 ;
  assign n33749 = n14678 ^ n5723 ^ n2047 ;
  assign n33750 = ~n30114 & n33749 ;
  assign n33751 = n33750 ^ n26541 ^ 1'b0 ;
  assign n33753 = n15361 ^ n14917 ^ n13407 ;
  assign n33752 = n28707 ^ n17699 ^ n610 ;
  assign n33754 = n33753 ^ n33752 ^ n31232 ;
  assign n33755 = n4869 | n33754 ;
  assign n33756 = n33755 ^ n2809 ^ 1'b0 ;
  assign n33757 = n2379 ^ n1605 ^ n1465 ;
  assign n33758 = n32150 ^ n27013 ^ n23662 ;
  assign n33759 = n8386 & ~n33758 ;
  assign n33760 = n25698 ^ n1811 ^ 1'b0 ;
  assign n33761 = n8011 | n33760 ;
  assign n33762 = n33761 ^ n29372 ^ n15534 ;
  assign n33773 = n1112 & ~n15632 ;
  assign n33763 = ( n11702 & n19017 ) | ( n11702 & n20094 ) | ( n19017 & n20094 ) ;
  assign n33767 = ( n1428 & n3267 ) | ( n1428 & n8581 ) | ( n3267 & n8581 ) ;
  assign n33768 = n19266 ^ n12146 ^ 1'b0 ;
  assign n33769 = n33767 & n33768 ;
  assign n33765 = n1572 & n3458 ;
  assign n33764 = n744 & ~n9113 ;
  assign n33766 = n33765 ^ n33764 ^ 1'b0 ;
  assign n33770 = n33769 ^ n33766 ^ n8486 ;
  assign n33771 = ( ~n10683 & n18994 ) | ( ~n10683 & n33770 ) | ( n18994 & n33770 ) ;
  assign n33772 = ( n1838 & n33763 ) | ( n1838 & n33771 ) | ( n33763 & n33771 ) ;
  assign n33774 = n33773 ^ n33772 ^ 1'b0 ;
  assign n33775 = n33762 | n33774 ;
  assign n33776 = ( n2552 & n14237 ) | ( n2552 & ~n31211 ) | ( n14237 & ~n31211 ) ;
  assign n33777 = ~n5654 & n33776 ;
  assign n33778 = ~n11216 & n33777 ;
  assign n33779 = n33778 ^ n7054 ^ 1'b0 ;
  assign n33780 = n26459 ^ n4415 ^ 1'b0 ;
  assign n33781 = n28473 ^ n21497 ^ 1'b0 ;
  assign n33782 = n33781 ^ n12852 ^ n6336 ;
  assign n33783 = ~n12975 & n27094 ;
  assign n33784 = ( ~n2465 & n14616 ) | ( ~n2465 & n18372 ) | ( n14616 & n18372 ) ;
  assign n33785 = ( n4427 & n6095 ) | ( n4427 & n8840 ) | ( n6095 & n8840 ) ;
  assign n33786 = n7301 ^ n5660 ^ 1'b0 ;
  assign n33787 = n33785 & ~n33786 ;
  assign n33788 = n33787 ^ n22017 ^ 1'b0 ;
  assign n33789 = n28525 & ~n33788 ;
  assign n33790 = n33789 ^ n10875 ^ 1'b0 ;
  assign n33791 = ( n26924 & n28861 ) | ( n26924 & n33790 ) | ( n28861 & n33790 ) ;
  assign n33792 = n1381 & n10167 ;
  assign n33793 = n5058 & n33792 ;
  assign n33794 = ( n8870 & n14815 ) | ( n8870 & ~n33793 ) | ( n14815 & ~n33793 ) ;
  assign n33795 = n24760 ^ n21411 ^ n7409 ;
  assign n33796 = n14465 ^ n3846 ^ 1'b0 ;
  assign n33797 = n17745 ^ n16415 ^ 1'b0 ;
  assign n33798 = n3094 & ~n33797 ;
  assign n33799 = ( n3926 & n12016 ) | ( n3926 & ~n17324 ) | ( n12016 & ~n17324 ) ;
  assign n33800 = n33799 ^ n29873 ^ n28895 ;
  assign n33801 = ( n3896 & n33798 ) | ( n3896 & ~n33800 ) | ( n33798 & ~n33800 ) ;
  assign n33802 = n7018 ^ n2323 ^ 1'b0 ;
  assign n33805 = n14202 & n17130 ;
  assign n33806 = n33805 ^ n9292 ^ n4381 ;
  assign n33803 = ( ~n3377 & n5421 ) | ( ~n3377 & n25148 ) | ( n5421 & n25148 ) ;
  assign n33804 = n33803 ^ n19256 ^ n6249 ;
  assign n33807 = n33806 ^ n33804 ^ n2802 ;
  assign n33808 = n583 & ~n33807 ;
  assign n33809 = n16267 & n33808 ;
  assign n33810 = n2631 | n4848 ;
  assign n33811 = ( ~n7781 & n13069 ) | ( ~n7781 & n33810 ) | ( n13069 & n33810 ) ;
  assign n33814 = n3927 & ~n27775 ;
  assign n33815 = n33814 ^ n4004 ^ 1'b0 ;
  assign n33813 = n15935 & ~n18542 ;
  assign n33816 = n33815 ^ n33813 ^ 1'b0 ;
  assign n33812 = n18431 ^ n15919 ^ n12618 ;
  assign n33817 = n33816 ^ n33812 ^ n11542 ;
  assign n33818 = n7989 | n11565 ;
  assign n33819 = n33818 ^ n17962 ^ 1'b0 ;
  assign n33820 = ~n4478 & n8869 ;
  assign n33823 = n23409 ^ n13356 ^ n3512 ;
  assign n33824 = n33823 ^ n13342 ^ n6672 ;
  assign n33821 = ( n4481 & n17294 ) | ( n4481 & ~n29893 ) | ( n17294 & ~n29893 ) ;
  assign n33822 = n33821 ^ n24254 ^ n5023 ;
  assign n33825 = n33824 ^ n33822 ^ n3877 ;
  assign n33826 = n24203 ^ n11524 ^ n10217 ;
  assign n33827 = n33826 ^ n8605 ^ 1'b0 ;
  assign n33830 = ( ~n7362 & n10723 ) | ( ~n7362 & n13607 ) | ( n10723 & n13607 ) ;
  assign n33828 = n15399 ^ n4983 ^ 1'b0 ;
  assign n33829 = ( n713 & n2662 ) | ( n713 & ~n33828 ) | ( n2662 & ~n33828 ) ;
  assign n33831 = n33830 ^ n33829 ^ n6093 ;
  assign n33832 = n21294 ^ n7267 ^ 1'b0 ;
  assign n33833 = n14790 & ~n33832 ;
  assign n33835 = n1450 | n4175 ;
  assign n33836 = n33835 ^ n5261 ^ 1'b0 ;
  assign n33837 = ( n4594 & n10439 ) | ( n4594 & ~n33836 ) | ( n10439 & ~n33836 ) ;
  assign n33834 = ~n5961 & n14097 ;
  assign n33838 = n33837 ^ n33834 ^ 1'b0 ;
  assign n33839 = n11532 | n33838 ;
  assign n33840 = n1258 & ~n33839 ;
  assign n33846 = n8301 ^ n594 ^ 1'b0 ;
  assign n33843 = n9293 & ~n10100 ;
  assign n33844 = n33843 ^ n9733 ^ n6785 ;
  assign n33841 = ~n519 & n2365 ;
  assign n33842 = n33841 ^ n570 ^ 1'b0 ;
  assign n33845 = n33844 ^ n33842 ^ n19783 ;
  assign n33847 = n33846 ^ n33845 ^ n6754 ;
  assign n33848 = n5373 ^ n4454 ^ n1620 ;
  assign n33849 = n19523 ^ n12010 ^ n9321 ;
  assign n33850 = n24572 | n25342 ;
  assign n33851 = n9597 & ~n33850 ;
  assign n33852 = n1134 | n33851 ;
  assign n33853 = n15392 | n33852 ;
  assign n33854 = n33853 ^ n12411 ^ 1'b0 ;
  assign n33855 = ( n33848 & n33849 ) | ( n33848 & n33854 ) | ( n33849 & n33854 ) ;
  assign n33856 = n13918 & n17557 ;
  assign n33857 = n22941 ^ n18110 ^ n7888 ;
  assign n33858 = ( n8403 & n33856 ) | ( n8403 & n33857 ) | ( n33856 & n33857 ) ;
  assign n33859 = n14680 & ~n25827 ;
  assign n33860 = ( n2660 & ~n22597 ) | ( n2660 & n33859 ) | ( ~n22597 & n33859 ) ;
  assign n33861 = n33860 ^ n5611 ^ n1202 ;
  assign n33862 = n3429 & ~n16726 ;
  assign n33863 = n28917 ^ n23187 ^ n17302 ;
  assign n33864 = ( n15341 & n19884 ) | ( n15341 & ~n27163 ) | ( n19884 & ~n27163 ) ;
  assign n33865 = ( n16520 & n17558 ) | ( n16520 & n29989 ) | ( n17558 & n29989 ) ;
  assign n33866 = n13711 ^ n13153 ^ n823 ;
  assign n33867 = ( n10960 & n18238 ) | ( n10960 & n33866 ) | ( n18238 & n33866 ) ;
  assign n33868 = n16752 ^ n15477 ^ 1'b0 ;
  assign n33869 = n13548 | n20612 ;
  assign n33871 = n13105 ^ n8848 ^ n3351 ;
  assign n33872 = n33871 ^ n17101 ^ n6820 ;
  assign n33873 = n16381 & ~n33872 ;
  assign n33874 = ~n14569 & n33873 ;
  assign n33870 = n21262 ^ n13610 ^ x80 ;
  assign n33875 = n33874 ^ n33870 ^ n3474 ;
  assign n33878 = n17042 ^ n7627 ^ 1'b0 ;
  assign n33876 = n13717 | n28905 ;
  assign n33877 = n33876 ^ n2787 ^ 1'b0 ;
  assign n33879 = n33878 ^ n33877 ^ n20539 ;
  assign n33880 = n28674 ^ n22213 ^ n5246 ;
  assign n33881 = n22714 & ~n33880 ;
  assign n33882 = ( n8501 & n16896 ) | ( n8501 & ~n19943 ) | ( n16896 & ~n19943 ) ;
  assign n33883 = n17572 & n33882 ;
  assign n33884 = n33883 ^ n30008 ^ 1'b0 ;
  assign n33885 = ~n8126 & n15317 ;
  assign n33886 = n33885 ^ n6264 ^ n4389 ;
  assign n33887 = ( n8456 & ~n28483 ) | ( n8456 & n33886 ) | ( ~n28483 & n33886 ) ;
  assign n33888 = n13737 ^ n1670 ^ 1'b0 ;
  assign n33889 = n33888 ^ n16598 ^ 1'b0 ;
  assign n33890 = n5637 | n33889 ;
  assign n33891 = n22044 | n33890 ;
  assign n33892 = ( n13577 & ~n17112 ) | ( n13577 & n29099 ) | ( ~n17112 & n29099 ) ;
  assign n33893 = n11205 & ~n22762 ;
  assign n33894 = ( n1156 & n1942 ) | ( n1156 & n12403 ) | ( n1942 & n12403 ) ;
  assign n33896 = ~n19043 & n19110 ;
  assign n33897 = n2197 & n33896 ;
  assign n33898 = n33897 ^ n9177 ^ n7925 ;
  assign n33895 = n20454 & ~n26098 ;
  assign n33899 = n33898 ^ n33895 ^ n6118 ;
  assign n33900 = ~n744 & n33899 ;
  assign n33901 = n847 | n1476 ;
  assign n33902 = n33901 ^ n14564 ^ 1'b0 ;
  assign n33903 = n20025 ^ n17752 ^ n2170 ;
  assign n33904 = n33903 ^ n3743 ^ 1'b0 ;
  assign n33905 = ~n1491 & n22899 ;
  assign n33906 = n3566 & n33905 ;
  assign n33907 = ~n3156 & n33906 ;
  assign n33908 = n33907 ^ n13891 ^ 1'b0 ;
  assign n33909 = n19387 & ~n33908 ;
  assign n33910 = n25773 ^ n20222 ^ n13715 ;
  assign n33911 = n27962 ^ n16154 ^ n1164 ;
  assign n33912 = ( ~n1773 & n18461 ) | ( ~n1773 & n33911 ) | ( n18461 & n33911 ) ;
  assign n33913 = n33910 & n33912 ;
  assign n33914 = n10300 ^ n2570 ^ x11 ;
  assign n33917 = ( ~n1484 & n5529 ) | ( ~n1484 & n15412 ) | ( n5529 & n15412 ) ;
  assign n33915 = n7968 ^ n6394 ^ 1'b0 ;
  assign n33916 = n25514 & ~n33915 ;
  assign n33918 = n33917 ^ n33916 ^ n12436 ;
  assign n33919 = ( n1902 & ~n5409 ) | ( n1902 & n9534 ) | ( ~n5409 & n9534 ) ;
  assign n33920 = n678 & ~n8831 ;
  assign n33921 = ( n9134 & ~n20373 ) | ( n9134 & n33920 ) | ( ~n20373 & n33920 ) ;
  assign n33922 = n2455 & n10268 ;
  assign n33923 = n2134 ^ n890 ^ 1'b0 ;
  assign n33924 = ~n22071 & n33923 ;
  assign n33925 = n33846 ^ n14929 ^ n3002 ;
  assign n33926 = n29062 ^ n7491 ^ n7162 ;
  assign n33927 = n28691 & ~n33926 ;
  assign n33928 = n33927 ^ n25149 ^ 1'b0 ;
  assign n33929 = n33925 & ~n33928 ;
  assign n33930 = n10405 | n13205 ;
  assign n33931 = n2319 | n9686 ;
  assign n33932 = n33931 ^ n31489 ^ n13325 ;
  assign n33933 = n33932 ^ n19937 ^ n7715 ;
  assign n33934 = ( n12863 & n33930 ) | ( n12863 & n33933 ) | ( n33930 & n33933 ) ;
  assign n33935 = ( n2589 & ~n5373 ) | ( n2589 & n19888 ) | ( ~n5373 & n19888 ) ;
  assign n33936 = n33935 ^ n19382 ^ 1'b0 ;
  assign n33937 = n6873 & ~n33936 ;
  assign n33938 = ~n10676 & n33937 ;
  assign n33939 = n15986 & ~n33938 ;
  assign n33940 = n16700 ^ n7475 ^ 1'b0 ;
  assign n33941 = n7039 | n33940 ;
  assign n33942 = ~n20415 & n33941 ;
  assign n33943 = n8722 ^ n7558 ^ n4820 ;
  assign n33944 = n21954 & ~n33943 ;
  assign n33945 = n33944 ^ n8517 ^ 1'b0 ;
  assign n33946 = n12898 ^ n3607 ^ 1'b0 ;
  assign n33947 = ~n14998 & n33946 ;
  assign n33950 = n23835 ^ n12518 ^ n12032 ;
  assign n33948 = n18409 | n24862 ;
  assign n33949 = n5974 | n33948 ;
  assign n33951 = n33950 ^ n33949 ^ n2302 ;
  assign n33957 = ( ~n14660 & n15145 ) | ( ~n14660 & n17793 ) | ( n15145 & n17793 ) ;
  assign n33955 = n27688 ^ n3345 ^ x88 ;
  assign n33952 = n16395 ^ n4383 ^ 1'b0 ;
  assign n33953 = ( n7335 & n7763 ) | ( n7335 & ~n33952 ) | ( n7763 & ~n33952 ) ;
  assign n33954 = n33953 ^ n9382 ^ n8182 ;
  assign n33956 = n33955 ^ n33954 ^ n9730 ;
  assign n33958 = n33957 ^ n33956 ^ n9529 ;
  assign n33959 = n24418 ^ n7673 ^ n942 ;
  assign n33960 = ( n11304 & n17795 ) | ( n11304 & ~n20908 ) | ( n17795 & ~n20908 ) ;
  assign n33962 = n13903 ^ n11919 ^ n9191 ;
  assign n33961 = x78 & ~n10945 ;
  assign n33963 = n33962 ^ n33961 ^ 1'b0 ;
  assign n33964 = n33960 & n33963 ;
  assign n33965 = n29942 ^ n2027 ^ 1'b0 ;
  assign n33966 = n33964 & n33965 ;
  assign n33967 = ( x248 & n20354 ) | ( x248 & n33966 ) | ( n20354 & n33966 ) ;
  assign n33968 = n33967 ^ n25366 ^ n549 ;
  assign n33969 = ( n2819 & ~n3018 ) | ( n2819 & n5888 ) | ( ~n3018 & n5888 ) ;
  assign n33973 = ( ~n4081 & n6664 ) | ( ~n4081 & n13555 ) | ( n6664 & n13555 ) ;
  assign n33970 = n5561 & n18551 ;
  assign n33971 = n5630 & n33970 ;
  assign n33972 = n14992 & ~n33971 ;
  assign n33974 = n33973 ^ n33972 ^ 1'b0 ;
  assign n33975 = n33974 ^ n20088 ^ 1'b0 ;
  assign n33976 = n33969 | n33975 ;
  assign n33977 = ~n7348 & n20174 ;
  assign n33980 = n1369 | n1582 ;
  assign n33981 = n2305 & ~n33980 ;
  assign n33982 = n33981 ^ n26728 ^ n13469 ;
  assign n33978 = n4501 & n29123 ;
  assign n33979 = n7487 & n33978 ;
  assign n33983 = n33982 ^ n33979 ^ 1'b0 ;
  assign n33985 = n1747 | n8949 ;
  assign n33986 = n25413 & ~n33985 ;
  assign n33984 = ( n2926 & ~n5251 ) | ( n2926 & n22263 ) | ( ~n5251 & n22263 ) ;
  assign n33987 = n33986 ^ n33984 ^ n9446 ;
  assign n33988 = n5224 & ~n6587 ;
  assign n33989 = n3708 & n33988 ;
  assign n33990 = n16510 & n21662 ;
  assign n33991 = n29842 ^ n28793 ^ n13231 ;
  assign n33992 = ( n1124 & n5532 ) | ( n1124 & ~n13586 ) | ( n5532 & ~n13586 ) ;
  assign n33993 = ( n17479 & ~n25050 ) | ( n17479 & n33992 ) | ( ~n25050 & n33992 ) ;
  assign n33994 = ( ~x160 & n26255 ) | ( ~x160 & n33993 ) | ( n26255 & n33993 ) ;
  assign n33996 = ( n4196 & n8560 ) | ( n4196 & n12593 ) | ( n8560 & n12593 ) ;
  assign n33995 = n21140 ^ n7582 ^ n1680 ;
  assign n33997 = n33996 ^ n33995 ^ n11207 ;
  assign n33998 = ( n407 & n2678 ) | ( n407 & ~n18820 ) | ( n2678 & ~n18820 ) ;
  assign n33999 = n33998 ^ n18972 ^ n501 ;
  assign n34000 = ( ~n30123 & n33997 ) | ( ~n30123 & n33999 ) | ( n33997 & n33999 ) ;
  assign n34001 = ( ~n696 & n2512 ) | ( ~n696 & n4635 ) | ( n2512 & n4635 ) ;
  assign n34002 = n34001 ^ n33031 ^ 1'b0 ;
  assign n34003 = n4399 & ~n16539 ;
  assign n34004 = n34003 ^ n23776 ^ n23134 ;
  assign n34005 = n3980 & ~n21377 ;
  assign n34006 = n34005 ^ n7105 ^ 1'b0 ;
  assign n34007 = n34006 ^ n25767 ^ 1'b0 ;
  assign n34008 = n10228 | n19244 ;
  assign n34009 = n3459 | n34008 ;
  assign n34010 = ~n15245 & n26518 ;
  assign n34011 = n34010 ^ n22314 ^ 1'b0 ;
  assign n34012 = ( n13397 & n34009 ) | ( n13397 & n34011 ) | ( n34009 & n34011 ) ;
  assign n34013 = ( n14375 & n17899 ) | ( n14375 & ~n31177 ) | ( n17899 & ~n31177 ) ;
  assign n34014 = n18452 ^ n807 ^ 1'b0 ;
  assign n34015 = n5648 | n34014 ;
  assign n34018 = n25432 ^ n18318 ^ n6453 ;
  assign n34016 = n2905 & n9812 ;
  assign n34017 = n17784 | n34016 ;
  assign n34019 = n34018 ^ n34017 ^ 1'b0 ;
  assign n34020 = ~n1204 & n7607 ;
  assign n34021 = n34020 ^ n16612 ^ 1'b0 ;
  assign n34022 = n34021 ^ n20756 ^ n18306 ;
  assign n34023 = ( n31334 & n31925 ) | ( n31334 & ~n34022 ) | ( n31925 & ~n34022 ) ;
  assign n34024 = n10727 | n18733 ;
  assign n34025 = n34024 ^ n28734 ^ 1'b0 ;
  assign n34026 = n34025 ^ n31912 ^ n10146 ;
  assign n34027 = n4110 & n13322 ;
  assign n34028 = ~n19728 & n34027 ;
  assign n34029 = n16982 & ~n34028 ;
  assign n34030 = n7582 & n17667 ;
  assign n34031 = n34030 ^ n20124 ^ 1'b0 ;
  assign n34032 = n9125 & n13933 ;
  assign n34033 = ~n33017 & n34032 ;
  assign n34034 = n29285 | n34033 ;
  assign n34035 = n34034 ^ n8375 ^ 1'b0 ;
  assign n34036 = n22422 ^ n20808 ^ n19459 ;
  assign n34037 = ( ~n2962 & n27242 ) | ( ~n2962 & n34036 ) | ( n27242 & n34036 ) ;
  assign n34038 = n4049 | n34037 ;
  assign n34040 = n32087 ^ n16870 ^ 1'b0 ;
  assign n34039 = n2603 | n4069 ;
  assign n34041 = n34040 ^ n34039 ^ 1'b0 ;
  assign n34042 = n4147 | n34041 ;
  assign n34043 = n15367 | n24576 ;
  assign n34044 = n34043 ^ n12708 ^ 1'b0 ;
  assign n34045 = ( n15660 & ~n21739 ) | ( n15660 & n34044 ) | ( ~n21739 & n34044 ) ;
  assign n34051 = n4323 & ~n15947 ;
  assign n34046 = ~n15821 & n16255 ;
  assign n34047 = n34046 ^ n22549 ^ n13489 ;
  assign n34048 = n11747 & ~n34047 ;
  assign n34049 = n21722 ^ n7817 ^ 1'b0 ;
  assign n34050 = ( ~n7045 & n34048 ) | ( ~n7045 & n34049 ) | ( n34048 & n34049 ) ;
  assign n34052 = n34051 ^ n34050 ^ n16401 ;
  assign n34053 = n31301 ^ n19472 ^ n2325 ;
  assign n34054 = n4976 | n8339 ;
  assign n34055 = ( ~n8332 & n20539 ) | ( ~n8332 & n34054 ) | ( n20539 & n34054 ) ;
  assign n34057 = n25431 ^ n22716 ^ n20673 ;
  assign n34056 = n6905 & n19645 ;
  assign n34058 = n34057 ^ n34056 ^ 1'b0 ;
  assign n34059 = ( n16170 & n29707 ) | ( n16170 & ~n34058 ) | ( n29707 & ~n34058 ) ;
  assign n34060 = n13493 ^ n11823 ^ n11152 ;
  assign n34062 = n2539 ^ n812 ^ 1'b0 ;
  assign n34063 = n1156 | n34062 ;
  assign n34061 = ( ~n6869 & n22996 ) | ( ~n6869 & n25101 ) | ( n22996 & n25101 ) ;
  assign n34064 = n34063 ^ n34061 ^ n2315 ;
  assign n34065 = n15015 ^ n6951 ^ n864 ;
  assign n34066 = n34065 ^ n10525 ^ 1'b0 ;
  assign n34067 = n21907 & n34066 ;
  assign n34068 = ( ~n2471 & n8851 ) | ( ~n2471 & n11362 ) | ( n8851 & n11362 ) ;
  assign n34069 = n33248 ^ n26076 ^ 1'b0 ;
  assign n34070 = n16083 ^ n12205 ^ n5095 ;
  assign n34071 = n24961 ^ n7861 ^ n7245 ;
  assign n34072 = n469 & n34071 ;
  assign n34073 = n10497 ^ n9167 ^ 1'b0 ;
  assign n34074 = x73 | n6226 ;
  assign n34075 = n10634 | n34074 ;
  assign n34076 = n8779 | n34075 ;
  assign n34077 = ( n34072 & ~n34073 ) | ( n34072 & n34076 ) | ( ~n34073 & n34076 ) ;
  assign n34078 = n14620 ^ n5055 ^ 1'b0 ;
  assign n34079 = ~n942 & n34078 ;
  assign n34080 = n17480 & n34079 ;
  assign n34081 = n32745 ^ n4769 ^ 1'b0 ;
  assign n34082 = ( n6239 & ~n10486 ) | ( n6239 & n15448 ) | ( ~n10486 & n15448 ) ;
  assign n34083 = ~n18488 & n24779 ;
  assign n34084 = ~n9855 & n34083 ;
  assign n34085 = n34082 & ~n34084 ;
  assign n34086 = n34081 & n34085 ;
  assign n34090 = n6217 ^ n4909 ^ 1'b0 ;
  assign n34087 = ~n3522 & n11107 ;
  assign n34088 = ~n4893 & n20130 ;
  assign n34089 = n34087 & n34088 ;
  assign n34091 = n34090 ^ n34089 ^ n17334 ;
  assign n34092 = ( n1327 & n3084 ) | ( n1327 & n34091 ) | ( n3084 & n34091 ) ;
  assign n34093 = ~n4269 & n18405 ;
  assign n34094 = ( n2174 & ~n24176 ) | ( n2174 & n34093 ) | ( ~n24176 & n34093 ) ;
  assign n34095 = n18364 ^ n801 ^ 1'b0 ;
  assign n34096 = ( n10670 & ~n17125 ) | ( n10670 & n34095 ) | ( ~n17125 & n34095 ) ;
  assign n34104 = n13266 ^ n2617 ^ 1'b0 ;
  assign n34105 = n4906 | n34104 ;
  assign n34101 = ( ~n12952 & n22556 ) | ( ~n12952 & n31612 ) | ( n22556 & n31612 ) ;
  assign n34102 = n34101 ^ n20641 ^ n13286 ;
  assign n34103 = n34102 ^ n30848 ^ n7139 ;
  assign n34097 = n27953 ^ n10547 ^ 1'b0 ;
  assign n34098 = n16007 | n28790 ;
  assign n34099 = ~n26697 & n34098 ;
  assign n34100 = ~n34097 & n34099 ;
  assign n34106 = n34105 ^ n34103 ^ n34100 ;
  assign n34107 = ( ~x168 & n4578 ) | ( ~x168 & n10216 ) | ( n4578 & n10216 ) ;
  assign n34108 = ~n8229 & n34107 ;
  assign n34109 = ( ~n1200 & n20868 ) | ( ~n1200 & n30788 ) | ( n20868 & n30788 ) ;
  assign n34110 = ( n3538 & n25631 ) | ( n3538 & ~n32829 ) | ( n25631 & ~n32829 ) ;
  assign n34111 = ~n34109 & n34110 ;
  assign n34112 = n34111 ^ n25792 ^ 1'b0 ;
  assign n34113 = n34112 ^ n27270 ^ n27054 ;
  assign n34114 = n28808 ^ n11244 ^ n3333 ;
  assign n34115 = ( n5892 & ~n8979 ) | ( n5892 & n21628 ) | ( ~n8979 & n21628 ) ;
  assign n34116 = n34115 ^ n28556 ^ n10930 ;
  assign n34117 = n32702 ^ n12508 ^ 1'b0 ;
  assign n34118 = n19960 & n34117 ;
  assign n34119 = x137 & ~n5959 ;
  assign n34120 = n34119 ^ n13584 ^ 1'b0 ;
  assign n34121 = n34120 ^ n29586 ^ n13546 ;
  assign n34122 = ( n26084 & n34118 ) | ( n26084 & n34121 ) | ( n34118 & n34121 ) ;
  assign n34123 = ( n8426 & n13028 ) | ( n8426 & n16531 ) | ( n13028 & n16531 ) ;
  assign n34124 = n14543 | n27609 ;
  assign n34125 = n34124 ^ n6915 ^ 1'b0 ;
  assign n34127 = ( n1068 & n9995 ) | ( n1068 & ~n14007 ) | ( n9995 & ~n14007 ) ;
  assign n34126 = n5491 | n13808 ;
  assign n34128 = n34127 ^ n34126 ^ n15838 ;
  assign n34129 = n25982 & n32099 ;
  assign n34130 = ~n34128 & n34129 ;
  assign n34131 = n2472 & n21975 ;
  assign n34132 = n453 | n12609 ;
  assign n34133 = n30807 & ~n34132 ;
  assign n34134 = n13639 ^ n11800 ^ 1'b0 ;
  assign n34135 = n31201 & ~n34134 ;
  assign n34136 = ( n6732 & n7780 ) | ( n6732 & n34135 ) | ( n7780 & n34135 ) ;
  assign n34137 = ( n14081 & ~n16926 ) | ( n14081 & n34136 ) | ( ~n16926 & n34136 ) ;
  assign n34138 = ( n29285 & ~n34133 ) | ( n29285 & n34137 ) | ( ~n34133 & n34137 ) ;
  assign n34139 = n34138 ^ n6207 ^ 1'b0 ;
  assign n34140 = n24092 ^ n18982 ^ 1'b0 ;
  assign n34141 = n24120 ^ n4698 ^ 1'b0 ;
  assign n34142 = ~n34140 & n34141 ;
  assign n34143 = n31202 ^ n14458 ^ 1'b0 ;
  assign n34144 = ( ~n525 & n771 ) | ( ~n525 & n3275 ) | ( n771 & n3275 ) ;
  assign n34145 = n1827 & n11564 ;
  assign n34146 = n34145 ^ n12012 ^ 1'b0 ;
  assign n34147 = n34146 ^ n5632 ^ 1'b0 ;
  assign n34148 = n34147 ^ n28621 ^ 1'b0 ;
  assign n34149 = n34144 & ~n34148 ;
  assign n34150 = n24743 | n28821 ;
  assign n34151 = ( n27984 & ~n32122 ) | ( n27984 & n34150 ) | ( ~n32122 & n34150 ) ;
  assign n34152 = n3659 & n11293 ;
  assign n34153 = ~n12592 & n16423 ;
  assign n34154 = x52 & ~n3911 ;
  assign n34155 = n18115 & n34154 ;
  assign n34156 = n24431 ^ n1434 ^ 1'b0 ;
  assign n34157 = ~n34155 & n34156 ;
  assign n34158 = n19969 ^ n14660 ^ 1'b0 ;
  assign n34159 = n15362 & n34158 ;
  assign n34160 = n24523 ^ n22665 ^ n13981 ;
  assign n34161 = n21347 ^ n9988 ^ 1'b0 ;
  assign n34162 = n13941 & ~n34161 ;
  assign n34166 = ( ~n288 & n7451 ) | ( ~n288 & n9063 ) | ( n7451 & n9063 ) ;
  assign n34164 = n8463 ^ n5542 ^ n2703 ;
  assign n34163 = ~n5910 & n8285 ;
  assign n34165 = n34164 ^ n34163 ^ n14455 ;
  assign n34167 = n34166 ^ n34165 ^ n28847 ;
  assign n34168 = ( ~n6987 & n34162 ) | ( ~n6987 & n34167 ) | ( n34162 & n34167 ) ;
  assign n34169 = ( n2807 & n4354 ) | ( n2807 & n5382 ) | ( n4354 & n5382 ) ;
  assign n34170 = n34169 ^ n19726 ^ n5108 ;
  assign n34171 = ( n3253 & ~n20333 ) | ( n3253 & n24382 ) | ( ~n20333 & n24382 ) ;
  assign n34172 = n2230 & n34171 ;
  assign n34173 = ~n19811 & n34172 ;
  assign n34174 = n4154 & n22727 ;
  assign n34175 = n34174 ^ n15562 ^ 1'b0 ;
  assign n34176 = ~n9396 & n34175 ;
  assign n34177 = n34176 ^ n24383 ^ 1'b0 ;
  assign n34178 = n5189 & ~n6546 ;
  assign n34179 = ~n6998 & n34178 ;
  assign n34180 = n9663 | n34179 ;
  assign n34181 = n34180 ^ n4992 ^ 1'b0 ;
  assign n34182 = n10306 ^ n4899 ^ 1'b0 ;
  assign n34183 = n1247 & n34182 ;
  assign n34184 = n34183 ^ n15264 ^ 1'b0 ;
  assign n34185 = n34184 ^ n12248 ^ n8190 ;
  assign n34194 = n11862 ^ n4433 ^ n789 ;
  assign n34192 = n10219 ^ n5107 ^ 1'b0 ;
  assign n34193 = ~n14783 & n34192 ;
  assign n34190 = n5754 ^ n5563 ^ 1'b0 ;
  assign n34191 = n20356 | n34190 ;
  assign n34195 = n34194 ^ n34193 ^ n34191 ;
  assign n34186 = ( n715 & n9959 ) | ( n715 & n13130 ) | ( n9959 & n13130 ) ;
  assign n34187 = n34186 ^ n31759 ^ 1'b0 ;
  assign n34188 = n16803 & n34187 ;
  assign n34189 = n34188 ^ n2827 ^ 1'b0 ;
  assign n34196 = n34195 ^ n34189 ^ n9697 ;
  assign n34197 = n30744 ^ n12542 ^ x70 ;
  assign n34198 = n21185 ^ n7289 ^ 1'b0 ;
  assign n34199 = ( ~n14772 & n18649 ) | ( ~n14772 & n24301 ) | ( n18649 & n24301 ) ;
  assign n34200 = n34199 ^ x210 ^ 1'b0 ;
  assign n34201 = ~n10888 & n10933 ;
  assign n34202 = ( n15780 & n16590 ) | ( n15780 & n34201 ) | ( n16590 & n34201 ) ;
  assign n34203 = ( ~n3811 & n34200 ) | ( ~n3811 & n34202 ) | ( n34200 & n34202 ) ;
  assign n34204 = ( n4177 & ~n9293 ) | ( n4177 & n15876 ) | ( ~n9293 & n15876 ) ;
  assign n34205 = ( n4096 & ~n9716 ) | ( n4096 & n34204 ) | ( ~n9716 & n34204 ) ;
  assign n34206 = n34205 ^ n13419 ^ 1'b0 ;
  assign n34207 = n34206 ^ n20460 ^ 1'b0 ;
  assign n34208 = n34203 | n34207 ;
  assign n34209 = ( n9150 & ~n34198 ) | ( n9150 & n34208 ) | ( ~n34198 & n34208 ) ;
  assign n34210 = ~n3335 & n7281 ;
  assign n34211 = ~n32679 & n34210 ;
  assign n34212 = n849 & n22742 ;
  assign n34213 = ( ~n12330 & n14379 ) | ( ~n12330 & n32197 ) | ( n14379 & n32197 ) ;
  assign n34214 = n1372 & n11924 ;
  assign n34215 = n34214 ^ n32875 ^ n25122 ;
  assign n34216 = ( n12313 & n15903 ) | ( n12313 & n34215 ) | ( n15903 & n34215 ) ;
  assign n34217 = n13110 ^ n6764 ^ 1'b0 ;
  assign n34218 = n15556 & n34217 ;
  assign n34219 = ( n2964 & n9048 ) | ( n2964 & ~n34218 ) | ( n9048 & ~n34218 ) ;
  assign n34220 = ( ~n1553 & n12513 ) | ( ~n1553 & n17751 ) | ( n12513 & n17751 ) ;
  assign n34221 = ( n17792 & ~n33137 ) | ( n17792 & n34220 ) | ( ~n33137 & n34220 ) ;
  assign n34222 = n6778 & ~n6796 ;
  assign n34223 = n34222 ^ n15450 ^ 1'b0 ;
  assign n34224 = ~n26627 & n34223 ;
  assign n34225 = n2189 ^ n370 ^ 1'b0 ;
  assign n34226 = n2854 & ~n34225 ;
  assign n34228 = n33563 ^ n30618 ^ 1'b0 ;
  assign n34227 = n20336 | n22849 ;
  assign n34229 = n34228 ^ n34227 ^ 1'b0 ;
  assign n34230 = n34226 & ~n34229 ;
  assign n34231 = n34230 ^ n19429 ^ 1'b0 ;
  assign n34233 = n21819 ^ n12732 ^ 1'b0 ;
  assign n34232 = n6239 ^ n4621 ^ n3664 ;
  assign n34234 = n34233 ^ n34232 ^ n22534 ;
  assign n34235 = n5899 ^ n5210 ^ 1'b0 ;
  assign n34236 = ~n12686 & n34235 ;
  assign n34237 = ( n19244 & ~n30513 ) | ( n19244 & n34236 ) | ( ~n30513 & n34236 ) ;
  assign n34238 = n32986 ^ n31002 ^ n7156 ;
  assign n34239 = n9371 ^ x212 ^ 1'b0 ;
  assign n34240 = n34239 ^ n14396 ^ 1'b0 ;
  assign n34241 = n28722 & ~n34240 ;
  assign n34243 = n1165 & ~n21583 ;
  assign n34242 = ( n7804 & n9115 ) | ( n7804 & n17254 ) | ( n9115 & n17254 ) ;
  assign n34244 = n34243 ^ n34242 ^ 1'b0 ;
  assign n34245 = n31997 & ~n34244 ;
  assign n34246 = ( n11643 & n16881 ) | ( n11643 & n20651 ) | ( n16881 & n20651 ) ;
  assign n34247 = n24424 ^ n11611 ^ n6635 ;
  assign n34248 = n34247 ^ n20158 ^ 1'b0 ;
  assign n34249 = n34248 ^ n32819 ^ n24179 ;
  assign n34250 = n9330 ^ n7925 ^ n1897 ;
  assign n34251 = n12112 ^ n10898 ^ n364 ;
  assign n34252 = n17939 | n34251 ;
  assign n34253 = n10394 & ~n34252 ;
  assign n34254 = n34253 ^ n18117 ^ 1'b0 ;
  assign n34255 = ~n9001 & n19451 ;
  assign n34256 = ( n34250 & n34254 ) | ( n34250 & n34255 ) | ( n34254 & n34255 ) ;
  assign n34257 = ( n1949 & n4667 ) | ( n1949 & n12366 ) | ( n4667 & n12366 ) ;
  assign n34258 = n34257 ^ n30464 ^ 1'b0 ;
  assign n34259 = n13940 ^ n13264 ^ n3985 ;
  assign n34260 = n7245 & n30920 ;
  assign n34261 = n34259 & n34260 ;
  assign n34262 = ( ~n11751 & n19015 ) | ( ~n11751 & n34261 ) | ( n19015 & n34261 ) ;
  assign n34263 = n34262 ^ n24443 ^ n20158 ;
  assign n34264 = n17686 ^ n10727 ^ 1'b0 ;
  assign n34265 = n29645 & n34264 ;
  assign n34266 = n15100 & ~n21142 ;
  assign n34267 = n34266 ^ n9677 ^ 1'b0 ;
  assign n34268 = n8688 | n9012 ;
  assign n34269 = n34268 ^ n28246 ^ 1'b0 ;
  assign n34270 = ( n7386 & n12307 ) | ( n7386 & ~n15449 ) | ( n12307 & ~n15449 ) ;
  assign n34271 = n25118 ^ n23229 ^ n12547 ;
  assign n34272 = n34271 ^ n13508 ^ 1'b0 ;
  assign n34273 = ( n2441 & n22850 ) | ( n2441 & ~n23364 ) | ( n22850 & ~n23364 ) ;
  assign n34274 = n29474 ^ n21506 ^ 1'b0 ;
  assign n34275 = ( n15841 & n31832 ) | ( n15841 & ~n34274 ) | ( n31832 & ~n34274 ) ;
  assign n34276 = ( ~n23478 & n25614 ) | ( ~n23478 & n34275 ) | ( n25614 & n34275 ) ;
  assign n34277 = n5051 ^ n4022 ^ n3185 ;
  assign n34278 = ( n2830 & n34276 ) | ( n2830 & n34277 ) | ( n34276 & n34277 ) ;
  assign n34279 = n7865 & ~n15377 ;
  assign n34280 = ( n640 & n3937 ) | ( n640 & ~n7007 ) | ( n3937 & ~n7007 ) ;
  assign n34281 = ( n29914 & n34279 ) | ( n29914 & n34280 ) | ( n34279 & n34280 ) ;
  assign n34283 = n4715 & n21101 ;
  assign n34284 = n7895 & n34283 ;
  assign n34282 = n4342 & n18406 ;
  assign n34285 = n34284 ^ n34282 ^ 1'b0 ;
  assign n34286 = n424 & ~n7809 ;
  assign n34287 = n34286 ^ n29668 ^ 1'b0 ;
  assign n34288 = n21261 ^ n7540 ^ 1'b0 ;
  assign n34289 = n5418 | n34288 ;
  assign n34290 = n34289 ^ n17370 ^ 1'b0 ;
  assign n34291 = n19508 ^ n3206 ^ n2733 ;
  assign n34292 = n34291 ^ n19158 ^ 1'b0 ;
  assign n34293 = x208 & n34292 ;
  assign n34294 = n34293 ^ n27654 ^ n2240 ;
  assign n34295 = ( n11410 & n34290 ) | ( n11410 & n34294 ) | ( n34290 & n34294 ) ;
  assign n34297 = ( n4373 & n7354 ) | ( n4373 & n29241 ) | ( n7354 & n29241 ) ;
  assign n34296 = ( n1719 & ~n4939 ) | ( n1719 & n11408 ) | ( ~n4939 & n11408 ) ;
  assign n34298 = n34297 ^ n34296 ^ n23981 ;
  assign n34299 = n10651 | n16349 ;
  assign n34300 = n6370 ^ n3962 ^ 1'b0 ;
  assign n34301 = ~n2920 & n34300 ;
  assign n34302 = n16998 | n34301 ;
  assign n34303 = n34302 ^ n21771 ^ n14679 ;
  assign n34304 = n21500 & n34303 ;
  assign n34305 = ~n28317 & n34304 ;
  assign n34306 = ( n5599 & n11183 ) | ( n5599 & ~n26941 ) | ( n11183 & ~n26941 ) ;
  assign n34307 = n9269 | n34306 ;
  assign n34308 = ( n1794 & ~n5560 ) | ( n1794 & n11075 ) | ( ~n5560 & n11075 ) ;
  assign n34309 = ( n8307 & ~n10615 ) | ( n8307 & n34308 ) | ( ~n10615 & n34308 ) ;
  assign n34310 = n3667 & ~n14673 ;
  assign n34311 = ~n31502 & n34310 ;
  assign n34312 = n34309 & ~n34311 ;
  assign n34313 = ~n3352 & n34312 ;
  assign n34314 = ( n17084 & ~n28264 ) | ( n17084 & n34313 ) | ( ~n28264 & n34313 ) ;
  assign n34315 = ( n1062 & n22075 ) | ( n1062 & ~n31016 ) | ( n22075 & ~n31016 ) ;
  assign n34316 = n14941 ^ n10647 ^ n7251 ;
  assign n34317 = ( ~n9279 & n30172 ) | ( ~n9279 & n34316 ) | ( n30172 & n34316 ) ;
  assign n34318 = n34315 & ~n34317 ;
  assign n34320 = n664 & n2862 ;
  assign n34319 = n16455 ^ n13461 ^ n5558 ;
  assign n34321 = n34320 ^ n34319 ^ 1'b0 ;
  assign n34322 = n13540 ^ n433 ^ 1'b0 ;
  assign n34323 = ~n3000 & n34322 ;
  assign n34324 = n13889 & n34323 ;
  assign n34325 = n34324 ^ n15941 ^ 1'b0 ;
  assign n34326 = n34325 ^ n27068 ^ 1'b0 ;
  assign n34327 = n7709 | n34326 ;
  assign n34328 = ( n15884 & n22549 ) | ( n15884 & n34327 ) | ( n22549 & n34327 ) ;
  assign n34331 = n22676 & n28129 ;
  assign n34332 = n34331 ^ n27443 ^ n16422 ;
  assign n34329 = ~n2283 & n26138 ;
  assign n34330 = n34329 ^ n14231 ^ 1'b0 ;
  assign n34333 = n34332 ^ n34330 ^ n24898 ;
  assign n34337 = n19817 ^ n18626 ^ n8391 ;
  assign n34334 = ( n4518 & n9899 ) | ( n4518 & ~n18207 ) | ( n9899 & ~n18207 ) ;
  assign n34335 = n25725 ^ n24593 ^ 1'b0 ;
  assign n34336 = n34334 & ~n34335 ;
  assign n34338 = n34337 ^ n34336 ^ 1'b0 ;
  assign n34339 = n22907 ^ n1536 ^ 1'b0 ;
  assign n34340 = n29247 & ~n34327 ;
  assign n34341 = ( n6182 & n13234 ) | ( n6182 & ~n18760 ) | ( n13234 & ~n18760 ) ;
  assign n34342 = n16591 & n34341 ;
  assign n34343 = n9351 & n34342 ;
  assign n34344 = n15434 | n18882 ;
  assign n34345 = n9601 | n34344 ;
  assign n34346 = n33729 ^ n5348 ^ n2115 ;
  assign n34347 = ( ~n33299 & n34345 ) | ( ~n33299 & n34346 ) | ( n34345 & n34346 ) ;
  assign n34348 = n574 & ~n34347 ;
  assign n34349 = ~n26111 & n34348 ;
  assign n34350 = n17363 ^ n14605 ^ n8764 ;
  assign n34351 = n34350 ^ n21015 ^ n11236 ;
  assign n34353 = ( ~n7347 & n8288 ) | ( ~n7347 & n10690 ) | ( n8288 & n10690 ) ;
  assign n34352 = n23722 ^ n17140 ^ n14010 ;
  assign n34354 = n34353 ^ n34352 ^ n15337 ;
  assign n34355 = n15002 ^ n1477 ^ 1'b0 ;
  assign n34356 = ~n15601 & n34355 ;
  assign n34357 = ( x232 & n14625 ) | ( x232 & n34356 ) | ( n14625 & n34356 ) ;
  assign n34358 = ( ~n1266 & n12521 ) | ( ~n1266 & n34357 ) | ( n12521 & n34357 ) ;
  assign n34359 = n15650 & ~n34358 ;
  assign n34360 = n34359 ^ n32618 ^ n19568 ;
  assign n34361 = n23745 ^ n22755 ^ n17339 ;
  assign n34362 = n607 & n11285 ;
  assign n34363 = n20882 & n34362 ;
  assign n34364 = n34363 ^ n22470 ^ 1'b0 ;
  assign n34365 = n17284 | n34364 ;
  assign n34366 = n34365 ^ n22812 ^ 1'b0 ;
  assign n34367 = n25212 ^ n9908 ^ 1'b0 ;
  assign n34368 = n34367 ^ n32008 ^ n17155 ;
  assign n34369 = n5027 & n6618 ;
  assign n34370 = n34369 ^ n24447 ^ n12956 ;
  assign n34371 = ( n1293 & n25570 ) | ( n1293 & n34370 ) | ( n25570 & n34370 ) ;
  assign n34372 = n24033 ^ n21679 ^ 1'b0 ;
  assign n34373 = ( ~n13511 & n31474 ) | ( ~n13511 & n34372 ) | ( n31474 & n34372 ) ;
  assign n34374 = n8086 ^ n1830 ^ 1'b0 ;
  assign n34375 = ( n945 & n3961 ) | ( n945 & ~n21253 ) | ( n3961 & ~n21253 ) ;
  assign n34376 = n20162 | n32572 ;
  assign n34377 = n15112 & ~n34376 ;
  assign n34378 = n28214 ^ n8524 ^ 1'b0 ;
  assign n34379 = n34378 ^ n12574 ^ n4510 ;
  assign n34380 = n12663 ^ n3126 ^ n2538 ;
  assign n34381 = n8102 & n17753 ;
  assign n34382 = n5294 & n34381 ;
  assign n34383 = n34382 ^ n30520 ^ 1'b0 ;
  assign n34384 = ( n34379 & n34380 ) | ( n34379 & n34383 ) | ( n34380 & n34383 ) ;
  assign n34385 = ( n17822 & n19248 ) | ( n17822 & n28999 ) | ( n19248 & n28999 ) ;
  assign n34386 = n33943 ^ n6401 ^ x136 ;
  assign n34387 = ( n27889 & n34385 ) | ( n27889 & n34386 ) | ( n34385 & n34386 ) ;
  assign n34388 = ~n4915 & n34387 ;
  assign n34389 = n34388 ^ n13712 ^ 1'b0 ;
  assign n34390 = ( n3492 & n26111 ) | ( n3492 & n34389 ) | ( n26111 & n34389 ) ;
  assign n34391 = ( n8153 & n15000 ) | ( n8153 & ~n22263 ) | ( n15000 & ~n22263 ) ;
  assign n34392 = n34391 ^ n21789 ^ n17566 ;
  assign n34393 = n26967 ^ n23221 ^ n19093 ;
  assign n34395 = ( n5906 & n16389 ) | ( n5906 & n25640 ) | ( n16389 & n25640 ) ;
  assign n34394 = n28908 | n29225 ;
  assign n34396 = n34395 ^ n34394 ^ n1309 ;
  assign n34397 = n33728 ^ n25274 ^ 1'b0 ;
  assign n34398 = ( n1181 & n21187 ) | ( n1181 & n34397 ) | ( n21187 & n34397 ) ;
  assign n34399 = n23507 ^ n14680 ^ n1446 ;
  assign n34401 = n16156 ^ n8971 ^ n7890 ;
  assign n34402 = n8547 ^ n5118 ^ n2292 ;
  assign n34403 = n7151 & n34402 ;
  assign n34404 = ( n3378 & n16538 ) | ( n3378 & n34403 ) | ( n16538 & n34403 ) ;
  assign n34405 = n34404 ^ n13307 ^ n10161 ;
  assign n34406 = ( n14197 & n34401 ) | ( n14197 & ~n34405 ) | ( n34401 & ~n34405 ) ;
  assign n34400 = n8276 & n30752 ;
  assign n34407 = n34406 ^ n34400 ^ 1'b0 ;
  assign n34408 = n11455 | n19726 ;
  assign n34409 = n34408 ^ n12906 ^ 1'b0 ;
  assign n34410 = n33971 ^ n5916 ^ 1'b0 ;
  assign n34411 = ( n3039 & n5687 ) | ( n3039 & ~n7802 ) | ( n5687 & ~n7802 ) ;
  assign n34412 = ( n14603 & n27006 ) | ( n14603 & ~n34411 ) | ( n27006 & ~n34411 ) ;
  assign n34413 = n21129 | n34412 ;
  assign n34414 = ( n11970 & n16824 ) | ( n11970 & ~n34413 ) | ( n16824 & ~n34413 ) ;
  assign n34415 = n23962 ^ n9352 ^ n341 ;
  assign n34416 = ~n12192 & n16807 ;
  assign n34417 = n34416 ^ n17241 ^ 1'b0 ;
  assign n34418 = n34417 ^ n26940 ^ n14699 ;
  assign n34419 = ~n2051 & n8345 ;
  assign n34420 = n34419 ^ n4135 ^ 1'b0 ;
  assign n34421 = n18512 | n34420 ;
  assign n34422 = n19608 ^ n6310 ^ 1'b0 ;
  assign n34423 = n19503 & ~n34422 ;
  assign n34424 = ( n12456 & n25101 ) | ( n12456 & ~n26892 ) | ( n25101 & ~n26892 ) ;
  assign n34425 = n23849 | n34424 ;
  assign n34434 = n16951 ^ n10225 ^ 1'b0 ;
  assign n34431 = n5882 | n13597 ;
  assign n34432 = n34431 ^ n6168 ^ 1'b0 ;
  assign n34426 = n830 & n7957 ;
  assign n34427 = ~n4379 & n34426 ;
  assign n34428 = n34427 ^ n16531 ^ 1'b0 ;
  assign n34429 = ~n11580 & n34428 ;
  assign n34430 = n34429 ^ n30552 ^ n4477 ;
  assign n34433 = n34432 ^ n34430 ^ n752 ;
  assign n34435 = n34434 ^ n34433 ^ n20025 ;
  assign n34436 = ( n1179 & n1868 ) | ( n1179 & ~n32595 ) | ( n1868 & ~n32595 ) ;
  assign n34437 = ( n2182 & n10040 ) | ( n2182 & n15694 ) | ( n10040 & n15694 ) ;
  assign n34438 = ( n3293 & n32293 ) | ( n3293 & n34437 ) | ( n32293 & n34437 ) ;
  assign n34439 = n5737 & n22923 ;
  assign n34440 = ~n6561 & n34439 ;
  assign n34441 = n34440 ^ n19916 ^ n18348 ;
  assign n34442 = ( n9812 & ~n20493 ) | ( n9812 & n34441 ) | ( ~n20493 & n34441 ) ;
  assign n34443 = ( n1603 & n1933 ) | ( n1603 & n2315 ) | ( n1933 & n2315 ) ;
  assign n34444 = n34443 ^ n24344 ^ n13993 ;
  assign n34445 = n7783 & n34444 ;
  assign n34446 = n34445 ^ n29619 ^ 1'b0 ;
  assign n34447 = n15591 & n34446 ;
  assign n34448 = n17323 | n29961 ;
  assign n34449 = n9775 & ~n34448 ;
  assign n34450 = n17891 & ~n34449 ;
  assign n34458 = n31382 ^ n18946 ^ n6867 ;
  assign n34452 = ( n3411 & n8948 ) | ( n3411 & n21667 ) | ( n8948 & n21667 ) ;
  assign n34453 = n34452 ^ n5566 ^ n2393 ;
  assign n34454 = ( n15895 & n20724 ) | ( n15895 & ~n34453 ) | ( n20724 & ~n34453 ) ;
  assign n34455 = n34454 ^ n17816 ^ 1'b0 ;
  assign n34456 = ~n26290 & n34455 ;
  assign n34451 = ( n1530 & ~n12040 ) | ( n1530 & n15171 ) | ( ~n12040 & n15171 ) ;
  assign n34457 = n34456 ^ n34451 ^ n23106 ;
  assign n34459 = n34458 ^ n34457 ^ 1'b0 ;
  assign n34460 = n28962 ^ n26766 ^ n17569 ;
  assign n34461 = ~n9217 & n34460 ;
  assign n34462 = ~n8827 & n34461 ;
  assign n34463 = n5581 & ~n26951 ;
  assign n34464 = n34462 & n34463 ;
  assign n34465 = n3538 & ~n26874 ;
  assign n34466 = n34465 ^ n5596 ^ 1'b0 ;
  assign n34468 = n29281 ^ n10574 ^ 1'b0 ;
  assign n34469 = n16331 & n34468 ;
  assign n34470 = ~n11320 & n34469 ;
  assign n34471 = ( n5829 & ~n18853 ) | ( n5829 & n34470 ) | ( ~n18853 & n34470 ) ;
  assign n34467 = n1137 & n11199 ;
  assign n34472 = n34471 ^ n34467 ^ n15968 ;
  assign n34475 = n7187 ^ n7135 ^ n4279 ;
  assign n34476 = ( ~n7890 & n21702 ) | ( ~n7890 & n34475 ) | ( n21702 & n34475 ) ;
  assign n34477 = ( n12928 & ~n16029 ) | ( n12928 & n34476 ) | ( ~n16029 & n34476 ) ;
  assign n34473 = n4984 ^ x230 ^ 1'b0 ;
  assign n34474 = n4104 | n34473 ;
  assign n34478 = n34477 ^ n34474 ^ 1'b0 ;
  assign n34479 = ( n21910 & n24882 ) | ( n21910 & ~n30375 ) | ( n24882 & ~n30375 ) ;
  assign n34480 = n18901 ^ n2514 ^ n2170 ;
  assign n34481 = n18368 & ~n34480 ;
  assign n34482 = n34481 ^ n26581 ^ 1'b0 ;
  assign n34483 = n11424 ^ n3542 ^ 1'b0 ;
  assign n34484 = n5860 & n23183 ;
  assign n34485 = ~n2524 & n34484 ;
  assign n34486 = n4201 & ~n15880 ;
  assign n34487 = n34486 ^ n11825 ^ 1'b0 ;
  assign n34488 = ( n4030 & ~n7010 ) | ( n4030 & n34487 ) | ( ~n7010 & n34487 ) ;
  assign n34490 = n10660 & n29135 ;
  assign n34489 = n28604 ^ n21179 ^ 1'b0 ;
  assign n34491 = n34490 ^ n34489 ^ n12270 ;
  assign n34492 = n7084 & n11245 ;
  assign n34493 = n3699 & n34492 ;
  assign n34494 = n8613 & n20645 ;
  assign n34495 = n34494 ^ n28906 ^ 1'b0 ;
  assign n34496 = ~n34493 & n34495 ;
  assign n34497 = n34496 ^ n15056 ^ n5690 ;
  assign n34498 = ~n12690 & n18738 ;
  assign n34499 = ( n5860 & n21201 ) | ( n5860 & n34498 ) | ( n21201 & n34498 ) ;
  assign n34500 = ~n20835 & n34499 ;
  assign n34501 = ~n29409 & n34500 ;
  assign n34502 = n12059 ^ n4239 ^ 1'b0 ;
  assign n34503 = n20359 | n34502 ;
  assign n34504 = ( ~n15316 & n20400 ) | ( ~n15316 & n34412 ) | ( n20400 & n34412 ) ;
  assign n34505 = n13248 & n15194 ;
  assign n34506 = n17869 & ~n34505 ;
  assign n34509 = ( ~n1454 & n1498 ) | ( ~n1454 & n9331 ) | ( n1498 & n9331 ) ;
  assign n34510 = ( n3137 & n19070 ) | ( n3137 & ~n34509 ) | ( n19070 & ~n34509 ) ;
  assign n34507 = n10303 ^ n1717 ^ n1611 ;
  assign n34508 = ~n32294 & n34507 ;
  assign n34511 = n34510 ^ n34508 ^ n18642 ;
  assign n34512 = n6394 ^ n690 ^ 1'b0 ;
  assign n34513 = n23439 | n34512 ;
  assign n34514 = n7325 & ~n11209 ;
  assign n34515 = ~n5578 & n34514 ;
  assign n34516 = n22557 ^ n2849 ^ 1'b0 ;
  assign n34517 = n34515 | n34516 ;
  assign n34518 = ( n4406 & ~n6429 ) | ( n4406 & n26287 ) | ( ~n6429 & n26287 ) ;
  assign n34519 = ( n5770 & n6767 ) | ( n5770 & ~n33109 ) | ( n6767 & ~n33109 ) ;
  assign n34520 = n22960 ^ n11291 ^ n10049 ;
  assign n34521 = n30366 ^ n4425 ^ 1'b0 ;
  assign n34522 = ( ~n23085 & n26927 ) | ( ~n23085 & n34521 ) | ( n26927 & n34521 ) ;
  assign n34523 = ~n8082 & n30651 ;
  assign n34524 = n32574 & n34523 ;
  assign n34525 = ( n27660 & n34522 ) | ( n27660 & n34524 ) | ( n34522 & n34524 ) ;
  assign n34526 = ( ~n15725 & n17407 ) | ( ~n15725 & n21819 ) | ( n17407 & n21819 ) ;
  assign n34527 = n33106 ^ n28351 ^ n7973 ;
  assign n34528 = ( n5285 & ~n34526 ) | ( n5285 & n34527 ) | ( ~n34526 & n34527 ) ;
  assign n34529 = n9692 ^ n8944 ^ n1599 ;
  assign n34530 = n1309 & n5179 ;
  assign n34531 = ( ~n17803 & n30219 ) | ( ~n17803 & n34530 ) | ( n30219 & n34530 ) ;
  assign n34532 = n28228 ^ n2011 ^ 1'b0 ;
  assign n34533 = n34531 | n34532 ;
  assign n34534 = ( n9486 & n13794 ) | ( n9486 & n22087 ) | ( n13794 & n22087 ) ;
  assign n34535 = n25305 & ~n34534 ;
  assign n34536 = ~n6577 & n23136 ;
  assign n34537 = ( n17803 & n25510 ) | ( n17803 & ~n31063 ) | ( n25510 & ~n31063 ) ;
  assign n34538 = ( ~n8673 & n13566 ) | ( ~n8673 & n24821 ) | ( n13566 & n24821 ) ;
  assign n34539 = n34538 ^ n22192 ^ n6709 ;
  assign n34540 = n6366 ^ n3710 ^ 1'b0 ;
  assign n34546 = n24283 ^ n20744 ^ n6075 ;
  assign n34543 = n357 & n8415 ;
  assign n34544 = ~n10250 & n34543 ;
  assign n34545 = ( n15870 & ~n17383 ) | ( n15870 & n34544 ) | ( ~n17383 & n34544 ) ;
  assign n34541 = n12686 ^ n9792 ^ 1'b0 ;
  assign n34542 = n34541 ^ n22524 ^ n19878 ;
  assign n34547 = n34546 ^ n34545 ^ n34542 ;
  assign n34548 = ( n2584 & n10007 ) | ( n2584 & n19715 ) | ( n10007 & n19715 ) ;
  assign n34549 = ( n1967 & ~n16898 ) | ( n1967 & n34548 ) | ( ~n16898 & n34548 ) ;
  assign n34550 = n18304 ^ n3217 ^ 1'b0 ;
  assign n34551 = ( n26219 & n33754 ) | ( n26219 & ~n34550 ) | ( n33754 & ~n34550 ) ;
  assign n34552 = ( n3889 & n5279 ) | ( n3889 & n14930 ) | ( n5279 & n14930 ) ;
  assign n34553 = n31759 ^ n10363 ^ n661 ;
  assign n34554 = n34553 ^ n20420 ^ 1'b0 ;
  assign n34555 = n1768 & ~n34554 ;
  assign n34556 = ( n8529 & ~n15333 ) | ( n8529 & n22935 ) | ( ~n15333 & n22935 ) ;
  assign n34557 = n34556 ^ n23276 ^ n6600 ;
  assign n34558 = n6221 ^ n2778 ^ 1'b0 ;
  assign n34559 = n34557 & ~n34558 ;
  assign n34560 = ( n6612 & n15254 ) | ( n6612 & ~n22180 ) | ( n15254 & ~n22180 ) ;
  assign n34561 = n1981 & n17257 ;
  assign n34562 = ~n20645 & n34561 ;
  assign n34563 = n10338 ^ n9028 ^ n4890 ;
  assign n34564 = ( ~n815 & n7221 ) | ( ~n815 & n34563 ) | ( n7221 & n34563 ) ;
  assign n34565 = n34564 ^ n33986 ^ n20942 ;
  assign n34566 = ( n1266 & n3973 ) | ( n1266 & ~n23268 ) | ( n3973 & ~n23268 ) ;
  assign n34567 = n34566 ^ n8880 ^ n6260 ;
  assign n34568 = ~n7866 & n24711 ;
  assign n34569 = n34568 ^ n16819 ^ 1'b0 ;
  assign n34570 = n34569 ^ n10776 ^ n9646 ;
  assign n34572 = n7337 & n22742 ;
  assign n34573 = n4352 & n34572 ;
  assign n34571 = n16425 ^ n13744 ^ n7292 ;
  assign n34574 = n34573 ^ n34571 ^ n22860 ;
  assign n34577 = ~n22250 & n25887 ;
  assign n34575 = n2382 & ~n9859 ;
  assign n34576 = n10815 & ~n34575 ;
  assign n34578 = n34577 ^ n34576 ^ n1851 ;
  assign n34579 = n26206 ^ n17863 ^ 1'b0 ;
  assign n34580 = n31076 ^ n11031 ^ 1'b0 ;
  assign n34581 = n30392 ^ n1272 ^ 1'b0 ;
  assign n34582 = ~n17111 & n34581 ;
  assign n34583 = n34582 ^ n23354 ^ n10027 ;
  assign n34584 = ( ~n11579 & n34580 ) | ( ~n11579 & n34583 ) | ( n34580 & n34583 ) ;
  assign n34585 = n30896 ^ n17903 ^ n15980 ;
  assign n34586 = n6265 ^ n2678 ^ 1'b0 ;
  assign n34587 = ( n5206 & n12827 ) | ( n5206 & ~n22278 ) | ( n12827 & ~n22278 ) ;
  assign n34588 = n3383 | n34587 ;
  assign n34589 = n33012 ^ n2835 ^ 1'b0 ;
  assign n34590 = n32287 ^ n1526 ^ 1'b0 ;
  assign n34591 = ( ~n755 & n31211 ) | ( ~n755 & n34590 ) | ( n31211 & n34590 ) ;
  assign n34592 = n10500 & ~n18038 ;
  assign n34593 = n8685 ^ n6596 ^ 1'b0 ;
  assign n34594 = ~n9883 & n34593 ;
  assign n34595 = n34594 ^ n11550 ^ n2039 ;
  assign n34596 = n34595 ^ n4017 ^ n1196 ;
  assign n34597 = n34596 ^ n21674 ^ 1'b0 ;
  assign n34598 = n9310 & n34597 ;
  assign n34600 = n33024 ^ n21473 ^ 1'b0 ;
  assign n34599 = n17966 ^ n8929 ^ n1955 ;
  assign n34601 = n34600 ^ n34599 ^ n3163 ;
  assign n34602 = ( n20190 & n24597 ) | ( n20190 & ~n34601 ) | ( n24597 & ~n34601 ) ;
  assign n34603 = n6936 & ~n34602 ;
  assign n34604 = ~n19811 & n34603 ;
  assign n34605 = ( n7794 & n23691 ) | ( n7794 & ~n23904 ) | ( n23691 & ~n23904 ) ;
  assign n34606 = ~n9722 & n21479 ;
  assign n34607 = n10188 & ~n13778 ;
  assign n34608 = n34607 ^ n17302 ^ 1'b0 ;
  assign n34609 = n34608 ^ n24442 ^ 1'b0 ;
  assign n34610 = ( n705 & n8606 ) | ( n705 & n10644 ) | ( n8606 & n10644 ) ;
  assign n34611 = ( n9467 & n26994 ) | ( n9467 & ~n34610 ) | ( n26994 & ~n34610 ) ;
  assign n34612 = n3853 & ~n10907 ;
  assign n34613 = n2852 & n34612 ;
  assign n34614 = n34613 ^ n16476 ^ n12998 ;
  assign n34615 = n34614 ^ n25586 ^ n1031 ;
  assign n34616 = n2974 & ~n13604 ;
  assign n34617 = ~n17985 & n34616 ;
  assign n34619 = x5 & ~n12263 ;
  assign n34620 = n34619 ^ n27848 ^ 1'b0 ;
  assign n34621 = ( n8089 & ~n25906 ) | ( n8089 & n34620 ) | ( ~n25906 & n34620 ) ;
  assign n34618 = n8087 ^ n1852 ^ n975 ;
  assign n34622 = n34621 ^ n34618 ^ n2173 ;
  assign n34623 = ( ~n4296 & n9716 ) | ( ~n4296 & n13191 ) | ( n9716 & n13191 ) ;
  assign n34624 = n34623 ^ n12733 ^ n11851 ;
  assign n34625 = n25433 & n34624 ;
  assign n34626 = ( n25179 & n34622 ) | ( n25179 & n34625 ) | ( n34622 & n34625 ) ;
  assign n34627 = n25938 & n34626 ;
  assign n34628 = ( ~n12946 & n34617 ) | ( ~n12946 & n34627 ) | ( n34617 & n34627 ) ;
  assign n34629 = n6747 | n30660 ;
  assign n34630 = n13546 | n34629 ;
  assign n34631 = ( ~n3406 & n21549 ) | ( ~n3406 & n34630 ) | ( n21549 & n34630 ) ;
  assign n34632 = n34631 ^ n22860 ^ 1'b0 ;
  assign n34633 = ( n21508 & ~n26255 ) | ( n21508 & n34632 ) | ( ~n26255 & n34632 ) ;
  assign n34634 = n6352 ^ n2452 ^ n1823 ;
  assign n34635 = n34634 ^ n10807 ^ n4589 ;
  assign n34636 = ( n10929 & n31776 ) | ( n10929 & ~n33145 ) | ( n31776 & ~n33145 ) ;
  assign n34637 = n13887 & ~n26553 ;
  assign n34638 = n34637 ^ n1785 ^ 1'b0 ;
  assign n34639 = ( n1130 & n25506 ) | ( n1130 & n26311 ) | ( n25506 & n26311 ) ;
  assign n34640 = ( n19314 & n34638 ) | ( n19314 & ~n34639 ) | ( n34638 & ~n34639 ) ;
  assign n34641 = n11075 ^ n4324 ^ 1'b0 ;
  assign n34642 = n18025 ^ n11115 ^ 1'b0 ;
  assign n34643 = n34641 & ~n34642 ;
  assign n34644 = n34643 ^ n10777 ^ 1'b0 ;
  assign n34645 = ( n8669 & n12780 ) | ( n8669 & ~n13100 ) | ( n12780 & ~n13100 ) ;
  assign n34646 = n34645 ^ n21411 ^ 1'b0 ;
  assign n34647 = ~n34644 & n34646 ;
  assign n34648 = n30784 ^ n30490 ^ n3951 ;
  assign n34649 = n34648 ^ n10189 ^ 1'b0 ;
  assign n34650 = n11316 | n34649 ;
  assign n34651 = ( n1826 & ~n2934 ) | ( n1826 & n6708 ) | ( ~n2934 & n6708 ) ;
  assign n34652 = n25858 ^ n15616 ^ 1'b0 ;
  assign n34654 = n31730 ^ n15434 ^ n8949 ;
  assign n34653 = ( n8435 & ~n13645 ) | ( n8435 & n18741 ) | ( ~n13645 & n18741 ) ;
  assign n34655 = n34654 ^ n34653 ^ n24366 ;
  assign n34656 = n20556 ^ n3866 ^ 1'b0 ;
  assign n34657 = ( n1064 & ~n6105 ) | ( n1064 & n34656 ) | ( ~n6105 & n34656 ) ;
  assign n34658 = n16824 & n21836 ;
  assign n34659 = n9380 & n34658 ;
  assign n34661 = n7521 & n11719 ;
  assign n34662 = n34661 ^ n6971 ^ 1'b0 ;
  assign n34660 = n1860 & n2641 ;
  assign n34663 = n34662 ^ n34660 ^ 1'b0 ;
  assign n34664 = n6138 & ~n21376 ;
  assign n34665 = n12909 ^ n8697 ^ n5884 ;
  assign n34666 = ( ~n1865 & n32072 ) | ( ~n1865 & n33236 ) | ( n32072 & n33236 ) ;
  assign n34667 = ~n34665 & n34666 ;
  assign n34668 = n34667 ^ n3486 ^ 1'b0 ;
  assign n34669 = ( n1332 & ~n12669 ) | ( n1332 & n14582 ) | ( ~n12669 & n14582 ) ;
  assign n34670 = n33601 | n34669 ;
  assign n34671 = n34670 ^ n20909 ^ 1'b0 ;
  assign n34672 = ( n3263 & ~n9439 ) | ( n3263 & n26814 ) | ( ~n9439 & n26814 ) ;
  assign n34673 = n34672 ^ n21816 ^ 1'b0 ;
  assign n34674 = n34673 ^ n7155 ^ 1'b0 ;
  assign n34675 = ~n2164 & n2367 ;
  assign n34676 = n5911 & ~n24051 ;
  assign n34677 = n21512 & n34676 ;
  assign n34678 = n34677 ^ n28221 ^ n2133 ;
  assign n34679 = ( n7597 & n15114 ) | ( n7597 & ~n25518 ) | ( n15114 & ~n25518 ) ;
  assign n34680 = ( n18715 & n24882 ) | ( n18715 & ~n34679 ) | ( n24882 & ~n34679 ) ;
  assign n34681 = n5416 | n34680 ;
  assign n34682 = n34681 ^ n30570 ^ 1'b0 ;
  assign n34683 = n29721 ^ n10140 ^ n4161 ;
  assign n34684 = n34683 ^ n10033 ^ n3889 ;
  assign n34685 = n34684 ^ n28159 ^ n26988 ;
  assign n34686 = n25610 | n27486 ;
  assign n34687 = n14733 | n22634 ;
  assign n34688 = n20885 ^ n15141 ^ n11067 ;
  assign n34689 = n4172 | n32222 ;
  assign n34690 = n15186 | n24426 ;
  assign n34691 = n15056 & ~n34690 ;
  assign n34693 = ( n3164 & n13739 ) | ( n3164 & n30889 ) | ( n13739 & n30889 ) ;
  assign n34694 = n34693 ^ n4832 ^ n492 ;
  assign n34692 = n10792 ^ n6085 ^ n5674 ;
  assign n34695 = n34694 ^ n34692 ^ x214 ;
  assign n34696 = n34695 ^ n7021 ^ n4526 ;
  assign n34697 = ~n1595 & n1761 ;
  assign n34698 = n34697 ^ n1974 ^ 1'b0 ;
  assign n34699 = ( n7889 & ~n8147 ) | ( n7889 & n34698 ) | ( ~n8147 & n34698 ) ;
  assign n34700 = n25936 ^ n5367 ^ 1'b0 ;
  assign n34701 = n34700 ^ n19259 ^ 1'b0 ;
  assign n34702 = n8688 | n34701 ;
  assign n34703 = ( n30904 & ~n34699 ) | ( n30904 & n34702 ) | ( ~n34699 & n34702 ) ;
  assign n34704 = n34703 ^ n19677 ^ 1'b0 ;
  assign n34705 = n34696 | n34704 ;
  assign n34706 = n20839 ^ n2445 ^ 1'b0 ;
  assign n34707 = n12241 ^ n5911 ^ 1'b0 ;
  assign n34708 = n34707 ^ n24227 ^ n8931 ;
  assign n34709 = n34708 ^ n9579 ^ 1'b0 ;
  assign n34710 = n34709 ^ n33146 ^ n5134 ;
  assign n34711 = n8374 ^ n4479 ^ 1'b0 ;
  assign n34712 = ~n15314 & n34711 ;
  assign n34713 = n34712 ^ n12850 ^ n7658 ;
  assign n34715 = n5444 ^ n1784 ^ n501 ;
  assign n34714 = ~n14996 & n29481 ;
  assign n34716 = n34715 ^ n34714 ^ 1'b0 ;
  assign n34717 = ( n6109 & n21025 ) | ( n6109 & ~n25529 ) | ( n21025 & ~n25529 ) ;
  assign n34718 = n32459 ^ n15316 ^ n10545 ;
  assign n34719 = ( n8520 & n19424 ) | ( n8520 & ~n34718 ) | ( n19424 & ~n34718 ) ;
  assign n34720 = n9525 | n18679 ;
  assign n34721 = n34720 ^ n34587 ^ n2452 ;
  assign n34722 = n25769 ^ n9358 ^ n2232 ;
  assign n34723 = n2586 | n7792 ;
  assign n34724 = n4939 | n34723 ;
  assign n34725 = n3914 & ~n34724 ;
  assign n34726 = n34725 ^ n10236 ^ n7434 ;
  assign n34727 = n4774 ^ n3885 ^ 1'b0 ;
  assign n34728 = ~n34726 & n34727 ;
  assign n34729 = n23827 ^ n22443 ^ 1'b0 ;
  assign n34730 = n13709 & ~n34729 ;
  assign n34732 = n1634 | n10384 ;
  assign n34733 = n25497 | n34732 ;
  assign n34731 = n19461 ^ n16612 ^ n10981 ;
  assign n34734 = n34733 ^ n34731 ^ n28339 ;
  assign n34735 = ( n4588 & n20924 ) | ( n4588 & ~n22224 ) | ( n20924 & ~n22224 ) ;
  assign n34736 = n7776 ^ n3526 ^ 1'b0 ;
  assign n34737 = n8756 & ~n34736 ;
  assign n34738 = n9028 ^ n6868 ^ 1'b0 ;
  assign n34739 = ~n30383 & n34738 ;
  assign n34740 = ( n3309 & n17148 ) | ( n3309 & ~n30552 ) | ( n17148 & ~n30552 ) ;
  assign n34741 = n7417 ^ n4391 ^ 1'b0 ;
  assign n34742 = ~n15994 & n34741 ;
  assign n34743 = n4741 & n34742 ;
  assign n34744 = n34740 & n34743 ;
  assign n34745 = n24890 ^ n18432 ^ n17745 ;
  assign n34746 = ( n8357 & n34453 ) | ( n8357 & n34745 ) | ( n34453 & n34745 ) ;
  assign n34747 = n13576 ^ n4198 ^ x77 ;
  assign n34748 = n13964 | n34747 ;
  assign n34751 = n28065 ^ n17190 ^ n9605 ;
  assign n34749 = n22787 ^ n19792 ^ n275 ;
  assign n34750 = n34749 ^ n10036 ^ 1'b0 ;
  assign n34752 = n34751 ^ n34750 ^ 1'b0 ;
  assign n34753 = n11791 & n16806 ;
  assign n34754 = n34753 ^ n20844 ^ n408 ;
  assign n34755 = ( n9840 & n18882 ) | ( n9840 & n34754 ) | ( n18882 & n34754 ) ;
  assign n34757 = n9318 ^ n5915 ^ n2797 ;
  assign n34758 = ~n3068 & n34757 ;
  assign n34759 = n34758 ^ n1484 ^ 1'b0 ;
  assign n34760 = ( n4769 & ~n13631 ) | ( n4769 & n34759 ) | ( ~n13631 & n34759 ) ;
  assign n34756 = n23598 ^ n9042 ^ 1'b0 ;
  assign n34761 = n34760 ^ n34756 ^ n5432 ;
  assign n34762 = n17978 & n32395 ;
  assign n34763 = ( n5626 & n15681 ) | ( n5626 & n34762 ) | ( n15681 & n34762 ) ;
  assign n34764 = ( n5274 & n17775 ) | ( n5274 & ~n34763 ) | ( n17775 & ~n34763 ) ;
  assign n34765 = n29491 ^ n15270 ^ n9580 ;
  assign n34766 = ( n9450 & n19684 ) | ( n9450 & ~n34765 ) | ( n19684 & ~n34765 ) ;
  assign n34767 = n30468 ^ n20794 ^ 1'b0 ;
  assign n34768 = ( n25138 & ~n34406 ) | ( n25138 & n34767 ) | ( ~n34406 & n34767 ) ;
  assign n34769 = n9373 | n21079 ;
  assign n34770 = n17905 | n34769 ;
  assign n34771 = n34770 ^ n28450 ^ 1'b0 ;
  assign n34772 = n6396 ^ n2125 ^ 1'b0 ;
  assign n34773 = n975 | n6434 ;
  assign n34774 = n15154 | n34773 ;
  assign n34775 = n11878 ^ n3986 ^ 1'b0 ;
  assign n34776 = n34775 ^ n11817 ^ 1'b0 ;
  assign n34777 = n34776 ^ n13556 ^ n10509 ;
  assign n34778 = n34777 ^ n30600 ^ 1'b0 ;
  assign n34779 = ( n15145 & ~n16979 ) | ( n15145 & n20943 ) | ( ~n16979 & n20943 ) ;
  assign n34780 = n10338 ^ n5208 ^ 1'b0 ;
  assign n34781 = n22448 | n26682 ;
  assign n34782 = n34780 & ~n34781 ;
  assign n34783 = n34782 ^ n16188 ^ n8513 ;
  assign n34784 = n16248 ^ n3207 ^ 1'b0 ;
  assign n34785 = n27708 ^ n11602 ^ n2852 ;
  assign n34786 = n3707 & ~n5452 ;
  assign n34787 = ( n5211 & n34785 ) | ( n5211 & n34786 ) | ( n34785 & n34786 ) ;
  assign n34788 = n34787 ^ n1965 ^ 1'b0 ;
  assign n34789 = n18837 & ~n34788 ;
  assign n34790 = ( n2450 & n11540 ) | ( n2450 & n19248 ) | ( n11540 & n19248 ) ;
  assign n34791 = n17387 ^ n8707 ^ n8438 ;
  assign n34792 = n32653 ^ n14158 ^ x114 ;
  assign n34793 = ~n4148 & n17853 ;
  assign n34794 = n34793 ^ n4036 ^ 1'b0 ;
  assign n34795 = n22280 | n25266 ;
  assign n34796 = n31727 ^ n26669 ^ 1'b0 ;
  assign n34797 = ( n6702 & ~n21910 ) | ( n6702 & n26738 ) | ( ~n21910 & n26738 ) ;
  assign n34798 = n34797 ^ n8255 ^ 1'b0 ;
  assign n34799 = n905 | n13057 ;
  assign n34800 = n34799 ^ n6030 ^ 1'b0 ;
  assign n34801 = ( n29634 & n33973 ) | ( n29634 & n34800 ) | ( n33973 & n34800 ) ;
  assign n34802 = ( n10150 & ~n28602 ) | ( n10150 & n31920 ) | ( ~n28602 & n31920 ) ;
  assign n34803 = ~n1760 & n12339 ;
  assign n34804 = n29671 ^ n13706 ^ n10800 ;
  assign n34805 = n6480 | n18592 ;
  assign n34806 = n34805 ^ n15056 ^ 1'b0 ;
  assign n34807 = n34806 ^ n23904 ^ n3103 ;
  assign n34808 = ~n32211 & n34807 ;
  assign n34809 = n34808 ^ n2892 ^ 1'b0 ;
  assign n34810 = n2085 | n12714 ;
  assign n34811 = n34809 | n34810 ;
  assign n34812 = ~n16462 & n18472 ;
  assign n34813 = n2390 | n2646 ;
  assign n34814 = n34813 ^ n7754 ^ 1'b0 ;
  assign n34815 = ~n268 & n5237 ;
  assign n34816 = n7293 & n34815 ;
  assign n34817 = n11359 & ~n34816 ;
  assign n34818 = n34817 ^ n4894 ^ 1'b0 ;
  assign n34819 = ( n11341 & n13327 ) | ( n11341 & ~n34818 ) | ( n13327 & ~n34818 ) ;
  assign n34820 = ( n16669 & n24080 ) | ( n16669 & n34819 ) | ( n24080 & n34819 ) ;
  assign n34821 = n34820 ^ n25699 ^ 1'b0 ;
  assign n34822 = n25413 ^ n3229 ^ 1'b0 ;
  assign n34823 = n34821 | n34822 ;
  assign n34824 = n11339 ^ n6114 ^ 1'b0 ;
  assign n34825 = n9072 | n34824 ;
  assign n34826 = n34823 & ~n34825 ;
  assign n34827 = ( ~n8360 & n34814 ) | ( ~n8360 & n34826 ) | ( n34814 & n34826 ) ;
  assign n34828 = ( n16582 & ~n25550 ) | ( n16582 & n33452 ) | ( ~n25550 & n33452 ) ;
  assign n34829 = ~n2752 & n10734 ;
  assign n34830 = n28295 & n34829 ;
  assign n34831 = ( n14560 & ~n34828 ) | ( n14560 & n34830 ) | ( ~n34828 & n34830 ) ;
  assign n34832 = n17053 ^ n12680 ^ n6470 ;
  assign n34833 = n23873 ^ n3456 ^ n581 ;
  assign n34834 = n32308 ^ n1991 ^ 1'b0 ;
  assign n34835 = n34833 & ~n34834 ;
  assign n34836 = ( n21976 & ~n23368 ) | ( n21976 & n23914 ) | ( ~n23368 & n23914 ) ;
  assign n34837 = n34836 ^ n15157 ^ n4517 ;
  assign n34838 = n34837 ^ n23256 ^ n21269 ;
  assign n34839 = n2408 & ~n3016 ;
  assign n34840 = ( n6947 & n34838 ) | ( n6947 & ~n34839 ) | ( n34838 & ~n34839 ) ;
  assign n34841 = ( ~n31736 & n34835 ) | ( ~n31736 & n34840 ) | ( n34835 & n34840 ) ;
  assign n34842 = n7857 & n15756 ;
  assign n34843 = ( n20878 & n30651 ) | ( n20878 & n34842 ) | ( n30651 & n34842 ) ;
  assign n34844 = n24752 & n34303 ;
  assign n34845 = ( n7324 & n26072 ) | ( n7324 & n32442 ) | ( n26072 & n32442 ) ;
  assign n34847 = ( n287 & n3597 ) | ( n287 & ~n13113 ) | ( n3597 & ~n13113 ) ;
  assign n34848 = ( n4570 & n5700 ) | ( n4570 & n20446 ) | ( n5700 & n20446 ) ;
  assign n34849 = ( n1505 & n34847 ) | ( n1505 & n34848 ) | ( n34847 & n34848 ) ;
  assign n34846 = n15697 & n21400 ;
  assign n34850 = n34849 ^ n34846 ^ 1'b0 ;
  assign n34851 = ( n11908 & n18251 ) | ( n11908 & n30997 ) | ( n18251 & n30997 ) ;
  assign n34852 = ( n1679 & ~n21060 ) | ( n1679 & n34851 ) | ( ~n21060 & n34851 ) ;
  assign n34853 = ~n7371 & n7942 ;
  assign n34854 = ( ~n1046 & n4116 ) | ( ~n1046 & n34853 ) | ( n4116 & n34853 ) ;
  assign n34855 = n34854 ^ n30128 ^ n3853 ;
  assign n34856 = n22935 ^ n6218 ^ 1'b0 ;
  assign n34857 = n11592 & n34856 ;
  assign n34858 = n34857 ^ n18596 ^ n14720 ;
  assign n34859 = n1232 & n12363 ;
  assign n34860 = n34859 ^ n22666 ^ 1'b0 ;
  assign n34863 = n2934 | n21854 ;
  assign n34864 = n968 & ~n34863 ;
  assign n34861 = n14681 ^ n11152 ^ 1'b0 ;
  assign n34862 = n34861 ^ n7080 ^ n2728 ;
  assign n34865 = n34864 ^ n34862 ^ n25734 ;
  assign n34866 = n1455 & ~n34865 ;
  assign n34867 = ~n19352 & n34866 ;
  assign n34868 = n34867 ^ n15515 ^ n3064 ;
  assign n34870 = n5075 ^ n3949 ^ 1'b0 ;
  assign n34871 = n17066 & n34870 ;
  assign n34869 = ( x177 & n4089 ) | ( x177 & ~n10410 ) | ( n4089 & ~n10410 ) ;
  assign n34872 = n34871 ^ n34869 ^ x239 ;
  assign n34873 = n34872 ^ n6413 ^ n5815 ;
  assign n34874 = n28934 ^ n6294 ^ 1'b0 ;
  assign n34875 = n12901 | n34874 ;
  assign n34876 = n30021 ^ n6404 ^ 1'b0 ;
  assign n34877 = ( n12217 & n34819 ) | ( n12217 & ~n34876 ) | ( n34819 & ~n34876 ) ;
  assign n34878 = n34877 ^ n5498 ^ 1'b0 ;
  assign n34879 = n34878 ^ n29600 ^ n9969 ;
  assign n34880 = n12774 ^ n7293 ^ 1'b0 ;
  assign n34881 = n34880 ^ n33547 ^ n29899 ;
  assign n34882 = ( n6073 & ~n28908 ) | ( n6073 & n34569 ) | ( ~n28908 & n34569 ) ;
  assign n34883 = n18237 ^ n10930 ^ 1'b0 ;
  assign n34884 = ( n5685 & n7709 ) | ( n5685 & n34883 ) | ( n7709 & n34883 ) ;
  assign n34885 = n34884 ^ n31255 ^ n1087 ;
  assign n34886 = n34885 ^ n11065 ^ n2974 ;
  assign n34887 = n34867 ^ n16379 ^ n13551 ;
  assign n34888 = n34887 ^ n22167 ^ n11115 ;
  assign n34889 = n994 & ~n2311 ;
  assign n34890 = n8630 & n34889 ;
  assign n34893 = n9380 ^ n7322 ^ x227 ;
  assign n34894 = n34893 ^ n614 ^ 1'b0 ;
  assign n34891 = ( n11704 & n24149 ) | ( n11704 & n32851 ) | ( n24149 & n32851 ) ;
  assign n34892 = n9784 | n34891 ;
  assign n34895 = n34894 ^ n34892 ^ 1'b0 ;
  assign n34896 = n31127 ^ n26188 ^ 1'b0 ;
  assign n34897 = ~n10075 & n34896 ;
  assign n34898 = ~n12476 & n34897 ;
  assign n34899 = n5309 | n13448 ;
  assign n34900 = n34898 & ~n34899 ;
  assign n34901 = ( n10007 & n31572 ) | ( n10007 & ~n31919 ) | ( n31572 & ~n31919 ) ;
  assign n34902 = n6616 | n8226 ;
  assign n34903 = n29919 ^ n10597 ^ n2018 ;
  assign n34904 = ( n2854 & ~n4170 ) | ( n2854 & n34903 ) | ( ~n4170 & n34903 ) ;
  assign n34905 = n15919 ^ n12234 ^ n9822 ;
  assign n34906 = n34905 ^ n23478 ^ n15422 ;
  assign n34909 = n20032 ^ n7471 ^ 1'b0 ;
  assign n34910 = n34101 & n34909 ;
  assign n34907 = ( n11061 & n12955 ) | ( n11061 & ~n32999 ) | ( n12955 & ~n32999 ) ;
  assign n34908 = ~n9097 & n34907 ;
  assign n34911 = n34910 ^ n34908 ^ 1'b0 ;
  assign n34913 = n17508 ^ n6687 ^ n6682 ;
  assign n34912 = n11731 & ~n17343 ;
  assign n34914 = n34913 ^ n34912 ^ 1'b0 ;
  assign n34918 = n16355 ^ n12620 ^ n363 ;
  assign n34919 = n30061 | n34918 ;
  assign n34920 = n19439 | n34919 ;
  assign n34915 = ~n4422 & n20623 ;
  assign n34916 = n34915 ^ n5178 ^ 1'b0 ;
  assign n34917 = n1846 & n34916 ;
  assign n34921 = n34920 ^ n34917 ^ 1'b0 ;
  assign n34922 = ( n6527 & n14682 ) | ( n6527 & ~n16344 ) | ( n14682 & ~n16344 ) ;
  assign n34923 = n34922 ^ n12803 ^ 1'b0 ;
  assign n34924 = n7984 ^ n4901 ^ 1'b0 ;
  assign n34925 = n34924 ^ n4311 ^ n3128 ;
  assign n34926 = n34925 ^ n23687 ^ x109 ;
  assign n34927 = n27313 ^ n859 ^ 1'b0 ;
  assign n34928 = ~n26404 & n34927 ;
  assign n34929 = ( ~n621 & n16411 ) | ( ~n621 & n20595 ) | ( n16411 & n20595 ) ;
  assign n34930 = n34929 ^ n15814 ^ n5796 ;
  assign n34931 = n34930 ^ n21503 ^ 1'b0 ;
  assign n34932 = n21471 & n34931 ;
  assign n34935 = n10202 & n20741 ;
  assign n34936 = n34935 ^ n18735 ^ 1'b0 ;
  assign n34933 = n22869 ^ n15473 ^ 1'b0 ;
  assign n34934 = n28821 & ~n34933 ;
  assign n34937 = n34936 ^ n34934 ^ n12231 ;
  assign n34938 = n28357 ^ n21734 ^ n2097 ;
  assign n34939 = n17348 ^ n6224 ^ 1'b0 ;
  assign n34940 = ~n22235 & n34939 ;
  assign n34941 = ( ~n3493 & n7535 ) | ( ~n3493 & n19240 ) | ( n7535 & n19240 ) ;
  assign n34942 = ( n11824 & ~n34940 ) | ( n11824 & n34941 ) | ( ~n34940 & n34941 ) ;
  assign n34943 = n31760 ^ n22449 ^ n12931 ;
  assign n34944 = n15136 ^ n1241 ^ 1'b0 ;
  assign n34945 = ~n20521 & n34944 ;
  assign n34946 = ( n16091 & n16606 ) | ( n16091 & n34945 ) | ( n16606 & n34945 ) ;
  assign n34947 = ( n8938 & ~n9012 ) | ( n8938 & n34946 ) | ( ~n9012 & n34946 ) ;
  assign n34948 = n27446 ^ n602 ^ 1'b0 ;
  assign n34949 = n34947 & ~n34948 ;
  assign n34950 = n28301 ^ n25569 ^ n13104 ;
  assign n34951 = n750 | n21431 ;
  assign n34953 = ( ~n2868 & n20310 ) | ( ~n2868 & n33901 ) | ( n20310 & n33901 ) ;
  assign n34954 = n34953 ^ n21831 ^ n19518 ;
  assign n34952 = n11408 ^ n9473 ^ n2631 ;
  assign n34955 = n34954 ^ n34952 ^ 1'b0 ;
  assign n34956 = n5309 ^ n2649 ^ 1'b0 ;
  assign n34957 = ( n291 & n20006 ) | ( n291 & n34956 ) | ( n20006 & n34956 ) ;
  assign n34958 = n12219 ^ n4476 ^ 1'b0 ;
  assign n34959 = n24003 & n34958 ;
  assign n34960 = n18414 ^ n6048 ^ 1'b0 ;
  assign n34961 = ( n9131 & n25533 ) | ( n9131 & ~n34960 ) | ( n25533 & ~n34960 ) ;
  assign n34962 = n17727 ^ n13751 ^ n3205 ;
  assign n34963 = ( n13205 & n15814 ) | ( n13205 & ~n21289 ) | ( n15814 & ~n21289 ) ;
  assign n34964 = n34963 ^ n27263 ^ n14320 ;
  assign n34965 = ~n22046 & n34964 ;
  assign n34966 = n8983 | n20533 ;
  assign n34967 = ( n34048 & n34437 ) | ( n34048 & ~n34966 ) | ( n34437 & ~n34966 ) ;
  assign n34968 = ( ~n621 & n644 ) | ( ~n621 & n13294 ) | ( n644 & n13294 ) ;
  assign n34969 = ( n2914 & n14524 ) | ( n2914 & n34968 ) | ( n14524 & n34968 ) ;
  assign n34970 = n32978 & ~n34969 ;
  assign n34971 = ~n22446 & n34970 ;
  assign n34972 = ( n8535 & n12606 ) | ( n8535 & n21040 ) | ( n12606 & n21040 ) ;
  assign n34973 = n26077 ^ n10023 ^ 1'b0 ;
  assign n34974 = n9007 & n34973 ;
  assign n34975 = ( n16289 & n34972 ) | ( n16289 & n34974 ) | ( n34972 & n34974 ) ;
  assign n34976 = n27859 ^ n7753 ^ 1'b0 ;
  assign n34977 = n34976 ^ n30317 ^ n2522 ;
  assign n34978 = n19225 & ~n34977 ;
  assign n34979 = n34975 & n34978 ;
  assign n34980 = n23796 ^ n10627 ^ 1'b0 ;
  assign n34981 = n34979 | n34980 ;
  assign n34982 = n13759 & n17694 ;
  assign n34984 = n21263 ^ n15042 ^ n5874 ;
  assign n34985 = n2468 | n14941 ;
  assign n34986 = n9093 & ~n34985 ;
  assign n34987 = n18119 | n34986 ;
  assign n34988 = n34984 & ~n34987 ;
  assign n34983 = n5689 & n27016 ;
  assign n34989 = n34988 ^ n34983 ^ n10771 ;
  assign n34990 = n24234 ^ n14571 ^ n5032 ;
  assign n34991 = ~n4238 & n20256 ;
  assign n34992 = n34990 & n34991 ;
  assign n34993 = n365 & n14895 ;
  assign n34994 = ( ~n7741 & n32510 ) | ( ~n7741 & n33132 ) | ( n32510 & n33132 ) ;
  assign n34995 = n34994 ^ n2738 ^ n1367 ;
  assign n34996 = n34995 ^ n25139 ^ n8569 ;
  assign n34997 = n7761 ^ n1587 ^ 1'b0 ;
  assign n34998 = ~n14649 & n24335 ;
  assign n34999 = n2278 & ~n29178 ;
  assign n35000 = n31441 & n34999 ;
  assign n35001 = n5412 & ~n19564 ;
  assign n35002 = n35001 ^ n24317 ^ 1'b0 ;
  assign n35003 = n32713 & n35002 ;
  assign n35004 = ~n10476 & n35003 ;
  assign n35005 = ( n9372 & n35000 ) | ( n9372 & ~n35004 ) | ( n35000 & ~n35004 ) ;
  assign n35006 = n12926 & ~n21622 ;
  assign n35007 = ( n2027 & ~n10796 ) | ( n2027 & n15845 ) | ( ~n10796 & n15845 ) ;
  assign n35008 = n10271 | n21021 ;
  assign n35009 = n35007 | n35008 ;
  assign n35010 = n15825 ^ n14305 ^ n12599 ;
  assign n35011 = n23786 ^ n18882 ^ 1'b0 ;
  assign n35012 = n35011 ^ n14063 ^ 1'b0 ;
  assign n35013 = ( n18899 & ~n21126 ) | ( n18899 & n29482 ) | ( ~n21126 & n29482 ) ;
  assign n35014 = n35013 ^ n15594 ^ n10657 ;
  assign n35015 = ~n883 & n23893 ;
  assign n35017 = ~n3261 & n6752 ;
  assign n35016 = ( n10247 & n21789 ) | ( n10247 & n29385 ) | ( n21789 & n29385 ) ;
  assign n35018 = n35017 ^ n35016 ^ n13460 ;
  assign n35019 = n15050 | n35018 ;
  assign n35020 = ( n10923 & ~n15768 ) | ( n10923 & n35019 ) | ( ~n15768 & n35019 ) ;
  assign n35021 = ( n1927 & ~n4012 ) | ( n1927 & n4603 ) | ( ~n4012 & n4603 ) ;
  assign n35022 = n23455 | n35021 ;
  assign n35023 = n6676 & ~n35022 ;
  assign n35024 = ( ~n8534 & n9808 ) | ( ~n8534 & n11882 ) | ( n9808 & n11882 ) ;
  assign n35025 = n35024 ^ n31707 ^ n10270 ;
  assign n35026 = ( n19271 & n35023 ) | ( n19271 & n35025 ) | ( n35023 & n35025 ) ;
  assign n35027 = n1549 & n9276 ;
  assign n35028 = n35027 ^ n5974 ^ 1'b0 ;
  assign n35029 = n29563 ^ n17150 ^ n17105 ;
  assign n35030 = n13803 & n35029 ;
  assign n35034 = n28688 ^ n18093 ^ n9656 ;
  assign n35031 = ( ~n2550 & n4044 ) | ( ~n2550 & n16069 ) | ( n4044 & n16069 ) ;
  assign n35032 = n35031 ^ n33695 ^ 1'b0 ;
  assign n35033 = n5552 & n35032 ;
  assign n35035 = n35034 ^ n35033 ^ n35024 ;
  assign n35036 = ( n1497 & n3012 ) | ( n1497 & n9460 ) | ( n3012 & n9460 ) ;
  assign n35037 = ( n8822 & n10896 ) | ( n8822 & n26950 ) | ( n10896 & n26950 ) ;
  assign n35038 = ( n17278 & ~n35036 ) | ( n17278 & n35037 ) | ( ~n35036 & n35037 ) ;
  assign n35042 = n28905 ^ n23641 ^ n7227 ;
  assign n35039 = n31723 ^ n10980 ^ n3024 ;
  assign n35040 = n19802 & ~n34786 ;
  assign n35041 = n35039 | n35040 ;
  assign n35043 = n35042 ^ n35041 ^ 1'b0 ;
  assign n35044 = n18764 ^ n9901 ^ n9460 ;
  assign n35045 = n10513 & n35044 ;
  assign n35046 = ~n9326 & n35045 ;
  assign n35047 = ~n12998 & n35046 ;
  assign n35048 = n13907 & ~n24013 ;
  assign n35049 = ~n13358 & n35048 ;
  assign n35050 = ~n18060 & n35049 ;
  assign n35051 = ( n7196 & n16500 ) | ( n7196 & n30714 ) | ( n16500 & n30714 ) ;
  assign n35053 = ( n2530 & ~n14995 ) | ( n2530 & n15483 ) | ( ~n14995 & n15483 ) ;
  assign n35054 = n4093 & ~n35053 ;
  assign n35055 = n35054 ^ n10267 ^ 1'b0 ;
  assign n35052 = n2648 & n9782 ;
  assign n35056 = n35055 ^ n35052 ^ n15352 ;
  assign n35057 = n5318 & ~n7571 ;
  assign n35058 = n35057 ^ n12401 ^ 1'b0 ;
  assign n35059 = n20095 ^ n18069 ^ n8030 ;
  assign n35060 = n22415 ^ n1241 ^ 1'b0 ;
  assign n35061 = ( ~x78 & n35059 ) | ( ~x78 & n35060 ) | ( n35059 & n35060 ) ;
  assign n35062 = ( n4092 & ~n4651 ) | ( n4092 & n10235 ) | ( ~n4651 & n10235 ) ;
  assign n35063 = n35062 ^ n19674 ^ n16604 ;
  assign n35064 = ( n11102 & n17918 ) | ( n11102 & ~n35063 ) | ( n17918 & ~n35063 ) ;
  assign n35065 = n35064 ^ n5187 ^ 1'b0 ;
  assign n35066 = n3371 & n35065 ;
  assign n35067 = ~n13431 & n25017 ;
  assign n35068 = n35067 ^ n29873 ^ 1'b0 ;
  assign n35069 = n28238 ^ n22869 ^ n1375 ;
  assign n35070 = n26688 | n35069 ;
  assign n35071 = n35070 ^ n32185 ^ 1'b0 ;
  assign n35072 = n35071 ^ n27976 ^ 1'b0 ;
  assign n35073 = n7594 & ~n35072 ;
  assign n35078 = ( n3524 & n8451 ) | ( n3524 & n20395 ) | ( n8451 & n20395 ) ;
  assign n35074 = n11011 | n19699 ;
  assign n35075 = n35074 ^ n3915 ^ 1'b0 ;
  assign n35076 = ~n30223 & n35075 ;
  assign n35077 = n18049 & n35076 ;
  assign n35079 = n35078 ^ n35077 ^ 1'b0 ;
  assign n35080 = n33611 ^ n13996 ^ n8881 ;
  assign n35081 = n9195 | n33097 ;
  assign n35082 = n10372 ^ n6153 ^ n802 ;
  assign n35083 = n35082 ^ n14189 ^ 1'b0 ;
  assign n35084 = n1232 & n35083 ;
  assign n35085 = n35084 ^ n17710 ^ n13100 ;
  assign n35086 = ~n6513 & n10821 ;
  assign n35087 = ~n28263 & n35086 ;
  assign n35088 = n2126 & n24683 ;
  assign n35089 = n2728 & n35088 ;
  assign n35090 = n18325 ^ n4998 ^ 1'b0 ;
  assign n35091 = n31045 | n35090 ;
  assign n35092 = ( n7366 & n7573 ) | ( n7366 & ~n16513 ) | ( n7573 & ~n16513 ) ;
  assign n35093 = n35092 ^ n21233 ^ 1'b0 ;
  assign n35094 = n33180 & n35093 ;
  assign n35095 = n15728 ^ n14332 ^ n5253 ;
  assign n35096 = ( ~n32127 & n35094 ) | ( ~n32127 & n35095 ) | ( n35094 & n35095 ) ;
  assign n35097 = ( n398 & ~n2401 ) | ( n398 & n6626 ) | ( ~n2401 & n6626 ) ;
  assign n35098 = n6662 ^ n5056 ^ n277 ;
  assign n35099 = n13546 ^ n11213 ^ 1'b0 ;
  assign n35100 = n18131 | n20412 ;
  assign n35101 = n35099 & ~n35100 ;
  assign n35102 = n4540 | n6851 ;
  assign n35103 = n22606 | n35102 ;
  assign n35104 = n10659 ^ n9383 ^ n4437 ;
  assign n35105 = n33089 ^ n25538 ^ n20071 ;
  assign n35106 = ~n19800 & n35105 ;
  assign n35107 = ~n35104 & n35106 ;
  assign n35108 = n14044 | n35107 ;
  assign n35109 = n16050 & n21550 ;
  assign n35110 = n35109 ^ n9822 ^ 1'b0 ;
  assign n35111 = ( ~n6054 & n6602 ) | ( ~n6054 & n22286 ) | ( n6602 & n22286 ) ;
  assign n35112 = ( n8714 & ~n31112 ) | ( n8714 & n35111 ) | ( ~n31112 & n35111 ) ;
  assign n35113 = ~n29719 & n35112 ;
  assign n35114 = n9217 | n21945 ;
  assign n35115 = n942 & ~n35114 ;
  assign n35116 = n4944 & n14209 ;
  assign n35117 = n18573 & n35116 ;
  assign n35118 = n8293 & ~n35117 ;
  assign n35119 = ~n8231 & n35118 ;
  assign n35120 = n35119 ^ n1694 ^ n1101 ;
  assign n35121 = ( ~n31626 & n35115 ) | ( ~n31626 & n35120 ) | ( n35115 & n35120 ) ;
  assign n35124 = n12232 & n14334 ;
  assign n35122 = n5842 ^ n2690 ^ n1247 ;
  assign n35123 = n35122 ^ n24321 ^ n13891 ;
  assign n35125 = n35124 ^ n35123 ^ n9629 ;
  assign n35126 = n11653 | n21109 ;
  assign n35127 = ( ~n6642 & n13726 ) | ( ~n6642 & n33467 ) | ( n13726 & n33467 ) ;
  assign n35128 = ( ~n18135 & n19920 ) | ( ~n18135 & n30788 ) | ( n19920 & n30788 ) ;
  assign n35129 = ( n16145 & ~n19115 ) | ( n16145 & n28406 ) | ( ~n19115 & n28406 ) ;
  assign n35130 = ( n4285 & n6697 ) | ( n4285 & ~n30713 ) | ( n6697 & ~n30713 ) ;
  assign n35131 = ( ~n27801 & n31503 ) | ( ~n27801 & n35130 ) | ( n31503 & n35130 ) ;
  assign n35132 = n35131 ^ n6053 ^ 1'b0 ;
  assign n35133 = n19699 & ~n35132 ;
  assign n35138 = n21951 ^ n19558 ^ n7322 ;
  assign n35139 = n35138 ^ n19123 ^ n9988 ;
  assign n35134 = n30557 ^ n7113 ^ n2583 ;
  assign n35135 = n11754 | n23783 ;
  assign n35136 = n13596 | n35135 ;
  assign n35137 = n35134 & n35136 ;
  assign n35140 = n35139 ^ n35137 ^ n7355 ;
  assign n35141 = ( n4541 & n5360 ) | ( n4541 & ~n17985 ) | ( n5360 & ~n17985 ) ;
  assign n35142 = ( x99 & ~n5619 ) | ( x99 & n35141 ) | ( ~n5619 & n35141 ) ;
  assign n35143 = n35142 ^ n29869 ^ n15410 ;
  assign n35144 = n21272 & ~n35143 ;
  assign n35145 = n9431 | n28009 ;
  assign n35146 = ( n6035 & ~n10948 ) | ( n6035 & n16390 ) | ( ~n10948 & n16390 ) ;
  assign n35150 = n10661 & ~n12422 ;
  assign n35151 = n35150 ^ n15891 ^ n3989 ;
  assign n35148 = n23506 ^ n16147 ^ n5736 ;
  assign n35147 = n16287 & ~n19539 ;
  assign n35149 = n35148 ^ n35147 ^ n23526 ;
  assign n35152 = n35151 ^ n35149 ^ n13584 ;
  assign n35153 = n19842 ^ n11696 ^ n382 ;
  assign n35154 = n22328 ^ n6575 ^ n4108 ;
  assign n35155 = n35154 ^ n23175 ^ n8349 ;
  assign n35156 = n12439 | n35155 ;
  assign n35157 = ~n35153 & n35156 ;
  assign n35158 = n27730 ^ n14702 ^ 1'b0 ;
  assign n35164 = n7532 & ~n28945 ;
  assign n35165 = n7344 & n35164 ;
  assign n35161 = n6979 | n14906 ;
  assign n35162 = n35161 ^ n11931 ^ 1'b0 ;
  assign n35159 = n31136 ^ n5693 ^ n570 ;
  assign n35160 = ( ~n19555 & n24781 ) | ( ~n19555 & n35159 ) | ( n24781 & n35159 ) ;
  assign n35163 = n35162 ^ n35160 ^ n19493 ;
  assign n35166 = n35165 ^ n35163 ^ n33063 ;
  assign n35167 = n11286 ^ n3377 ^ n1109 ;
  assign n35168 = n6271 | n19626 ;
  assign n35169 = ( n17457 & n35167 ) | ( n17457 & ~n35168 ) | ( n35167 & ~n35168 ) ;
  assign n35170 = n22672 ^ n11795 ^ 1'b0 ;
  assign n35171 = n14148 & ~n27685 ;
  assign n35172 = ~n35170 & n35171 ;
  assign n35173 = n11534 ^ n9684 ^ n7795 ;
  assign n35174 = n30287 ^ n9753 ^ 1'b0 ;
  assign n35175 = n28238 & n35174 ;
  assign n35176 = ( ~n3945 & n4645 ) | ( ~n3945 & n7013 ) | ( n4645 & n7013 ) ;
  assign n35177 = ~n16441 & n35176 ;
  assign n35178 = ( ~n1154 & n15583 ) | ( ~n1154 & n15895 ) | ( n15583 & n15895 ) ;
  assign n35179 = n35178 ^ n5635 ^ 1'b0 ;
  assign n35180 = n2809 ^ n2334 ^ 1'b0 ;
  assign n35181 = n30285 ^ n24903 ^ n6168 ;
  assign n35182 = ( n15140 & n32439 ) | ( n15140 & n35181 ) | ( n32439 & n35181 ) ;
  assign n35196 = n6930 & ~n18859 ;
  assign n35197 = n35196 ^ n19124 ^ n18489 ;
  assign n35190 = ~n1910 & n6697 ;
  assign n35191 = n10935 & n35190 ;
  assign n35192 = n35191 ^ n9926 ^ 1'b0 ;
  assign n35193 = ( n24343 & n27718 ) | ( n24343 & ~n35192 ) | ( n27718 & ~n35192 ) ;
  assign n35194 = n8379 & ~n35193 ;
  assign n35183 = n16862 ^ n1290 ^ 1'b0 ;
  assign n35186 = n13065 | n32222 ;
  assign n35187 = n35186 ^ n13219 ^ 1'b0 ;
  assign n35184 = n8486 ^ n5416 ^ n892 ;
  assign n35185 = n35184 ^ n20288 ^ 1'b0 ;
  assign n35188 = n35187 ^ n35185 ^ n14160 ;
  assign n35189 = n35183 | n35188 ;
  assign n35195 = n35194 ^ n35189 ^ 1'b0 ;
  assign n35198 = n35197 ^ n35195 ^ n7035 ;
  assign n35199 = ( n2098 & n9103 ) | ( n2098 & n10920 ) | ( n9103 & n10920 ) ;
  assign n35200 = n35199 ^ n13084 ^ n3365 ;
  assign n35201 = n35200 ^ n7722 ^ 1'b0 ;
  assign n35202 = n13443 | n35201 ;
  assign n35203 = n23486 ^ n430 ^ 1'b0 ;
  assign n35204 = n339 & n35203 ;
  assign n35205 = ( ~n2989 & n31557 ) | ( ~n2989 & n35204 ) | ( n31557 & n35204 ) ;
  assign n35206 = n31421 ^ n27599 ^ n11388 ;
  assign n35207 = n35205 & ~n35206 ;
  assign n35208 = n35207 ^ n6700 ^ 1'b0 ;
  assign n35209 = n35208 ^ n12319 ^ 1'b0 ;
  assign n35210 = ( ~n6212 & n27159 ) | ( ~n6212 & n27205 ) | ( n27159 & n27205 ) ;
  assign n35211 = ( n3530 & n4606 ) | ( n3530 & ~n21343 ) | ( n4606 & ~n21343 ) ;
  assign n35212 = n31127 ^ n24585 ^ n6036 ;
  assign n35213 = n35212 ^ n31980 ^ n10201 ;
  assign n35214 = ~n656 & n2659 ;
  assign n35215 = ~n5224 & n35214 ;
  assign n35216 = n35215 ^ n30049 ^ x112 ;
  assign n35217 = n35216 ^ n19106 ^ 1'b0 ;
  assign n35218 = n25227 & n35217 ;
  assign n35219 = ~n15927 & n17045 ;
  assign n35220 = ~n4652 & n35219 ;
  assign n35221 = ( n1006 & n3682 ) | ( n1006 & ~n27352 ) | ( n3682 & ~n27352 ) ;
  assign n35222 = n35221 ^ n20972 ^ x133 ;
  assign n35224 = n3690 ^ n389 ^ 1'b0 ;
  assign n35225 = n11520 | n35224 ;
  assign n35223 = ( n4605 & n15850 ) | ( n4605 & ~n24067 ) | ( n15850 & ~n24067 ) ;
  assign n35226 = n35225 ^ n35223 ^ n17171 ;
  assign n35227 = ( ~n6786 & n27708 ) | ( ~n6786 & n32011 ) | ( n27708 & n32011 ) ;
  assign n35228 = ( n6690 & ~n15504 ) | ( n6690 & n35227 ) | ( ~n15504 & n35227 ) ;
  assign n35229 = n35228 ^ n10032 ^ 1'b0 ;
  assign n35233 = ( n4950 & n6105 ) | ( n4950 & n8062 ) | ( n6105 & n8062 ) ;
  assign n35232 = n23464 ^ n11757 ^ n6523 ;
  assign n35234 = n35233 ^ n35232 ^ n23234 ;
  assign n35230 = n13550 | n27256 ;
  assign n35231 = n35230 ^ n14452 ^ 1'b0 ;
  assign n35235 = n35234 ^ n35231 ^ 1'b0 ;
  assign n35236 = n9298 | n10154 ;
  assign n35237 = n6977 | n35236 ;
  assign n35238 = ~n18938 & n19200 ;
  assign n35239 = ~n35237 & n35238 ;
  assign n35240 = n7829 & n33245 ;
  assign n35241 = ~n24123 & n35240 ;
  assign n35242 = n31869 ^ n27603 ^ 1'b0 ;
  assign n35243 = n21105 ^ n19548 ^ 1'b0 ;
  assign n35244 = n25985 ^ n24178 ^ n13304 ;
  assign n35245 = ( n7805 & n11439 ) | ( n7805 & n35244 ) | ( n11439 & n35244 ) ;
  assign n35255 = ( n6092 & ~n8282 ) | ( n6092 & n19148 ) | ( ~n8282 & n19148 ) ;
  assign n35246 = ~n2022 & n33145 ;
  assign n35247 = n35246 ^ n12000 ^ 1'b0 ;
  assign n35248 = n35247 ^ n21586 ^ 1'b0 ;
  assign n35249 = n16016 & n35248 ;
  assign n35250 = ~n1365 & n9034 ;
  assign n35251 = ~n25785 & n35250 ;
  assign n35252 = ~n35249 & n35251 ;
  assign n35253 = n11461 & ~n35252 ;
  assign n35254 = ~n19908 & n35253 ;
  assign n35256 = n35255 ^ n35254 ^ n6104 ;
  assign n35257 = n16293 ^ n13342 ^ n10858 ;
  assign n35258 = n35257 ^ n19078 ^ n7504 ;
  assign n35259 = n8342 & ~n23601 ;
  assign n35260 = n14783 & n35259 ;
  assign n35261 = n3706 | n28031 ;
  assign n35262 = n35261 ^ n32633 ^ 1'b0 ;
  assign n35263 = n23353 ^ n10187 ^ n6582 ;
  assign n35264 = n5789 | n35263 ;
  assign n35265 = n25209 & ~n35264 ;
  assign n35266 = n7424 ^ n5827 ^ n781 ;
  assign n35268 = n7913 ^ n3356 ^ 1'b0 ;
  assign n35269 = n15836 & ~n35268 ;
  assign n35267 = n8165 & ~n13436 ;
  assign n35270 = n35269 ^ n35267 ^ 1'b0 ;
  assign n35271 = ( n5642 & ~n26820 ) | ( n5642 & n35270 ) | ( ~n26820 & n35270 ) ;
  assign n35273 = n26587 ^ n22676 ^ x183 ;
  assign n35272 = ~n15383 & n24150 ;
  assign n35274 = n35273 ^ n35272 ^ n25408 ;
  assign n35275 = n29151 ^ n26903 ^ n7306 ;
  assign n35276 = n19158 ^ n4657 ^ 1'b0 ;
  assign n35277 = ( ~n3921 & n14911 ) | ( ~n3921 & n23420 ) | ( n14911 & n23420 ) ;
  assign n35278 = n1149 | n35277 ;
  assign n35279 = n35278 ^ n20239 ^ 1'b0 ;
  assign n35292 = n6845 & n8286 ;
  assign n35293 = ( ~n7613 & n23340 ) | ( ~n7613 & n35292 ) | ( n23340 & n35292 ) ;
  assign n35287 = ~n2085 & n5972 ;
  assign n35288 = n35287 ^ n3006 ^ 1'b0 ;
  assign n35289 = n35288 ^ n27996 ^ n23333 ;
  assign n35290 = n24139 & n35289 ;
  assign n35291 = n35290 ^ n24488 ^ 1'b0 ;
  assign n35294 = n35293 ^ n35291 ^ n9191 ;
  assign n35295 = n35294 ^ n5008 ^ 1'b0 ;
  assign n35296 = ( n606 & n20341 ) | ( n606 & n25579 ) | ( n20341 & n25579 ) ;
  assign n35297 = ( n4322 & n33388 ) | ( n4322 & ~n35296 ) | ( n33388 & ~n35296 ) ;
  assign n35298 = n35295 & n35297 ;
  assign n35280 = n17553 ^ n7566 ^ n361 ;
  assign n35281 = n26878 ^ n19354 ^ n4570 ;
  assign n35282 = n35281 ^ n9531 ^ 1'b0 ;
  assign n35283 = n7664 & n35282 ;
  assign n35284 = n26219 & n35283 ;
  assign n35285 = n35284 ^ n22856 ^ 1'b0 ;
  assign n35286 = n35280 | n35285 ;
  assign n35299 = n35298 ^ n35286 ^ 1'b0 ;
  assign n35301 = ( n1711 & n10370 ) | ( n1711 & n15232 ) | ( n10370 & n15232 ) ;
  assign n35300 = n14206 ^ n8384 ^ n2892 ;
  assign n35302 = n35301 ^ n35300 ^ n12102 ;
  assign n35303 = n19695 ^ n15455 ^ n5918 ;
  assign n35304 = n35303 ^ n32636 ^ n23413 ;
  assign n35305 = ( ~x34 & n34236 ) | ( ~x34 & n35304 ) | ( n34236 & n35304 ) ;
  assign n35306 = n35305 ^ n33353 ^ n13608 ;
  assign n35309 = n22690 ^ n6439 ^ 1'b0 ;
  assign n35310 = ( n21321 & n31388 ) | ( n21321 & ~n35309 ) | ( n31388 & ~n35309 ) ;
  assign n35307 = n21748 ^ n19570 ^ n4781 ;
  assign n35308 = ( n11919 & n19633 ) | ( n11919 & ~n35307 ) | ( n19633 & ~n35307 ) ;
  assign n35311 = n35310 ^ n35308 ^ n602 ;
  assign n35312 = n22606 ^ n9711 ^ 1'b0 ;
  assign n35313 = n1455 & ~n35312 ;
  assign n35314 = n5973 & ~n35313 ;
  assign n35315 = x18 & ~n11428 ;
  assign n35316 = n35315 ^ n14769 ^ 1'b0 ;
  assign n35317 = n35316 ^ n14002 ^ n9692 ;
  assign n35318 = n24125 | n35317 ;
  assign n35319 = ( n2031 & n2598 ) | ( n2031 & ~n6927 ) | ( n2598 & ~n6927 ) ;
  assign n35320 = ~n20940 & n35319 ;
  assign n35321 = n35320 ^ n14546 ^ 1'b0 ;
  assign n35322 = ( n6518 & n14310 ) | ( n6518 & n35321 ) | ( n14310 & n35321 ) ;
  assign n35323 = n6759 & ~n9258 ;
  assign n35325 = n4352 ^ n2382 ^ 1'b0 ;
  assign n35324 = ( n1164 & ~n27083 ) | ( n1164 & n27457 ) | ( ~n27083 & n27457 ) ;
  assign n35326 = n35325 ^ n35324 ^ x23 ;
  assign n35327 = n6473 ^ n3899 ^ 1'b0 ;
  assign n35328 = n17918 ^ n2402 ^ 1'b0 ;
  assign n35329 = ( n24084 & ~n28558 ) | ( n24084 & n35328 ) | ( ~n28558 & n35328 ) ;
  assign n35330 = n33458 ^ n28793 ^ 1'b0 ;
  assign n35331 = n35330 ^ n14652 ^ 1'b0 ;
  assign n35332 = n35329 | n35331 ;
  assign n35333 = ( n7503 & n7512 ) | ( n7503 & n8861 ) | ( n7512 & n8861 ) ;
  assign n35334 = ( n2299 & n19599 ) | ( n2299 & ~n35333 ) | ( n19599 & ~n35333 ) ;
  assign n35335 = ( ~n8482 & n22213 ) | ( ~n8482 & n35334 ) | ( n22213 & n35334 ) ;
  assign n35336 = ( n1413 & ~n14800 ) | ( n1413 & n20244 ) | ( ~n14800 & n20244 ) ;
  assign n35338 = n11182 ^ n11088 ^ n6500 ;
  assign n35337 = n7491 | n10466 ;
  assign n35339 = n35338 ^ n35337 ^ 1'b0 ;
  assign n35343 = n18171 ^ n13875 ^ n9602 ;
  assign n35340 = n29705 ^ n16480 ^ n15828 ;
  assign n35341 = n34412 & n35340 ;
  assign n35342 = n19767 & n35341 ;
  assign n35344 = n35343 ^ n35342 ^ 1'b0 ;
  assign n35345 = ( n790 & ~n13275 ) | ( n790 & n33124 ) | ( ~n13275 & n33124 ) ;
  assign n35346 = n29935 ^ n25171 ^ n899 ;
  assign n35347 = n35346 ^ n34672 ^ n9007 ;
  assign n35348 = n5579 & ~n35347 ;
  assign n35349 = n3554 & n35348 ;
  assign n35350 = ( x134 & ~n10492 ) | ( x134 & n28065 ) | ( ~n10492 & n28065 ) ;
  assign n35351 = n35350 ^ n10395 ^ n9441 ;
  assign n35352 = ( ~n19395 & n21620 ) | ( ~n19395 & n32510 ) | ( n21620 & n32510 ) ;
  assign n35353 = ( ~n8870 & n24808 ) | ( ~n8870 & n27588 ) | ( n24808 & n27588 ) ;
  assign n35354 = n35353 ^ n28854 ^ n25752 ;
  assign n35355 = n14967 | n30234 ;
  assign n35356 = n35355 ^ n30403 ^ 1'b0 ;
  assign n35357 = n35356 ^ n18167 ^ n15421 ;
  assign n35358 = n31098 ^ n21565 ^ 1'b0 ;
  assign n35359 = n35357 & ~n35358 ;
  assign n35361 = ( ~n8187 & n11006 ) | ( ~n8187 & n13992 ) | ( n11006 & n13992 ) ;
  assign n35360 = n14840 & n21246 ;
  assign n35362 = n35361 ^ n35360 ^ 1'b0 ;
  assign n35363 = ~n12140 & n35362 ;
  assign n35364 = n11764 & n35363 ;
  assign n35365 = ~n11883 & n35364 ;
  assign n35366 = n1165 & ~n1713 ;
  assign n35367 = n271 & ~n14510 ;
  assign n35368 = n35367 ^ n17790 ^ 1'b0 ;
  assign n35369 = n35368 ^ n23099 ^ 1'b0 ;
  assign n35370 = n16749 | n35369 ;
  assign n35371 = n35370 ^ n21402 ^ 1'b0 ;
  assign n35372 = ~n20041 & n35371 ;
  assign n35373 = n35372 ^ n23967 ^ n7452 ;
  assign n35374 = n35373 ^ n20441 ^ n6184 ;
  assign n35375 = n29803 ^ n21058 ^ n1315 ;
  assign n35376 = ~n23824 & n31477 ;
  assign n35378 = n6356 ^ n4520 ^ n1085 ;
  assign n35377 = n32128 ^ n12108 ^ 1'b0 ;
  assign n35379 = n35378 ^ n35377 ^ n13909 ;
  assign n35380 = n35379 ^ n24892 ^ 1'b0 ;
  assign n35381 = ( ~x159 & n321 ) | ( ~x159 & n16097 ) | ( n321 & n16097 ) ;
  assign n35382 = n35381 ^ n30967 ^ 1'b0 ;
  assign n35383 = ( n7043 & n17394 ) | ( n7043 & n18078 ) | ( n17394 & n18078 ) ;
  assign n35384 = ~n33226 & n35383 ;
  assign n35385 = n35382 & n35384 ;
  assign n35386 = x186 & ~n29315 ;
  assign n35387 = n35386 ^ n1976 ^ 1'b0 ;
  assign n35388 = ~n16454 & n19917 ;
  assign n35389 = n30032 & n35388 ;
  assign n35390 = n35389 ^ n26669 ^ 1'b0 ;
  assign n35391 = n13677 | n35390 ;
  assign n35392 = n21620 ^ n11475 ^ n3322 ;
  assign n35393 = n25114 ^ n20312 ^ n9908 ;
  assign n35394 = ~n19131 & n35393 ;
  assign n35395 = n33597 ^ n7197 ^ n3748 ;
  assign n35396 = n35395 ^ n1433 ^ 1'b0 ;
  assign n35397 = n17392 & n21619 ;
  assign n35398 = n35397 ^ n6946 ^ 1'b0 ;
  assign n35399 = ( n5593 & ~n20998 ) | ( n5593 & n35398 ) | ( ~n20998 & n35398 ) ;
  assign n35400 = ~n35396 & n35399 ;
  assign n35401 = n35400 ^ n19219 ^ 1'b0 ;
  assign n35402 = n3794 & ~n4896 ;
  assign n35403 = ( ~n21426 & n34332 ) | ( ~n21426 & n35402 ) | ( n34332 & n35402 ) ;
  assign n35404 = x236 & ~n4717 ;
  assign n35405 = ~n35403 & n35404 ;
  assign n35406 = n28856 ^ n16214 ^ 1'b0 ;
  assign n35407 = n29105 ^ n3920 ^ n471 ;
  assign n35408 = n12239 | n33859 ;
  assign n35409 = n26184 ^ n22209 ^ n4072 ;
  assign n35411 = ( n12163 & ~n22682 ) | ( n12163 & n31769 ) | ( ~n22682 & n31769 ) ;
  assign n35410 = n35356 ^ n29628 ^ n1886 ;
  assign n35412 = n35411 ^ n35410 ^ 1'b0 ;
  assign n35413 = ~n17687 & n35096 ;
  assign n35414 = n35412 & n35413 ;
  assign n35415 = n19863 ^ n9148 ^ n967 ;
  assign n35416 = n1459 & ~n35415 ;
  assign n35417 = n28512 ^ n23829 ^ 1'b0 ;
  assign n35418 = n35416 | n35417 ;
  assign n35419 = n12828 & ~n21683 ;
  assign n35420 = ~n14267 & n35419 ;
  assign n35421 = n15177 ^ n15171 ^ n5037 ;
  assign n35422 = n35421 ^ n18751 ^ n14887 ;
  assign n35423 = n35422 ^ n32861 ^ n3562 ;
  assign n35424 = n35415 ^ n13742 ^ n4967 ;
  assign n35425 = n33156 & n35424 ;
  assign n35426 = ( n694 & ~n25194 ) | ( n694 & n35425 ) | ( ~n25194 & n35425 ) ;
  assign n35427 = n13172 & ~n30660 ;
  assign n35428 = n5466 | n20145 ;
  assign n35429 = ( n15795 & n33650 ) | ( n15795 & n35428 ) | ( n33650 & n35428 ) ;
  assign n35430 = n15071 ^ n3938 ^ n2625 ;
  assign n35431 = ( n8922 & n29942 ) | ( n8922 & n35430 ) | ( n29942 & n35430 ) ;
  assign n35432 = n830 & ~n3601 ;
  assign n35433 = n35432 ^ n847 ^ 1'b0 ;
  assign n35434 = n35433 ^ n31742 ^ n15684 ;
  assign n35435 = n17218 & n35434 ;
  assign n35436 = ~n16779 & n35435 ;
  assign n35437 = n35436 ^ n13455 ^ 1'b0 ;
  assign n35438 = ~n13925 & n29941 ;
  assign n35439 = n20947 & n35438 ;
  assign n35440 = n14364 & n16881 ;
  assign n35441 = n35440 ^ n1594 ^ 1'b0 ;
  assign n35442 = n35441 ^ n13935 ^ 1'b0 ;
  assign n35443 = n12563 ^ n6889 ^ n4782 ;
  assign n35444 = n35443 ^ n25823 ^ n8917 ;
  assign n35445 = n7881 | n17941 ;
  assign n35446 = n35445 ^ n5636 ^ 1'b0 ;
  assign n35447 = ~n14007 & n20826 ;
  assign n35448 = n14313 & n35447 ;
  assign n35449 = n3536 & ~n35448 ;
  assign n35450 = ~n14492 & n35449 ;
  assign n35451 = ( n7878 & n10992 ) | ( n7878 & ~n23846 ) | ( n10992 & ~n23846 ) ;
  assign n35452 = n2961 & n10169 ;
  assign n35453 = n35452 ^ n13083 ^ 1'b0 ;
  assign n35454 = n35453 ^ n34872 ^ n9318 ;
  assign n35455 = ( n15293 & n28714 ) | ( n15293 & ~n35454 ) | ( n28714 & ~n35454 ) ;
  assign n35456 = n30884 ^ n8157 ^ 1'b0 ;
  assign n35457 = n22928 ^ n2930 ^ n1897 ;
  assign n35458 = n35457 ^ n3113 ^ x83 ;
  assign n35459 = n17418 & n18030 ;
  assign n35460 = n35459 ^ n9718 ^ 1'b0 ;
  assign n35461 = n23316 & ~n35460 ;
  assign n35462 = n35461 ^ n20437 ^ 1'b0 ;
  assign n35463 = ( n5398 & ~n14215 ) | ( n5398 & n21707 ) | ( ~n14215 & n21707 ) ;
  assign n35464 = n11478 ^ n4877 ^ n4642 ;
  assign n35465 = ( ~n21931 & n35463 ) | ( ~n21931 & n35464 ) | ( n35463 & n35464 ) ;
  assign n35466 = n5151 & n5705 ;
  assign n35467 = n2350 & ~n35466 ;
  assign n35468 = n26146 & ~n32581 ;
  assign n35469 = n35468 ^ n18732 ^ 1'b0 ;
  assign n35470 = n35469 ^ n15604 ^ n13349 ;
  assign n35472 = n32685 ^ n21917 ^ 1'b0 ;
  assign n35471 = ( ~x109 & n8303 ) | ( ~x109 & n33682 ) | ( n8303 & n33682 ) ;
  assign n35473 = n35472 ^ n35471 ^ n310 ;
  assign n35474 = n28141 ^ n6716 ^ n3693 ;
  assign n35475 = ( n13047 & n15143 ) | ( n13047 & n27503 ) | ( n15143 & n27503 ) ;
  assign n35476 = n35475 ^ n29302 ^ n13880 ;
  assign n35481 = n25311 ^ n13792 ^ 1'b0 ;
  assign n35478 = n7608 & n27350 ;
  assign n35479 = ~n8308 & n35478 ;
  assign n35477 = ( ~n15446 & n19965 ) | ( ~n15446 & n29882 ) | ( n19965 & n29882 ) ;
  assign n35480 = n35479 ^ n35477 ^ 1'b0 ;
  assign n35482 = n35481 ^ n35480 ^ 1'b0 ;
  assign n35485 = n24725 ^ n8562 ^ n813 ;
  assign n35483 = n28929 ^ n19607 ^ n16607 ;
  assign n35484 = n3232 & ~n35483 ;
  assign n35486 = n35485 ^ n35484 ^ 1'b0 ;
  assign n35487 = n16866 | n24542 ;
  assign n35488 = n35487 ^ n4066 ^ 1'b0 ;
  assign n35489 = n35488 ^ n1820 ^ 1'b0 ;
  assign n35490 = ~n15438 & n35489 ;
  assign n35491 = n31549 ^ n30554 ^ 1'b0 ;
  assign n35492 = ( ~n4411 & n13732 ) | ( ~n4411 & n25943 ) | ( n13732 & n25943 ) ;
  assign n35493 = n35492 ^ n20190 ^ 1'b0 ;
  assign n35494 = n21357 ^ n12533 ^ x6 ;
  assign n35495 = n35494 ^ n27304 ^ n6037 ;
  assign n35496 = n18226 ^ n4293 ^ n3949 ;
  assign n35497 = n12291 ^ n7855 ^ 1'b0 ;
  assign n35498 = x121 & n35497 ;
  assign n35499 = n22271 & n35498 ;
  assign n35500 = ( n8338 & ~n33571 ) | ( n8338 & n35499 ) | ( ~n33571 & n35499 ) ;
  assign n35501 = ( ~n1942 & n4230 ) | ( ~n1942 & n15858 ) | ( n4230 & n15858 ) ;
  assign n35502 = n35501 ^ n32036 ^ 1'b0 ;
  assign n35503 = n7275 & ~n35502 ;
  assign n35504 = n23164 & n35503 ;
  assign n35505 = n8316 & ~n35504 ;
  assign n35506 = n23802 ^ n12715 ^ 1'b0 ;
  assign n35507 = n10415 & n35506 ;
  assign n35508 = ~n18204 & n21007 ;
  assign n35509 = n15089 ^ n11039 ^ n8166 ;
  assign n35510 = ( ~n12559 & n15456 ) | ( ~n12559 & n17288 ) | ( n15456 & n17288 ) ;
  assign n35511 = ( ~n13859 & n28448 ) | ( ~n13859 & n35510 ) | ( n28448 & n35510 ) ;
  assign n35512 = n35511 ^ n3217 ^ n897 ;
  assign n35513 = ( n30006 & n35509 ) | ( n30006 & n35512 ) | ( n35509 & n35512 ) ;
  assign n35514 = n5602 & n9992 ;
  assign n35515 = n3722 & n35514 ;
  assign n35516 = n35515 ^ n20834 ^ 1'b0 ;
  assign n35517 = n25897 ^ n18331 ^ 1'b0 ;
  assign n35519 = n20124 ^ n17903 ^ 1'b0 ;
  assign n35520 = n8731 | n35519 ;
  assign n35518 = n26501 ^ n17056 ^ n257 ;
  assign n35521 = n35520 ^ n35518 ^ 1'b0 ;
  assign n35522 = n29668 & ~n35521 ;
  assign n35523 = n35522 ^ n5687 ^ 1'b0 ;
  assign n35524 = n33191 ^ n17256 ^ 1'b0 ;
  assign n35525 = n10708 | n33141 ;
  assign n35526 = n35524 | n35525 ;
  assign n35527 = n20152 ^ n13238 ^ 1'b0 ;
  assign n35528 = ( n3654 & n26514 ) | ( n3654 & n35527 ) | ( n26514 & n35527 ) ;
  assign n35529 = n31002 ^ n19998 ^ n12255 ;
  assign n35534 = n9634 ^ n2763 ^ 1'b0 ;
  assign n35532 = n3096 & n12561 ;
  assign n35533 = n35532 ^ n16533 ^ x220 ;
  assign n35530 = ( n9946 & n13166 ) | ( n9946 & ~n20244 ) | ( n13166 & ~n20244 ) ;
  assign n35531 = n30131 | n35530 ;
  assign n35535 = n35534 ^ n35533 ^ n35531 ;
  assign n35536 = n26184 | n33616 ;
  assign n35537 = ( n5285 & n6767 ) | ( n5285 & ~n12010 ) | ( n6767 & ~n12010 ) ;
  assign n35538 = ( n4426 & n14175 ) | ( n4426 & n35537 ) | ( n14175 & n35537 ) ;
  assign n35539 = ( n4396 & ~n9326 ) | ( n4396 & n14632 ) | ( ~n9326 & n14632 ) ;
  assign n35540 = ( ~n9279 & n18050 ) | ( ~n9279 & n35539 ) | ( n18050 & n35539 ) ;
  assign n35541 = n552 & n29175 ;
  assign n35543 = ~n325 & n27120 ;
  assign n35544 = n11487 & n35543 ;
  assign n35542 = n3305 & n4635 ;
  assign n35545 = n35544 ^ n35542 ^ 1'b0 ;
  assign n35546 = ( n11803 & n21954 ) | ( n11803 & n35545 ) | ( n21954 & n35545 ) ;
  assign n35547 = n9235 & n33337 ;
  assign n35548 = n35547 ^ n31621 ^ 1'b0 ;
  assign n35549 = ~n3733 & n21884 ;
  assign n35550 = n35549 ^ n20469 ^ 1'b0 ;
  assign n35551 = n33917 & n35550 ;
  assign n35552 = n22125 ^ n10065 ^ 1'b0 ;
  assign n35553 = ~n14215 & n35552 ;
  assign n35556 = n20272 ^ n5513 ^ n3784 ;
  assign n35554 = n943 ^ n890 ^ 1'b0 ;
  assign n35555 = ~n21523 & n35554 ;
  assign n35557 = n35556 ^ n35555 ^ n26987 ;
  assign n35558 = n35557 ^ n26711 ^ n23698 ;
  assign n35559 = n31365 ^ n18159 ^ 1'b0 ;
  assign n35561 = n8364 & ~n9267 ;
  assign n35560 = n9444 ^ n1473 ^ 1'b0 ;
  assign n35562 = n35561 ^ n35560 ^ n8140 ;
  assign n35563 = n2622 | n16010 ;
  assign n35564 = n16749 | n35563 ;
  assign n35565 = n13370 | n35564 ;
  assign n35566 = n35565 ^ n35451 ^ 1'b0 ;
  assign n35567 = n35562 | n35566 ;
  assign n35568 = n5878 & n10146 ;
  assign n35569 = n35568 ^ n3789 ^ 1'b0 ;
  assign n35570 = n31832 ^ n27567 ^ n947 ;
  assign n35571 = n35570 ^ n21185 ^ n5484 ;
  assign n35572 = n19778 ^ n1598 ^ 1'b0 ;
  assign n35573 = n6130 & ~n35572 ;
  assign n35574 = n35573 ^ n9372 ^ x170 ;
  assign n35575 = ( ~n1207 & n5648 ) | ( ~n1207 & n7681 ) | ( n5648 & n7681 ) ;
  assign n35576 = n35575 ^ n18225 ^ n13236 ;
  assign n35577 = n10187 ^ n9269 ^ n5842 ;
  assign n35578 = ( n1433 & n24565 ) | ( n1433 & n35577 ) | ( n24565 & n35577 ) ;
  assign n35579 = n22336 ^ n18013 ^ n1753 ;
  assign n35580 = ( n5107 & n25514 ) | ( n5107 & ~n27376 ) | ( n25514 & ~n27376 ) ;
  assign n35581 = ( n28373 & n35579 ) | ( n28373 & ~n35580 ) | ( n35579 & ~n35580 ) ;
  assign n35582 = ( ~x215 & n3546 ) | ( ~x215 & n13518 ) | ( n3546 & n13518 ) ;
  assign n35583 = n35582 ^ n26697 ^ 1'b0 ;
  assign n35585 = n9843 ^ n2729 ^ 1'b0 ;
  assign n35586 = n2208 | n35585 ;
  assign n35587 = n35586 ^ n16614 ^ 1'b0 ;
  assign n35588 = n18195 & ~n35587 ;
  assign n35584 = n20636 ^ n12874 ^ n12581 ;
  assign n35589 = n35588 ^ n35584 ^ 1'b0 ;
  assign n35590 = n2676 ^ n1448 ^ 1'b0 ;
  assign n35591 = n35590 ^ n35298 ^ n7881 ;
  assign n35592 = n9948 & ~n12260 ;
  assign n35593 = n28503 ^ n14719 ^ 1'b0 ;
  assign n35594 = ( n15035 & n16933 ) | ( n15035 & ~n35593 ) | ( n16933 & ~n35593 ) ;
  assign n35595 = n20620 ^ n10415 ^ n5087 ;
  assign n35596 = n35595 ^ n12191 ^ 1'b0 ;
  assign n35597 = ( x49 & n10124 ) | ( x49 & ~n27261 ) | ( n10124 & ~n27261 ) ;
  assign n35598 = n7940 ^ n4792 ^ n3130 ;
  assign n35599 = n35598 ^ n13524 ^ n4256 ;
  assign n35600 = n8230 & n35599 ;
  assign n35601 = ~n10589 & n35600 ;
  assign n35602 = n30917 ^ n2076 ^ 1'b0 ;
  assign n35603 = n4788 & n35602 ;
  assign n35604 = n8648 & ~n16732 ;
  assign n35605 = ( n6316 & n35603 ) | ( n6316 & n35604 ) | ( n35603 & n35604 ) ;
  assign n35606 = n5649 & ~n7653 ;
  assign n35607 = ~n35605 & n35606 ;
  assign n35608 = n16809 ^ n15701 ^ n1858 ;
  assign n35609 = ( ~n5813 & n10574 ) | ( ~n5813 & n16823 ) | ( n10574 & n16823 ) ;
  assign n35610 = ( n6864 & n29826 ) | ( n6864 & n31697 ) | ( n29826 & n31697 ) ;
  assign n35611 = n35610 ^ n6042 ^ 1'b0 ;
  assign n35612 = ( n7171 & n15311 ) | ( n7171 & ~n35611 ) | ( n15311 & ~n35611 ) ;
  assign n35613 = ~n9105 & n33235 ;
  assign n35614 = ( ~n7529 & n15786 ) | ( ~n7529 & n24864 ) | ( n15786 & n24864 ) ;
  assign n35615 = ( n24888 & n25599 ) | ( n24888 & n35614 ) | ( n25599 & n35614 ) ;
  assign n35617 = n28221 ^ n6014 ^ n1453 ;
  assign n35616 = n11936 ^ n3542 ^ 1'b0 ;
  assign n35618 = n35617 ^ n35616 ^ 1'b0 ;
  assign n35619 = ~n35615 & n35618 ;
  assign n35620 = ( n2047 & ~n4013 ) | ( n2047 & n11361 ) | ( ~n4013 & n11361 ) ;
  assign n35621 = n35620 ^ n16004 ^ 1'b0 ;
  assign n35622 = n8504 | n35621 ;
  assign n35623 = n23898 ^ n16257 ^ n12322 ;
  assign n35625 = n7886 | n13162 ;
  assign n35626 = n14772 & ~n35625 ;
  assign n35624 = ~n9898 & n24516 ;
  assign n35627 = n35626 ^ n35624 ^ n34271 ;
  assign n35628 = ( ~n9812 & n27054 ) | ( ~n9812 & n35627 ) | ( n27054 & n35627 ) ;
  assign n35629 = n1183 ^ x154 ^ 1'b0 ;
  assign n35630 = ( n2777 & n7303 ) | ( n2777 & ~n13531 ) | ( n7303 & ~n13531 ) ;
  assign n35631 = n15393 ^ n6788 ^ 1'b0 ;
  assign n35632 = ~n35630 & n35631 ;
  assign n35633 = n21185 ^ n12620 ^ n2454 ;
  assign n35634 = n35633 ^ n8066 ^ 1'b0 ;
  assign n35635 = ~n6698 & n35634 ;
  assign n35636 = n13072 & n21678 ;
  assign n35637 = n35636 ^ n13554 ^ n8352 ;
  assign n35638 = ( n3502 & ~n6771 ) | ( n3502 & n26168 ) | ( ~n6771 & n26168 ) ;
  assign n35639 = n35638 ^ n21839 ^ n3328 ;
  assign n35640 = n35639 ^ n22373 ^ n19163 ;
  assign n35641 = ( n7149 & ~n17812 ) | ( n7149 & n26999 ) | ( ~n17812 & n26999 ) ;
  assign n35642 = ~n30611 & n35641 ;
  assign n35643 = n15765 ^ n14105 ^ 1'b0 ;
  assign n35646 = n3697 | n11910 ;
  assign n35647 = n35646 ^ n18322 ^ n4697 ;
  assign n35648 = n9130 | n35647 ;
  assign n35649 = n33728 ^ n31428 ^ 1'b0 ;
  assign n35650 = ( n16515 & n25457 ) | ( n16515 & ~n35649 ) | ( n25457 & ~n35649 ) ;
  assign n35651 = ( ~n5021 & n35648 ) | ( ~n5021 & n35650 ) | ( n35648 & n35650 ) ;
  assign n35652 = n2414 & ~n35651 ;
  assign n35644 = n19167 ^ n13759 ^ n1818 ;
  assign n35645 = ( n1873 & ~n10089 ) | ( n1873 & n35644 ) | ( ~n10089 & n35644 ) ;
  assign n35653 = n35652 ^ n35645 ^ n7290 ;
  assign n35654 = ( n25142 & ~n35643 ) | ( n25142 & n35653 ) | ( ~n35643 & n35653 ) ;
  assign n35655 = n22635 ^ n17022 ^ 1'b0 ;
  assign n35656 = n19604 & n35655 ;
  assign n35657 = n23493 ^ n19269 ^ 1'b0 ;
  assign n35658 = n35657 ^ n3306 ^ n2528 ;
  assign n35659 = n21512 ^ n3200 ^ 1'b0 ;
  assign n35660 = n35659 ^ n6323 ^ n5886 ;
  assign n35661 = n26473 ^ n23998 ^ n19550 ;
  assign n35662 = ( n10504 & n21788 ) | ( n10504 & n35661 ) | ( n21788 & n35661 ) ;
  assign n35663 = ( n1591 & ~n1636 ) | ( n1591 & n33459 ) | ( ~n1636 & n33459 ) ;
  assign n35664 = ( n740 & ~n3078 ) | ( n740 & n19590 ) | ( ~n3078 & n19590 ) ;
  assign n35665 = n35664 ^ n14030 ^ n3484 ;
  assign n35666 = n33013 | n35665 ;
  assign n35667 = n26151 & ~n35666 ;
  assign n35668 = ~n14129 & n24280 ;
  assign n35669 = n34760 | n35668 ;
  assign n35670 = ( n4858 & ~n6882 ) | ( n4858 & n21522 ) | ( ~n6882 & n21522 ) ;
  assign n35671 = n35670 ^ n35411 ^ n22979 ;
  assign n35672 = n35671 ^ n33133 ^ 1'b0 ;
  assign n35673 = n32405 & n35672 ;
  assign n35674 = n32899 ^ n11342 ^ 1'b0 ;
  assign n35675 = ( n4747 & ~n28366 ) | ( n4747 & n35674 ) | ( ~n28366 & n35674 ) ;
  assign n35676 = n35590 ^ n15057 ^ 1'b0 ;
  assign n35677 = n21191 ^ n17790 ^ n11693 ;
  assign n35678 = ( n6294 & n7286 ) | ( n6294 & ~n35677 ) | ( n7286 & ~n35677 ) ;
  assign n35679 = n5137 & ~n12332 ;
  assign n35680 = n23125 & n35679 ;
  assign n35681 = n35680 ^ n7038 ^ 1'b0 ;
  assign n35682 = n2689 & ~n35681 ;
  assign n35683 = n35682 ^ n27466 ^ 1'b0 ;
  assign n35684 = ( ~n5322 & n7492 ) | ( ~n5322 & n35683 ) | ( n7492 & n35683 ) ;
  assign n35687 = n26627 ^ n4365 ^ n1446 ;
  assign n35688 = ( ~n4705 & n11639 ) | ( ~n4705 & n35687 ) | ( n11639 & n35687 ) ;
  assign n35689 = n5225 & n35688 ;
  assign n35685 = n28688 ^ n27832 ^ n12228 ;
  assign n35686 = n35685 ^ n23535 ^ 1'b0 ;
  assign n35690 = n35689 ^ n35686 ^ n34642 ;
  assign n35691 = ( n16104 & n24953 ) | ( n16104 & ~n31782 ) | ( n24953 & ~n31782 ) ;
  assign n35692 = n35691 ^ n9254 ^ n3561 ;
  assign n35693 = n31499 ^ n29774 ^ n21642 ;
  assign n35694 = n6923 ^ n6768 ^ 1'b0 ;
  assign n35695 = n18180 | n35694 ;
  assign n35696 = n35693 & ~n35695 ;
  assign n35697 = n35696 ^ n21038 ^ n4022 ;
  assign n35698 = ( ~n7531 & n10907 ) | ( ~n7531 & n12806 ) | ( n10907 & n12806 ) ;
  assign n35699 = n6144 & n20425 ;
  assign n35700 = n25757 & n35699 ;
  assign n35701 = n35698 | n35700 ;
  assign n35702 = ( n6701 & n10600 ) | ( n6701 & n35701 ) | ( n10600 & n35701 ) ;
  assign n35703 = n28235 ^ n20550 ^ n9971 ;
  assign n35704 = n26174 & n33079 ;
  assign n35705 = x115 & n12328 ;
  assign n35706 = n35705 ^ n21552 ^ 1'b0 ;
  assign n35707 = n34006 ^ n30185 ^ n20685 ;
  assign n35708 = ( n719 & n12738 ) | ( n719 & n29097 ) | ( n12738 & n29097 ) ;
  assign n35709 = n20163 ^ n18414 ^ 1'b0 ;
  assign n35710 = n17519 ^ n16503 ^ n11402 ;
  assign n35711 = n10504 | n35710 ;
  assign n35712 = n35711 ^ n20077 ^ 1'b0 ;
  assign n35713 = ~n11643 & n20669 ;
  assign n35714 = n12858 ^ n6424 ^ 1'b0 ;
  assign n35715 = n906 & n35714 ;
  assign n35719 = n22138 ^ n16601 ^ n15619 ;
  assign n35720 = ( n1808 & n3423 ) | ( n1808 & n35719 ) | ( n3423 & n35719 ) ;
  assign n35716 = ~n6015 & n33441 ;
  assign n35717 = n35206 & n35716 ;
  assign n35718 = n32916 | n35717 ;
  assign n35721 = n35720 ^ n35718 ^ 1'b0 ;
  assign n35722 = ( n2631 & n27621 ) | ( n2631 & n35721 ) | ( n27621 & n35721 ) ;
  assign n35723 = ( ~n20872 & n28261 ) | ( ~n20872 & n30116 ) | ( n28261 & n30116 ) ;
  assign n35724 = n481 & n5886 ;
  assign n35725 = n22111 & n35724 ;
  assign n35726 = ( ~n4523 & n20834 ) | ( ~n4523 & n35725 ) | ( n20834 & n35725 ) ;
  assign n35727 = n12794 ^ n6005 ^ 1'b0 ;
  assign n35728 = n34179 | n35727 ;
  assign n35729 = n19461 | n35728 ;
  assign n35730 = n35729 ^ n9114 ^ 1'b0 ;
  assign n35731 = n30570 ^ n20736 ^ 1'b0 ;
  assign n35732 = n12386 | n35731 ;
  assign n35734 = ( n3059 & n5922 ) | ( n3059 & ~n27511 ) | ( n5922 & ~n27511 ) ;
  assign n35733 = n4794 ^ n2139 ^ n883 ;
  assign n35735 = n35734 ^ n35733 ^ 1'b0 ;
  assign n35736 = ~n35732 & n35735 ;
  assign n35737 = n24711 ^ n12142 ^ 1'b0 ;
  assign n35738 = ( ~n4389 & n33896 ) | ( ~n4389 & n35737 ) | ( n33896 & n35737 ) ;
  assign n35739 = n17102 & ~n35738 ;
  assign n35740 = n25323 ^ n22425 ^ n2408 ;
  assign n35741 = n33256 ^ n13762 ^ n12544 ;
  assign n35742 = n35741 ^ n14074 ^ n3538 ;
  assign n35743 = n4873 & ~n10319 ;
  assign n35744 = n8113 ^ n1117 ^ 1'b0 ;
  assign n35746 = ( ~n3966 & n21762 ) | ( ~n3966 & n30420 ) | ( n21762 & n30420 ) ;
  assign n35747 = ( n13719 & n19335 ) | ( n13719 & ~n35746 ) | ( n19335 & ~n35746 ) ;
  assign n35745 = ( n11590 & ~n23085 ) | ( n11590 & n27564 ) | ( ~n23085 & n27564 ) ;
  assign n35748 = n35747 ^ n35745 ^ n22423 ;
  assign n35749 = n15264 ^ n11046 ^ n6444 ;
  assign n35750 = n35749 ^ n3745 ^ 1'b0 ;
  assign n35751 = n35748 & ~n35750 ;
  assign n35752 = ~n15830 & n22603 ;
  assign n35753 = ~n8064 & n11579 ;
  assign n35754 = n35753 ^ n328 ^ 1'b0 ;
  assign n35758 = n3049 & n4442 ;
  assign n35759 = n35758 ^ n8714 ^ 1'b0 ;
  assign n35755 = ( n9596 & ~n16057 ) | ( n9596 & n24140 ) | ( ~n16057 & n24140 ) ;
  assign n35756 = n35755 ^ n7072 ^ 1'b0 ;
  assign n35757 = ~n33425 & n35756 ;
  assign n35760 = n35759 ^ n35757 ^ n1320 ;
  assign n35761 = n34835 ^ n13148 ^ n1670 ;
  assign n35762 = x173 | n7272 ;
  assign n35763 = n4939 ^ n598 ^ 1'b0 ;
  assign n35764 = n35762 | n35763 ;
  assign n35765 = n17552 | n35764 ;
  assign n35766 = n35765 ^ n31574 ^ 1'b0 ;
  assign n35767 = n4245 | n27136 ;
  assign n35768 = n35767 ^ n31400 ^ 1'b0 ;
  assign n35769 = ( n5902 & ~n24135 ) | ( n5902 & n35768 ) | ( ~n24135 & n35768 ) ;
  assign n35770 = n32930 ^ n10209 ^ 1'b0 ;
  assign n35771 = ~n8316 & n35770 ;
  assign n35778 = n8126 | n11140 ;
  assign n35777 = ( n287 & n20345 ) | ( n287 & ~n32027 ) | ( n20345 & ~n32027 ) ;
  assign n35779 = n35778 ^ n35777 ^ n1665 ;
  assign n35772 = n8102 & n12409 ;
  assign n35773 = n35772 ^ n23292 ^ 1'b0 ;
  assign n35774 = ~n4069 & n35773 ;
  assign n35775 = n18432 & n35774 ;
  assign n35776 = n35775 ^ n33845 ^ n7186 ;
  assign n35780 = n35779 ^ n35776 ^ n15937 ;
  assign n35781 = ( n11585 & ~n14031 ) | ( n11585 & n17749 ) | ( ~n14031 & n17749 ) ;
  assign n35782 = n10346 & ~n14723 ;
  assign n35783 = n26665 & n35782 ;
  assign n35784 = n6162 | n35783 ;
  assign n35785 = n35784 ^ n22861 ^ n11962 ;
  assign n35786 = n18369 ^ n10092 ^ 1'b0 ;
  assign n35787 = n30431 ^ n21822 ^ 1'b0 ;
  assign n35788 = ( n35254 & ~n35786 ) | ( n35254 & n35787 ) | ( ~n35786 & n35787 ) ;
  assign n35789 = n2926 & ~n5220 ;
  assign n35790 = n8651 | n21352 ;
  assign n35791 = n19175 & ~n35790 ;
  assign n35792 = ~n7438 & n10513 ;
  assign n35793 = n35792 ^ n5464 ^ 1'b0 ;
  assign n35794 = n18517 ^ n495 ^ 1'b0 ;
  assign n35795 = n15408 | n35794 ;
  assign n35796 = n2015 | n9910 ;
  assign n35797 = n3517 | n35796 ;
  assign n35798 = ( ~n7006 & n33799 ) | ( ~n7006 & n35797 ) | ( n33799 & n35797 ) ;
  assign n35799 = ( n6766 & ~n9783 ) | ( n6766 & n10430 ) | ( ~n9783 & n10430 ) ;
  assign n35800 = ~n13639 & n35799 ;
  assign n35801 = ~n9945 & n35800 ;
  assign n35802 = n7690 ^ n2648 ^ 1'b0 ;
  assign n35803 = ~n9895 & n35802 ;
  assign n35804 = ( ~x25 & n35801 ) | ( ~x25 & n35803 ) | ( n35801 & n35803 ) ;
  assign n35805 = n35804 ^ n33141 ^ 1'b0 ;
  assign n35806 = n22614 ^ n6778 ^ 1'b0 ;
  assign n35807 = ~n20652 & n35806 ;
  assign n35808 = ( ~n17752 & n19606 ) | ( ~n17752 & n35807 ) | ( n19606 & n35807 ) ;
  assign n35809 = n12274 ^ n12047 ^ 1'b0 ;
  assign n35812 = ( n19539 & n28530 ) | ( n19539 & n28929 ) | ( n28530 & n28929 ) ;
  assign n35813 = ( n13969 & n17551 ) | ( n13969 & ~n35812 ) | ( n17551 & ~n35812 ) ;
  assign n35810 = n28707 ^ n19789 ^ 1'b0 ;
  assign n35811 = n6207 | n35810 ;
  assign n35814 = n35813 ^ n35811 ^ n19288 ;
  assign n35817 = ( ~n10530 & n12212 ) | ( ~n10530 & n15537 ) | ( n12212 & n15537 ) ;
  assign n35815 = n8830 ^ n2939 ^ n717 ;
  assign n35816 = n6283 & n35815 ;
  assign n35818 = n35817 ^ n35816 ^ 1'b0 ;
  assign n35819 = n33532 ^ n12614 ^ n9754 ;
  assign n35820 = n35819 ^ n21494 ^ 1'b0 ;
  assign n35821 = n6663 & ~n35820 ;
  assign n35824 = n16998 ^ n5449 ^ n2767 ;
  assign n35825 = n35824 ^ n22623 ^ n20571 ;
  assign n35822 = n31705 ^ n476 ^ 1'b0 ;
  assign n35823 = ~n1706 & n35822 ;
  assign n35826 = n35825 ^ n35823 ^ 1'b0 ;
  assign n35827 = n5300 & ~n13532 ;
  assign n35828 = n35827 ^ n27573 ^ 1'b0 ;
  assign n35829 = n18636 | n35828 ;
  assign n35830 = n28384 ^ n27599 ^ n17423 ;
  assign n35831 = ( n1282 & n14398 ) | ( n1282 & n21696 ) | ( n14398 & n21696 ) ;
  assign n35832 = n35831 ^ n29919 ^ n19625 ;
  assign n35835 = ( n3050 & n12659 ) | ( n3050 & n30193 ) | ( n12659 & n30193 ) ;
  assign n35833 = ( n14558 & n20391 ) | ( n14558 & ~n21025 ) | ( n20391 & ~n21025 ) ;
  assign n35834 = ( n32847 & n34188 ) | ( n32847 & ~n35833 ) | ( n34188 & ~n35833 ) ;
  assign n35836 = n35835 ^ n35834 ^ n15852 ;
  assign n35837 = ( n6355 & n6825 ) | ( n6355 & ~n13258 ) | ( n6825 & ~n13258 ) ;
  assign n35838 = ( n3222 & n33222 ) | ( n3222 & n35837 ) | ( n33222 & n35837 ) ;
  assign n35839 = ( n1056 & n21537 ) | ( n1056 & ~n32218 ) | ( n21537 & ~n32218 ) ;
  assign n35840 = n7567 | n12518 ;
  assign n35841 = ( n7254 & ~n18197 ) | ( n7254 & n35840 ) | ( ~n18197 & n35840 ) ;
  assign n35842 = n35841 ^ n20207 ^ n1292 ;
  assign n35843 = ~n14388 & n23478 ;
  assign n35844 = ~n29099 & n35843 ;
  assign n35845 = n35844 ^ n26425 ^ 1'b0 ;
  assign n35846 = n35845 ^ n12848 ^ 1'b0 ;
  assign n35847 = n19812 ^ n11324 ^ 1'b0 ;
  assign n35848 = n35846 | n35847 ;
  assign n35849 = n22195 ^ n16255 ^ n1740 ;
  assign n35850 = n35849 ^ n22930 ^ 1'b0 ;
  assign n35851 = n21220 & ~n35850 ;
  assign n35852 = n30106 ^ n23753 ^ n280 ;
  assign n35853 = n35852 ^ n34164 ^ 1'b0 ;
  assign n35854 = n5415 & n35853 ;
  assign n35855 = ( n26456 & n32610 ) | ( n26456 & n35854 ) | ( n32610 & n35854 ) ;
  assign n35856 = n31345 ^ n25485 ^ x6 ;
  assign n35857 = n27109 ^ n20943 ^ n1548 ;
  assign n35858 = ( ~n983 & n3038 ) | ( ~n983 & n25649 ) | ( n3038 & n25649 ) ;
  assign n35861 = ~n24485 & n35381 ;
  assign n35859 = n346 & n4380 ;
  assign n35860 = n35859 ^ n1379 ^ 1'b0 ;
  assign n35862 = n35861 ^ n35860 ^ n20411 ;
  assign n35863 = n3638 & ~n12991 ;
  assign n35864 = n21367 & ~n33132 ;
  assign n35865 = ~n35863 & n35864 ;
  assign n35866 = n35865 ^ n29701 ^ n2856 ;
  assign n35867 = n35862 & ~n35866 ;
  assign n35868 = n11539 & n13958 ;
  assign n35869 = ~n18879 & n35868 ;
  assign n35870 = n35869 ^ n19387 ^ 1'b0 ;
  assign n35871 = n23183 & ~n28147 ;
  assign n35872 = n3508 & ~n18364 ;
  assign n35873 = ( ~n14309 & n17542 ) | ( ~n14309 & n35872 ) | ( n17542 & n35872 ) ;
  assign n35874 = n16881 & n28063 ;
  assign n35875 = n35874 ^ n33805 ^ 1'b0 ;
  assign n35876 = n4026 & n35875 ;
  assign n35877 = n18589 | n20787 ;
  assign n35878 = n10497 | n35877 ;
  assign n35879 = n35878 ^ n10976 ^ 1'b0 ;
  assign n35880 = n12997 & ~n35879 ;
  assign n35881 = n34406 ^ n12065 ^ 1'b0 ;
  assign n35882 = n30911 & n35881 ;
  assign n35883 = n13869 ^ n3679 ^ 1'b0 ;
  assign n35884 = n10345 | n35883 ;
  assign n35885 = n20175 & n30128 ;
  assign n35886 = n35885 ^ n14355 ^ 1'b0 ;
  assign n35887 = ( ~n1466 & n19624 ) | ( ~n1466 & n35886 ) | ( n19624 & n35886 ) ;
  assign n35888 = n35887 ^ n18804 ^ n3005 ;
  assign n35889 = n6918 & ~n25235 ;
  assign n35890 = n35889 ^ n6869 ^ n664 ;
  assign n35891 = n5335 & n12462 ;
  assign n35892 = ( n14502 & n15880 ) | ( n14502 & ~n35891 ) | ( n15880 & ~n35891 ) ;
  assign n35896 = ~n1746 & n6209 ;
  assign n35897 = n35896 ^ n18369 ^ 1'b0 ;
  assign n35898 = ( n3313 & ~n13351 ) | ( n3313 & n35897 ) | ( ~n13351 & n35897 ) ;
  assign n35893 = n17552 | n29872 ;
  assign n35894 = n35893 ^ n2759 ^ 1'b0 ;
  assign n35895 = n10939 & ~n35894 ;
  assign n35899 = n35898 ^ n35895 ^ 1'b0 ;
  assign n35900 = n27737 ^ n574 ^ 1'b0 ;
  assign n35901 = n19506 & ~n35900 ;
  assign n35902 = n9959 & n12247 ;
  assign n35903 = n9789 & n35902 ;
  assign n35904 = n35903 ^ n27980 ^ n22705 ;
  assign n35905 = n6138 & ~n35904 ;
  assign n35906 = ~n35901 & n35905 ;
  assign n35907 = n20328 ^ n4656 ^ n2676 ;
  assign n35908 = ( n17770 & n29264 ) | ( n17770 & ~n35907 ) | ( n29264 & ~n35907 ) ;
  assign n35909 = x183 & n16689 ;
  assign n35910 = ~n11066 & n35909 ;
  assign n35911 = n35910 ^ n22592 ^ 1'b0 ;
  assign n35912 = n28481 ^ n17362 ^ 1'b0 ;
  assign n35913 = ( n18423 & n21198 ) | ( n18423 & n22923 ) | ( n21198 & n22923 ) ;
  assign n35914 = ~n25663 & n32559 ;
  assign n35915 = n12463 ^ n10931 ^ 1'b0 ;
  assign n35916 = n35914 | n35915 ;
  assign n35917 = n17058 ^ n9287 ^ n7172 ;
  assign n35918 = n25765 | n35917 ;
  assign n35919 = n9376 & n35918 ;
  assign n35920 = n35916 & n35919 ;
  assign n35921 = n11320 & ~n12432 ;
  assign n35922 = ~n34057 & n35921 ;
  assign n35923 = ~n11633 & n15774 ;
  assign n35924 = n35923 ^ n8971 ^ 1'b0 ;
  assign n35925 = ( ~n5628 & n13223 ) | ( ~n5628 & n18469 ) | ( n13223 & n18469 ) ;
  assign n35926 = n13801 & ~n35925 ;
  assign n35927 = ( n15813 & n16176 ) | ( n15813 & ~n35926 ) | ( n16176 & ~n35926 ) ;
  assign n35928 = n30043 ^ n20221 ^ n896 ;
  assign n35929 = ( n22277 & n35927 ) | ( n22277 & ~n35928 ) | ( n35927 & ~n35928 ) ;
  assign n35930 = n19063 ^ n14722 ^ n2289 ;
  assign n35931 = ( n20178 & n24518 ) | ( n20178 & ~n35930 ) | ( n24518 & ~n35930 ) ;
  assign n35932 = n8486 | n35931 ;
  assign n35933 = n35932 ^ n21394 ^ 1'b0 ;
  assign n35934 = n4144 & ~n25387 ;
  assign n35935 = n6106 | n12377 ;
  assign n35936 = n21292 | n35935 ;
  assign n35937 = n20664 & n35936 ;
  assign n35938 = n32425 & n35937 ;
  assign n35939 = n35938 ^ n24505 ^ n1295 ;
  assign n35940 = ( ~n13875 & n20044 ) | ( ~n13875 & n35939 ) | ( n20044 & n35939 ) ;
  assign n35941 = n13687 ^ n5100 ^ 1'b0 ;
  assign n35942 = n9594 | n35941 ;
  assign n35943 = n2784 | n12319 ;
  assign n35944 = ( n21435 & n31577 ) | ( n21435 & ~n35943 ) | ( n31577 & ~n35943 ) ;
  assign n35948 = n14030 ^ n11772 ^ n1703 ;
  assign n35949 = n35948 ^ n6150 ^ 1'b0 ;
  assign n35945 = n18802 ^ n12987 ^ 1'b0 ;
  assign n35946 = n16520 & n35945 ;
  assign n35947 = n35946 ^ n11220 ^ 1'b0 ;
  assign n35950 = n35949 ^ n35947 ^ n20553 ;
  assign n35951 = n35950 ^ n27587 ^ n9774 ;
  assign n35952 = ~n8019 & n8128 ;
  assign n35953 = n24811 ^ n14074 ^ n12685 ;
  assign n35954 = ( n1572 & n6722 ) | ( n1572 & n9959 ) | ( n6722 & n9959 ) ;
  assign n35955 = n35954 ^ n9554 ^ 1'b0 ;
  assign n35956 = ( n6482 & n35953 ) | ( n6482 & n35955 ) | ( n35953 & n35955 ) ;
  assign n35957 = ( n4467 & n30552 ) | ( n4467 & ~n35956 ) | ( n30552 & ~n35956 ) ;
  assign n35958 = n29472 ^ n20941 ^ n18358 ;
  assign n35961 = n2964 | n15231 ;
  assign n35962 = n35961 ^ n14498 ^ 1'b0 ;
  assign n35963 = n6252 & ~n35962 ;
  assign n35959 = n1729 & ~n3578 ;
  assign n35960 = ~n17020 & n35959 ;
  assign n35964 = n35963 ^ n35960 ^ n18781 ;
  assign n35965 = n35310 ^ n16940 ^ 1'b0 ;
  assign n35966 = ( n5888 & n34206 ) | ( n5888 & n35965 ) | ( n34206 & n35965 ) ;
  assign n35967 = n31549 ^ n23741 ^ n9406 ;
  assign n35968 = ( n2148 & n6028 ) | ( n2148 & n6954 ) | ( n6028 & n6954 ) ;
  assign n35969 = n34087 ^ n19493 ^ n15545 ;
  assign n35970 = n11928 ^ n4156 ^ n1672 ;
  assign n35971 = ( ~n10708 & n35969 ) | ( ~n10708 & n35970 ) | ( n35969 & n35970 ) ;
  assign n35972 = n35971 ^ n15092 ^ 1'b0 ;
  assign n35973 = n30596 ^ n12131 ^ n2520 ;
  assign n35974 = n35973 ^ n28791 ^ n8829 ;
  assign n35975 = n2443 & n25173 ;
  assign n35976 = n6042 & n35975 ;
  assign n35977 = ( n26246 & ~n29669 ) | ( n26246 & n35976 ) | ( ~n29669 & n35976 ) ;
  assign n35978 = n35977 ^ n12598 ^ n2648 ;
  assign n35980 = n4420 | n10974 ;
  assign n35979 = n3671 & ~n17537 ;
  assign n35981 = n35980 ^ n35979 ^ 1'b0 ;
  assign n35982 = n35981 ^ n16749 ^ n16147 ;
  assign n35983 = ( n2818 & n8163 ) | ( n2818 & n11962 ) | ( n8163 & n11962 ) ;
  assign n35987 = n8845 ^ n3798 ^ 1'b0 ;
  assign n35988 = n12563 & ~n35987 ;
  assign n35985 = n25752 ^ n16756 ^ n4610 ;
  assign n35984 = n1076 ^ n859 ^ 1'b0 ;
  assign n35986 = n35985 ^ n35984 ^ 1'b0 ;
  assign n35989 = n35988 ^ n35986 ^ n13869 ;
  assign n35990 = n17519 & n22617 ;
  assign n35991 = n12458 & ~n35990 ;
  assign n35992 = n35991 ^ n34564 ^ n17185 ;
  assign n35993 = n4151 | n6985 ;
  assign n35994 = n35993 ^ n26731 ^ n12029 ;
  assign n35995 = n15213 ^ n5182 ^ 1'b0 ;
  assign n35996 = n35994 & n35995 ;
  assign n35997 = n31254 ^ n12206 ^ n8177 ;
  assign n35998 = ( n16500 & n16607 ) | ( n16500 & ~n17897 ) | ( n16607 & ~n17897 ) ;
  assign n35999 = ( ~n8700 & n14601 ) | ( ~n8700 & n28707 ) | ( n14601 & n28707 ) ;
  assign n36000 = n12053 ^ n3461 ^ n2356 ;
  assign n36001 = ( ~n16669 & n17121 ) | ( ~n16669 & n36000 ) | ( n17121 & n36000 ) ;
  assign n36002 = ( n17829 & ~n22644 ) | ( n17829 & n33222 ) | ( ~n22644 & n33222 ) ;
  assign n36003 = ( n26949 & ~n36001 ) | ( n26949 & n36002 ) | ( ~n36001 & n36002 ) ;
  assign n36004 = ( n1558 & ~n21107 ) | ( n1558 & n36003 ) | ( ~n21107 & n36003 ) ;
  assign n36005 = n35819 ^ n11143 ^ n7089 ;
  assign n36006 = n10976 | n36005 ;
  assign n36007 = ( n5192 & n8782 ) | ( n5192 & n17008 ) | ( n8782 & n17008 ) ;
  assign n36008 = n36007 ^ n1437 ^ 1'b0 ;
  assign n36009 = ~n31224 & n36008 ;
  assign n36010 = n9714 & n33297 ;
  assign n36011 = n36010 ^ n33430 ^ 1'b0 ;
  assign n36012 = n23726 ^ n18153 ^ n12675 ;
  assign n36013 = ~n4537 & n14999 ;
  assign n36014 = n25182 ^ n8813 ^ 1'b0 ;
  assign n36015 = ( n12335 & n33127 ) | ( n12335 & ~n36014 ) | ( n33127 & ~n36014 ) ;
  assign n36016 = ( n9923 & n11565 ) | ( n9923 & n36015 ) | ( n11565 & n36015 ) ;
  assign n36017 = n3871 | n20908 ;
  assign n36018 = n36017 ^ n24511 ^ 1'b0 ;
  assign n36019 = n7101 & ~n28290 ;
  assign n36020 = n36019 ^ n22109 ^ n16581 ;
  assign n36021 = n13858 & n17767 ;
  assign n36023 = ( n15881 & n17387 ) | ( n15881 & ~n28638 ) | ( n17387 & ~n28638 ) ;
  assign n36022 = ( n5618 & ~n11754 ) | ( n5618 & n24187 ) | ( ~n11754 & n24187 ) ;
  assign n36024 = n36023 ^ n36022 ^ n984 ;
  assign n36025 = ( n11400 & n17659 ) | ( n11400 & ~n21443 ) | ( n17659 & ~n21443 ) ;
  assign n36026 = n36025 ^ n3381 ^ 1'b0 ;
  assign n36027 = n24980 ^ n7185 ^ n5238 ;
  assign n36028 = n36027 ^ n12157 ^ n591 ;
  assign n36029 = ( n12712 & ~n27518 ) | ( n12712 & n36028 ) | ( ~n27518 & n36028 ) ;
  assign n36030 = n36029 ^ n31863 ^ n4330 ;
  assign n36031 = ( n13490 & ~n36026 ) | ( n13490 & n36030 ) | ( ~n36026 & n36030 ) ;
  assign n36032 = ( n1866 & n4093 ) | ( n1866 & ~n8340 ) | ( n4093 & ~n8340 ) ;
  assign n36033 = n6633 & ~n15967 ;
  assign n36034 = n36032 & n36033 ;
  assign n36035 = ( n17547 & ~n21653 ) | ( n17547 & n30319 ) | ( ~n21653 & n30319 ) ;
  assign n36036 = n36035 ^ n830 ^ 1'b0 ;
  assign n36037 = ~n1718 & n5326 ;
  assign n36038 = ~n9079 & n36037 ;
  assign n36039 = n36038 ^ n23493 ^ 1'b0 ;
  assign n36040 = n861 & n36039 ;
  assign n36041 = n36040 ^ n25239 ^ n6118 ;
  assign n36042 = ~n36036 & n36041 ;
  assign n36043 = n15084 ^ n8148 ^ n7878 ;
  assign n36044 = n36043 ^ n20257 ^ n19978 ;
  assign n36045 = n11689 ^ n9583 ^ n2939 ;
  assign n36046 = ~n1855 & n36045 ;
  assign n36047 = n19656 ^ n8790 ^ n6689 ;
  assign n36048 = n36047 ^ n7149 ^ 1'b0 ;
  assign n36049 = n10091 & n31993 ;
  assign n36051 = n2564 ^ n2088 ^ n1134 ;
  assign n36052 = n711 & n36051 ;
  assign n36053 = n36052 ^ n4275 ^ 1'b0 ;
  assign n36050 = n6199 & ~n20562 ;
  assign n36054 = n36053 ^ n36050 ^ 1'b0 ;
  assign n36055 = n36054 ^ n5928 ^ 1'b0 ;
  assign n36056 = ~n854 & n14246 ;
  assign n36057 = n20913 ^ n5648 ^ x141 ;
  assign n36058 = ( ~n602 & n36056 ) | ( ~n602 & n36057 ) | ( n36056 & n36057 ) ;
  assign n36059 = n8413 ^ n4406 ^ n1716 ;
  assign n36060 = n36059 ^ n13226 ^ n6917 ;
  assign n36062 = n21497 ^ n8061 ^ 1'b0 ;
  assign n36061 = n19572 ^ n4636 ^ 1'b0 ;
  assign n36063 = n36062 ^ n36061 ^ n27810 ;
  assign n36064 = ~n9385 & n36063 ;
  assign n36065 = ( n6712 & n13286 ) | ( n6712 & ~n27746 ) | ( n13286 & ~n27746 ) ;
  assign n36066 = n29069 ^ n11591 ^ n9176 ;
  assign n36067 = n4009 | n27585 ;
  assign n36068 = ( n36065 & n36066 ) | ( n36065 & ~n36067 ) | ( n36066 & ~n36067 ) ;
  assign n36069 = ( ~n27624 & n32459 ) | ( ~n27624 & n36068 ) | ( n32459 & n36068 ) ;
  assign n36070 = n6050 & ~n36069 ;
  assign n36071 = n15878 & n36070 ;
  assign n36072 = n16964 ^ n13686 ^ n9843 ;
  assign n36073 = n17765 | n19248 ;
  assign n36074 = ( n6676 & ~n7183 ) | ( n6676 & n36073 ) | ( ~n7183 & n36073 ) ;
  assign n36083 = n11206 | n12813 ;
  assign n36084 = n36083 ^ n19526 ^ 1'b0 ;
  assign n36085 = ~n23042 & n36084 ;
  assign n36086 = n18592 & n36085 ;
  assign n36078 = n16533 & ~n23226 ;
  assign n36079 = n11845 & n36078 ;
  assign n36080 = ~n6314 & n36079 ;
  assign n36075 = n18960 ^ n16304 ^ 1'b0 ;
  assign n36076 = n9754 & n36075 ;
  assign n36077 = n12817 & n36076 ;
  assign n36081 = n36080 ^ n36077 ^ n26933 ;
  assign n36082 = n36081 ^ n22783 ^ 1'b0 ;
  assign n36087 = n36086 ^ n36082 ^ n22025 ;
  assign n36088 = n24571 ^ n13654 ^ 1'b0 ;
  assign n36089 = n36088 ^ n28166 ^ n1561 ;
  assign n36090 = ( n740 & n2275 ) | ( n740 & ~n7286 ) | ( n2275 & ~n7286 ) ;
  assign n36091 = n7769 & ~n36090 ;
  assign n36092 = n5326 & ~n18946 ;
  assign n36093 = ~n36091 & n36092 ;
  assign n36094 = ( n8047 & n9707 ) | ( n8047 & ~n14593 ) | ( n9707 & ~n14593 ) ;
  assign n36095 = x227 & ~n36094 ;
  assign n36096 = n36095 ^ n4300 ^ 1'b0 ;
  assign n36097 = n33743 ^ n7218 ^ 1'b0 ;
  assign n36098 = n36097 ^ n10056 ^ 1'b0 ;
  assign n36099 = n3789 | n18409 ;
  assign n36100 = n36099 ^ n23087 ^ n22868 ;
  assign n36101 = n29165 ^ x224 ^ 1'b0 ;
  assign n36102 = n36101 ^ n27216 ^ n9222 ;
  assign n36103 = ( ~n5611 & n15833 ) | ( ~n5611 & n36102 ) | ( n15833 & n36102 ) ;
  assign n36104 = n13875 & n30641 ;
  assign n36105 = n11572 ^ n11230 ^ n5926 ;
  assign n36106 = n36105 ^ n7015 ^ n5799 ;
  assign n36107 = n36104 & n36106 ;
  assign n36110 = n33692 ^ n23680 ^ n1206 ;
  assign n36108 = n6927 ^ n6221 ^ n2553 ;
  assign n36109 = ~n11442 & n36108 ;
  assign n36111 = n36110 ^ n36109 ^ n9963 ;
  assign n36112 = ( n35872 & n36107 ) | ( n35872 & n36111 ) | ( n36107 & n36111 ) ;
  assign n36113 = ( n10500 & n11843 ) | ( n10500 & n16397 ) | ( n11843 & n16397 ) ;
  assign n36114 = n29924 ^ n2629 ^ x192 ;
  assign n36117 = ( n1903 & n5166 ) | ( n1903 & n16256 ) | ( n5166 & n16256 ) ;
  assign n36115 = n34673 ^ n27777 ^ n15034 ;
  assign n36116 = n36115 ^ n18940 ^ n4404 ;
  assign n36118 = n36117 ^ n36116 ^ n4823 ;
  assign n36119 = n36118 ^ n7378 ^ 1'b0 ;
  assign n36121 = ( n6234 & n10742 ) | ( n6234 & n14787 ) | ( n10742 & n14787 ) ;
  assign n36120 = n3124 | n14012 ;
  assign n36122 = n36121 ^ n36120 ^ n10600 ;
  assign n36123 = n36122 ^ n3316 ^ 1'b0 ;
  assign n36124 = n21587 ^ n13589 ^ 1'b0 ;
  assign n36125 = ~n7147 & n36124 ;
  assign n36126 = n24894 ^ n8934 ^ 1'b0 ;
  assign n36127 = ( ~n20770 & n36125 ) | ( ~n20770 & n36126 ) | ( n36125 & n36126 ) ;
  assign n36128 = n2020 & n36127 ;
  assign n36129 = n36128 ^ n8577 ^ 1'b0 ;
  assign n36135 = n36002 ^ n32880 ^ n29183 ;
  assign n36132 = n23270 ^ n14643 ^ n1054 ;
  assign n36130 = ( n311 & ~n12947 ) | ( n311 & n20206 ) | ( ~n12947 & n20206 ) ;
  assign n36131 = n36130 ^ n20396 ^ n2192 ;
  assign n36133 = n36132 ^ n36131 ^ n7547 ;
  assign n36134 = n36133 ^ n17840 ^ n7137 ;
  assign n36136 = n36135 ^ n36134 ^ 1'b0 ;
  assign n36137 = ( n6871 & n10317 ) | ( n6871 & n12070 ) | ( n10317 & n12070 ) ;
  assign n36138 = ( n1168 & ~n20097 ) | ( n1168 & n32264 ) | ( ~n20097 & n32264 ) ;
  assign n36139 = n3242 & ~n16310 ;
  assign n36140 = n36139 ^ n1349 ^ 1'b0 ;
  assign n36141 = n36140 ^ n15893 ^ n1426 ;
  assign n36142 = n35163 ^ n7473 ^ n5929 ;
  assign n36143 = n19205 ^ n8866 ^ n5661 ;
  assign n36144 = n36143 ^ n22797 ^ n2041 ;
  assign n36145 = ( n1195 & ~n8817 ) | ( n1195 & n12455 ) | ( ~n8817 & n12455 ) ;
  assign n36146 = n24227 ^ n4314 ^ 1'b0 ;
  assign n36147 = n36145 & ~n36146 ;
  assign n36148 = ~n24365 & n36147 ;
  assign n36149 = n36148 ^ n7975 ^ 1'b0 ;
  assign n36150 = n36149 ^ n31552 ^ n12385 ;
  assign n36151 = n8990 ^ n540 ^ 1'b0 ;
  assign n36152 = n11072 & ~n36151 ;
  assign n36153 = ~n36150 & n36152 ;
  assign n36154 = n2627 & n12464 ;
  assign n36155 = n21888 ^ n20173 ^ 1'b0 ;
  assign n36156 = n36155 ^ n9159 ^ 1'b0 ;
  assign n36157 = n36156 ^ n19613 ^ n10727 ;
  assign n36158 = ( ~n3859 & n8371 ) | ( ~n3859 & n20280 ) | ( n8371 & n20280 ) ;
  assign n36159 = n13247 ^ n7127 ^ n2068 ;
  assign n36160 = ( n13030 & ~n18051 ) | ( n13030 & n36159 ) | ( ~n18051 & n36159 ) ;
  assign n36161 = n27503 ^ n24219 ^ n7912 ;
  assign n36162 = ( n10799 & n14306 ) | ( n10799 & ~n36161 ) | ( n14306 & ~n36161 ) ;
  assign n36164 = ( n7844 & n21030 ) | ( n7844 & n25678 ) | ( n21030 & n25678 ) ;
  assign n36163 = n5418 | n34582 ;
  assign n36165 = n36164 ^ n36163 ^ n30583 ;
  assign n36168 = ( ~x163 & n8750 ) | ( ~x163 & n24118 ) | ( n8750 & n24118 ) ;
  assign n36166 = n33019 ^ n8022 ^ 1'b0 ;
  assign n36167 = n22066 | n36166 ;
  assign n36169 = n36168 ^ n36167 ^ n1806 ;
  assign n36170 = n7405 ^ x227 ^ 1'b0 ;
  assign n36171 = ( n5390 & n13921 ) | ( n5390 & n17349 ) | ( n13921 & n17349 ) ;
  assign n36172 = ( n27204 & ~n30552 ) | ( n27204 & n36171 ) | ( ~n30552 & n36171 ) ;
  assign n36173 = ( n9486 & n22408 ) | ( n9486 & ~n28620 ) | ( n22408 & ~n28620 ) ;
  assign n36174 = n10381 | n18716 ;
  assign n36175 = ( n2183 & n10016 ) | ( n2183 & ~n36174 ) | ( n10016 & ~n36174 ) ;
  assign n36176 = ( ~n14648 & n16194 ) | ( ~n14648 & n35925 ) | ( n16194 & n35925 ) ;
  assign n36177 = n36176 ^ n8574 ^ n5503 ;
  assign n36178 = n33915 ^ n12239 ^ n5045 ;
  assign n36179 = n28172 ^ n20442 ^ 1'b0 ;
  assign n36180 = n11545 & n36179 ;
  assign n36181 = ( n1408 & n6602 ) | ( n1408 & ~n11803 ) | ( n6602 & ~n11803 ) ;
  assign n36182 = ~n26590 & n36181 ;
  assign n36183 = n36182 ^ n21109 ^ n12954 ;
  assign n36184 = n28581 ^ n22841 ^ n13730 ;
  assign n36185 = ( n7153 & ~n10703 ) | ( n7153 & n36184 ) | ( ~n10703 & n36184 ) ;
  assign n36189 = ~n3311 & n6556 ;
  assign n36187 = n3056 ^ n1452 ^ 1'b0 ;
  assign n36188 = n12246 & n36187 ;
  assign n36186 = n10240 | n17056 ;
  assign n36190 = n36189 ^ n36188 ^ n36186 ;
  assign n36191 = n17142 | n18512 ;
  assign n36192 = n36191 ^ n15245 ^ 1'b0 ;
  assign n36193 = n22844 | n36192 ;
  assign n36194 = n23343 ^ n12463 ^ n4404 ;
  assign n36195 = n3191 & ~n19502 ;
  assign n36196 = ~x222 & n20466 ;
  assign n36197 = n36196 ^ n13264 ^ n843 ;
  assign n36198 = ( n8606 & n32472 ) | ( n8606 & ~n36197 ) | ( n32472 & ~n36197 ) ;
  assign n36199 = ( ~n14031 & n16070 ) | ( ~n14031 & n16099 ) | ( n16070 & n16099 ) ;
  assign n36200 = ( n8659 & n8819 ) | ( n8659 & n12374 ) | ( n8819 & n12374 ) ;
  assign n36201 = ( n2696 & n4866 ) | ( n2696 & ~n33478 ) | ( n4866 & ~n33478 ) ;
  assign n36202 = n3212 & ~n20958 ;
  assign n36203 = ( n10547 & ~n15699 ) | ( n10547 & n36202 ) | ( ~n15699 & n36202 ) ;
  assign n36204 = n14175 | n18840 ;
  assign n36205 = n22257 ^ n11034 ^ n8010 ;
  assign n36206 = ( ~n2694 & n23188 ) | ( ~n2694 & n36205 ) | ( n23188 & n36205 ) ;
  assign n36207 = ( n3561 & n15030 ) | ( n3561 & ~n34140 ) | ( n15030 & ~n34140 ) ;
  assign n36208 = ( n4405 & n10368 ) | ( n4405 & n15573 ) | ( n10368 & n15573 ) ;
  assign n36209 = n36208 ^ n24211 ^ 1'b0 ;
  assign n36210 = ( n4712 & n6064 ) | ( n4712 & n36209 ) | ( n6064 & n36209 ) ;
  assign n36211 = ( ~n19572 & n25368 ) | ( ~n19572 & n31762 ) | ( n25368 & n31762 ) ;
  assign n36212 = n2377 & n33430 ;
  assign n36213 = n26681 ^ n19752 ^ 1'b0 ;
  assign n36214 = n36212 & ~n36213 ;
  assign n36215 = ~n1962 & n3550 ;
  assign n36216 = n18126 | n36215 ;
  assign n36217 = n5403 | n34317 ;
  assign n36218 = n35835 ^ n27370 ^ 1'b0 ;
  assign n36219 = n32273 | n36218 ;
  assign n36220 = ( n6613 & ~n7051 ) | ( n6613 & n21589 ) | ( ~n7051 & n21589 ) ;
  assign n36221 = n36220 ^ n15968 ^ 1'b0 ;
  assign n36222 = n30961 ^ n28330 ^ n20727 ;
  assign n36223 = n33570 ^ n10790 ^ 1'b0 ;
  assign n36224 = ( ~n3051 & n21346 ) | ( ~n3051 & n36223 ) | ( n21346 & n36223 ) ;
  assign n36225 = ( x43 & n11524 ) | ( x43 & ~n36224 ) | ( n11524 & ~n36224 ) ;
  assign n36226 = ( n5745 & n9922 ) | ( n5745 & n29473 ) | ( n9922 & n29473 ) ;
  assign n36227 = n17568 & n17706 ;
  assign n36228 = n20029 | n23364 ;
  assign n36229 = n36228 ^ n13821 ^ 1'b0 ;
  assign n36230 = n36229 ^ n4459 ^ 1'b0 ;
  assign n36231 = n20652 ^ n13758 ^ n8178 ;
  assign n36232 = n1139 & ~n3483 ;
  assign n36233 = n36232 ^ n24086 ^ 1'b0 ;
  assign n36234 = n36233 ^ n22700 ^ 1'b0 ;
  assign n36235 = ( n523 & n23281 ) | ( n523 & n36234 ) | ( n23281 & n36234 ) ;
  assign n36236 = n24137 ^ n23134 ^ n5811 ;
  assign n36237 = n25101 ^ n12396 ^ 1'b0 ;
  assign n36238 = n19526 ^ n12213 ^ n8426 ;
  assign n36239 = n36238 ^ n30021 ^ n13514 ;
  assign n36240 = ~n36237 & n36239 ;
  assign n36241 = ( ~n29814 & n36236 ) | ( ~n29814 & n36240 ) | ( n36236 & n36240 ) ;
  assign n36242 = n34165 ^ n23893 ^ n21667 ;
  assign n36243 = n36242 ^ n33433 ^ n31581 ;
  assign n36248 = ( ~n3546 & n5944 ) | ( ~n3546 & n9195 ) | ( n5944 & n9195 ) ;
  assign n36246 = ~n6986 & n8549 ;
  assign n36247 = n36246 ^ n3759 ^ 1'b0 ;
  assign n36249 = n36248 ^ n36247 ^ 1'b0 ;
  assign n36244 = ~n24016 & n33145 ;
  assign n36245 = n36244 ^ n11837 ^ 1'b0 ;
  assign n36250 = n36249 ^ n36245 ^ n7101 ;
  assign n36251 = ( x173 & ~n27650 ) | ( x173 & n36250 ) | ( ~n27650 & n36250 ) ;
  assign n36252 = ~n24502 & n27247 ;
  assign n36253 = ~n9575 & n36252 ;
  assign n36254 = n30542 ^ n24418 ^ 1'b0 ;
  assign n36255 = n23145 | n36254 ;
  assign n36256 = ( n19802 & n29059 ) | ( n19802 & n36255 ) | ( n29059 & n36255 ) ;
  assign n36262 = ( ~n3122 & n12988 ) | ( ~n3122 & n15882 ) | ( n12988 & n15882 ) ;
  assign n36259 = n13850 ^ n10951 ^ n3142 ;
  assign n36258 = n1448 | n3768 ;
  assign n36260 = n36259 ^ n36258 ^ 1'b0 ;
  assign n36257 = ~n22240 & n23878 ;
  assign n36261 = n36260 ^ n36257 ^ n11497 ;
  assign n36263 = n36262 ^ n36261 ^ n33912 ;
  assign n36264 = n23349 ^ n18162 ^ n6915 ;
  assign n36265 = n29635 ^ n28170 ^ 1'b0 ;
  assign n36266 = ( ~n24241 & n27186 ) | ( ~n24241 & n36265 ) | ( n27186 & n36265 ) ;
  assign n36267 = n3525 & ~n9278 ;
  assign n36268 = n23256 ^ n22358 ^ n11724 ;
  assign n36269 = ( n31343 & n36267 ) | ( n31343 & n36268 ) | ( n36267 & n36268 ) ;
  assign n36270 = ( n13749 & ~n26751 ) | ( n13749 & n36269 ) | ( ~n26751 & n36269 ) ;
  assign n36271 = ~n8122 & n17946 ;
  assign n36272 = ~n30626 & n36271 ;
  assign n36273 = ( n6126 & n19121 ) | ( n6126 & ~n24778 ) | ( n19121 & ~n24778 ) ;
  assign n36274 = n22657 & ~n36273 ;
  assign n36275 = n36274 ^ n6465 ^ 1'b0 ;
  assign n36276 = ( ~n4070 & n19590 ) | ( ~n4070 & n34331 ) | ( n19590 & n34331 ) ;
  assign n36278 = n27150 ^ n7881 ^ 1'b0 ;
  assign n36277 = n27188 ^ n9877 ^ 1'b0 ;
  assign n36279 = n36278 ^ n36277 ^ n35610 ;
  assign n36280 = n8924 | n10008 ;
  assign n36281 = ( n2684 & n26602 ) | ( n2684 & n30551 ) | ( n26602 & n30551 ) ;
  assign n36282 = ( n31817 & n34097 ) | ( n31817 & ~n36281 ) | ( n34097 & ~n36281 ) ;
  assign n36283 = ( n1972 & n32405 ) | ( n1972 & n34327 ) | ( n32405 & n34327 ) ;
  assign n36284 = ( ~n2989 & n5249 ) | ( ~n2989 & n14212 ) | ( n5249 & n14212 ) ;
  assign n36285 = n36284 ^ n31010 ^ 1'b0 ;
  assign n36286 = n24412 ^ n12707 ^ n7926 ;
  assign n36287 = ( n264 & n21178 ) | ( n264 & ~n24197 ) | ( n21178 & ~n24197 ) ;
  assign n36288 = n4196 ^ n3292 ^ 1'b0 ;
  assign n36289 = n36287 & ~n36288 ;
  assign n36290 = n18222 & ~n36289 ;
  assign n36291 = ~n400 & n6275 ;
  assign n36292 = n36291 ^ n2719 ^ 1'b0 ;
  assign n36293 = n13830 & ~n14008 ;
  assign n36294 = n36293 ^ n15572 ^ 1'b0 ;
  assign n36295 = n18797 & ~n23143 ;
  assign n36296 = n36294 & n36295 ;
  assign n36297 = n2370 | n36296 ;
  assign n36298 = n36297 ^ n31847 ^ 1'b0 ;
  assign n36300 = n11206 ^ n7907 ^ n6834 ;
  assign n36301 = n36300 ^ n15227 ^ 1'b0 ;
  assign n36302 = n24479 ^ n8370 ^ 1'b0 ;
  assign n36303 = n5024 & n36302 ;
  assign n36304 = n7189 | n36303 ;
  assign n36305 = ( n14702 & n36301 ) | ( n14702 & n36304 ) | ( n36301 & n36304 ) ;
  assign n36299 = n24584 ^ n17332 ^ 1'b0 ;
  assign n36306 = n36305 ^ n36299 ^ 1'b0 ;
  assign n36307 = ~n17829 & n36306 ;
  assign n36308 = n13815 & n27405 ;
  assign n36309 = ~n13647 & n36308 ;
  assign n36310 = n12697 & n22553 ;
  assign n36311 = n20184 & n36310 ;
  assign n36312 = n36311 ^ n20325 ^ n6812 ;
  assign n36313 = n36312 ^ n21707 ^ 1'b0 ;
  assign n36314 = n36313 ^ n35454 ^ n4594 ;
  assign n36319 = ( n6338 & ~n6992 ) | ( n6338 & n15839 ) | ( ~n6992 & n15839 ) ;
  assign n36318 = ~n1502 & n7188 ;
  assign n36315 = n1005 & n7937 ;
  assign n36316 = ~n9525 & n36315 ;
  assign n36317 = ( n20753 & n23592 ) | ( n20753 & n36316 ) | ( n23592 & n36316 ) ;
  assign n36320 = n36319 ^ n36318 ^ n36317 ;
  assign n36321 = n27570 ^ n14632 ^ n1896 ;
  assign n36322 = n36321 ^ n22169 ^ 1'b0 ;
  assign n36323 = ~n1595 & n36322 ;
  assign n36324 = n36323 ^ n17855 ^ 1'b0 ;
  assign n36326 = n6966 ^ n4720 ^ 1'b0 ;
  assign n36327 = n7103 | n36326 ;
  assign n36325 = ( n9955 & n22518 ) | ( n9955 & n24572 ) | ( n22518 & n24572 ) ;
  assign n36328 = n36327 ^ n36325 ^ n12678 ;
  assign n36329 = n3792 & n3814 ;
  assign n36330 = ~n21154 & n36329 ;
  assign n36331 = n36330 ^ n20145 ^ n8603 ;
  assign n36332 = n23128 & ~n31135 ;
  assign n36333 = ~n3230 & n14688 ;
  assign n36334 = n36333 ^ n12894 ^ 1'b0 ;
  assign n36335 = n36334 ^ n19250 ^ n4376 ;
  assign n36336 = n11898 & n36335 ;
  assign n36337 = ~n2886 & n36336 ;
  assign n36338 = n36337 ^ n22118 ^ n10912 ;
  assign n36339 = n14014 ^ n11918 ^ n1787 ;
  assign n36340 = n8216 & ~n16863 ;
  assign n36341 = n36339 & n36340 ;
  assign n36342 = n36341 ^ n18416 ^ n15986 ;
  assign n36343 = n20777 | n34273 ;
  assign n36344 = n8917 & ~n36343 ;
  assign n36345 = n4438 & n9873 ;
  assign n36346 = ~n26911 & n36345 ;
  assign n36347 = n25167 ^ n6537 ^ 1'b0 ;
  assign n36348 = n19564 ^ n7992 ^ n2101 ;
  assign n36349 = ( n2828 & ~n26032 ) | ( n2828 & n36348 ) | ( ~n26032 & n36348 ) ;
  assign n36350 = n36349 ^ n21867 ^ 1'b0 ;
  assign n36351 = n7632 ^ n5275 ^ n691 ;
  assign n36352 = n30393 ^ n4779 ^ 1'b0 ;
  assign n36353 = n31278 & ~n36352 ;
  assign n36354 = n36353 ^ n32730 ^ n520 ;
  assign n36355 = ( n19848 & n20050 ) | ( n19848 & n30340 ) | ( n20050 & n30340 ) ;
  assign n36356 = n3098 ^ n1579 ^ n1477 ;
  assign n36357 = ( n1910 & n24297 ) | ( n1910 & ~n34291 ) | ( n24297 & ~n34291 ) ;
  assign n36358 = ( n11137 & ~n12786 ) | ( n11137 & n29505 ) | ( ~n12786 & n29505 ) ;
  assign n36359 = ( n36356 & n36357 ) | ( n36356 & n36358 ) | ( n36357 & n36358 ) ;
  assign n36362 = n18176 ^ n11667 ^ 1'b0 ;
  assign n36363 = n13788 & n36362 ;
  assign n36360 = n24054 ^ n19002 ^ n17787 ;
  assign n36361 = n23170 & ~n36360 ;
  assign n36364 = n36363 ^ n36361 ^ 1'b0 ;
  assign n36365 = ( n6960 & ~n7730 ) | ( n6960 & n13969 ) | ( ~n7730 & n13969 ) ;
  assign n36366 = n17589 ^ n1397 ^ 1'b0 ;
  assign n36367 = n36365 & n36366 ;
  assign n36368 = n10140 ^ n5948 ^ n2735 ;
  assign n36369 = ( n719 & n2254 ) | ( n719 & n36368 ) | ( n2254 & n36368 ) ;
  assign n36370 = n36369 ^ n18185 ^ n13272 ;
  assign n36371 = ( n1115 & n1799 ) | ( n1115 & ~n20526 ) | ( n1799 & ~n20526 ) ;
  assign n36372 = ( n883 & ~n36370 ) | ( n883 & n36371 ) | ( ~n36370 & n36371 ) ;
  assign n36376 = ( n10612 & ~n12928 ) | ( n10612 & n14314 ) | ( ~n12928 & n14314 ) ;
  assign n36373 = n24525 ^ n8939 ^ n7327 ;
  assign n36374 = n36373 ^ n10391 ^ n7163 ;
  assign n36375 = n36374 ^ n24083 ^ n6667 ;
  assign n36377 = n36376 ^ n36375 ^ n27540 ;
  assign n36378 = n20223 ^ n5374 ^ 1'b0 ;
  assign n36379 = ~n5352 & n36378 ;
  assign n36380 = n20698 ^ n13345 ^ n2105 ;
  assign n36381 = ( ~n5105 & n36379 ) | ( ~n5105 & n36380 ) | ( n36379 & n36380 ) ;
  assign n36382 = n21804 ^ n16718 ^ n9867 ;
  assign n36383 = ( n2732 & n24169 ) | ( n2732 & ~n32116 ) | ( n24169 & ~n32116 ) ;
  assign n36384 = ( n3270 & ~n19590 ) | ( n3270 & n36383 ) | ( ~n19590 & n36383 ) ;
  assign n36385 = n14521 ^ n11415 ^ n4229 ;
  assign n36386 = n12860 | n30627 ;
  assign n36387 = n12108 ^ n4780 ^ 1'b0 ;
  assign n36388 = n36387 ^ n19655 ^ n5402 ;
  assign n36389 = n35488 ^ n19363 ^ 1'b0 ;
  assign n36390 = n35467 ^ n24822 ^ 1'b0 ;
  assign n36391 = n852 & ~n13460 ;
  assign n36392 = n36391 ^ n7531 ^ 1'b0 ;
  assign n36393 = n1968 | n12136 ;
  assign n36394 = n36392 | n36393 ;
  assign n36395 = n3715 ^ n3340 ^ 1'b0 ;
  assign n36396 = n8419 & n36395 ;
  assign n36397 = ( n1980 & n17082 ) | ( n1980 & ~n28284 ) | ( n17082 & ~n28284 ) ;
  assign n36398 = n7352 ^ n1287 ^ 1'b0 ;
  assign n36399 = n34952 & n36398 ;
  assign n36400 = n36399 ^ n35824 ^ n13403 ;
  assign n36404 = n15370 ^ n9756 ^ 1'b0 ;
  assign n36405 = n2864 & n36404 ;
  assign n36401 = n20378 ^ n10488 ^ 1'b0 ;
  assign n36402 = n19804 ^ n19512 ^ n18385 ;
  assign n36403 = ( ~n17205 & n36401 ) | ( ~n17205 & n36402 ) | ( n36401 & n36402 ) ;
  assign n36406 = n36405 ^ n36403 ^ n25996 ;
  assign n36407 = n34627 ^ n24000 ^ n2306 ;
  assign n36408 = n32376 ^ n29390 ^ n7123 ;
  assign n36409 = n21542 ^ n11300 ^ 1'b0 ;
  assign n36410 = n30672 ^ n23201 ^ n11792 ;
  assign n36416 = ( n2190 & n11626 ) | ( n2190 & ~n13678 ) | ( n11626 & ~n13678 ) ;
  assign n36417 = ( n9283 & n31440 ) | ( n9283 & n36416 ) | ( n31440 & n36416 ) ;
  assign n36418 = ( n7442 & ~n30641 ) | ( n7442 & n36417 ) | ( ~n30641 & n36417 ) ;
  assign n36413 = n8986 ^ n7654 ^ 1'b0 ;
  assign n36414 = n3338 & n36413 ;
  assign n36411 = n16518 ^ n6671 ^ n2798 ;
  assign n36412 = n36411 ^ n11892 ^ n7713 ;
  assign n36415 = n36414 ^ n36412 ^ n15997 ;
  assign n36419 = n36418 ^ n36415 ^ n11320 ;
  assign n36420 = n29985 ^ n23982 ^ n2429 ;
  assign n36421 = ~n2801 & n36420 ;
  assign n36422 = ( n3549 & n7127 ) | ( n3549 & ~n21748 ) | ( n7127 & ~n21748 ) ;
  assign n36423 = n8177 | n26332 ;
  assign n36424 = n36422 | n36423 ;
  assign n36425 = ( ~n6560 & n24170 ) | ( ~n6560 & n28554 ) | ( n24170 & n28554 ) ;
  assign n36426 = n2188 & n36425 ;
  assign n36427 = n36426 ^ n10663 ^ 1'b0 ;
  assign n36428 = n3203 & ~n29733 ;
  assign n36429 = n26003 | n35990 ;
  assign n36430 = n33481 & ~n36429 ;
  assign n36431 = n22620 & ~n36430 ;
  assign n36432 = n36428 & n36431 ;
  assign n36433 = n23950 ^ n11365 ^ 1'b0 ;
  assign n36434 = n10020 | n36433 ;
  assign n36435 = n31260 ^ n15581 ^ n8182 ;
  assign n36436 = n34913 ^ n18186 ^ n15490 ;
  assign n36437 = n21357 ^ n18746 ^ n13418 ;
  assign n36438 = n26162 & n30019 ;
  assign n36439 = n1055 & n26971 ;
  assign n36440 = n5705 ^ n3517 ^ n1882 ;
  assign n36441 = n36440 ^ n32265 ^ 1'b0 ;
  assign n36442 = n25130 ^ n22472 ^ n2905 ;
  assign n36443 = ( ~n15964 & n28054 ) | ( ~n15964 & n36442 ) | ( n28054 & n36442 ) ;
  assign n36444 = ( n5724 & n13360 ) | ( n5724 & n24060 ) | ( n13360 & n24060 ) ;
  assign n36445 = ( ~n2461 & n23901 ) | ( ~n2461 & n25803 ) | ( n23901 & n25803 ) ;
  assign n36446 = n32742 ^ n20627 ^ 1'b0 ;
  assign n36447 = n8336 | n36446 ;
  assign n36448 = n28817 | n36447 ;
  assign n36449 = ( ~n36444 & n36445 ) | ( ~n36444 & n36448 ) | ( n36445 & n36448 ) ;
  assign n36450 = n20381 ^ n14568 ^ 1'b0 ;
  assign n36451 = n8143 & ~n21944 ;
  assign n36452 = ~n34394 & n36451 ;
  assign n36453 = n36452 ^ n25883 ^ n20940 ;
  assign n36454 = n8172 ^ n652 ^ 1'b0 ;
  assign n36455 = n36454 ^ n29955 ^ n5209 ;
  assign n36456 = n36455 ^ n28133 ^ n23260 ;
  assign n36457 = ( n13232 & ~n14405 ) | ( n13232 & n36379 ) | ( ~n14405 & n36379 ) ;
  assign n36458 = ( n6730 & ~n12194 ) | ( n6730 & n36457 ) | ( ~n12194 & n36457 ) ;
  assign n36459 = n18453 ^ n7965 ^ 1'b0 ;
  assign n36460 = n36459 ^ n33367 ^ n7020 ;
  assign n36461 = n3669 | n6765 ;
  assign n36462 = n36461 ^ n4925 ^ n4880 ;
  assign n36463 = n16841 | n36462 ;
  assign n36464 = ( n7107 & n36460 ) | ( n7107 & n36463 ) | ( n36460 & n36463 ) ;
  assign n36465 = ( n8279 & n15725 ) | ( n8279 & n15852 ) | ( n15725 & n15852 ) ;
  assign n36466 = ( ~n11743 & n30296 ) | ( ~n11743 & n36465 ) | ( n30296 & n36465 ) ;
  assign n36467 = n11553 & n18906 ;
  assign n36468 = n3077 & n16331 ;
  assign n36469 = n4832 & n9896 ;
  assign n36470 = n18847 ^ n5490 ^ 1'b0 ;
  assign n36471 = n12735 & n36470 ;
  assign n36472 = ~n36469 & n36471 ;
  assign n36473 = ( n3083 & n28923 ) | ( n3083 & n31141 ) | ( n28923 & n31141 ) ;
  assign n36474 = n4677 | n8762 ;
  assign n36475 = n36474 ^ n9880 ^ n2187 ;
  assign n36476 = n32291 ^ n30121 ^ n16916 ;
  assign n36477 = n33070 ^ n28465 ^ n9350 ;
  assign n36478 = ( ~n16378 & n31949 ) | ( ~n16378 & n33447 ) | ( n31949 & n33447 ) ;
  assign n36479 = n27360 ^ n21642 ^ n8472 ;
  assign n36480 = n32290 ^ n19520 ^ n1576 ;
  assign n36481 = ( n3879 & ~n14528 ) | ( n3879 & n36480 ) | ( ~n14528 & n36480 ) ;
  assign n36482 = ( n6516 & ~n24686 ) | ( n6516 & n36481 ) | ( ~n24686 & n36481 ) ;
  assign n36483 = n35208 ^ n23687 ^ n1752 ;
  assign n36484 = n32832 ^ n31956 ^ n15017 ;
  assign n36485 = ( n2749 & n8438 ) | ( n2749 & n9222 ) | ( n8438 & n9222 ) ;
  assign n36486 = n1237 & n1713 ;
  assign n36487 = n36486 ^ n26349 ^ 1'b0 ;
  assign n36488 = n36487 ^ n15178 ^ 1'b0 ;
  assign n36489 = n36485 | n36488 ;
  assign n36490 = n672 ^ x97 ^ 1'b0 ;
  assign n36491 = n14608 ^ n3474 ^ x161 ;
  assign n36492 = n36491 ^ n6006 ^ 1'b0 ;
  assign n36493 = n36073 & ~n36492 ;
  assign n36494 = ( ~n24281 & n36490 ) | ( ~n24281 & n36493 ) | ( n36490 & n36493 ) ;
  assign n36496 = ~n2985 & n11424 ;
  assign n36497 = ~n34698 & n36496 ;
  assign n36495 = n27244 ^ n6263 ^ n2321 ;
  assign n36498 = n36497 ^ n36495 ^ n35504 ;
  assign n36501 = n13775 & ~n18625 ;
  assign n36499 = ( n668 & n11768 ) | ( n668 & ~n36105 ) | ( n11768 & ~n36105 ) ;
  assign n36500 = n36499 ^ n8730 ^ 1'b0 ;
  assign n36502 = n36501 ^ n36500 ^ n27314 ;
  assign n36503 = n23099 ^ n19144 ^ n5577 ;
  assign n36504 = n2892 | n20488 ;
  assign n36505 = n32066 | n36504 ;
  assign n36506 = ( n4812 & n36503 ) | ( n4812 & ~n36505 ) | ( n36503 & ~n36505 ) ;
  assign n36507 = n323 | n2641 ;
  assign n36508 = n33276 & ~n36507 ;
  assign n36509 = n6963 | n16011 ;
  assign n36510 = n36509 ^ n14094 ^ n1258 ;
  assign n36513 = n760 & n9352 ;
  assign n36511 = n10012 & ~n28907 ;
  assign n36512 = n36511 ^ n11022 ^ 1'b0 ;
  assign n36514 = n36513 ^ n36512 ^ n8285 ;
  assign n36515 = n14043 & n36514 ;
  assign n36516 = n36510 & n36515 ;
  assign n36517 = n32022 ^ n1963 ^ 1'b0 ;
  assign n36518 = ~n28972 & n36517 ;
  assign n36519 = n14313 ^ n12588 ^ n5502 ;
  assign n36520 = n36519 ^ n34006 ^ n10054 ;
  assign n36521 = n36520 ^ n22250 ^ n12545 ;
  assign n36522 = ( n10448 & n18930 ) | ( n10448 & ~n36521 ) | ( n18930 & ~n36521 ) ;
  assign n36523 = ( n4824 & n20763 ) | ( n4824 & ~n36522 ) | ( n20763 & ~n36522 ) ;
  assign n36524 = ( n3450 & n4541 ) | ( n3450 & n10836 ) | ( n4541 & n10836 ) ;
  assign n36525 = n3156 & ~n35746 ;
  assign n36526 = ( n5411 & n36524 ) | ( n5411 & ~n36525 ) | ( n36524 & ~n36525 ) ;
  assign n36527 = ( n814 & n3601 ) | ( n814 & ~n18966 ) | ( n3601 & ~n18966 ) ;
  assign n36528 = n36527 ^ n13144 ^ n12766 ;
  assign n36530 = n5839 & n8076 ;
  assign n36531 = n36530 ^ n11665 ^ 1'b0 ;
  assign n36532 = n36531 ^ n27352 ^ n12781 ;
  assign n36529 = n21217 | n22534 ;
  assign n36533 = n36532 ^ n36529 ^ n33115 ;
  assign n36534 = ( n11722 & n36528 ) | ( n11722 & ~n36533 ) | ( n36528 & ~n36533 ) ;
  assign n36535 = n2160 & ~n35433 ;
  assign n36536 = n19823 | n22481 ;
  assign n36537 = n36536 ^ n32807 ^ 1'b0 ;
  assign n36538 = n29208 ^ n16237 ^ 1'b0 ;
  assign n36539 = n13079 & ~n36538 ;
  assign n36540 = n36539 ^ n5870 ^ n2206 ;
  assign n36541 = n36540 ^ n29889 ^ n2101 ;
  assign n36542 = n1645 | n21056 ;
  assign n36543 = n36542 ^ n8824 ^ n8522 ;
  assign n36544 = n12387 ^ n12152 ^ n8173 ;
  assign n36548 = ( ~n341 & n9289 ) | ( ~n341 & n20584 ) | ( n9289 & n20584 ) ;
  assign n36547 = n21945 ^ n15572 ^ n10920 ;
  assign n36545 = ( n10759 & n10957 ) | ( n10759 & n14398 ) | ( n10957 & n14398 ) ;
  assign n36546 = ~n5627 & n36545 ;
  assign n36549 = n36548 ^ n36547 ^ n36546 ;
  assign n36550 = n28239 ^ n17369 ^ n17169 ;
  assign n36551 = ( n24510 & n36549 ) | ( n24510 & ~n36550 ) | ( n36549 & ~n36550 ) ;
  assign n36552 = n10390 & ~n13317 ;
  assign n36553 = n36552 ^ n20630 ^ 1'b0 ;
  assign n36554 = n36553 ^ n22458 ^ 1'b0 ;
  assign n36557 = n21209 ^ n4802 ^ n3395 ;
  assign n36555 = n1708 & ~n23435 ;
  assign n36556 = n8346 & n36555 ;
  assign n36558 = n36557 ^ n36556 ^ n29687 ;
  assign n36559 = n8450 & ~n21854 ;
  assign n36560 = ( ~x123 & n11171 ) | ( ~x123 & n33822 ) | ( n11171 & n33822 ) ;
  assign n36561 = n36560 ^ n33622 ^ 1'b0 ;
  assign n36562 = n16739 | n36561 ;
  assign n36563 = ( n26902 & n36559 ) | ( n26902 & ~n36562 ) | ( n36559 & ~n36562 ) ;
  assign n36564 = ( n13840 & ~n16660 ) | ( n13840 & n19760 ) | ( ~n16660 & n19760 ) ;
  assign n36565 = n21872 ^ n3170 ^ n3056 ;
  assign n36566 = n26665 ^ n20468 ^ 1'b0 ;
  assign n36567 = ~n15636 & n22393 ;
  assign n36568 = n36567 ^ n30874 ^ 1'b0 ;
  assign n36569 = n30804 ^ n8743 ^ n2128 ;
  assign n36570 = ~n17534 & n18581 ;
  assign n36571 = n36570 ^ n24320 ^ n15903 ;
  assign n36572 = n36571 ^ n8230 ^ 1'b0 ;
  assign n36575 = n31301 ^ n29040 ^ n4189 ;
  assign n36573 = ( n1770 & n16790 ) | ( n1770 & n22526 ) | ( n16790 & n22526 ) ;
  assign n36574 = n36573 ^ n34417 ^ n23929 ;
  assign n36576 = n36575 ^ n36574 ^ n6112 ;
  assign n36577 = ~n3953 & n5515 ;
  assign n36578 = n12374 ^ n11840 ^ 1'b0 ;
  assign n36579 = n5119 & ~n36578 ;
  assign n36580 = n36579 ^ n26996 ^ n20732 ;
  assign n36581 = n19369 ^ n13563 ^ n5106 ;
  assign n36582 = n3044 & ~n3334 ;
  assign n36583 = ~n36581 & n36582 ;
  assign n36584 = n36583 ^ n27455 ^ n24880 ;
  assign n36585 = n13754 & n36584 ;
  assign n36586 = n36585 ^ n32698 ^ 1'b0 ;
  assign n36587 = ( n4931 & n10268 ) | ( n4931 & n29685 ) | ( n10268 & n29685 ) ;
  assign n36588 = n33491 & ~n36587 ;
  assign n36589 = ~n19424 & n36588 ;
  assign n36590 = n17217 & n23671 ;
  assign n36591 = n13425 & ~n36590 ;
  assign n36592 = n36591 ^ n1730 ^ 1'b0 ;
  assign n36593 = n4793 & ~n36592 ;
  assign n36594 = n25614 | n36593 ;
  assign n36595 = n36594 ^ n14089 ^ 1'b0 ;
  assign n36596 = n36595 ^ n32939 ^ n6857 ;
  assign n36597 = ~n1280 & n36596 ;
  assign n36598 = n14021 ^ n9498 ^ n6728 ;
  assign n36599 = ( n28444 & n33750 ) | ( n28444 & ~n36598 ) | ( n33750 & ~n36598 ) ;
  assign n36600 = n2952 & n3824 ;
  assign n36601 = n36600 ^ n12685 ^ 1'b0 ;
  assign n36602 = n36601 ^ n29685 ^ 1'b0 ;
  assign n36603 = n23854 ^ n20931 ^ n280 ;
  assign n36604 = ~n7009 & n36603 ;
  assign n36605 = n36604 ^ n33538 ^ n28500 ;
  assign n36606 = n10979 | n28854 ;
  assign n36607 = n11328 & ~n36606 ;
  assign n36608 = ( n2704 & n7504 ) | ( n2704 & ~n24103 ) | ( n7504 & ~n24103 ) ;
  assign n36609 = n36608 ^ n10664 ^ 1'b0 ;
  assign n36610 = n18373 ^ n16931 ^ n4886 ;
  assign n36611 = n23395 ^ n5229 ^ 1'b0 ;
  assign n36612 = n36611 ^ n19901 ^ n7153 ;
  assign n36613 = ( n14386 & n21292 ) | ( n14386 & n25130 ) | ( n21292 & n25130 ) ;
  assign n36614 = ( ~n1796 & n1939 ) | ( ~n1796 & n17605 ) | ( n1939 & n17605 ) ;
  assign n36615 = n6883 & ~n36614 ;
  assign n36616 = n36615 ^ n23511 ^ 1'b0 ;
  assign n36617 = n19266 | n24487 ;
  assign n36618 = n25819 ^ n15560 ^ 1'b0 ;
  assign n36619 = n36618 ^ n18479 ^ n6253 ;
  assign n36623 = n18364 ^ n4038 ^ 1'b0 ;
  assign n36624 = ~n275 & n8010 ;
  assign n36625 = n29697 & ~n36624 ;
  assign n36626 = ( ~n3298 & n36623 ) | ( ~n3298 & n36625 ) | ( n36623 & n36625 ) ;
  assign n36620 = n4362 & ~n6047 ;
  assign n36621 = n13390 & ~n36620 ;
  assign n36622 = ( n10125 & ~n18149 ) | ( n10125 & n36621 ) | ( ~n18149 & n36621 ) ;
  assign n36627 = n36626 ^ n36622 ^ n13189 ;
  assign n36628 = ( n25560 & n33297 ) | ( n25560 & n34179 ) | ( n33297 & n34179 ) ;
  assign n36629 = n21911 ^ n17611 ^ n13789 ;
  assign n36630 = ( n766 & n842 ) | ( n766 & n21994 ) | ( n842 & n21994 ) ;
  assign n36631 = n4610 ^ n677 ^ 1'b0 ;
  assign n36632 = ~n3914 & n13307 ;
  assign n36633 = ~n9125 & n36632 ;
  assign n36634 = n36633 ^ n35988 ^ n2791 ;
  assign n36635 = n36634 ^ n22219 ^ 1'b0 ;
  assign n36636 = n16521 ^ x48 ^ 1'b0 ;
  assign n36637 = n1095 & ~n16137 ;
  assign n36638 = n36637 ^ n18930 ^ x124 ;
  assign n36639 = n18246 ^ n544 ^ 1'b0 ;
  assign n36640 = n14233 | n36639 ;
  assign n36641 = n20588 | n22249 ;
  assign n36642 = n26665 ^ n825 ^ n290 ;
  assign n36643 = ( n16631 & n28366 ) | ( n16631 & ~n36642 ) | ( n28366 & ~n36642 ) ;
  assign n36652 = n25539 ^ n14347 ^ n11227 ;
  assign n36653 = n36652 ^ n6267 ^ n5277 ;
  assign n36644 = n2896 | n10536 ;
  assign n36645 = ( n4174 & n18765 ) | ( n4174 & n19194 ) | ( n18765 & n19194 ) ;
  assign n36646 = n15955 & n36645 ;
  assign n36647 = n36646 ^ n6980 ^ 1'b0 ;
  assign n36648 = n12831 & ~n29697 ;
  assign n36649 = n16595 & n36648 ;
  assign n36650 = ( ~n14930 & n25522 ) | ( ~n14930 & n36649 ) | ( n25522 & n36649 ) ;
  assign n36651 = ( n36644 & n36647 ) | ( n36644 & ~n36650 ) | ( n36647 & ~n36650 ) ;
  assign n36654 = n36653 ^ n36651 ^ 1'b0 ;
  assign n36655 = ( ~n8133 & n9750 ) | ( ~n8133 & n25384 ) | ( n9750 & n25384 ) ;
  assign n36656 = ( n770 & ~n2853 ) | ( n770 & n12360 ) | ( ~n2853 & n12360 ) ;
  assign n36657 = n2583 & ~n36656 ;
  assign n36658 = n23203 & ~n36657 ;
  assign n36659 = n28065 & n36658 ;
  assign n36661 = ( n1909 & n8813 ) | ( n1909 & ~n10152 ) | ( n8813 & ~n10152 ) ;
  assign n36660 = n16231 & n19917 ;
  assign n36662 = n36661 ^ n36660 ^ 1'b0 ;
  assign n36663 = n29126 ^ n11205 ^ n9534 ;
  assign n36664 = n16727 ^ n2876 ^ 1'b0 ;
  assign n36665 = n36663 | n36664 ;
  assign n36666 = ( n2032 & n27117 ) | ( n2032 & ~n36665 ) | ( n27117 & ~n36665 ) ;
  assign n36667 = n14691 ^ n5014 ^ n4447 ;
  assign n36668 = n13210 ^ n10737 ^ n7183 ;
  assign n36669 = n35488 ^ n3708 ^ n2586 ;
  assign n36670 = n36669 ^ n36109 ^ n2457 ;
  assign n36671 = n36668 & n36670 ;
  assign n36672 = ( ~n1900 & n23479 ) | ( ~n1900 & n34222 ) | ( n23479 & n34222 ) ;
  assign n36673 = ( ~n13407 & n20095 ) | ( ~n13407 & n28498 ) | ( n20095 & n28498 ) ;
  assign n36674 = n36673 ^ n16319 ^ 1'b0 ;
  assign n36675 = n8723 ^ n5055 ^ n1060 ;
  assign n36676 = ~n14769 & n36675 ;
  assign n36677 = n36676 ^ n2506 ^ 1'b0 ;
  assign n36678 = n1179 & n36677 ;
  assign n36679 = ~n16850 & n36678 ;
  assign n36685 = n6797 ^ x101 ^ 1'b0 ;
  assign n36680 = ~n8496 & n9467 ;
  assign n36681 = n36680 ^ n20042 ^ 1'b0 ;
  assign n36682 = n35031 ^ n29345 ^ n6978 ;
  assign n36683 = n36682 ^ n31079 ^ 1'b0 ;
  assign n36684 = ~n36681 & n36683 ;
  assign n36686 = n36685 ^ n36684 ^ n31490 ;
  assign n36687 = n15026 | n18684 ;
  assign n36688 = x208 | n36687 ;
  assign n36691 = n2530 | n8747 ;
  assign n36692 = n36691 ^ n2173 ^ 1'b0 ;
  assign n36689 = n14279 | n14766 ;
  assign n36690 = n36689 ^ n1419 ^ 1'b0 ;
  assign n36693 = n36692 ^ n36690 ^ n35142 ;
  assign n36694 = ( n31474 & ~n36688 ) | ( n31474 & n36693 ) | ( ~n36688 & n36693 ) ;
  assign n36695 = n15715 ^ n12517 ^ n10514 ;
  assign n36696 = ( n6111 & ~n36661 ) | ( n6111 & n36695 ) | ( ~n36661 & n36695 ) ;
  assign n36697 = ( n1933 & ~n22279 ) | ( n1933 & n24716 ) | ( ~n22279 & n24716 ) ;
  assign n36698 = n4715 & n14898 ;
  assign n36699 = n22249 ^ n18663 ^ n17851 ;
  assign n36700 = n36699 ^ n7659 ^ 1'b0 ;
  assign n36701 = n17363 | n36700 ;
  assign n36704 = n1243 & ~n16434 ;
  assign n36705 = ~n29984 & n36704 ;
  assign n36703 = n18738 & n33640 ;
  assign n36706 = n36705 ^ n36703 ^ 1'b0 ;
  assign n36702 = n10802 | n12498 ;
  assign n36707 = n36706 ^ n36702 ^ 1'b0 ;
  assign n36708 = n18613 ^ n12066 ^ n8036 ;
  assign n36709 = n12198 ^ n7856 ^ 1'b0 ;
  assign n36710 = ( n10951 & n16714 ) | ( n10951 & n32914 ) | ( n16714 & n32914 ) ;
  assign n36711 = ( ~n10892 & n14050 ) | ( ~n10892 & n32125 ) | ( n14050 & n32125 ) ;
  assign n36712 = ( x6 & n36710 ) | ( x6 & n36711 ) | ( n36710 & n36711 ) ;
  assign n36716 = n5580 ^ n2443 ^ 1'b0 ;
  assign n36717 = n13596 & ~n36716 ;
  assign n36713 = n10292 ^ n4529 ^ n317 ;
  assign n36714 = n27394 ^ n22389 ^ 1'b0 ;
  assign n36715 = n36713 & ~n36714 ;
  assign n36718 = n36717 ^ n36715 ^ n28068 ;
  assign n36719 = n5304 ^ n3485 ^ 1'b0 ;
  assign n36720 = n36719 ^ n35153 ^ n23322 ;
  assign n36721 = n2176 & ~n22907 ;
  assign n36722 = n20212 ^ n5453 ^ n742 ;
  assign n36723 = n36722 ^ n16574 ^ n880 ;
  assign n36724 = n36722 ^ n30322 ^ n12088 ;
  assign n36725 = n36724 ^ n10728 ^ n2124 ;
  assign n36726 = ( ~n27840 & n28424 ) | ( ~n27840 & n36725 ) | ( n28424 & n36725 ) ;
  assign n36727 = ( ~n3298 & n7822 ) | ( ~n3298 & n11499 ) | ( n7822 & n11499 ) ;
  assign n36728 = n16985 & ~n24664 ;
  assign n36729 = ~n36727 & n36728 ;
  assign n36730 = n869 | n36729 ;
  assign n36731 = n3376 | n36730 ;
  assign n36732 = n35181 ^ n6905 ^ n2583 ;
  assign n36733 = n3279 | n7889 ;
  assign n36734 = n25983 | n36733 ;
  assign n36735 = ( ~n9847 & n18865 ) | ( ~n9847 & n36734 ) | ( n18865 & n36734 ) ;
  assign n36736 = n1186 | n14494 ;
  assign n36737 = n1910 | n4469 ;
  assign n36738 = n36737 ^ n30665 ^ 1'b0 ;
  assign n36739 = ( n13393 & ~n36736 ) | ( n13393 & n36738 ) | ( ~n36736 & n36738 ) ;
  assign n36740 = n19355 | n36739 ;
  assign n36741 = n16718 ^ n15112 ^ n14316 ;
  assign n36742 = n7819 | n36575 ;
  assign n36743 = n36742 ^ n34986 ^ 1'b0 ;
  assign n36744 = n34554 ^ n9773 ^ 1'b0 ;
  assign n36745 = n13689 | n36744 ;
  assign n36746 = n7979 & n21220 ;
  assign n36747 = n36746 ^ n2114 ^ 1'b0 ;
  assign n36748 = n36747 ^ n12526 ^ 1'b0 ;
  assign n36749 = n22253 ^ n17395 ^ n11082 ;
  assign n36751 = n1060 & ~n7946 ;
  assign n36750 = n24957 ^ n2956 ^ n2456 ;
  assign n36752 = n36751 ^ n36750 ^ n1287 ;
  assign n36753 = n11724 ^ n2296 ^ n1133 ;
  assign n36754 = n36753 ^ n24562 ^ n17655 ;
  assign n36755 = ( ~n2663 & n17047 ) | ( ~n2663 & n22716 ) | ( n17047 & n22716 ) ;
  assign n36756 = n25969 ^ n21789 ^ n8869 ;
  assign n36758 = n36065 ^ n14788 ^ n9861 ;
  assign n36757 = n33018 ^ n3196 ^ 1'b0 ;
  assign n36759 = n36758 ^ n36757 ^ n5039 ;
  assign n36760 = n11696 | n36759 ;
  assign n36761 = n36760 ^ n18686 ^ 1'b0 ;
  assign n36762 = ( ~n2245 & n3272 ) | ( ~n2245 & n14535 ) | ( n3272 & n14535 ) ;
  assign n36763 = n36762 ^ n32597 ^ n30778 ;
  assign n36764 = n34167 ^ n11596 ^ 1'b0 ;
  assign n36765 = n4796 & n36764 ;
  assign n36766 = n36765 ^ n11304 ^ n8845 ;
  assign n36767 = ( n13474 & n19462 ) | ( n13474 & n36766 ) | ( n19462 & n36766 ) ;
  assign n36768 = n19455 ^ n4062 ^ 1'b0 ;
  assign n36769 = n1002 & ~n36768 ;
  assign n36770 = ( n14535 & n25533 ) | ( n14535 & n36769 ) | ( n25533 & n36769 ) ;
  assign n36771 = n4881 & ~n31255 ;
  assign n36772 = n18265 ^ n15285 ^ 1'b0 ;
  assign n36773 = ~n36771 & n36772 ;
  assign n36774 = n36773 ^ n346 ^ 1'b0 ;
  assign n36775 = ~n10781 & n36774 ;
  assign n36776 = ~n4012 & n25032 ;
  assign n36777 = n36776 ^ n36509 ^ 1'b0 ;
  assign n36778 = ( n6030 & n7228 ) | ( n6030 & ~n30991 ) | ( n7228 & ~n30991 ) ;
  assign n36779 = n17106 | n36778 ;
  assign n36780 = n18781 ^ n14222 ^ n645 ;
  assign n36781 = ( ~n24703 & n27799 ) | ( ~n24703 & n36780 ) | ( n27799 & n36780 ) ;
  assign n36782 = ( n7451 & n22462 ) | ( n7451 & ~n36781 ) | ( n22462 & ~n36781 ) ;
  assign n36783 = ( n13474 & n14250 ) | ( n13474 & ~n15016 ) | ( n14250 & ~n15016 ) ;
  assign n36784 = n36783 ^ n2742 ^ 1'b0 ;
  assign n36785 = n36784 ^ n34594 ^ n20354 ;
  assign n36786 = ( n7106 & ~n8776 ) | ( n7106 & n30711 ) | ( ~n8776 & n30711 ) ;
  assign n36787 = ( n18544 & n19298 ) | ( n18544 & n36786 ) | ( n19298 & n36786 ) ;
  assign n36788 = n17161 ^ n6202 ^ 1'b0 ;
  assign n36789 = ( n21074 & n33376 ) | ( n21074 & ~n36788 ) | ( n33376 & ~n36788 ) ;
  assign n36790 = n20353 ^ n19136 ^ n7928 ;
  assign n36791 = ( n36787 & n36789 ) | ( n36787 & ~n36790 ) | ( n36789 & ~n36790 ) ;
  assign n36792 = n33211 ^ n24811 ^ n2918 ;
  assign n36793 = n24608 | n32354 ;
  assign n36794 = ~n15305 & n36793 ;
  assign n36795 = n30461 & n36794 ;
  assign n36796 = n3653 ^ n2658 ^ n1588 ;
  assign n36797 = n26980 ^ n6237 ^ 1'b0 ;
  assign n36798 = ~n23636 & n23691 ;
  assign n36799 = n29662 & n36798 ;
  assign n36800 = ( n23161 & ~n36797 ) | ( n23161 & n36799 ) | ( ~n36797 & n36799 ) ;
  assign n36801 = n22940 ^ n21236 ^ n14651 ;
  assign n36802 = n36801 ^ n21048 ^ n19936 ;
  assign n36803 = n36802 ^ n22325 ^ n19349 ;
  assign n36804 = ( n12689 & ~n15402 ) | ( n12689 & n18783 ) | ( ~n15402 & n18783 ) ;
  assign n36805 = n26915 ^ n9202 ^ 1'b0 ;
  assign n36806 = x151 & ~n36805 ;
  assign n36807 = ( n29264 & ~n36804 ) | ( n29264 & n36806 ) | ( ~n36804 & n36806 ) ;
  assign n36808 = n5794 & ~n33381 ;
  assign n36809 = ~n28147 & n36808 ;
  assign n36810 = n12020 & n36809 ;
  assign n36811 = n3703 ^ n2767 ^ 1'b0 ;
  assign n36812 = ( ~n11731 & n13357 ) | ( ~n11731 & n14433 ) | ( n13357 & n14433 ) ;
  assign n36813 = n36812 ^ n18228 ^ n11667 ;
  assign n36814 = n18240 ^ x227 ^ 1'b0 ;
  assign n36815 = n36814 ^ n18414 ^ n5824 ;
  assign n36816 = n30179 ^ n20138 ^ n1154 ;
  assign n36817 = ( n15382 & ~n27826 ) | ( n15382 & n29567 ) | ( ~n27826 & n29567 ) ;
  assign n36818 = n36817 ^ n22317 ^ n17335 ;
  assign n36819 = n11819 ^ n4603 ^ 1'b0 ;
  assign n36820 = n35728 | n36819 ;
  assign n36821 = n30113 ^ n18741 ^ 1'b0 ;
  assign n36822 = ~n24271 & n36821 ;
  assign n36823 = n11280 & ~n20838 ;
  assign n36824 = n36823 ^ n36390 ^ 1'b0 ;
  assign n36825 = n12065 ^ n6023 ^ n2133 ;
  assign n36826 = n1436 | n10690 ;
  assign n36827 = n14020 ^ n7475 ^ 1'b0 ;
  assign n36828 = n36826 | n36827 ;
  assign n36829 = ( n1413 & n18620 ) | ( n1413 & n36828 ) | ( n18620 & n36828 ) ;
  assign n36830 = ( x203 & ~n19432 ) | ( x203 & n25311 ) | ( ~n19432 & n25311 ) ;
  assign n36831 = ~n9883 & n36830 ;
  assign n36832 = n1214 | n1218 ;
  assign n36833 = n36832 ^ n12193 ^ 1'b0 ;
  assign n36835 = ( ~n5554 & n5575 ) | ( ~n5554 & n15329 ) | ( n5575 & n15329 ) ;
  assign n36836 = n36835 ^ n26394 ^ n22614 ;
  assign n36834 = n12416 & n17785 ;
  assign n36837 = n36836 ^ n36834 ^ 1'b0 ;
  assign n36838 = x222 | n1368 ;
  assign n36839 = ( n1716 & n14067 ) | ( n1716 & ~n27070 ) | ( n14067 & ~n27070 ) ;
  assign n36840 = ( x7 & n11264 ) | ( x7 & n36839 ) | ( n11264 & n36839 ) ;
  assign n36841 = ( n34229 & ~n36838 ) | ( n34229 & n36840 ) | ( ~n36838 & n36840 ) ;
  assign n36842 = n34272 ^ n20779 ^ 1'b0 ;
  assign n36843 = ( n4886 & n10745 ) | ( n4886 & n29424 ) | ( n10745 & n29424 ) ;
  assign n36844 = n26947 ^ n8732 ^ n2434 ;
  assign n36845 = ( n1686 & n11833 ) | ( n1686 & ~n20902 ) | ( n11833 & ~n20902 ) ;
  assign n36847 = ~n8115 & n11406 ;
  assign n36848 = n24777 & n36847 ;
  assign n36846 = n27179 ^ n2045 ^ 1'b0 ;
  assign n36849 = n36848 ^ n36846 ^ n2802 ;
  assign n36850 = n36849 ^ n18501 ^ n4568 ;
  assign n36851 = n21854 | n27249 ;
  assign n36852 = n36850 | n36851 ;
  assign n36853 = n11882 & n19692 ;
  assign n36854 = ~n27719 & n36853 ;
  assign n36855 = ( n22082 & n29293 ) | ( n22082 & n35936 ) | ( n29293 & n35936 ) ;
  assign n36856 = n36855 ^ n3214 ^ 1'b0 ;
  assign n36857 = ( ~n10173 & n32037 ) | ( ~n10173 & n33444 ) | ( n32037 & n33444 ) ;
  assign n36858 = ( n3336 & n20416 ) | ( n3336 & ~n36857 ) | ( n20416 & ~n36857 ) ;
  assign n36860 = n11663 ^ n7113 ^ 1'b0 ;
  assign n36859 = n24258 ^ n16426 ^ n3188 ;
  assign n36861 = n36860 ^ n36859 ^ 1'b0 ;
  assign n36862 = n14856 ^ n8462 ^ 1'b0 ;
  assign n36863 = n18167 ^ n14452 ^ n10566 ;
  assign n36864 = ( ~n6211 & n17029 ) | ( ~n6211 & n36863 ) | ( n17029 & n36863 ) ;
  assign n36866 = ( n11842 & ~n16652 ) | ( n11842 & n28065 ) | ( ~n16652 & n28065 ) ;
  assign n36867 = ( n4649 & ~n17739 ) | ( n4649 & n36866 ) | ( ~n17739 & n36866 ) ;
  assign n36868 = ( n1454 & ~n36801 ) | ( n1454 & n36867 ) | ( ~n36801 & n36867 ) ;
  assign n36865 = n34155 ^ n33826 ^ n5194 ;
  assign n36869 = n36868 ^ n36865 ^ n12947 ;
  assign n36870 = n4341 & ~n7443 ;
  assign n36871 = n36870 ^ n18257 ^ n12361 ;
  assign n36872 = n34624 ^ n18287 ^ 1'b0 ;
  assign n36873 = ~n36871 & n36872 ;
  assign n36874 = n10204 ^ n8095 ^ 1'b0 ;
  assign n36875 = n11975 ^ n6127 ^ 1'b0 ;
  assign n36876 = ~n2521 & n36875 ;
  assign n36877 = ( n24155 & ~n36874 ) | ( n24155 & n36876 ) | ( ~n36874 & n36876 ) ;
  assign n36878 = n36877 ^ n33752 ^ n13510 ;
  assign n36879 = ~n3940 & n36878 ;
  assign n36880 = n34672 & n36879 ;
  assign n36881 = n9134 ^ n1302 ^ 1'b0 ;
  assign n36882 = n23662 ^ n9711 ^ 1'b0 ;
  assign n36883 = n22290 & ~n36882 ;
  assign n36884 = n5600 | n36883 ;
  assign n36885 = n6854 ^ n3330 ^ 1'b0 ;
  assign n36886 = ~n4156 & n36885 ;
  assign n36887 = ( n5044 & n7115 ) | ( n5044 & n36886 ) | ( n7115 & n36886 ) ;
  assign n36888 = ( n7577 & n17368 ) | ( n7577 & n36887 ) | ( n17368 & n36887 ) ;
  assign n36889 = ( n2139 & n6833 ) | ( n2139 & ~n24935 ) | ( n6833 & ~n24935 ) ;
  assign n36890 = ( n12598 & n29270 ) | ( n12598 & ~n30284 ) | ( n29270 & ~n30284 ) ;
  assign n36891 = ( n14184 & n36889 ) | ( n14184 & n36890 ) | ( n36889 & n36890 ) ;
  assign n36892 = n36888 & ~n36891 ;
  assign n36893 = n36892 ^ n4498 ^ 1'b0 ;
  assign n36894 = n28040 & n35378 ;
  assign n36895 = ( n14123 & ~n15222 ) | ( n14123 & n16625 ) | ( ~n15222 & n16625 ) ;
  assign n36896 = n27270 & ~n30295 ;
  assign n36897 = ~n31016 & n36896 ;
  assign n36898 = n28076 ^ n13360 ^ 1'b0 ;
  assign n36899 = ~n9047 & n36898 ;
  assign n36900 = n18902 ^ n18041 ^ n16228 ;
  assign n36901 = n36900 ^ n29778 ^ 1'b0 ;
  assign n36902 = n15067 ^ n4301 ^ 1'b0 ;
  assign n36903 = n36902 ^ n3318 ^ n2043 ;
  assign n36904 = n3106 & ~n14497 ;
  assign n36905 = n15857 & n36904 ;
  assign n36906 = n790 | n17093 ;
  assign n36907 = n16418 | n36906 ;
  assign n36908 = n4113 & ~n23370 ;
  assign n36909 = n32926 ^ n27938 ^ n20033 ;
  assign n36910 = ( n2729 & n20585 ) | ( n2729 & ~n33859 ) | ( n20585 & ~n33859 ) ;
  assign n36911 = n7757 ^ n7558 ^ 1'b0 ;
  assign n36912 = ~n15687 & n36911 ;
  assign n36913 = n36912 ^ n34128 ^ 1'b0 ;
  assign n36914 = ~n19477 & n26106 ;
  assign n36915 = ( ~n3014 & n11068 ) | ( ~n3014 & n11210 ) | ( n11068 & n11210 ) ;
  assign n36916 = n24006 ^ n13172 ^ 1'b0 ;
  assign n36917 = ( ~n25097 & n36915 ) | ( ~n25097 & n36916 ) | ( n36915 & n36916 ) ;
  assign n36918 = n19349 ^ n2889 ^ 1'b0 ;
  assign n36919 = n3331 & n36918 ;
  assign n36920 = n36919 ^ n8261 ^ 1'b0 ;
  assign n36921 = ( n13406 & ~n14623 ) | ( n13406 & n36920 ) | ( ~n14623 & n36920 ) ;
  assign n36922 = ( ~n9888 & n17466 ) | ( ~n9888 & n17551 ) | ( n17466 & n17551 ) ;
  assign n36923 = ~n6240 & n36922 ;
  assign n36924 = n8717 ^ n2160 ^ n1633 ;
  assign n36925 = n36924 ^ n28498 ^ n13345 ;
  assign n36926 = n13603 ^ n12219 ^ n5084 ;
  assign n36927 = n36926 ^ n17045 ^ 1'b0 ;
  assign n36928 = n12891 & n36927 ;
  assign n36929 = n10999 & n36928 ;
  assign n36930 = ~n2017 & n36929 ;
  assign n36931 = n23685 ^ n6364 ^ 1'b0 ;
  assign n36932 = ~n27353 & n36931 ;
  assign n36933 = ~n20861 & n36932 ;
  assign n36934 = ~n1109 & n20157 ;
  assign n36935 = n15561 | n36934 ;
  assign n36936 = ( ~n7522 & n8803 ) | ( ~n7522 & n20064 ) | ( n8803 & n20064 ) ;
  assign n36937 = n36936 ^ n13244 ^ n9774 ;
  assign n36938 = n36937 ^ n33202 ^ n23114 ;
  assign n36939 = ( ~n666 & n14564 ) | ( ~n666 & n22690 ) | ( n14564 & n22690 ) ;
  assign n36940 = ( n10133 & n26345 ) | ( n10133 & n29830 ) | ( n26345 & n29830 ) ;
  assign n36941 = ( ~n13789 & n21191 ) | ( ~n13789 & n27334 ) | ( n21191 & n27334 ) ;
  assign n36942 = ~n6833 & n25123 ;
  assign n36943 = n33804 ^ n23324 ^ 1'b0 ;
  assign n36944 = n19256 & n36943 ;
  assign n36945 = ( n3936 & n12260 ) | ( n3936 & ~n15405 ) | ( n12260 & ~n15405 ) ;
  assign n36946 = n36945 ^ n33003 ^ n4330 ;
  assign n36947 = ( n20475 & ~n36061 ) | ( n20475 & n36946 ) | ( ~n36061 & n36946 ) ;
  assign n36948 = ( n981 & n4533 ) | ( n981 & n36947 ) | ( n4533 & n36947 ) ;
  assign n36949 = n3097 ^ n2757 ^ 1'b0 ;
  assign n36952 = ( n3113 & ~n6657 ) | ( n3113 & n28137 ) | ( ~n6657 & n28137 ) ;
  assign n36950 = n1503 & ~n24417 ;
  assign n36951 = n36950 ^ n18010 ^ 1'b0 ;
  assign n36953 = n36952 ^ n36951 ^ 1'b0 ;
  assign n36954 = n12463 ^ n3621 ^ n434 ;
  assign n36955 = n8588 & n36954 ;
  assign n36956 = n36955 ^ x119 ^ 1'b0 ;
  assign n36957 = ( n13031 & n13788 ) | ( n13031 & n36956 ) | ( n13788 & n36956 ) ;
  assign n36958 = ~n19148 & n36957 ;
  assign n36959 = n12616 & ~n23746 ;
  assign n36961 = n28463 & n30665 ;
  assign n36960 = n36601 ^ n35289 ^ 1'b0 ;
  assign n36962 = n36961 ^ n36960 ^ n27550 ;
  assign n36963 = ~n6004 & n34226 ;
  assign n36964 = ~n11075 & n36963 ;
  assign n36965 = ( n19194 & n28243 ) | ( n19194 & ~n36964 ) | ( n28243 & ~n36964 ) ;
  assign n36966 = n25614 ^ n5935 ^ 1'b0 ;
  assign n36967 = n9775 ^ n7792 ^ n5233 ;
  assign n36968 = ( n14684 & n20669 ) | ( n14684 & n20822 ) | ( n20669 & n20822 ) ;
  assign n36969 = ( n29699 & ~n36967 ) | ( n29699 & n36968 ) | ( ~n36967 & n36968 ) ;
  assign n36970 = n1345 | n1763 ;
  assign n36971 = n18257 | n36970 ;
  assign n36972 = n36971 ^ n30535 ^ n12948 ;
  assign n36973 = n27323 & ~n34663 ;
  assign n36974 = n781 | n17036 ;
  assign n36975 = n9922 | n36974 ;
  assign n36976 = n19917 & ~n36975 ;
  assign n36977 = n6139 ^ n615 ^ x70 ;
  assign n36978 = n36977 ^ n19467 ^ n4014 ;
  assign n36979 = n23808 & n36978 ;
  assign n36980 = n36979 ^ n3136 ^ 1'b0 ;
  assign n36981 = ~n3488 & n23505 ;
  assign n36982 = ( ~n6311 & n20012 ) | ( ~n6311 & n36981 ) | ( n20012 & n36981 ) ;
  assign n36983 = n36982 ^ n23032 ^ 1'b0 ;
  assign n36984 = ( ~n18399 & n19820 ) | ( ~n18399 & n35872 ) | ( n19820 & n35872 ) ;
  assign n36985 = n24647 ^ n17230 ^ n16949 ;
  assign n36986 = ( n33050 & n36984 ) | ( n33050 & n36985 ) | ( n36984 & n36985 ) ;
  assign n36987 = n11034 ^ n10762 ^ 1'b0 ;
  assign n36988 = ~n10624 & n36987 ;
  assign n36989 = ( ~n16181 & n23752 ) | ( ~n16181 & n36988 ) | ( n23752 & n36988 ) ;
  assign n36996 = n27632 ^ n18552 ^ 1'b0 ;
  assign n36992 = ( n3741 & ~n7229 ) | ( n3741 & n11382 ) | ( ~n7229 & n11382 ) ;
  assign n36993 = ( ~n3044 & n5847 ) | ( ~n3044 & n36992 ) | ( n5847 & n36992 ) ;
  assign n36994 = n36993 ^ n12291 ^ 1'b0 ;
  assign n36995 = ~n23664 & n36994 ;
  assign n36990 = ( n4630 & n26014 ) | ( n4630 & n29814 ) | ( n26014 & n29814 ) ;
  assign n36991 = n36990 ^ n32574 ^ n1541 ;
  assign n36997 = n36996 ^ n36995 ^ n36991 ;
  assign n36998 = n12699 & n24818 ;
  assign n36999 = ~n17020 & n36998 ;
  assign n37000 = ~n34877 & n36999 ;
  assign n37001 = n22101 ^ n8468 ^ 1'b0 ;
  assign n37002 = n37001 ^ n26314 ^ 1'b0 ;
  assign n37003 = n37000 | n37002 ;
  assign n37004 = n9413 | n27268 ;
  assign n37005 = n31588 & ~n37004 ;
  assign n37006 = n16436 ^ n9494 ^ 1'b0 ;
  assign n37007 = n37006 ^ n30335 ^ n23686 ;
  assign n37008 = n37007 ^ n2570 ^ 1'b0 ;
  assign n37009 = ~n37005 & n37008 ;
  assign n37011 = ( n8163 & ~n16148 ) | ( n8163 & n21423 ) | ( ~n16148 & n21423 ) ;
  assign n37012 = ~n33824 & n34136 ;
  assign n37013 = ~n37011 & n37012 ;
  assign n37010 = ( n18167 & n28837 ) | ( n18167 & n36311 ) | ( n28837 & n36311 ) ;
  assign n37014 = n37013 ^ n37010 ^ n4243 ;
  assign n37015 = n1115 & ~n23501 ;
  assign n37016 = n21457 ^ n3065 ^ 1'b0 ;
  assign n37017 = ( ~n10492 & n12029 ) | ( ~n10492 & n17775 ) | ( n12029 & n17775 ) ;
  assign n37018 = n12524 & n37017 ;
  assign n37019 = n37018 ^ n5578 ^ 1'b0 ;
  assign n37020 = n8036 | n37019 ;
  assign n37021 = n37020 ^ n12526 ^ 1'b0 ;
  assign n37022 = n24475 ^ n10982 ^ 1'b0 ;
  assign n37023 = ( n10004 & n22472 ) | ( n10004 & n37022 ) | ( n22472 & n37022 ) ;
  assign n37024 = n37023 ^ n15582 ^ n4379 ;
  assign n37025 = n25773 & ~n37024 ;
  assign n37026 = n37025 ^ n381 ^ 1'b0 ;
  assign n37027 = n10595 & n24505 ;
  assign n37028 = ~n16896 & n37027 ;
  assign n37029 = n35181 ^ n33132 ^ 1'b0 ;
  assign n37030 = ( n19014 & ~n20807 ) | ( n19014 & n27550 ) | ( ~n20807 & n27550 ) ;
  assign n37031 = ( n15760 & ~n24163 ) | ( n15760 & n27764 ) | ( ~n24163 & n27764 ) ;
  assign n37032 = n37031 ^ n17583 ^ n2568 ;
  assign n37033 = ( n7078 & ~n31073 ) | ( n7078 & n37032 ) | ( ~n31073 & n37032 ) ;
  assign n37034 = n3816 ^ n3601 ^ n1930 ;
  assign n37035 = n37034 ^ n18471 ^ n13964 ;
  assign n37044 = n17727 & n19483 ;
  assign n37041 = n12464 ^ n1344 ^ 1'b0 ;
  assign n37042 = n37041 ^ n25756 ^ n14767 ;
  assign n37037 = n8973 ^ n1574 ^ 1'b0 ;
  assign n37038 = ~n7209 & n37037 ;
  assign n37039 = ( n17987 & n30809 ) | ( n17987 & n37038 ) | ( n30809 & n37038 ) ;
  assign n37036 = n11941 ^ n5557 ^ n5077 ;
  assign n37040 = n37039 ^ n37036 ^ n24212 ;
  assign n37043 = n37042 ^ n37040 ^ n11470 ;
  assign n37045 = n37044 ^ n37043 ^ 1'b0 ;
  assign n37046 = n26065 & n33444 ;
  assign n37047 = n37046 ^ n16846 ^ 1'b0 ;
  assign n37048 = n30956 ^ n12753 ^ x226 ;
  assign n37049 = ( n7994 & n35292 ) | ( n7994 & n37048 ) | ( n35292 & n37048 ) ;
  assign n37050 = ( n2306 & n30217 ) | ( n2306 & ~n30437 ) | ( n30217 & ~n30437 ) ;
  assign n37051 = n30390 ^ n10485 ^ 1'b0 ;
  assign n37052 = n37050 & n37051 ;
  assign n37053 = n1924 & n37052 ;
  assign n37054 = n37049 & n37053 ;
  assign n37055 = n9808 & ~n19705 ;
  assign n37056 = n37055 ^ n28994 ^ n28815 ;
  assign n37057 = n25809 ^ n9854 ^ 1'b0 ;
  assign n37058 = ~n13432 & n37057 ;
  assign n37059 = n37058 ^ n10447 ^ n2941 ;
  assign n37060 = n19718 ^ n1546 ^ 1'b0 ;
  assign n37061 = n15311 & n37060 ;
  assign n37062 = n18527 | n31315 ;
  assign n37063 = n7365 | n28194 ;
  assign n37064 = ( n5504 & ~n13055 ) | ( n5504 & n20708 ) | ( ~n13055 & n20708 ) ;
  assign n37065 = n30669 | n37064 ;
  assign n37066 = ~n17484 & n37065 ;
  assign n37067 = ~n37063 & n37066 ;
  assign n37068 = ( n37061 & ~n37062 ) | ( n37061 & n37067 ) | ( ~n37062 & n37067 ) ;
  assign n37069 = n25098 ^ n20368 ^ 1'b0 ;
  assign n37070 = n37069 ^ n7525 ^ 1'b0 ;
  assign n37071 = n27933 & ~n36295 ;
  assign n37072 = n37071 ^ n12444 ^ 1'b0 ;
  assign n37073 = ( n1672 & ~n2626 ) | ( n1672 & n11747 ) | ( ~n2626 & n11747 ) ;
  assign n37074 = n25261 & n36915 ;
  assign n37075 = ~n37073 & n37074 ;
  assign n37076 = n1756 & ~n37075 ;
  assign n37077 = n37076 ^ n29988 ^ 1'b0 ;
  assign n37078 = ( n3077 & n22025 ) | ( n3077 & n29479 ) | ( n22025 & n29479 ) ;
  assign n37079 = ~n2376 & n2923 ;
  assign n37080 = ~n1189 & n37079 ;
  assign n37081 = n37080 ^ n30364 ^ n2527 ;
  assign n37082 = n32935 ^ n21316 ^ n4358 ;
  assign n37083 = ( n26720 & n36233 ) | ( n26720 & n37082 ) | ( n36233 & n37082 ) ;
  assign n37084 = n37083 ^ n32423 ^ n4810 ;
  assign n37085 = n5286 & ~n33368 ;
  assign n37086 = n4064 & n22506 ;
  assign n37087 = ~n35052 & n37086 ;
  assign n37089 = n7483 ^ n3833 ^ 1'b0 ;
  assign n37090 = n18045 & n37089 ;
  assign n37088 = n14497 & ~n35570 ;
  assign n37091 = n37090 ^ n37088 ^ n25161 ;
  assign n37092 = n11668 ^ n11645 ^ n3573 ;
  assign n37093 = ( n11300 & ~n22740 ) | ( n11300 & n37092 ) | ( ~n22740 & n37092 ) ;
  assign n37094 = n1886 & n34144 ;
  assign n37095 = ( n6281 & n37093 ) | ( n6281 & ~n37094 ) | ( n37093 & ~n37094 ) ;
  assign n37096 = ~n3706 & n34700 ;
  assign n37097 = n37096 ^ n18738 ^ n17118 ;
  assign n37098 = n3051 & n15968 ;
  assign n37099 = n8956 & ~n34215 ;
  assign n37100 = n34548 ^ n34493 ^ n26761 ;
  assign n37101 = ( n10936 & n18335 ) | ( n10936 & ~n36850 ) | ( n18335 & ~n36850 ) ;
  assign n37102 = n17531 ^ n14849 ^ n7671 ;
  assign n37103 = ( ~n12213 & n15950 ) | ( ~n12213 & n37102 ) | ( n15950 & n37102 ) ;
  assign n37104 = n13927 ^ n687 ^ 1'b0 ;
  assign n37105 = ~n37103 & n37104 ;
  assign n37106 = x201 & n19200 ;
  assign n37107 = n37106 ^ n10534 ^ 1'b0 ;
  assign n37108 = n5040 & n37107 ;
  assign n37109 = n11639 & n37108 ;
  assign n37110 = ( ~n1304 & n30470 ) | ( ~n1304 & n30799 ) | ( n30470 & n30799 ) ;
  assign n37111 = n17299 ^ n16013 ^ n6794 ;
  assign n37112 = ( ~n15158 & n29774 ) | ( ~n15158 & n37111 ) | ( n29774 & n37111 ) ;
  assign n37113 = n37112 ^ n20979 ^ n6557 ;
  assign n37114 = n37113 ^ n34037 ^ n859 ;
  assign n37115 = ( n1337 & n11164 ) | ( n1337 & ~n20190 ) | ( n11164 & ~n20190 ) ;
  assign n37116 = n15072 ^ n418 ^ 1'b0 ;
  assign n37117 = ~n17517 & n37116 ;
  assign n37118 = ~n6170 & n33596 ;
  assign n37119 = ~n24416 & n37118 ;
  assign n37120 = n6455 | n14851 ;
  assign n37121 = n37120 ^ n22416 ^ n2228 ;
  assign n37122 = n24346 ^ n5673 ^ 1'b0 ;
  assign n37123 = ( x47 & ~n12126 ) | ( x47 & n15144 ) | ( ~n12126 & n15144 ) ;
  assign n37124 = ( ~n9640 & n9994 ) | ( ~n9640 & n37123 ) | ( n9994 & n37123 ) ;
  assign n37125 = ( n4279 & n5158 ) | ( n4279 & n37124 ) | ( n5158 & n37124 ) ;
  assign n37126 = ( n37121 & n37122 ) | ( n37121 & ~n37125 ) | ( n37122 & ~n37125 ) ;
  assign n37127 = n19399 ^ n16829 ^ n14629 ;
  assign n37128 = ~n8916 & n12411 ;
  assign n37129 = n37128 ^ n6024 ^ 1'b0 ;
  assign n37130 = ( ~n15042 & n21015 ) | ( ~n15042 & n37129 ) | ( n21015 & n37129 ) ;
  assign n37131 = n10022 ^ x144 ^ 1'b0 ;
  assign n37132 = n37131 ^ n5926 ^ n4732 ;
  assign n37133 = ( n1017 & n11587 ) | ( n1017 & n12551 ) | ( n11587 & n12551 ) ;
  assign n37134 = ( n2838 & n8892 ) | ( n2838 & ~n17099 ) | ( n8892 & ~n17099 ) ;
  assign n37135 = n9684 ^ n4215 ^ 1'b0 ;
  assign n37136 = n25445 ^ n22487 ^ 1'b0 ;
  assign n37137 = ( n3785 & ~n6670 ) | ( n3785 & n9040 ) | ( ~n6670 & n9040 ) ;
  assign n37138 = n1360 & n37137 ;
  assign n37139 = ( n11728 & n37136 ) | ( n11728 & ~n37138 ) | ( n37136 & ~n37138 ) ;
  assign n37144 = n36669 ^ n35755 ^ n31162 ;
  assign n37140 = n11303 ^ n7611 ^ n4005 ;
  assign n37141 = ~n14924 & n37140 ;
  assign n37142 = n1698 & n37141 ;
  assign n37143 = n17634 | n37142 ;
  assign n37145 = n37144 ^ n37143 ^ 1'b0 ;
  assign n37147 = n2318 | n14933 ;
  assign n37148 = n3888 & ~n37147 ;
  assign n37146 = n7746 & n19271 ;
  assign n37149 = n37148 ^ n37146 ^ 1'b0 ;
  assign n37155 = n31899 ^ n12917 ^ n3309 ;
  assign n37156 = n27505 | n37155 ;
  assign n37157 = n37156 ^ n14044 ^ 1'b0 ;
  assign n37158 = n6915 | n37157 ;
  assign n37153 = n12325 | n18484 ;
  assign n37154 = n37153 ^ n19771 ^ 1'b0 ;
  assign n37150 = n12732 ^ n5243 ^ 1'b0 ;
  assign n37151 = n7764 | n37150 ;
  assign n37152 = n37151 ^ n8839 ^ 1'b0 ;
  assign n37159 = n37158 ^ n37154 ^ n37152 ;
  assign n37160 = n8088 ^ n4450 ^ n871 ;
  assign n37161 = n26884 | n37160 ;
  assign n37162 = ( n5448 & n24719 ) | ( n5448 & n34745 ) | ( n24719 & n34745 ) ;
  assign n37163 = n11284 ^ n4599 ^ 1'b0 ;
  assign n37164 = n9709 & n37163 ;
  assign n37165 = n431 | n8780 ;
  assign n37166 = n37165 ^ n1927 ^ 1'b0 ;
  assign n37167 = ( x209 & n31291 ) | ( x209 & n37166 ) | ( n31291 & n37166 ) ;
  assign n37168 = n7570 | n10370 ;
  assign n37169 = n37167 | n37168 ;
  assign n37170 = n31384 ^ n17042 ^ n14350 ;
  assign n37171 = n15976 & ~n22942 ;
  assign n37172 = ( n2089 & n12158 ) | ( n2089 & ~n18820 ) | ( n12158 & ~n18820 ) ;
  assign n37173 = ( n17330 & ~n27959 ) | ( n17330 & n37172 ) | ( ~n27959 & n37172 ) ;
  assign n37174 = ( n22249 & n37171 ) | ( n22249 & ~n37173 ) | ( n37171 & ~n37173 ) ;
  assign n37175 = n4793 & ~n18054 ;
  assign n37176 = n37175 ^ n5540 ^ 1'b0 ;
  assign n37177 = n37176 ^ n26554 ^ n26287 ;
  assign n37178 = n29771 ^ n10399 ^ 1'b0 ;
  assign n37179 = n10948 ^ n6841 ^ n4701 ;
  assign n37180 = ( ~n5863 & n27940 ) | ( ~n5863 & n33033 ) | ( n27940 & n33033 ) ;
  assign n37181 = ( n24070 & n37179 ) | ( n24070 & ~n37180 ) | ( n37179 & ~n37180 ) ;
  assign n37182 = ( n5159 & n14219 ) | ( n5159 & ~n23211 ) | ( n14219 & ~n23211 ) ;
  assign n37183 = n37182 ^ n19288 ^ n12483 ;
  assign n37184 = ~n27429 & n37183 ;
  assign n37185 = ~n11854 & n37184 ;
  assign n37186 = n4917 | n7727 ;
  assign n37187 = n20904 & ~n37186 ;
  assign n37188 = ( n12328 & n19492 ) | ( n12328 & ~n20047 ) | ( n19492 & ~n20047 ) ;
  assign n37189 = n8041 ^ n7091 ^ n6593 ;
  assign n37190 = ( n9872 & n19052 ) | ( n9872 & ~n29703 ) | ( n19052 & ~n29703 ) ;
  assign n37191 = n2839 ^ n791 ^ 1'b0 ;
  assign n37192 = n11989 & n37191 ;
  assign n37193 = n14033 & ~n37192 ;
  assign n37194 = n724 & n33326 ;
  assign n37195 = n37194 ^ n5318 ^ 1'b0 ;
  assign n37196 = ( ~n20502 & n23028 ) | ( ~n20502 & n37195 ) | ( n23028 & n37195 ) ;
  assign n37197 = n3999 & ~n7283 ;
  assign n37198 = ~n37196 & n37197 ;
  assign n37199 = n13798 ^ n4894 ^ 1'b0 ;
  assign n37200 = n37199 ^ n17835 ^ n720 ;
  assign n37201 = n3597 | n37200 ;
  assign n37202 = n1133 & ~n37201 ;
  assign n37203 = n37202 ^ n5459 ^ 1'b0 ;
  assign n37204 = n37203 ^ n17004 ^ 1'b0 ;
  assign n37205 = n21406 & ~n37204 ;
  assign n37206 = ( ~n11251 & n19157 ) | ( ~n11251 & n37205 ) | ( n19157 & n37205 ) ;
  assign n37207 = ( n16047 & n16589 ) | ( n16047 & ~n22562 ) | ( n16589 & ~n22562 ) ;
  assign n37208 = n35868 & n37207 ;
  assign n37209 = ( n9502 & n14540 ) | ( n9502 & ~n37208 ) | ( n14540 & ~n37208 ) ;
  assign n37210 = ( ~n12258 & n16073 ) | ( ~n12258 & n20753 ) | ( n16073 & n20753 ) ;
  assign n37211 = n18840 ^ n1198 ^ 1'b0 ;
  assign n37212 = n22030 ^ n18019 ^ n17346 ;
  assign n37213 = ~n21495 & n37212 ;
  assign n37214 = ~n32620 & n37213 ;
  assign n37215 = n31985 ^ n24391 ^ 1'b0 ;
  assign n37216 = n33260 & n37215 ;
  assign n37217 = n28384 ^ n2397 ^ 1'b0 ;
  assign n37220 = n28310 ^ n13847 ^ n7641 ;
  assign n37218 = ( n2715 & n10434 ) | ( n2715 & n24423 ) | ( n10434 & n24423 ) ;
  assign n37219 = n37218 ^ n18608 ^ n18502 ;
  assign n37221 = n37220 ^ n37219 ^ n14573 ;
  assign n37222 = n35379 ^ n18541 ^ n18153 ;
  assign n37223 = n16495 ^ n2752 ^ 1'b0 ;
  assign n37224 = n8762 ^ n5119 ^ 1'b0 ;
  assign n37225 = n16608 & n32674 ;
  assign n37226 = n34105 ^ n33806 ^ n32745 ;
  assign n37227 = ( ~n2104 & n6490 ) | ( ~n2104 & n13356 ) | ( n6490 & n13356 ) ;
  assign n37228 = ( ~n4449 & n31580 ) | ( ~n4449 & n37227 ) | ( n31580 & n37227 ) ;
  assign n37229 = ( n16726 & n37226 ) | ( n16726 & n37228 ) | ( n37226 & n37228 ) ;
  assign n37230 = ~n4142 & n28848 ;
  assign n37231 = n37230 ^ n31725 ^ 1'b0 ;
  assign n37232 = n20365 | n37231 ;
  assign n37233 = n37232 ^ n11591 ^ 1'b0 ;
  assign n37234 = n25329 & n37233 ;
  assign n37235 = ( n5657 & n10209 ) | ( n5657 & ~n10557 ) | ( n10209 & ~n10557 ) ;
  assign n37236 = n4096 & ~n12257 ;
  assign n37237 = n10990 & n37236 ;
  assign n37238 = n19240 | n35230 ;
  assign n37239 = n37238 ^ n34214 ^ 1'b0 ;
  assign n37240 = ( ~n4692 & n24067 ) | ( ~n4692 & n28779 ) | ( n24067 & n28779 ) ;
  assign n37241 = n11408 | n16609 ;
  assign n37242 = n4538 | n17425 ;
  assign n37243 = ~n35296 & n37242 ;
  assign n37244 = n37243 ^ n8495 ^ 1'b0 ;
  assign n37245 = n15624 ^ n9165 ^ 1'b0 ;
  assign n37246 = n19964 & ~n37245 ;
  assign n37247 = n12181 ^ n8621 ^ 1'b0 ;
  assign n37248 = n13718 | n37247 ;
  assign n37249 = ( ~n23753 & n26070 ) | ( ~n23753 & n37248 ) | ( n26070 & n37248 ) ;
  assign n37250 = n32827 & n37249 ;
  assign n37251 = n37246 & n37250 ;
  assign n37255 = n1408 & n10583 ;
  assign n37256 = n37255 ^ n5725 ^ 1'b0 ;
  assign n37254 = n26936 ^ n25765 ^ n22166 ;
  assign n37252 = n18919 ^ n13730 ^ n11195 ;
  assign n37253 = ( n27447 & ~n31301 ) | ( n27447 & n37252 ) | ( ~n31301 & n37252 ) ;
  assign n37257 = n37256 ^ n37254 ^ n37253 ;
  assign n37259 = ~n9238 & n15033 ;
  assign n37258 = n32629 ^ n27618 ^ n2774 ;
  assign n37260 = n37259 ^ n37258 ^ n28320 ;
  assign n37261 = n32042 ^ n17454 ^ 1'b0 ;
  assign n37262 = n3846 & ~n37261 ;
  assign n37263 = n2240 | n33375 ;
  assign n37264 = n24160 ^ n4441 ^ 1'b0 ;
  assign n37265 = ~n37263 & n37264 ;
  assign n37266 = ~n3078 & n37265 ;
  assign n37267 = ~n12697 & n37266 ;
  assign n37268 = ( n10565 & ~n37262 ) | ( n10565 & n37267 ) | ( ~n37262 & n37267 ) ;
  assign n37269 = ~n19855 & n37268 ;
  assign n37270 = n37269 ^ n34411 ^ 1'b0 ;
  assign n37271 = n13232 ^ n9594 ^ 1'b0 ;
  assign n37272 = n25150 & ~n37271 ;
  assign n37273 = ( n4828 & ~n7123 ) | ( n4828 & n8237 ) | ( ~n7123 & n8237 ) ;
  assign n37274 = n37273 ^ n5707 ^ 1'b0 ;
  assign n37275 = n14136 ^ n9848 ^ n5458 ;
  assign n37276 = n17239 | n37275 ;
  assign n37277 = n13971 ^ n8784 ^ n3037 ;
  assign n37278 = n37277 ^ n35368 ^ 1'b0 ;
  assign n37279 = n13536 & n37278 ;
  assign n37280 = ( n31930 & n35350 ) | ( n31930 & n37279 ) | ( n35350 & n37279 ) ;
  assign n37281 = ( n4341 & n37276 ) | ( n4341 & n37280 ) | ( n37276 & n37280 ) ;
  assign n37282 = ~n25532 & n28170 ;
  assign n37283 = n30393 ^ n15276 ^ 1'b0 ;
  assign n37284 = n3517 & n6985 ;
  assign n37285 = ( n5675 & n16898 ) | ( n5675 & n37284 ) | ( n16898 & n37284 ) ;
  assign n37286 = n37285 ^ n6982 ^ n2969 ;
  assign n37287 = n21595 ^ n15311 ^ n909 ;
  assign n37288 = n3209 & n6669 ;
  assign n37289 = n28121 & n37288 ;
  assign n37291 = ~n5823 & n7121 ;
  assign n37292 = n37291 ^ n1755 ^ 1'b0 ;
  assign n37290 = n3583 & n20351 ;
  assign n37293 = n37292 ^ n37290 ^ n12911 ;
  assign n37294 = n9360 & n37293 ;
  assign n37295 = ( n1479 & n2382 ) | ( n1479 & n6920 ) | ( n2382 & n6920 ) ;
  assign n37296 = n1935 & ~n4418 ;
  assign n37297 = ~n37295 & n37296 ;
  assign n37298 = n30113 ^ n10612 ^ n2406 ;
  assign n37299 = n37298 ^ n7702 ^ 1'b0 ;
  assign n37300 = n8080 & ~n37299 ;
  assign n37301 = n34457 ^ n15046 ^ 1'b0 ;
  assign n37303 = ( n3628 & n11139 ) | ( n3628 & ~n12741 ) | ( n11139 & ~n12741 ) ;
  assign n37302 = n13272 | n21559 ;
  assign n37304 = n37303 ^ n37302 ^ 1'b0 ;
  assign n37305 = n13934 | n24627 ;
  assign n37306 = n37304 | n37305 ;
  assign n37307 = ~n1935 & n34301 ;
  assign n37308 = n37307 ^ n5267 ^ 1'b0 ;
  assign n37309 = ( n1382 & n13566 ) | ( n1382 & ~n37308 ) | ( n13566 & ~n37308 ) ;
  assign n37310 = ( ~n33174 & n37306 ) | ( ~n33174 & n37309 ) | ( n37306 & n37309 ) ;
  assign n37311 = n1934 & ~n9742 ;
  assign n37312 = n37310 & n37311 ;
  assign n37313 = n19671 ^ n16207 ^ n16097 ;
  assign n37314 = n25128 & ~n37313 ;
  assign n37315 = n26119 ^ n3048 ^ x254 ;
  assign n37316 = n9846 & n15709 ;
  assign n37317 = n37316 ^ n8885 ^ 1'b0 ;
  assign n37318 = ( n15091 & n37315 ) | ( n15091 & ~n37317 ) | ( n37315 & ~n37317 ) ;
  assign n37319 = ~n7910 & n8880 ;
  assign n37320 = n21245 & n37319 ;
  assign n37321 = n37320 ^ n20998 ^ 1'b0 ;
  assign n37322 = n37321 ^ n35878 ^ n16585 ;
  assign n37323 = ( n890 & ~n2517 ) | ( n890 & n8441 ) | ( ~n2517 & n8441 ) ;
  assign n37324 = n37323 ^ n15582 ^ n8760 ;
  assign n37325 = ~n20849 & n37324 ;
  assign n37326 = n12034 | n37325 ;
  assign n37327 = ~n2224 & n37326 ;
  assign n37328 = n37327 ^ n9796 ^ n2367 ;
  assign n37329 = ( n468 & n2193 ) | ( n468 & n9995 ) | ( n2193 & n9995 ) ;
  assign n37330 = n16121 & n17960 ;
  assign n37331 = n37330 ^ n2352 ^ 1'b0 ;
  assign n37332 = n28097 ^ n301 ^ 1'b0 ;
  assign n37333 = n34872 & ~n37332 ;
  assign n37334 = ( ~n3764 & n4893 ) | ( ~n3764 & n6836 ) | ( n4893 & n6836 ) ;
  assign n37335 = n26718 ^ n10841 ^ n7142 ;
  assign n37336 = ( ~n16949 & n37334 ) | ( ~n16949 & n37335 ) | ( n37334 & n37335 ) ;
  assign n37337 = n22992 ^ n310 ^ 1'b0 ;
  assign n37338 = ( n9866 & n12368 ) | ( n9866 & ~n37337 ) | ( n12368 & ~n37337 ) ;
  assign n37339 = n23863 ^ n22186 ^ n11140 ;
  assign n37340 = ( n26132 & n29422 ) | ( n26132 & ~n31274 ) | ( n29422 & ~n31274 ) ;
  assign n37341 = n7721 ^ n6943 ^ n4644 ;
  assign n37342 = n37341 ^ n32393 ^ n14443 ;
  assign n37343 = n15443 ^ n2640 ^ 1'b0 ;
  assign n37344 = n37342 | n37343 ;
  assign n37345 = ( n667 & n17872 ) | ( n667 & n37344 ) | ( n17872 & n37344 ) ;
  assign n37346 = ( n2242 & n2594 ) | ( n2242 & ~n5628 ) | ( n2594 & ~n5628 ) ;
  assign n37347 = n18553 ^ n14253 ^ 1'b0 ;
  assign n37348 = ( n9379 & n17564 ) | ( n9379 & ~n37347 ) | ( n17564 & ~n37347 ) ;
  assign n37349 = n25811 ^ n11078 ^ n10353 ;
  assign n37350 = n37349 ^ n3608 ^ 1'b0 ;
  assign n37351 = ( ~n6405 & n14432 ) | ( ~n6405 & n37350 ) | ( n14432 & n37350 ) ;
  assign n37352 = ~n16863 & n37351 ;
  assign n37353 = n8203 & ~n13558 ;
  assign n37354 = n37353 ^ n21201 ^ 1'b0 ;
  assign n37355 = n35082 ^ n32825 ^ n18691 ;
  assign n37356 = n11405 & ~n16784 ;
  assign n37357 = ~n10521 & n37356 ;
  assign n37358 = ~n17709 & n21498 ;
  assign n37359 = n13565 & n37358 ;
  assign n37360 = n37359 ^ n33061 ^ 1'b0 ;
  assign n37361 = n37357 | n37360 ;
  assign n37362 = ( n4108 & n9640 ) | ( n4108 & n22645 ) | ( n9640 & n22645 ) ;
  assign n37363 = n37362 ^ n28947 ^ 1'b0 ;
  assign n37364 = ( n1820 & n2480 ) | ( n1820 & n5961 ) | ( n2480 & n5961 ) ;
  assign n37365 = n37364 ^ n29433 ^ n2085 ;
  assign n37366 = n37365 ^ n12398 ^ 1'b0 ;
  assign n37367 = ~n18163 & n28022 ;
  assign n37368 = n37367 ^ n7970 ^ 1'b0 ;
  assign n37369 = n18595 ^ n7822 ^ x167 ;
  assign n37370 = n37369 ^ n14338 ^ 1'b0 ;
  assign n37371 = n1977 & n37370 ;
  assign n37372 = n11499 & n37371 ;
  assign n37373 = n23598 ^ n6175 ^ n4910 ;
  assign n37374 = ~n15443 & n37373 ;
  assign n37375 = ~n37372 & n37374 ;
  assign n37376 = n34001 ^ n17045 ^ 1'b0 ;
  assign n37377 = n37376 ^ n17210 ^ n5019 ;
  assign n37381 = n13883 ^ n9431 ^ n2435 ;
  assign n37378 = ~n4362 & n34446 ;
  assign n37379 = n37378 ^ n11189 ^ 1'b0 ;
  assign n37380 = n5124 | n37379 ;
  assign n37382 = n37381 ^ n37380 ^ 1'b0 ;
  assign n37383 = ( n34082 & n37377 ) | ( n34082 & ~n37382 ) | ( n37377 & ~n37382 ) ;
  assign n37384 = n10384 ^ n887 ^ 1'b0 ;
  assign n37385 = n8798 & n37384 ;
  assign n37386 = n37385 ^ n18797 ^ 1'b0 ;
  assign n37387 = n37386 ^ n23047 ^ 1'b0 ;
  assign n37388 = n17460 & n37387 ;
  assign n37389 = n10095 & n37388 ;
  assign n37390 = ( n6768 & ~n23939 ) | ( n6768 & n32312 ) | ( ~n23939 & n32312 ) ;
  assign n37391 = n17893 ^ n11307 ^ 1'b0 ;
  assign n37392 = n9569 & n37391 ;
  assign n37393 = n37392 ^ n27172 ^ n9853 ;
  assign n37394 = ( n3081 & ~n9510 ) | ( n3081 & n18904 ) | ( ~n9510 & n18904 ) ;
  assign n37395 = ( n24271 & n36804 ) | ( n24271 & n37394 ) | ( n36804 & n37394 ) ;
  assign n37396 = n9668 ^ n6396 ^ 1'b0 ;
  assign n37397 = n37396 ^ n16635 ^ 1'b0 ;
  assign n37398 = n450 & ~n37397 ;
  assign n37399 = ( n6624 & ~n15754 ) | ( n6624 & n31485 ) | ( ~n15754 & n31485 ) ;
  assign n37400 = ( n17975 & n26818 ) | ( n17975 & ~n33060 ) | ( n26818 & ~n33060 ) ;
  assign n37401 = n25113 ^ n17929 ^ n2437 ;
  assign n37402 = ~n4057 & n26122 ;
  assign n37403 = ~n16840 & n37402 ;
  assign n37404 = ( ~n16251 & n37401 ) | ( ~n16251 & n37403 ) | ( n37401 & n37403 ) ;
  assign n37405 = n25339 ^ n5524 ^ n380 ;
  assign n37406 = ( n4003 & n18767 ) | ( n4003 & n27237 ) | ( n18767 & n27237 ) ;
  assign n37407 = n37406 ^ n2912 ^ n1860 ;
  assign n37408 = ( n10667 & ~n11053 ) | ( n10667 & n37407 ) | ( ~n11053 & n37407 ) ;
  assign n37409 = ( n22181 & n30706 ) | ( n22181 & n33245 ) | ( n30706 & n33245 ) ;
  assign n37410 = x241 & n11710 ;
  assign n37411 = n37410 ^ n20591 ^ 1'b0 ;
  assign n37412 = n35977 ^ n20671 ^ 1'b0 ;
  assign n37413 = n33628 ^ n29972 ^ n8140 ;
  assign n37414 = n5267 ^ n3767 ^ 1'b0 ;
  assign n37415 = n37414 ^ n21292 ^ 1'b0 ;
  assign n37416 = ( n1960 & ~n18860 ) | ( n1960 & n37415 ) | ( ~n18860 & n37415 ) ;
  assign n37417 = n32468 ^ n7094 ^ 1'b0 ;
  assign n37418 = n25974 ^ n17360 ^ n6431 ;
  assign n37419 = n37418 ^ n28647 ^ n15047 ;
  assign n37420 = ( n21381 & ~n26535 ) | ( n21381 & n37419 ) | ( ~n26535 & n37419 ) ;
  assign n37421 = ~n1329 & n20619 ;
  assign n37422 = ~n3948 & n37421 ;
  assign n37423 = n37422 ^ n24829 ^ 1'b0 ;
  assign n37424 = n37423 ^ n25801 ^ n8793 ;
  assign n37425 = n34690 & n37424 ;
  assign n37426 = ~n10229 & n12168 ;
  assign n37427 = n37426 ^ n37342 ^ 1'b0 ;
  assign n37428 = x42 & ~n17988 ;
  assign n37429 = n17899 & n37428 ;
  assign n37430 = ~n2373 & n18718 ;
  assign n37431 = ~n36967 & n37430 ;
  assign n37432 = n24693 ^ n2572 ^ 1'b0 ;
  assign n37433 = n37432 ^ n11368 ^ n8488 ;
  assign n37434 = n15952 ^ n10967 ^ n10843 ;
  assign n37435 = n11152 & n16397 ;
  assign n37436 = n11631 & ~n32610 ;
  assign n37437 = ( n4406 & n5524 ) | ( n4406 & n24392 ) | ( n5524 & n24392 ) ;
  assign n37438 = n29893 & n37437 ;
  assign n37439 = ~n37436 & n37438 ;
  assign n37440 = n37435 & n37439 ;
  assign n37441 = ( n6292 & n19061 ) | ( n6292 & ~n22539 ) | ( n19061 & ~n22539 ) ;
  assign n37442 = n28547 ^ n5264 ^ 1'b0 ;
  assign n37447 = ( n6858 & n12841 ) | ( n6858 & ~n20477 ) | ( n12841 & ~n20477 ) ;
  assign n37445 = n33926 ^ n22243 ^ 1'b0 ;
  assign n37443 = n1673 | n15636 ;
  assign n37444 = n30806 & n37443 ;
  assign n37446 = n37445 ^ n37444 ^ 1'b0 ;
  assign n37448 = n37447 ^ n37446 ^ 1'b0 ;
  assign n37449 = ( n7647 & n9805 ) | ( n7647 & n18002 ) | ( n9805 & n18002 ) ;
  assign n37450 = ( n10698 & ~n20699 ) | ( n10698 & n37449 ) | ( ~n20699 & n37449 ) ;
  assign n37451 = ( n12640 & ~n21145 ) | ( n12640 & n24056 ) | ( ~n21145 & n24056 ) ;
  assign n37452 = ( ~n16585 & n22992 ) | ( ~n16585 & n24169 ) | ( n22992 & n24169 ) ;
  assign n37453 = ( n10049 & n27822 ) | ( n10049 & n36425 ) | ( n27822 & n36425 ) ;
  assign n37454 = n21664 ^ n13897 ^ 1'b0 ;
  assign n37455 = ( ~n4671 & n9727 ) | ( ~n4671 & n34454 ) | ( n9727 & n34454 ) ;
  assign n37456 = n16991 | n37455 ;
  assign n37457 = n1952 & ~n14084 ;
  assign n37459 = n36802 ^ n18492 ^ 1'b0 ;
  assign n37458 = n34440 ^ n24337 ^ n12321 ;
  assign n37460 = n37459 ^ n37458 ^ n25948 ;
  assign n37461 = ~n14494 & n16181 ;
  assign n37462 = n37461 ^ n28698 ^ 1'b0 ;
  assign n37463 = n8851 & ~n37462 ;
  assign n37464 = ( x93 & n20358 ) | ( x93 & ~n31899 ) | ( n20358 & ~n31899 ) ;
  assign n37465 = n5740 ^ n4322 ^ 1'b0 ;
  assign n37466 = n35325 & n37465 ;
  assign n37467 = n37466 ^ n11479 ^ 1'b0 ;
  assign n37468 = n909 ^ n336 ^ 1'b0 ;
  assign n37469 = n25308 ^ n5711 ^ 1'b0 ;
  assign n37470 = ( n4322 & ~n12059 ) | ( n4322 & n36945 ) | ( ~n12059 & n36945 ) ;
  assign n37471 = n37470 ^ n19052 ^ 1'b0 ;
  assign n37472 = ( n7676 & n17979 ) | ( n7676 & ~n26549 ) | ( n17979 & ~n26549 ) ;
  assign n37473 = ( n2103 & ~n13759 ) | ( n2103 & n37472 ) | ( ~n13759 & n37472 ) ;
  assign n37475 = n10821 & n13936 ;
  assign n37476 = ~n13051 & n37475 ;
  assign n37474 = ~n30098 & n32152 ;
  assign n37477 = n37476 ^ n37474 ^ 1'b0 ;
  assign n37478 = n31539 ^ n16148 ^ 1'b0 ;
  assign n37479 = n24458 & n37478 ;
  assign n37480 = n19097 ^ n16544 ^ n4207 ;
  assign n37481 = n5371 & ~n37480 ;
  assign n37482 = n37481 ^ n27658 ^ 1'b0 ;
  assign n37483 = n37482 ^ n5090 ^ n1439 ;
  assign n37484 = n9042 ^ n3740 ^ 1'b0 ;
  assign n37485 = n30950 & ~n37484 ;
  assign n37486 = n37483 & n37485 ;
  assign n37487 = n37486 ^ n26578 ^ n5035 ;
  assign n37488 = x161 & ~n1054 ;
  assign n37489 = n37488 ^ n22697 ^ 1'b0 ;
  assign n37490 = n37489 ^ n21490 ^ n14281 ;
  assign n37491 = n19800 | n30941 ;
  assign n37492 = n30859 ^ n25835 ^ n20504 ;
  assign n37493 = n37492 ^ n24318 ^ n2282 ;
  assign n37494 = n16763 ^ n16255 ^ n8523 ;
  assign n37495 = n18000 ^ n922 ^ 1'b0 ;
  assign n37496 = ( ~n482 & n1114 ) | ( ~n482 & n1632 ) | ( n1114 & n1632 ) ;
  assign n37497 = ( n8790 & n37495 ) | ( n8790 & n37496 ) | ( n37495 & n37496 ) ;
  assign n37498 = n7574 ^ n2373 ^ n2254 ;
  assign n37499 = n30241 & n37498 ;
  assign n37500 = n37497 & n37499 ;
  assign n37501 = n29075 ^ n10220 ^ n4628 ;
  assign n37502 = ( n5451 & ~n31042 ) | ( n5451 & n31395 ) | ( ~n31042 & n31395 ) ;
  assign n37503 = n37502 ^ n17915 ^ n3120 ;
  assign n37504 = n23274 ^ n15029 ^ 1'b0 ;
  assign n37505 = ~n12564 & n30159 ;
  assign n37506 = ~n20193 & n37505 ;
  assign n37507 = n24061 ^ n19658 ^ 1'b0 ;
  assign n37508 = ( ~n5607 & n26950 ) | ( ~n5607 & n29919 ) | ( n26950 & n29919 ) ;
  assign n37509 = ( n35215 & n36051 ) | ( n35215 & n37508 ) | ( n36051 & n37508 ) ;
  assign n37510 = ( n1490 & n28967 ) | ( n1490 & n37509 ) | ( n28967 & n37509 ) ;
  assign n37511 = ~n2952 & n14577 ;
  assign n37512 = n37511 ^ n23213 ^ n13055 ;
  assign n37513 = n17975 | n23057 ;
  assign n37514 = n27232 & ~n27406 ;
  assign n37515 = n37514 ^ n20960 ^ n9639 ;
  assign n37516 = ( n8549 & n37513 ) | ( n8549 & ~n37515 ) | ( n37513 & ~n37515 ) ;
  assign n37518 = n5789 | n12370 ;
  assign n37517 = n4855 ^ n2210 ^ 1'b0 ;
  assign n37519 = n37518 ^ n37517 ^ 1'b0 ;
  assign n37520 = ~n8168 & n37519 ;
  assign n37521 = ( n3773 & ~n17445 ) | ( n3773 & n17885 ) | ( ~n17445 & n17885 ) ;
  assign n37522 = n4749 & ~n28854 ;
  assign n37523 = n37521 & n37522 ;
  assign n37524 = ( n1309 & n8652 ) | ( n1309 & ~n26452 ) | ( n8652 & ~n26452 ) ;
  assign n37525 = ( n20036 & ~n37388 ) | ( n20036 & n37524 ) | ( ~n37388 & n37524 ) ;
  assign n37526 = n23521 ^ n17398 ^ n11816 ;
  assign n37527 = n19341 ^ n909 ^ 1'b0 ;
  assign n37528 = ~n37526 & n37527 ;
  assign n37529 = n12191 ^ n10694 ^ 1'b0 ;
  assign n37530 = ( n4896 & n13698 ) | ( n4896 & ~n37529 ) | ( n13698 & ~n37529 ) ;
  assign n37531 = n4621 & ~n37530 ;
  assign n37532 = ( n10265 & n23678 ) | ( n10265 & n33808 ) | ( n23678 & n33808 ) ;
  assign n37533 = n8472 | n29178 ;
  assign n37534 = n21449 | n37533 ;
  assign n37535 = n37534 ^ n35719 ^ 1'b0 ;
  assign n37536 = ( n1979 & n18388 ) | ( n1979 & ~n25594 ) | ( n18388 & ~n25594 ) ;
  assign n37537 = n37536 ^ n13510 ^ 1'b0 ;
  assign n37538 = n13348 ^ n1241 ^ 1'b0 ;
  assign n37539 = n37538 ^ n33964 ^ n31148 ;
  assign n37540 = n31073 ^ n15669 ^ 1'b0 ;
  assign n37541 = x173 | n37540 ;
  assign n37542 = n21476 ^ n2429 ^ 1'b0 ;
  assign n37543 = ~n37541 & n37542 ;
  assign n37544 = ( n10291 & n11613 ) | ( n10291 & ~n12603 ) | ( n11613 & ~n12603 ) ;
  assign n37545 = ~n33646 & n37544 ;
  assign n37546 = ~n37543 & n37545 ;
  assign n37547 = ( n1057 & n3160 ) | ( n1057 & ~n4875 ) | ( n3160 & ~n4875 ) ;
  assign n37548 = n37547 ^ n15883 ^ n2960 ;
  assign n37549 = n331 & n24088 ;
  assign n37550 = n32629 & n37549 ;
  assign n37551 = ( n29526 & n29921 ) | ( n29526 & n33859 ) | ( n29921 & n33859 ) ;
  assign n37552 = ( n18954 & n36379 ) | ( n18954 & ~n37551 ) | ( n36379 & ~n37551 ) ;
  assign n37553 = ( n37548 & n37550 ) | ( n37548 & ~n37552 ) | ( n37550 & ~n37552 ) ;
  assign n37554 = n36518 & ~n37553 ;
  assign n37555 = n28561 ^ n20974 ^ 1'b0 ;
  assign n37556 = ( ~n6907 & n7155 ) | ( ~n6907 & n10840 ) | ( n7155 & n10840 ) ;
  assign n37558 = n4762 ^ n2707 ^ 1'b0 ;
  assign n37559 = n870 & ~n37558 ;
  assign n37560 = ~n26356 & n37559 ;
  assign n37557 = n15064 & n35281 ;
  assign n37561 = n37560 ^ n37557 ^ 1'b0 ;
  assign n37562 = n33440 ^ n8732 ^ n678 ;
  assign n37563 = n37562 ^ n36045 ^ n18431 ;
  assign n37564 = ( n37556 & n37561 ) | ( n37556 & ~n37563 ) | ( n37561 & ~n37563 ) ;
  assign n37565 = n33367 ^ n6942 ^ n4366 ;
  assign n37566 = n1130 ^ n687 ^ 1'b0 ;
  assign n37567 = n37566 ^ n18646 ^ n15552 ;
  assign n37568 = ( n3888 & n6533 ) | ( n3888 & ~n16222 ) | ( n6533 & ~n16222 ) ;
  assign n37569 = ( ~n3119 & n19628 ) | ( ~n3119 & n22125 ) | ( n19628 & n22125 ) ;
  assign n37570 = n9265 ^ n8202 ^ n2091 ;
  assign n37571 = ( ~n1421 & n31801 ) | ( ~n1421 & n37570 ) | ( n31801 & n37570 ) ;
  assign n37572 = n37536 ^ n36121 ^ 1'b0 ;
  assign n37573 = n37572 ^ n9087 ^ n4445 ;
  assign n37574 = ( n3463 & n37571 ) | ( n3463 & n37573 ) | ( n37571 & n37573 ) ;
  assign n37575 = ( n37568 & n37569 ) | ( n37568 & ~n37574 ) | ( n37569 & ~n37574 ) ;
  assign n37576 = ( n6689 & ~n17699 ) | ( n6689 & n37575 ) | ( ~n17699 & n37575 ) ;
  assign n37577 = ( n2250 & n2800 ) | ( n2250 & n9554 ) | ( n2800 & n9554 ) ;
  assign n37578 = n27926 ^ n9533 ^ 1'b0 ;
  assign n37579 = ( ~n6238 & n37577 ) | ( ~n6238 & n37578 ) | ( n37577 & n37578 ) ;
  assign n37580 = n37579 ^ n18384 ^ 1'b0 ;
  assign n37581 = n16188 | n37580 ;
  assign n37582 = n34044 ^ n18661 ^ n17947 ;
  assign n37583 = ~n3481 & n18840 ;
  assign n37584 = n37583 ^ n28547 ^ n2864 ;
  assign n37585 = n13204 & n37584 ;
  assign n37586 = n37582 & n37585 ;
  assign n37587 = n36608 ^ n28079 ^ n17501 ;
  assign n37588 = n30311 & ~n37587 ;
  assign n37590 = n32660 ^ n30061 ^ n6246 ;
  assign n37589 = ( n15555 & n34820 ) | ( n15555 & n36199 ) | ( n34820 & n36199 ) ;
  assign n37591 = n37590 ^ n37589 ^ n3516 ;
  assign n37592 = ~n9410 & n24327 ;
  assign n37593 = ( ~n465 & n18163 ) | ( ~n465 & n37592 ) | ( n18163 & n37592 ) ;
  assign n37594 = n14292 & n29401 ;
  assign n37595 = n16161 ^ n12151 ^ n485 ;
  assign n37596 = n6301 | n37595 ;
  assign n37597 = n4496 | n37596 ;
  assign n37598 = n24413 ^ n11499 ^ n4889 ;
  assign n37599 = ( n13355 & ~n37597 ) | ( n13355 & n37598 ) | ( ~n37597 & n37598 ) ;
  assign n37600 = n37285 ^ n15390 ^ 1'b0 ;
  assign n37601 = n25813 & n37600 ;
  assign n37602 = n34763 ^ n29254 ^ n14012 ;
  assign n37603 = n37501 ^ n37292 ^ n6532 ;
  assign n37604 = n15742 ^ n1623 ^ 1'b0 ;
  assign n37605 = ( ~n2099 & n23156 ) | ( ~n2099 & n25465 ) | ( n23156 & n25465 ) ;
  assign n37606 = n37605 ^ n24596 ^ n19092 ;
  assign n37607 = n11614 ^ n2410 ^ 1'b0 ;
  assign n37608 = n37607 ^ n29740 ^ n6474 ;
  assign n37609 = n6922 ^ n5700 ^ 1'b0 ;
  assign n37612 = n9476 ^ n1061 ^ 1'b0 ;
  assign n37610 = n6681 ^ n2824 ^ n2480 ;
  assign n37611 = n3676 & ~n37610 ;
  assign n37613 = n37612 ^ n37611 ^ 1'b0 ;
  assign n37614 = n19943 ^ n16166 ^ 1'b0 ;
  assign n37615 = n37614 ^ n22451 ^ 1'b0 ;
  assign n37616 = n37613 & n37615 ;
  assign n37617 = ( n3226 & ~n37609 ) | ( n3226 & n37616 ) | ( ~n37609 & n37616 ) ;
  assign n37618 = n5330 & n8541 ;
  assign n37619 = n25663 & n37618 ;
  assign n37623 = ( n16645 & ~n22376 ) | ( n16645 & n29604 ) | ( ~n22376 & n29604 ) ;
  assign n37624 = ( n2011 & n7156 ) | ( n2011 & n37623 ) | ( n7156 & n37623 ) ;
  assign n37620 = ( n2250 & ~n2263 ) | ( n2250 & n17630 ) | ( ~n2263 & n17630 ) ;
  assign n37621 = n37620 ^ n4768 ^ 1'b0 ;
  assign n37622 = n37621 ^ n30956 ^ n15599 ;
  assign n37625 = n37624 ^ n37622 ^ n28133 ;
  assign n37626 = n7973 ^ n4245 ^ 1'b0 ;
  assign n37627 = n37626 ^ n19723 ^ n9851 ;
  assign n37628 = n21526 ^ n6063 ^ n3546 ;
  assign n37629 = n20590 ^ n13321 ^ n10081 ;
  assign n37630 = n20691 ^ n13599 ^ 1'b0 ;
  assign n37631 = ( n1816 & ~n3122 ) | ( n1816 & n26708 ) | ( ~n3122 & n26708 ) ;
  assign n37632 = ( n710 & ~n4113 ) | ( n710 & n13700 ) | ( ~n4113 & n13700 ) ;
  assign n37633 = ~n5866 & n7311 ;
  assign n37634 = ~n3265 & n26000 ;
  assign n37636 = n4803 | n6547 ;
  assign n37637 = n37636 ^ x246 ^ 1'b0 ;
  assign n37638 = ~x224 & n37637 ;
  assign n37635 = ( ~n1645 & n1884 ) | ( ~n1645 & n11679 ) | ( n1884 & n11679 ) ;
  assign n37639 = n37638 ^ n37635 ^ n37482 ;
  assign n37640 = n10794 | n31397 ;
  assign n37641 = n37640 ^ n11387 ^ x70 ;
  assign n37642 = n37641 ^ n22235 ^ 1'b0 ;
  assign n37643 = n36812 | n37642 ;
  assign n37647 = ~n8993 & n15541 ;
  assign n37648 = n37647 ^ n17011 ^ 1'b0 ;
  assign n37644 = n36623 ^ n13545 ^ 1'b0 ;
  assign n37645 = ( n10191 & ~n11802 ) | ( n10191 & n37644 ) | ( ~n11802 & n37644 ) ;
  assign n37646 = n37645 ^ n12529 ^ 1'b0 ;
  assign n37649 = n37648 ^ n37646 ^ n9078 ;
  assign n37650 = n37643 | n37649 ;
  assign n37651 = n37639 & ~n37650 ;
  assign n37652 = n34974 ^ n9029 ^ n871 ;
  assign n37653 = n14668 & ~n37566 ;
  assign n37654 = ~n37652 & n37653 ;
  assign n37655 = n37492 ^ n30933 ^ 1'b0 ;
  assign n37656 = n6376 & n19793 ;
  assign n37657 = n37656 ^ n2313 ^ 1'b0 ;
  assign n37658 = n17933 ^ n7097 ^ n4803 ;
  assign n37659 = n37657 | n37658 ;
  assign n37660 = n18577 ^ n1770 ^ n517 ;
  assign n37661 = n21920 ^ n19590 ^ n1719 ;
  assign n37662 = ( n22535 & ~n37660 ) | ( n22535 & n37661 ) | ( ~n37660 & n37661 ) ;
  assign n37663 = n34848 ^ n3030 ^ 1'b0 ;
  assign n37664 = ( ~n2113 & n10218 ) | ( ~n2113 & n29588 ) | ( n10218 & n29588 ) ;
  assign n37665 = n5719 ^ n1484 ^ 1'b0 ;
  assign n37666 = ~n5014 & n14250 ;
  assign n37667 = n37666 ^ n3808 ^ 1'b0 ;
  assign n37668 = n3555 & n4904 ;
  assign n37669 = ~n11205 & n37668 ;
  assign n37670 = n7462 ^ n6338 ^ n3412 ;
  assign n37671 = ~n37669 & n37670 ;
  assign n37672 = n37667 & n37671 ;
  assign n37673 = n7845 | n37672 ;
  assign n37674 = n12301 & ~n37673 ;
  assign n37675 = n9218 & ~n30011 ;
  assign n37676 = n37675 ^ n23995 ^ n13090 ;
  assign n37678 = n14017 ^ n9424 ^ n8783 ;
  assign n37677 = n3244 | n7072 ;
  assign n37679 = n37678 ^ n37677 ^ 1'b0 ;
  assign n37680 = n37679 ^ n16523 ^ n14145 ;
  assign n37681 = n32231 ^ n7447 ^ n5348 ;
  assign n37682 = n37681 ^ n18349 ^ x9 ;
  assign n37683 = n10694 | n18703 ;
  assign n37684 = n37683 ^ n4538 ^ 1'b0 ;
  assign n37685 = ( n5664 & n12057 ) | ( n5664 & ~n19364 ) | ( n12057 & ~n19364 ) ;
  assign n37686 = ( n2868 & n12762 ) | ( n2868 & n35544 ) | ( n12762 & n35544 ) ;
  assign n37687 = ( ~n37073 & n37685 ) | ( ~n37073 & n37686 ) | ( n37685 & n37686 ) ;
  assign n37688 = n37687 ^ n11021 ^ 1'b0 ;
  assign n37689 = ( n22599 & n26193 ) | ( n22599 & ~n37688 ) | ( n26193 & ~n37688 ) ;
  assign n37693 = ( n2318 & n18176 ) | ( n2318 & n25870 ) | ( n18176 & n25870 ) ;
  assign n37690 = n14057 ^ n5172 ^ n2306 ;
  assign n37691 = ( n5962 & n20995 ) | ( n5962 & ~n33724 ) | ( n20995 & ~n33724 ) ;
  assign n37692 = ( n2740 & ~n37690 ) | ( n2740 & n37691 ) | ( ~n37690 & n37691 ) ;
  assign n37694 = n37693 ^ n37692 ^ n697 ;
  assign n37695 = n12488 ^ n10007 ^ 1'b0 ;
  assign n37696 = n1497 | n37695 ;
  assign n37697 = ( ~n12526 & n18576 ) | ( ~n12526 & n37696 ) | ( n18576 & n37696 ) ;
  assign n37698 = n29974 ^ n4558 ^ 1'b0 ;
  assign n37699 = ( n1808 & n5720 ) | ( n1808 & ~n37698 ) | ( n5720 & ~n37698 ) ;
  assign n37700 = n3446 | n17169 ;
  assign n37701 = ~n11355 & n11720 ;
  assign n37702 = n37701 ^ n22312 ^ 1'b0 ;
  assign n37703 = ( n2471 & n4030 ) | ( n2471 & n10090 ) | ( n4030 & n10090 ) ;
  assign n37704 = n37703 ^ n8199 ^ n5673 ;
  assign n37705 = ( ~n1061 & n12848 ) | ( ~n1061 & n37704 ) | ( n12848 & n37704 ) ;
  assign n37706 = n10224 & ~n23151 ;
  assign n37707 = n21477 & ~n37706 ;
  assign n37708 = n1961 ^ n396 ^ 1'b0 ;
  assign n37709 = n6281 & ~n37708 ;
  assign n37710 = ( n19314 & ~n33846 ) | ( n19314 & n37709 ) | ( ~n33846 & n37709 ) ;
  assign n37711 = ( ~n37705 & n37707 ) | ( ~n37705 & n37710 ) | ( n37707 & n37710 ) ;
  assign n37712 = n4792 ^ n3622 ^ n710 ;
  assign n37713 = n37712 ^ n30263 ^ n25415 ;
  assign n37714 = ( ~n12112 & n12762 ) | ( ~n12112 & n37638 ) | ( n12762 & n37638 ) ;
  assign n37715 = n7901 ^ n4373 ^ 1'b0 ;
  assign n37716 = ~n18544 & n37715 ;
  assign n37717 = ( ~n2778 & n3899 ) | ( ~n2778 & n33326 ) | ( n3899 & n33326 ) ;
  assign n37718 = n37717 ^ n19723 ^ n7235 ;
  assign n37719 = ~n19502 & n37718 ;
  assign n37720 = ~n23679 & n37719 ;
  assign n37721 = ~n20888 & n35082 ;
  assign n37722 = n25538 ^ n1925 ^ 1'b0 ;
  assign n37723 = ( n1840 & n5711 ) | ( n1840 & ~n34194 ) | ( n5711 & ~n34194 ) ;
  assign n37724 = n12259 | n37723 ;
  assign n37725 = n9787 & ~n37724 ;
  assign n37726 = n37722 & ~n37725 ;
  assign n37727 = n28535 & n37726 ;
  assign n37728 = ( n1463 & n7058 ) | ( n1463 & n37727 ) | ( n7058 & n37727 ) ;
  assign n37729 = n34470 ^ n24111 ^ n6430 ;
  assign n37730 = n4828 & n23571 ;
  assign n37731 = ~n21048 & n37730 ;
  assign n37732 = ~n14698 & n37731 ;
  assign n37733 = n37732 ^ n8824 ^ n2306 ;
  assign n37734 = n10196 | n19767 ;
  assign n37735 = ( ~n1037 & n18051 ) | ( ~n1037 & n37734 ) | ( n18051 & n37734 ) ;
  assign n37736 = n7240 & ~n12444 ;
  assign n37737 = n37736 ^ n8307 ^ 1'b0 ;
  assign n37738 = n25886 ^ n2560 ^ 1'b0 ;
  assign n37739 = n37737 & ~n37738 ;
  assign n37740 = ( n27175 & n31326 ) | ( n27175 & ~n37739 ) | ( n31326 & ~n37739 ) ;
  assign n37741 = n37740 ^ n12940 ^ n7440 ;
  assign n37742 = n20071 ^ n8940 ^ 1'b0 ;
  assign n37743 = ~n9035 & n18002 ;
  assign n37744 = ~n6939 & n37743 ;
  assign n37745 = n12341 ^ n9686 ^ n9512 ;
  assign n37746 = n9303 ^ n1278 ^ n729 ;
  assign n37747 = n37746 ^ n1146 ^ 1'b0 ;
  assign n37748 = ~n19139 & n37747 ;
  assign n37749 = n37745 & n37748 ;
  assign n37750 = n8811 & n35233 ;
  assign n37751 = ~n12108 & n37750 ;
  assign n37752 = ( n17792 & ~n18589 ) | ( n17792 & n20090 ) | ( ~n18589 & n20090 ) ;
  assign n37753 = ( n4241 & ~n6404 ) | ( n4241 & n17608 ) | ( ~n6404 & n17608 ) ;
  assign n37754 = n37753 ^ n8951 ^ x195 ;
  assign n37755 = n29961 ^ n11676 ^ 1'b0 ;
  assign n37756 = n14105 & ~n37755 ;
  assign n37757 = n25167 ^ n15182 ^ 1'b0 ;
  assign n37759 = n22613 ^ n21526 ^ 1'b0 ;
  assign n37758 = ~n6465 & n29451 ;
  assign n37760 = n37759 ^ n37758 ^ 1'b0 ;
  assign n37761 = n6785 ^ n1672 ^ n1144 ;
  assign n37762 = n37761 ^ n24271 ^ n905 ;
  assign n37763 = ( n899 & n14341 ) | ( n899 & ~n37762 ) | ( n14341 & ~n37762 ) ;
  assign n37764 = ( ~n32637 & n37760 ) | ( ~n32637 & n37763 ) | ( n37760 & n37763 ) ;
  assign n37766 = ~n4102 & n9611 ;
  assign n37767 = n37766 ^ n299 ^ 1'b0 ;
  assign n37765 = n598 & n20932 ;
  assign n37768 = n37767 ^ n37765 ^ 1'b0 ;
  assign n37769 = n2270 & n7026 ;
  assign n37770 = n37769 ^ n21328 ^ 1'b0 ;
  assign n37771 = n37770 ^ n37424 ^ n3958 ;
  assign n37772 = n12430 & ~n37771 ;
  assign n37773 = n37772 ^ n4735 ^ 1'b0 ;
  assign n37774 = n37768 | n37773 ;
  assign n37775 = n8047 | n22655 ;
  assign n37776 = ( n9253 & n22922 ) | ( n9253 & n36789 ) | ( n22922 & n36789 ) ;
  assign n37777 = n25886 & ~n37776 ;
  assign n37778 = ( n25045 & ~n30172 ) | ( n25045 & n37777 ) | ( ~n30172 & n37777 ) ;
  assign n37779 = ( ~n7671 & n25244 ) | ( ~n7671 & n29553 ) | ( n25244 & n29553 ) ;
  assign n37780 = n37779 ^ n20415 ^ n19785 ;
  assign n37781 = n474 & ~n3429 ;
  assign n37782 = ( n21018 & n21817 ) | ( n21018 & n37781 ) | ( n21817 & n37781 ) ;
  assign n37783 = n37722 ^ n8544 ^ 1'b0 ;
  assign n37784 = n6944 ^ n6216 ^ n3674 ;
  assign n37785 = ( ~n2406 & n6444 ) | ( ~n2406 & n37784 ) | ( n6444 & n37784 ) ;
  assign n37786 = n37785 ^ n35089 ^ 1'b0 ;
  assign n37787 = ~n31692 & n37786 ;
  assign n37788 = n33723 ^ n24343 ^ 1'b0 ;
  assign n37789 = n37788 ^ n28176 ^ n12303 ;
  assign n37790 = n36738 ^ n16573 ^ n14341 ;
  assign n37791 = n24602 & ~n37790 ;
  assign n37792 = ~n37789 & n37791 ;
  assign n37793 = n16382 ^ n7374 ^ 1'b0 ;
  assign n37794 = n21245 ^ n6685 ^ 1'b0 ;
  assign n37795 = n37793 | n37794 ;
  assign n37796 = ( n30065 & ~n36421 ) | ( n30065 & n37795 ) | ( ~n36421 & n37795 ) ;
  assign n37797 = n36753 ^ n16152 ^ n14112 ;
  assign n37798 = n15065 & n17563 ;
  assign n37799 = ( n27790 & n37797 ) | ( n27790 & n37798 ) | ( n37797 & n37798 ) ;
  assign n37800 = n37799 ^ n34107 ^ n4421 ;
  assign n37801 = n37800 ^ n26522 ^ 1'b0 ;
  assign n37803 = ( n8703 & n9336 ) | ( n8703 & ~n13427 ) | ( n9336 & ~n13427 ) ;
  assign n37802 = n36392 ^ n15133 ^ n6317 ;
  assign n37804 = n37803 ^ n37802 ^ 1'b0 ;
  assign n37805 = n15173 ^ n8472 ^ 1'b0 ;
  assign n37806 = n37805 ^ n25228 ^ n1475 ;
  assign n37807 = n37806 ^ n1554 ^ 1'b0 ;
  assign n37808 = n37804 & n37807 ;
  assign n37809 = ( n1472 & n6639 ) | ( n1472 & ~n9067 ) | ( n6639 & ~n9067 ) ;
  assign n37810 = ( n735 & n9493 ) | ( n735 & n37809 ) | ( n9493 & n37809 ) ;
  assign n37811 = ~n33547 & n37810 ;
  assign n37812 = ( n12471 & n37808 ) | ( n12471 & ~n37811 ) | ( n37808 & ~n37811 ) ;
  assign n37813 = n12328 ^ n1197 ^ 1'b0 ;
  assign n37814 = n20351 ^ n18883 ^ 1'b0 ;
  assign n37815 = n3136 & ~n37814 ;
  assign n37816 = ( n4502 & ~n4687 ) | ( n4502 & n25342 ) | ( ~n4687 & n25342 ) ;
  assign n37817 = n37816 ^ n7171 ^ n4247 ;
  assign n37818 = n12089 ^ n2313 ^ 1'b0 ;
  assign n37819 = n37817 & n37818 ;
  assign n37820 = n11126 ^ n1175 ^ 1'b0 ;
  assign n37821 = ~n16145 & n37820 ;
  assign n37822 = ~n12326 & n37821 ;
  assign n37823 = n27793 & n37822 ;
  assign n37824 = n2296 | n19219 ;
  assign n37825 = n37824 ^ n18369 ^ n14246 ;
  assign n37826 = n34493 ^ n18612 ^ n2341 ;
  assign n37827 = ( n713 & ~n7321 ) | ( n713 & n17037 ) | ( ~n7321 & n17037 ) ;
  assign n37828 = n37827 ^ n7732 ^ n639 ;
  assign n37829 = ~n21693 & n37828 ;
  assign n37830 = n28881 ^ n5392 ^ 1'b0 ;
  assign n37831 = n3412 & ~n37830 ;
  assign n37832 = n26206 ^ n6653 ^ 1'b0 ;
  assign n37833 = n37831 & ~n37832 ;
  assign n37834 = n37833 ^ n36422 ^ n8760 ;
  assign n37835 = n28752 ^ n24509 ^ 1'b0 ;
  assign n37836 = ~n3820 & n36278 ;
  assign n37837 = n37836 ^ n22344 ^ 1'b0 ;
  assign n37838 = n2961 & n14715 ;
  assign n37839 = ~n10074 & n37838 ;
  assign n37840 = n37839 ^ n2687 ^ 1'b0 ;
  assign n37841 = n24799 ^ n10415 ^ n5294 ;
  assign n37842 = n37841 ^ n27299 ^ n10490 ;
  assign n37843 = ( n302 & ~n21908 ) | ( n302 & n32827 ) | ( ~n21908 & n32827 ) ;
  assign n37845 = ( n555 & ~n6673 ) | ( n555 & n29104 ) | ( ~n6673 & n29104 ) ;
  assign n37844 = n13957 | n31455 ;
  assign n37846 = n37845 ^ n37844 ^ n26951 ;
  assign n37847 = n17987 ^ n1360 ^ 1'b0 ;
  assign n37848 = ~n6146 & n37847 ;
  assign n37850 = n2221 & ~n12952 ;
  assign n37851 = n37850 ^ n15635 ^ 1'b0 ;
  assign n37849 = n12396 & n12680 ;
  assign n37852 = n37851 ^ n37849 ^ 1'b0 ;
  assign n37853 = n16739 & n32751 ;
  assign n37854 = ~n37852 & n37853 ;
  assign n37864 = n24845 ^ n20643 ^ 1'b0 ;
  assign n37858 = n5761 & n11072 ;
  assign n37859 = n37858 ^ n16900 ^ 1'b0 ;
  assign n37860 = ~n35861 & n37859 ;
  assign n37861 = ( n3268 & n19983 ) | ( n3268 & n37860 ) | ( n19983 & n37860 ) ;
  assign n37862 = ~n25869 & n37861 ;
  assign n37863 = n1844 & n37862 ;
  assign n37855 = n33761 ^ n24291 ^ n5323 ;
  assign n37856 = n37855 ^ n6621 ^ 1'b0 ;
  assign n37857 = n24440 & n37856 ;
  assign n37865 = n37864 ^ n37863 ^ n37857 ;
  assign n37866 = ( n2480 & n13666 ) | ( n2480 & ~n19210 ) | ( n13666 & ~n19210 ) ;
  assign n37867 = n3897 & n8799 ;
  assign n37868 = n37867 ^ n34242 ^ n23879 ;
  assign n37869 = n37868 ^ n30153 ^ n11073 ;
  assign n37870 = n30137 ^ n19156 ^ n14515 ;
  assign n37871 = ( n5863 & n6626 ) | ( n5863 & ~n6757 ) | ( n6626 & ~n6757 ) ;
  assign n37872 = n37871 ^ n14651 ^ n339 ;
  assign n37873 = ~n13797 & n37872 ;
  assign n37876 = ~n5913 & n25221 ;
  assign n37877 = n12632 & n37876 ;
  assign n37878 = ~n16588 & n35579 ;
  assign n37879 = n37877 & n37878 ;
  assign n37874 = n5380 | n15537 ;
  assign n37875 = ~n6664 & n37874 ;
  assign n37880 = n37879 ^ n37875 ^ 1'b0 ;
  assign n37881 = ( ~n2265 & n17150 ) | ( ~n2265 & n32874 ) | ( n17150 & n32874 ) ;
  assign n37882 = ( ~n12663 & n33986 ) | ( ~n12663 & n37881 ) | ( n33986 & n37881 ) ;
  assign n37883 = x223 & n14110 ;
  assign n37884 = n37883 ^ n3306 ^ 1'b0 ;
  assign n37885 = n37884 ^ n29719 ^ n1368 ;
  assign n37886 = n8167 & n37885 ;
  assign n37887 = n8749 ^ n5111 ^ 1'b0 ;
  assign n37888 = ~n16692 & n37887 ;
  assign n37889 = ( n8494 & n31630 ) | ( n8494 & ~n37888 ) | ( n31630 & ~n37888 ) ;
  assign n37890 = n11808 | n37889 ;
  assign n37891 = n1435 & ~n37890 ;
  assign n37892 = ( n7303 & n8543 ) | ( n7303 & n28960 ) | ( n8543 & n28960 ) ;
  assign n37893 = n37892 ^ n4721 ^ n833 ;
  assign n37895 = n29444 ^ n16355 ^ 1'b0 ;
  assign n37894 = n33585 ^ n18718 ^ n15204 ;
  assign n37896 = n37895 ^ n37894 ^ n1316 ;
  assign n37897 = ( ~n1116 & n13970 ) | ( ~n1116 & n37896 ) | ( n13970 & n37896 ) ;
  assign n37898 = n37897 ^ n27503 ^ 1'b0 ;
  assign n37899 = n5124 ^ n2717 ^ n526 ;
  assign n37900 = n3901 & ~n11489 ;
  assign n37901 = n6097 & n37900 ;
  assign n37902 = ( ~n20865 & n37899 ) | ( ~n20865 & n37901 ) | ( n37899 & n37901 ) ;
  assign n37903 = ~n18064 & n22242 ;
  assign n37904 = n9853 ^ n4960 ^ n648 ;
  assign n37905 = ~n7659 & n33905 ;
  assign n37906 = ( ~n10212 & n37904 ) | ( ~n10212 & n37905 ) | ( n37904 & n37905 ) ;
  assign n37907 = n27921 ^ n3449 ^ n2358 ;
  assign n37908 = n8285 & ~n37907 ;
  assign n37909 = ~n15043 & n37908 ;
  assign n37910 = n4851 & ~n37909 ;
  assign n37911 = ~n13876 & n37910 ;
  assign n37912 = n37329 | n37911 ;
  assign n37913 = n37906 | n37912 ;
  assign n37914 = n20256 ^ n1756 ^ 1'b0 ;
  assign n37915 = n37913 & n37914 ;
  assign n37916 = n34251 ^ n31368 ^ n30942 ;
  assign n37917 = n37916 ^ n27543 ^ n11855 ;
  assign n37918 = ( n13194 & ~n31972 ) | ( n13194 & n37917 ) | ( ~n31972 & n37917 ) ;
  assign n37919 = ( ~n15318 & n15674 ) | ( ~n15318 & n27758 ) | ( n15674 & n27758 ) ;
  assign n37920 = n5034 & ~n33872 ;
  assign n37921 = ~n2947 & n37920 ;
  assign n37922 = ( n1852 & n3418 ) | ( n1852 & ~n6210 ) | ( n3418 & ~n6210 ) ;
  assign n37923 = n37922 ^ n26119 ^ n1805 ;
  assign n37924 = ( n9011 & n33880 ) | ( n9011 & n37923 ) | ( n33880 & n37923 ) ;
  assign n37925 = n5480 & ~n37924 ;
  assign n37926 = ~n17844 & n37925 ;
  assign n37927 = ( ~n5632 & n37921 ) | ( ~n5632 & n37926 ) | ( n37921 & n37926 ) ;
  assign n37928 = ( n5165 & ~n37919 ) | ( n5165 & n37927 ) | ( ~n37919 & n37927 ) ;
  assign n37929 = ~n453 & n7671 ;
  assign n37930 = ~n12345 & n37929 ;
  assign n37931 = n37930 ^ n11904 ^ n1939 ;
  assign n37932 = n28029 ^ n3327 ^ 1'b0 ;
  assign n37933 = ( n19056 & n32093 ) | ( n19056 & ~n37932 ) | ( n32093 & ~n37932 ) ;
  assign n37934 = ( n15526 & ~n37931 ) | ( n15526 & n37933 ) | ( ~n37931 & n37933 ) ;
  assign n37935 = n6676 | n36390 ;
  assign n37936 = n4468 & ~n37935 ;
  assign n37937 = n30067 ^ n28536 ^ n2806 ;
  assign n37938 = n10516 ^ n8882 ^ 1'b0 ;
  assign n37939 = n37938 ^ n23479 ^ n10751 ;
  assign n37940 = n37939 ^ n34840 ^ n18212 ;
  assign n37941 = n7480 | n18772 ;
  assign n37942 = n20025 ^ n12930 ^ n6972 ;
  assign n37943 = n37942 ^ n25071 ^ n14641 ;
  assign n37944 = ( x112 & ~n37941 ) | ( x112 & n37943 ) | ( ~n37941 & n37943 ) ;
  assign n37945 = n24908 ^ n18772 ^ 1'b0 ;
  assign n37946 = n32350 ^ n15483 ^ n13221 ;
  assign n37947 = ( ~n3898 & n7196 ) | ( ~n3898 & n37946 ) | ( n7196 & n37946 ) ;
  assign n37948 = n31277 ^ n20851 ^ n14523 ;
  assign n37949 = n15577 ^ n3802 ^ 1'b0 ;
  assign n37950 = ~n574 & n37949 ;
  assign n37951 = ~n3051 & n26554 ;
  assign n37954 = ~n729 & n5612 ;
  assign n37955 = n37954 ^ n3811 ^ 1'b0 ;
  assign n37952 = ( n26480 & n27768 ) | ( n26480 & ~n30288 ) | ( n27768 & ~n30288 ) ;
  assign n37953 = ( ~n4104 & n26653 ) | ( ~n4104 & n37952 ) | ( n26653 & n37952 ) ;
  assign n37956 = n37955 ^ n37953 ^ 1'b0 ;
  assign n37957 = n29702 | n35986 ;
  assign n37958 = n14063 | n37957 ;
  assign n37959 = n21179 ^ n4368 ^ n1995 ;
  assign n37960 = n34968 ^ n13050 ^ n10705 ;
  assign n37963 = n5516 ^ n5264 ^ n2096 ;
  assign n37961 = n26987 ^ n1385 ^ n527 ;
  assign n37962 = n37961 ^ n6131 ^ 1'b0 ;
  assign n37964 = n37963 ^ n37962 ^ n36155 ;
  assign n37965 = n23408 ^ n358 ^ 1'b0 ;
  assign n37966 = n33041 & n37965 ;
  assign n37967 = n37966 ^ n22039 ^ 1'b0 ;
  assign n37968 = ( n8914 & ~n15583 ) | ( n8914 & n30875 ) | ( ~n15583 & n30875 ) ;
  assign n37969 = n11964 ^ n2741 ^ n905 ;
  assign n37970 = n6965 | n18600 ;
  assign n37971 = n37969 & ~n37970 ;
  assign n37972 = n23609 ^ n8826 ^ 1'b0 ;
  assign n37973 = n28770 & ~n37972 ;
  assign n37974 = ~n2472 & n5146 ;
  assign n37975 = n27949 & n37974 ;
  assign n37976 = ~n15157 & n37975 ;
  assign n37977 = ( x135 & ~n576 ) | ( x135 & n3947 ) | ( ~n576 & n3947 ) ;
  assign n37978 = n37977 ^ n26912 ^ n23150 ;
  assign n37979 = n37978 ^ n10924 ^ 1'b0 ;
  assign n37980 = n10958 ^ n10250 ^ n3284 ;
  assign n37981 = ( n360 & n37979 ) | ( n360 & n37980 ) | ( n37979 & n37980 ) ;
  assign n37982 = n28293 & ~n28815 ;
  assign n37983 = n8841 ^ n7968 ^ 1'b0 ;
  assign n37984 = n8099 | n37983 ;
  assign n37985 = ( n2848 & n23332 ) | ( n2848 & ~n37984 ) | ( n23332 & ~n37984 ) ;
  assign n37986 = n5293 ^ n2539 ^ 1'b0 ;
  assign n37987 = n30065 & n37986 ;
  assign n37988 = n37987 ^ n32036 ^ x65 ;
  assign n37989 = n32504 | n37988 ;
  assign n37990 = n37989 ^ n14591 ^ 1'b0 ;
  assign n37991 = n12101 & ~n18496 ;
  assign n37992 = n37991 ^ n5763 ^ 1'b0 ;
  assign n37993 = n13462 ^ n8166 ^ 1'b0 ;
  assign n37994 = n35223 | n37993 ;
  assign n37995 = n18917 ^ n14763 ^ n10885 ;
  assign n37996 = n37995 ^ n24161 ^ n11170 ;
  assign n37997 = ( n12409 & n18275 ) | ( n12409 & n34186 ) | ( n18275 & n34186 ) ;
  assign n37998 = n4404 ^ n994 ^ 1'b0 ;
  assign n37999 = n7698 | n37998 ;
  assign n38000 = n37999 ^ n17955 ^ 1'b0 ;
  assign n38001 = n15524 | n38000 ;
  assign n38002 = n10565 | n38001 ;
  assign n38003 = n2311 & n23234 ;
  assign n38004 = n12391 ^ n4851 ^ 1'b0 ;
  assign n38005 = ~n1154 & n38004 ;
  assign n38006 = n38005 ^ n18485 ^ 1'b0 ;
  assign n38007 = n12930 | n38006 ;
  assign n38008 = n32700 ^ n7359 ^ n661 ;
  assign n38009 = ( n17686 & n27432 ) | ( n17686 & ~n38008 ) | ( n27432 & ~n38008 ) ;
  assign n38010 = ( n5920 & ~n20834 ) | ( n5920 & n28193 ) | ( ~n20834 & n28193 ) ;
  assign n38011 = n23584 ^ n22392 ^ n9408 ;
  assign n38012 = n6340 & n8851 ;
  assign n38013 = n38012 ^ n37568 ^ 1'b0 ;
  assign n38014 = ( n1383 & n2632 ) | ( n1383 & ~n11075 ) | ( n2632 & ~n11075 ) ;
  assign n38015 = n13622 ^ n2825 ^ 1'b0 ;
  assign n38016 = ~n38014 & n38015 ;
  assign n38017 = n1936 & ~n34327 ;
  assign n38018 = n38017 ^ n4883 ^ 1'b0 ;
  assign n38019 = n38018 ^ n30538 ^ n11727 ;
  assign n38020 = n10656 ^ n3312 ^ 1'b0 ;
  assign n38021 = ( ~n12084 & n13145 ) | ( ~n12084 & n38020 ) | ( n13145 & n38020 ) ;
  assign n38023 = n37017 ^ n15356 ^ n1209 ;
  assign n38022 = n25433 ^ n11060 ^ n3369 ;
  assign n38024 = n38023 ^ n38022 ^ n25646 ;
  assign n38025 = n11663 ^ n5589 ^ 1'b0 ;
  assign n38026 = n12850 ^ n10358 ^ n3496 ;
  assign n38027 = n38026 ^ n16411 ^ n11332 ;
  assign n38028 = ( ~n5824 & n28536 ) | ( ~n5824 & n38027 ) | ( n28536 & n38027 ) ;
  assign n38029 = ( n36337 & ~n38025 ) | ( n36337 & n38028 ) | ( ~n38025 & n38028 ) ;
  assign n38030 = n10726 ^ n8247 ^ 1'b0 ;
  assign n38031 = n3793 & n38030 ;
  assign n38032 = n38031 ^ n18428 ^ n4527 ;
  assign n38033 = n29648 ^ n28821 ^ n9334 ;
  assign n38034 = ( n7637 & ~n13523 ) | ( n7637 & n16518 ) | ( ~n13523 & n16518 ) ;
  assign n38035 = n38034 ^ n37248 ^ n14474 ;
  assign n38036 = n38035 ^ n27599 ^ n14892 ;
  assign n38037 = ( n13267 & ~n24872 ) | ( n13267 & n37831 ) | ( ~n24872 & n37831 ) ;
  assign n38038 = n38037 ^ n18174 ^ n9474 ;
  assign n38039 = ( n8322 & ~n38036 ) | ( n8322 & n38038 ) | ( ~n38036 & n38038 ) ;
  assign n38040 = n31213 ^ n1737 ^ n1552 ;
  assign n38041 = n24151 ^ n19556 ^ n13498 ;
  assign n38042 = n24311 ^ n23995 ^ n21725 ;
  assign n38043 = ( n2164 & n20543 ) | ( n2164 & ~n38042 ) | ( n20543 & ~n38042 ) ;
  assign n38044 = ( n7153 & ~n28752 ) | ( n7153 & n38043 ) | ( ~n28752 & n38043 ) ;
  assign n38045 = n9677 ^ n1580 ^ 1'b0 ;
  assign n38046 = n8378 & n38045 ;
  assign n38047 = n7727 & n38046 ;
  assign n38048 = n38047 ^ n21986 ^ n17899 ;
  assign n38049 = n18801 | n28519 ;
  assign n38050 = ( n2914 & ~n9066 ) | ( n2914 & n25665 ) | ( ~n9066 & n25665 ) ;
  assign n38051 = n7635 ^ n358 ^ 1'b0 ;
  assign n38052 = ( n12949 & ~n15678 ) | ( n12949 & n38051 ) | ( ~n15678 & n38051 ) ;
  assign n38053 = n14366 ^ n5419 ^ 1'b0 ;
  assign n38054 = ( ~n16220 & n21665 ) | ( ~n16220 & n38053 ) | ( n21665 & n38053 ) ;
  assign n38055 = ( n12968 & n26027 ) | ( n12968 & ~n27730 ) | ( n26027 & ~n27730 ) ;
  assign n38056 = n27673 ^ n13595 ^ 1'b0 ;
  assign n38057 = n26307 ^ n21789 ^ n2004 ;
  assign n38058 = ( ~n22337 & n38056 ) | ( ~n22337 & n38057 ) | ( n38056 & n38057 ) ;
  assign n38059 = ( n1870 & n24184 ) | ( n1870 & n37583 ) | ( n24184 & n37583 ) ;
  assign n38060 = n38059 ^ n13854 ^ 1'b0 ;
  assign n38061 = n28247 ^ n12440 ^ n3811 ;
  assign n38062 = ( n21113 & ~n29347 ) | ( n21113 & n38061 ) | ( ~n29347 & n38061 ) ;
  assign n38063 = ( n3763 & ~n6052 ) | ( n3763 & n18986 ) | ( ~n6052 & n18986 ) ;
  assign n38064 = ( ~n29612 & n38062 ) | ( ~n29612 & n38063 ) | ( n38062 & n38063 ) ;
  assign n38065 = n1651 | n35493 ;
  assign n38066 = ~n7267 & n30990 ;
  assign n38067 = n25795 & n38066 ;
  assign n38068 = n2648 & ~n15059 ;
  assign n38069 = n38068 ^ n7393 ^ 1'b0 ;
  assign n38070 = ( n12065 & n31220 ) | ( n12065 & n38069 ) | ( n31220 & n38069 ) ;
  assign n38071 = n29457 ^ n9921 ^ n9371 ;
  assign n38072 = n33532 ^ n21259 ^ 1'b0 ;
  assign n38073 = n4890 | n38072 ;
  assign n38074 = n27632 ^ x235 ^ 1'b0 ;
  assign n38075 = n23712 & ~n38074 ;
  assign n38076 = n9947 ^ n1331 ^ 1'b0 ;
  assign n38077 = ~n12842 & n38076 ;
  assign n38078 = n38077 ^ n13594 ^ 1'b0 ;
  assign n38079 = n38075 & n38078 ;
  assign n38080 = n7903 ^ n5607 ^ n2025 ;
  assign n38081 = ~n35280 & n38080 ;
  assign n38082 = n18013 | n22267 ;
  assign n38083 = n36505 ^ n29348 ^ 1'b0 ;
  assign n38084 = ( n12212 & n24941 ) | ( n12212 & ~n33955 ) | ( n24941 & ~n33955 ) ;
  assign n38090 = n925 & ~n13052 ;
  assign n38086 = n18794 ^ n5970 ^ 1'b0 ;
  assign n38087 = n14397 | n38086 ;
  assign n38088 = n38087 ^ n770 ^ 1'b0 ;
  assign n38085 = ~n7647 & n13985 ;
  assign n38089 = n38088 ^ n38085 ^ n1337 ;
  assign n38091 = n38090 ^ n38089 ^ n35033 ;
  assign n38092 = n7349 & ~n10093 ;
  assign n38093 = n38092 ^ n15753 ^ n4077 ;
  assign n38094 = n33620 ^ n29183 ^ n9931 ;
  assign n38095 = n38094 ^ n28580 ^ 1'b0 ;
  assign n38096 = ( n6404 & ~n9146 ) | ( n6404 & n19928 ) | ( ~n9146 & n19928 ) ;
  assign n38097 = ( n20585 & n38095 ) | ( n20585 & ~n38096 ) | ( n38095 & ~n38096 ) ;
  assign n38098 = ~n956 & n6304 ;
  assign n38099 = n3894 & n38098 ;
  assign n38100 = n3969 ^ n1206 ^ 1'b0 ;
  assign n38101 = ~n598 & n38100 ;
  assign n38102 = n36754 & n38101 ;
  assign n38103 = n38102 ^ n11870 ^ 1'b0 ;
  assign n38104 = n7768 & n11515 ;
  assign n38105 = ~n3398 & n38104 ;
  assign n38106 = n31925 ^ n20088 ^ n5534 ;
  assign n38107 = n15891 ^ n5975 ^ 1'b0 ;
  assign n38108 = ( n10990 & n17124 ) | ( n10990 & n38107 ) | ( n17124 & n38107 ) ;
  assign n38109 = ( ~n18119 & n18257 ) | ( ~n18119 & n38108 ) | ( n18257 & n38108 ) ;
  assign n38110 = n38109 ^ n7168 ^ n390 ;
  assign n38111 = n13528 ^ n4885 ^ 1'b0 ;
  assign n38112 = ( n626 & n13097 ) | ( n626 & n19502 ) | ( n13097 & n19502 ) ;
  assign n38113 = ( n7613 & ~n38111 ) | ( n7613 & n38112 ) | ( ~n38111 & n38112 ) ;
  assign n38114 = n8885 & ~n26748 ;
  assign n38115 = n16076 & n38114 ;
  assign n38116 = n38115 ^ n33828 ^ 1'b0 ;
  assign n38119 = ( n463 & ~n5401 ) | ( n463 & n7273 ) | ( ~n5401 & n7273 ) ;
  assign n38118 = n21761 ^ n3384 ^ 1'b0 ;
  assign n38120 = n38119 ^ n38118 ^ n19497 ;
  assign n38117 = ~n13047 & n15475 ;
  assign n38121 = n38120 ^ n38117 ^ n26480 ;
  assign n38122 = n18930 ^ n18816 ^ 1'b0 ;
  assign n38123 = n16521 & ~n38122 ;
  assign n38124 = n24270 ^ n6783 ^ n1242 ;
  assign n38125 = ~n5994 & n24245 ;
  assign n38126 = ( n5655 & n7665 ) | ( n5655 & n8019 ) | ( n7665 & n8019 ) ;
  assign n38127 = ( n10725 & ~n10765 ) | ( n10725 & n38126 ) | ( ~n10765 & n38126 ) ;
  assign n38130 = n27036 ^ n14889 ^ n1828 ;
  assign n38128 = n19396 | n29935 ;
  assign n38129 = n13925 & ~n38128 ;
  assign n38131 = n38130 ^ n38129 ^ 1'b0 ;
  assign n38132 = n10987 | n38131 ;
  assign n38133 = n14745 ^ n5921 ^ 1'b0 ;
  assign n38134 = ~n38132 & n38133 ;
  assign n38135 = n35840 ^ n34814 ^ n6143 ;
  assign n38136 = n38135 ^ n28821 ^ 1'b0 ;
  assign n38137 = n14321 | n38136 ;
  assign n38138 = n38137 ^ n13462 ^ 1'b0 ;
  assign n38139 = ( n21102 & n28760 ) | ( n21102 & n38138 ) | ( n28760 & n38138 ) ;
  assign n38140 = ( ~n23147 & n23739 ) | ( ~n23147 & n29298 ) | ( n23739 & n29298 ) ;
  assign n38141 = ( n1519 & ~n16405 ) | ( n1519 & n22534 ) | ( ~n16405 & n22534 ) ;
  assign n38142 = n38141 ^ n22615 ^ 1'b0 ;
  assign n38143 = n5276 ^ n3039 ^ x203 ;
  assign n38144 = n21423 ^ n8481 ^ 1'b0 ;
  assign n38145 = ~n24898 & n38144 ;
  assign n38146 = n38145 ^ n28079 ^ 1'b0 ;
  assign n38147 = n38143 & n38146 ;
  assign n38148 = n30288 ^ n5459 ^ 1'b0 ;
  assign n38149 = ( ~n6796 & n8367 ) | ( ~n6796 & n38148 ) | ( n8367 & n38148 ) ;
  assign n38150 = ( n16326 & n22119 ) | ( n16326 & n38149 ) | ( n22119 & n38149 ) ;
  assign n38151 = ( n13298 & ~n25023 ) | ( n13298 & n38150 ) | ( ~n25023 & n38150 ) ;
  assign n38152 = n8611 ^ n6346 ^ 1'b0 ;
  assign n38153 = ( ~n408 & n4241 ) | ( ~n408 & n11696 ) | ( n4241 & n11696 ) ;
  assign n38154 = n38153 ^ n35025 ^ n15078 ;
  assign n38155 = ( n4213 & ~n29087 ) | ( n4213 & n38154 ) | ( ~n29087 & n38154 ) ;
  assign n38156 = ~n21489 & n38155 ;
  assign n38157 = ( n3096 & n24176 ) | ( n3096 & n26361 ) | ( n24176 & n26361 ) ;
  assign n38158 = n4692 ^ n4248 ^ 1'b0 ;
  assign n38159 = ( n3229 & ~n8701 ) | ( n3229 & n34204 ) | ( ~n8701 & n34204 ) ;
  assign n38160 = n3180 & ~n38159 ;
  assign n38161 = n38158 & n38160 ;
  assign n38162 = n23335 ^ x212 ^ 1'b0 ;
  assign n38163 = n6377 & ~n38162 ;
  assign n38164 = n32875 ^ n27653 ^ x44 ;
  assign n38165 = n20071 & ~n28360 ;
  assign n38166 = n19425 & n38165 ;
  assign n38167 = n33773 & ~n38166 ;
  assign n38168 = ( n7647 & n20876 ) | ( n7647 & n26358 ) | ( n20876 & n26358 ) ;
  assign n38169 = n3214 & ~n9653 ;
  assign n38170 = n38169 ^ n6523 ^ 1'b0 ;
  assign n38171 = n38170 ^ n23397 ^ n8973 ;
  assign n38172 = ~n7785 & n28051 ;
  assign n38173 = n38171 & n38172 ;
  assign n38174 = n21934 | n24138 ;
  assign n38175 = n32572 & ~n38174 ;
  assign n38176 = ( n7525 & n16866 ) | ( n7525 & n38175 ) | ( n16866 & n38175 ) ;
  assign n38177 = n12586 | n38176 ;
  assign n38178 = n10625 | n29268 ;
  assign n38179 = n12876 ^ n10650 ^ 1'b0 ;
  assign n38180 = ~n27059 & n38179 ;
  assign n38181 = n26208 ^ n20330 ^ 1'b0 ;
  assign n38182 = n38180 & n38181 ;
  assign n38183 = ~n3966 & n8340 ;
  assign n38184 = ~n17383 & n38183 ;
  assign n38185 = ( n1078 & n18044 ) | ( n1078 & ~n21870 ) | ( n18044 & ~n21870 ) ;
  assign n38186 = n38185 ^ n22304 ^ 1'b0 ;
  assign n38187 = n10268 ^ n6853 ^ n2785 ;
  assign n38188 = ( ~n12717 & n22029 ) | ( ~n12717 & n38187 ) | ( n22029 & n38187 ) ;
  assign n38189 = n25405 ^ n10618 ^ n9818 ;
  assign n38190 = ( n5735 & ~n18684 ) | ( n5735 & n38189 ) | ( ~n18684 & n38189 ) ;
  assign n38191 = n16373 ^ n12302 ^ n11597 ;
  assign n38192 = ( ~x29 & n6700 ) | ( ~x29 & n24245 ) | ( n6700 & n24245 ) ;
  assign n38193 = ~n8499 & n21705 ;
  assign n38194 = n38193 ^ x111 ^ 1'b0 ;
  assign n38195 = n21085 ^ n21054 ^ n20633 ;
  assign n38196 = ( n1820 & n8112 ) | ( n1820 & ~n12820 ) | ( n8112 & ~n12820 ) ;
  assign n38197 = ( n5797 & n7102 ) | ( n5797 & n38196 ) | ( n7102 & n38196 ) ;
  assign n38198 = ( n7346 & ~n38195 ) | ( n7346 & n38197 ) | ( ~n38195 & n38197 ) ;
  assign n38199 = n38194 | n38198 ;
  assign n38200 = n38199 ^ n12450 ^ 1'b0 ;
  assign n38201 = n838 & ~n22382 ;
  assign n38202 = ( ~n5566 & n8643 ) | ( ~n5566 & n38201 ) | ( n8643 & n38201 ) ;
  assign n38203 = ( n34336 & n38200 ) | ( n34336 & n38202 ) | ( n38200 & n38202 ) ;
  assign n38204 = ( n7057 & ~n16646 ) | ( n7057 & n17054 ) | ( ~n16646 & n17054 ) ;
  assign n38205 = n38204 ^ n24987 ^ n987 ;
  assign n38206 = ( ~n16233 & n22985 ) | ( ~n16233 & n36056 ) | ( n22985 & n36056 ) ;
  assign n38207 = ( n4749 & n14263 ) | ( n4749 & n23081 ) | ( n14263 & n23081 ) ;
  assign n38208 = ~n8532 & n34785 ;
  assign n38209 = n38208 ^ n831 ^ 1'b0 ;
  assign n38210 = n38209 ^ n11851 ^ n11016 ;
  assign n38211 = ( n9707 & ~n19121 ) | ( n9707 & n23871 ) | ( ~n19121 & n23871 ) ;
  assign n38212 = n17985 ^ n16238 ^ n12193 ;
  assign n38213 = n38212 ^ n12440 ^ 1'b0 ;
  assign n38214 = ( n3626 & n22326 ) | ( n3626 & n38213 ) | ( n22326 & n38213 ) ;
  assign n38215 = n3109 | n20931 ;
  assign n38216 = n38215 ^ n3800 ^ 1'b0 ;
  assign n38217 = n35141 ^ n13066 ^ 1'b0 ;
  assign n38218 = n2827 | n35783 ;
  assign n38219 = n14539 & ~n38218 ;
  assign n38220 = ( n10669 & n16661 ) | ( n10669 & n26846 ) | ( n16661 & n26846 ) ;
  assign n38221 = ( ~n8126 & n18086 ) | ( ~n8126 & n38220 ) | ( n18086 & n38220 ) ;
  assign n38222 = ( n38217 & n38219 ) | ( n38217 & ~n38221 ) | ( n38219 & ~n38221 ) ;
  assign n38223 = ( n37495 & n38216 ) | ( n37495 & n38222 ) | ( n38216 & n38222 ) ;
  assign n38225 = n7020 ^ n4194 ^ 1'b0 ;
  assign n38224 = ( n4181 & n7655 ) | ( n4181 & n10886 ) | ( n7655 & n10886 ) ;
  assign n38226 = n38225 ^ n38224 ^ n1003 ;
  assign n38227 = ~n12433 & n28874 ;
  assign n38228 = ( ~n5910 & n10123 ) | ( ~n5910 & n17872 ) | ( n10123 & n17872 ) ;
  assign n38229 = n38228 ^ n8072 ^ 1'b0 ;
  assign n38230 = n38227 | n38229 ;
  assign n38231 = ( n4169 & n38226 ) | ( n4169 & n38230 ) | ( n38226 & n38230 ) ;
  assign n38232 = n28678 ^ n17940 ^ 1'b0 ;
  assign n38233 = n15588 & ~n38232 ;
  assign n38234 = n1850 & ~n10359 ;
  assign n38235 = n16652 & n38234 ;
  assign n38236 = n12509 ^ n1424 ^ n984 ;
  assign n38237 = n38236 ^ n33138 ^ n13359 ;
  assign n38238 = n4904 & n15531 ;
  assign n38239 = n38238 ^ n15811 ^ 1'b0 ;
  assign n38240 = ( n5980 & n29071 ) | ( n5980 & n38239 ) | ( n29071 & n38239 ) ;
  assign n38241 = ( n17680 & ~n19114 ) | ( n17680 & n31173 ) | ( ~n19114 & n31173 ) ;
  assign n38242 = n38241 ^ n30486 ^ n12092 ;
  assign n38243 = n7823 & ~n38242 ;
  assign n38244 = n37458 ^ n27716 ^ n27091 ;
  assign n38245 = n20067 ^ n19439 ^ 1'b0 ;
  assign n38246 = n31878 | n38245 ;
  assign n38248 = n5402 ^ n2766 ^ n1143 ;
  assign n38247 = x34 & n16685 ;
  assign n38249 = n38248 ^ n38247 ^ 1'b0 ;
  assign n38250 = ( n17442 & ~n20071 ) | ( n17442 & n23564 ) | ( ~n20071 & n23564 ) ;
  assign n38251 = ( n7609 & n17218 ) | ( n7609 & ~n28035 ) | ( n17218 & ~n28035 ) ;
  assign n38252 = n16684 & n32943 ;
  assign n38253 = n38252 ^ n3406 ^ 1'b0 ;
  assign n38254 = n34848 ^ n33227 ^ n5511 ;
  assign n38255 = n6742 ^ n3495 ^ n1304 ;
  assign n38256 = n38255 ^ n35464 ^ n26624 ;
  assign n38257 = n33464 ^ n13618 ^ n4890 ;
  assign n38258 = ( x6 & n17388 ) | ( x6 & ~n38257 ) | ( n17388 & ~n38257 ) ;
  assign n38259 = n19829 ^ n9822 ^ n7652 ;
  assign n38260 = n27260 ^ n21742 ^ 1'b0 ;
  assign n38261 = n4299 | n38260 ;
  assign n38262 = n10499 | n38261 ;
  assign n38263 = n38259 & ~n38262 ;
  assign n38264 = n28236 ^ n3631 ^ 1'b0 ;
  assign n38265 = n5948 & n38264 ;
  assign n38267 = ( ~n2077 & n20833 ) | ( ~n2077 & n24794 ) | ( n20833 & n24794 ) ;
  assign n38266 = n4904 & n6292 ;
  assign n38268 = n38267 ^ n38266 ^ 1'b0 ;
  assign n38269 = n26998 | n37364 ;
  assign n38270 = n38269 ^ n15556 ^ n5705 ;
  assign n38271 = ( n17062 & n17548 ) | ( n17062 & ~n38270 ) | ( n17548 & ~n38270 ) ;
  assign n38272 = ( n8740 & n10312 ) | ( n8740 & n18384 ) | ( n10312 & n18384 ) ;
  assign n38273 = n38272 ^ n9749 ^ 1'b0 ;
  assign n38274 = n5000 ^ n351 ^ 1'b0 ;
  assign n38275 = n10912 ^ n9795 ^ 1'b0 ;
  assign n38276 = ( n8859 & n38274 ) | ( n8859 & ~n38275 ) | ( n38274 & ~n38275 ) ;
  assign n38277 = n38276 ^ n1897 ^ n1871 ;
  assign n38278 = n38277 ^ n16526 ^ 1'b0 ;
  assign n38279 = ( n16168 & n17205 ) | ( n16168 & n17224 ) | ( n17205 & n17224 ) ;
  assign n38280 = ( n33142 & n33969 ) | ( n33142 & ~n38279 ) | ( n33969 & ~n38279 ) ;
  assign n38281 = n4475 | n4832 ;
  assign n38282 = ( n9125 & ~n18889 ) | ( n9125 & n38281 ) | ( ~n18889 & n38281 ) ;
  assign n38283 = ( n2451 & n22067 ) | ( n2451 & ~n38282 ) | ( n22067 & ~n38282 ) ;
  assign n38284 = n23875 & n38283 ;
  assign n38285 = n38284 ^ n32921 ^ n32293 ;
  assign n38287 = n5513 & ~n17484 ;
  assign n38286 = n32438 ^ n2856 ^ 1'b0 ;
  assign n38288 = n38287 ^ n38286 ^ 1'b0 ;
  assign n38289 = n34046 ^ n26558 ^ n23886 ;
  assign n38290 = n6347 & n38289 ;
  assign n38291 = n30431 & n38290 ;
  assign n38292 = n25122 ^ n3931 ^ 1'b0 ;
  assign n38293 = n14917 | n38292 ;
  assign n38294 = ( n21101 & n22091 ) | ( n21101 & n28728 ) | ( n22091 & n28728 ) ;
  assign n38295 = ~n38293 & n38294 ;
  assign n38296 = ~n16485 & n38295 ;
  assign n38297 = ( n6882 & n10517 ) | ( n6882 & ~n11210 ) | ( n10517 & ~n11210 ) ;
  assign n38298 = ( ~n1465 & n9079 ) | ( ~n1465 & n19213 ) | ( n9079 & n19213 ) ;
  assign n38299 = n38297 & ~n38298 ;
  assign n38300 = n31568 & n38299 ;
  assign n38301 = n36944 ^ n6087 ^ 1'b0 ;
  assign n38302 = n35775 ^ n22593 ^ n2962 ;
  assign n38303 = n38302 ^ n28083 ^ n5591 ;
  assign n38304 = n23150 ^ n21630 ^ n615 ;
  assign n38305 = n38304 ^ n31872 ^ 1'b0 ;
  assign n38312 = n28600 ^ n14267 ^ 1'b0 ;
  assign n38306 = n22670 ^ n1127 ^ n378 ;
  assign n38307 = n38306 ^ n26613 ^ n12315 ;
  assign n38308 = n6750 ^ n555 ^ 1'b0 ;
  assign n38309 = ~n12521 & n38308 ;
  assign n38310 = ~n1807 & n38309 ;
  assign n38311 = ~n38307 & n38310 ;
  assign n38313 = n38312 ^ n38311 ^ n27503 ;
  assign n38314 = n9853 | n26399 ;
  assign n38315 = n28446 | n38314 ;
  assign n38316 = ( n12341 & n19688 ) | ( n12341 & n35656 ) | ( n19688 & n35656 ) ;
  assign n38317 = ( n3732 & n11303 ) | ( n3732 & n12812 ) | ( n11303 & n12812 ) ;
  assign n38318 = ~n6083 & n38317 ;
  assign n38319 = n38318 ^ n33925 ^ n951 ;
  assign n38320 = n5552 & ~n12900 ;
  assign n38321 = n4030 & n38320 ;
  assign n38322 = n6264 ^ n3316 ^ 1'b0 ;
  assign n38323 = ~n38321 & n38322 ;
  assign n38324 = ( ~n6569 & n7825 ) | ( ~n6569 & n17127 ) | ( n7825 & n17127 ) ;
  assign n38325 = n20974 | n33282 ;
  assign n38326 = ( n425 & ~n12135 ) | ( n425 & n27358 ) | ( ~n12135 & n27358 ) ;
  assign n38327 = n38326 ^ n22328 ^ n1487 ;
  assign n38328 = ( n7393 & n32362 ) | ( n7393 & n38327 ) | ( n32362 & n38327 ) ;
  assign n38329 = n14687 ^ n9450 ^ n2296 ;
  assign n38330 = n38329 ^ n27997 ^ n7611 ;
  assign n38331 = n38330 ^ n30237 ^ n11756 ;
  assign n38332 = n32020 ^ n19373 ^ 1'b0 ;
  assign n38333 = ( n19928 & n20118 ) | ( n19928 & n38332 ) | ( n20118 & n38332 ) ;
  assign n38334 = n35016 ^ n30903 ^ n22215 ;
  assign n38335 = ( n3340 & ~n21108 ) | ( n3340 & n37687 ) | ( ~n21108 & n37687 ) ;
  assign n38337 = n24872 ^ n22174 ^ 1'b0 ;
  assign n38336 = n37357 ^ n25020 ^ n4467 ;
  assign n38338 = n38337 ^ n38336 ^ n10721 ;
  assign n38339 = n24024 ^ n3490 ^ 1'b0 ;
  assign n38341 = n14757 ^ n1352 ^ n906 ;
  assign n38340 = n18614 ^ n7708 ^ n5165 ;
  assign n38342 = n38341 ^ n38340 ^ n10226 ;
  assign n38343 = ( ~n12701 & n21752 ) | ( ~n12701 & n33808 ) | ( n21752 & n33808 ) ;
  assign n38345 = n376 & ~n6982 ;
  assign n38344 = ~n28662 & n36903 ;
  assign n38346 = n38345 ^ n38344 ^ 1'b0 ;
  assign n38347 = n26274 ^ n15594 ^ 1'b0 ;
  assign n38348 = ( n15915 & n16439 ) | ( n15915 & ~n38347 ) | ( n16439 & ~n38347 ) ;
  assign n38349 = n7724 | n38348 ;
  assign n38350 = n10615 & ~n38349 ;
  assign n38351 = n6240 & ~n38350 ;
  assign n38352 = n32707 & n38351 ;
  assign n38353 = n25220 ^ n21769 ^ x14 ;
  assign n38354 = n35157 & ~n38353 ;
  assign n38355 = n14083 & ~n15157 ;
  assign n38356 = n9937 | n38355 ;
  assign n38357 = n38356 ^ n8734 ^ 1'b0 ;
  assign n38358 = ~n414 & n5113 ;
  assign n38359 = n11287 & n30642 ;
  assign n38360 = n38359 ^ n21994 ^ 1'b0 ;
  assign n38361 = ( ~n30552 & n38358 ) | ( ~n30552 & n38360 ) | ( n38358 & n38360 ) ;
  assign n38362 = ( n7027 & ~n35648 ) | ( n7027 & n37290 ) | ( ~n35648 & n37290 ) ;
  assign n38363 = ~n38361 & n38362 ;
  assign n38364 = n9872 & n38363 ;
  assign n38365 = ( n4597 & n24687 ) | ( n4597 & n33729 ) | ( n24687 & n33729 ) ;
  assign n38366 = n38365 ^ n8294 ^ n3670 ;
  assign n38367 = n36487 ^ n4597 ^ n3725 ;
  assign n38368 = n27218 ^ n24248 ^ n1175 ;
  assign n38369 = ( ~n15406 & n29897 ) | ( ~n15406 & n34021 ) | ( n29897 & n34021 ) ;
  assign n38370 = ~n27002 & n27862 ;
  assign n38371 = n823 | n38370 ;
  assign n38372 = ( n7348 & ~n28969 ) | ( n7348 & n38371 ) | ( ~n28969 & n38371 ) ;
  assign n38373 = n16836 & ~n18722 ;
  assign n38374 = n38373 ^ n29778 ^ 1'b0 ;
  assign n38377 = ~n12341 & n24265 ;
  assign n38375 = n12368 ^ n8352 ^ n5351 ;
  assign n38376 = ( n10574 & n23512 ) | ( n10574 & ~n38375 ) | ( n23512 & ~n38375 ) ;
  assign n38378 = n38377 ^ n38376 ^ 1'b0 ;
  assign n38379 = n29885 ^ n16260 ^ n15784 ;
  assign n38384 = n37443 ^ n7766 ^ 1'b0 ;
  assign n38382 = n17907 & n23395 ;
  assign n38383 = n34337 & n38382 ;
  assign n38380 = ( n2067 & n2896 ) | ( n2067 & ~n12024 ) | ( n2896 & ~n12024 ) ;
  assign n38381 = n38380 ^ n36503 ^ n26886 ;
  assign n38385 = n38384 ^ n38383 ^ n38381 ;
  assign n38386 = ( ~n1808 & n8971 ) | ( ~n1808 & n9675 ) | ( n8971 & n9675 ) ;
  assign n38387 = n8712 & n32547 ;
  assign n38388 = n38387 ^ n6336 ^ 1'b0 ;
  assign n38389 = ( n36069 & n38386 ) | ( n36069 & ~n38388 ) | ( n38386 & ~n38388 ) ;
  assign n38392 = n7764 | n14448 ;
  assign n38390 = n3740 & n10658 ;
  assign n38391 = n26465 & n38390 ;
  assign n38393 = n38392 ^ n38391 ^ n28246 ;
  assign n38394 = n17897 ^ n17441 ^ n11522 ;
  assign n38395 = ~n14772 & n28858 ;
  assign n38396 = n38394 & n38395 ;
  assign n38397 = n22801 ^ n13094 ^ 1'b0 ;
  assign n38398 = n4229 & ~n38397 ;
  assign n38399 = ( n12590 & ~n25853 ) | ( n12590 & n31698 ) | ( ~n25853 & n31698 ) ;
  assign n38400 = n19712 ^ n14940 ^ 1'b0 ;
  assign n38401 = n38400 ^ n7741 ^ 1'b0 ;
  assign n38402 = n12683 & ~n38401 ;
  assign n38403 = ( ~n7700 & n37966 ) | ( ~n7700 & n38402 ) | ( n37966 & n38402 ) ;
  assign n38404 = n12005 ^ n5800 ^ 1'b0 ;
  assign n38405 = n10493 ^ n8393 ^ 1'b0 ;
  assign n38406 = n24633 ^ n13079 ^ n8265 ;
  assign n38407 = n11471 ^ n3991 ^ 1'b0 ;
  assign n38408 = n38407 ^ n20342 ^ n5245 ;
  assign n38409 = n38408 ^ n11035 ^ n6465 ;
  assign n38410 = ~n10698 & n25163 ;
  assign n38411 = ( n5110 & n19730 ) | ( n5110 & n26259 ) | ( n19730 & n26259 ) ;
  assign n38412 = n29151 ^ n10824 ^ 1'b0 ;
  assign n38413 = ~n17249 & n38412 ;
  assign n38417 = n6556 ^ n1690 ^ 1'b0 ;
  assign n38414 = ~n4774 & n6905 ;
  assign n38415 = ~n4221 & n38414 ;
  assign n38416 = n10049 | n38415 ;
  assign n38418 = n38417 ^ n38416 ^ 1'b0 ;
  assign n38419 = n38413 & ~n38418 ;
  assign n38420 = n38419 ^ n28196 ^ n17490 ;
  assign n38421 = ( n13406 & ~n26713 ) | ( n13406 & n27428 ) | ( ~n26713 & n27428 ) ;
  assign n38422 = ( n24106 & n30385 ) | ( n24106 & n37923 ) | ( n30385 & n37923 ) ;
  assign n38423 = n38422 ^ n14386 ^ 1'b0 ;
  assign n38424 = ~n29433 & n38423 ;
  assign n38425 = ~n16125 & n20993 ;
  assign n38426 = n28161 ^ n2197 ^ 1'b0 ;
  assign n38427 = n3101 | n38426 ;
  assign n38429 = n32304 ^ n4380 ^ n1553 ;
  assign n38428 = ( n5358 & n7785 ) | ( n5358 & ~n8502 ) | ( n7785 & ~n8502 ) ;
  assign n38430 = n38429 ^ n38428 ^ n17677 ;
  assign n38431 = n38430 ^ n15148 ^ n4101 ;
  assign n38437 = n15399 ^ n8254 ^ n3048 ;
  assign n38432 = n29359 ^ n10217 ^ n3856 ;
  assign n38433 = n38432 ^ n27988 ^ n23246 ;
  assign n38434 = ( ~n10132 & n15133 ) | ( ~n10132 & n26702 ) | ( n15133 & n26702 ) ;
  assign n38435 = ( ~x154 & n2614 ) | ( ~x154 & n17878 ) | ( n2614 & n17878 ) ;
  assign n38436 = ( n38433 & n38434 ) | ( n38433 & ~n38435 ) | ( n38434 & ~n38435 ) ;
  assign n38438 = n38437 ^ n38436 ^ n32345 ;
  assign n38439 = n22149 ^ n19789 ^ 1'b0 ;
  assign n38442 = n2724 & ~n17454 ;
  assign n38443 = ~n865 & n38442 ;
  assign n38444 = n29503 ^ n17693 ^ 1'b0 ;
  assign n38445 = n38443 | n38444 ;
  assign n38446 = n29846 & n38445 ;
  assign n38440 = n820 & ~n10401 ;
  assign n38441 = ~x111 & n38440 ;
  assign n38447 = n38446 ^ n38441 ^ n17300 ;
  assign n38448 = n10209 & ~n26261 ;
  assign n38449 = n38448 ^ n11908 ^ 1'b0 ;
  assign n38450 = n4277 | n38449 ;
  assign n38451 = n38450 ^ n22783 ^ 1'b0 ;
  assign n38452 = n35125 | n38451 ;
  assign n38453 = n20648 & ~n38452 ;
  assign n38457 = ( ~n502 & n13131 ) | ( ~n502 & n21508 ) | ( n13131 & n21508 ) ;
  assign n38454 = n24963 ^ n14992 ^ 1'b0 ;
  assign n38455 = ~n14727 & n38454 ;
  assign n38456 = n38455 ^ n19027 ^ n16841 ;
  assign n38458 = n38457 ^ n38456 ^ n15689 ;
  assign n38459 = ~n34259 & n34554 ;
  assign n38460 = ( n1064 & n11217 ) | ( n1064 & ~n12746 ) | ( n11217 & ~n12746 ) ;
  assign n38461 = n25891 ^ n12307 ^ n5461 ;
  assign n38462 = ( ~n9351 & n38460 ) | ( ~n9351 & n38461 ) | ( n38460 & n38461 ) ;
  assign n38467 = n18479 ^ n4260 ^ n2210 ;
  assign n38468 = ~n23761 & n34512 ;
  assign n38469 = ( n11064 & n38467 ) | ( n11064 & ~n38468 ) | ( n38467 & ~n38468 ) ;
  assign n38463 = n38077 ^ n27057 ^ 1'b0 ;
  assign n38464 = n7302 & n38463 ;
  assign n38465 = n8014 ^ n6789 ^ 1'b0 ;
  assign n38466 = ( n35617 & ~n38464 ) | ( n35617 & n38465 ) | ( ~n38464 & n38465 ) ;
  assign n38470 = n38469 ^ n38466 ^ n28141 ;
  assign n38471 = n4056 ^ n2550 ^ 1'b0 ;
  assign n38472 = ( n17187 & n28384 ) | ( n17187 & ~n38471 ) | ( n28384 & ~n38471 ) ;
  assign n38473 = x197 & n7281 ;
  assign n38474 = n38473 ^ n29893 ^ 1'b0 ;
  assign n38475 = ~n18722 & n28765 ;
  assign n38476 = n34261 & n38475 ;
  assign n38477 = n38476 ^ n26892 ^ n5829 ;
  assign n38478 = n38474 | n38477 ;
  assign n38479 = n21944 ^ n12413 ^ n10659 ;
  assign n38480 = n14903 ^ n10967 ^ n4389 ;
  assign n38481 = n38480 ^ n17211 ^ n4067 ;
  assign n38482 = n22542 | n38481 ;
  assign n38483 = n38479 | n38482 ;
  assign n38484 = ( n15416 & ~n16803 ) | ( n15416 & n23889 ) | ( ~n16803 & n23889 ) ;
  assign n38485 = n13361 ^ n8127 ^ n4539 ;
  assign n38486 = ( n24433 & ~n30113 ) | ( n24433 & n38485 ) | ( ~n30113 & n38485 ) ;
  assign n38487 = n22391 & ~n32639 ;
  assign n38488 = n7122 ^ n1600 ^ 1'b0 ;
  assign n38489 = n1251 | n30654 ;
  assign n38490 = n38489 ^ n16186 ^ 1'b0 ;
  assign n38491 = ( n22385 & n38488 ) | ( n22385 & n38490 ) | ( n38488 & n38490 ) ;
  assign n38492 = ( n7467 & ~n14990 ) | ( n7467 & n16200 ) | ( ~n14990 & n16200 ) ;
  assign n38493 = n9014 & ~n38492 ;
  assign n38494 = ~n36971 & n38493 ;
  assign n38495 = n3781 & ~n24814 ;
  assign n38496 = n38495 ^ n24853 ^ 1'b0 ;
  assign n38497 = ~n35402 & n38496 ;
  assign n38498 = n4371 & n17501 ;
  assign n38499 = n36560 & n38498 ;
  assign n38500 = n34861 ^ n12795 ^ n4093 ;
  assign n38501 = n5108 & ~n14537 ;
  assign n38502 = n38501 ^ n5726 ^ 1'b0 ;
  assign n38503 = n28234 ^ n14847 ^ n9071 ;
  assign n38504 = ~n38502 & n38503 ;
  assign n38505 = n34918 ^ n12436 ^ n1451 ;
  assign n38506 = n24884 & ~n38505 ;
  assign n38507 = n33889 ^ n31912 ^ 1'b0 ;
  assign n38508 = ~n5745 & n17301 ;
  assign n38509 = n38508 ^ n23338 ^ 1'b0 ;
  assign n38510 = n15627 & n38509 ;
  assign n38511 = n34346 & n38510 ;
  assign n38512 = n38511 ^ n4744 ^ 1'b0 ;
  assign n38513 = n8414 & n24981 ;
  assign n38514 = n17509 & n18753 ;
  assign n38515 = n32734 ^ n30594 ^ 1'b0 ;
  assign n38516 = n38514 | n38515 ;
  assign n38517 = n24069 ^ n7315 ^ 1'b0 ;
  assign n38518 = n24823 ^ n21957 ^ n2853 ;
  assign n38519 = n38445 ^ n38167 ^ n18108 ;
  assign n38520 = n17429 ^ n15540 ^ n13387 ;
  assign n38521 = n9465 ^ n7881 ^ n4765 ;
  assign n38522 = n38521 ^ n21975 ^ 1'b0 ;
  assign n38523 = n32532 ^ n19902 ^ n18820 ;
  assign n38524 = ( n6642 & n20523 ) | ( n6642 & ~n24160 ) | ( n20523 & ~n24160 ) ;
  assign n38525 = ( ~n12226 & n21101 ) | ( ~n12226 & n38524 ) | ( n21101 & n38524 ) ;
  assign n38526 = n15145 ^ n8670 ^ 1'b0 ;
  assign n38527 = n30275 ^ n9707 ^ n7594 ;
  assign n38528 = ( ~n38525 & n38526 ) | ( ~n38525 & n38527 ) | ( n38526 & n38527 ) ;
  assign n38529 = n7466 & ~n9793 ;
  assign n38530 = n3115 & n38529 ;
  assign n38531 = n24497 ^ n19699 ^ 1'b0 ;
  assign n38532 = x61 & ~n38531 ;
  assign n38533 = ( n11368 & n15603 ) | ( n11368 & n36996 ) | ( n15603 & n36996 ) ;
  assign n38534 = ( n5637 & ~n7023 ) | ( n5637 & n38533 ) | ( ~n7023 & n38533 ) ;
  assign n38535 = n27505 ^ n25801 ^ n3617 ;
  assign n38536 = n38535 ^ n26165 ^ 1'b0 ;
  assign n38537 = ~n7005 & n38536 ;
  assign n38538 = n24507 ^ n11724 ^ 1'b0 ;
  assign n38539 = n8472 ^ n1241 ^ 1'b0 ;
  assign n38540 = n9499 | n38539 ;
  assign n38541 = ( n18907 & n33425 ) | ( n18907 & ~n38540 ) | ( n33425 & ~n38540 ) ;
  assign n38542 = n4400 ^ n2840 ^ 1'b0 ;
  assign n38543 = n38541 & ~n38542 ;
  assign n38544 = ~n31863 & n38543 ;
  assign n38545 = ~n38538 & n38544 ;
  assign n38546 = n17762 & n38545 ;
  assign n38547 = n21992 ^ n21461 ^ n19619 ;
  assign n38550 = n20741 & ~n22987 ;
  assign n38551 = n29604 & n38550 ;
  assign n38548 = n13486 ^ n11170 ^ 1'b0 ;
  assign n38549 = n18337 | n38548 ;
  assign n38552 = n38551 ^ n38549 ^ n36734 ;
  assign n38553 = ~n20067 & n30914 ;
  assign n38554 = ~n38552 & n38553 ;
  assign n38555 = n23569 ^ x163 ^ 1'b0 ;
  assign n38556 = n38555 ^ n14144 ^ 1'b0 ;
  assign n38557 = n37381 ^ n32286 ^ n15932 ;
  assign n38559 = n10325 & n30991 ;
  assign n38558 = n18917 ^ n12279 ^ n3128 ;
  assign n38560 = n38559 ^ n38558 ^ n27567 ;
  assign n38561 = ( n6710 & ~n15556 ) | ( n6710 & n38560 ) | ( ~n15556 & n38560 ) ;
  assign n38562 = n19555 ^ n15022 ^ 1'b0 ;
  assign n38563 = n8825 | n38562 ;
  assign n38564 = ( ~n4049 & n30426 ) | ( ~n4049 & n38563 ) | ( n30426 & n38563 ) ;
  assign n38565 = n38564 ^ n3387 ^ 1'b0 ;
  assign n38566 = n12702 ^ n7686 ^ n1495 ;
  assign n38567 = n10547 & n12344 ;
  assign n38568 = ( n5230 & n17121 ) | ( n5230 & ~n38567 ) | ( n17121 & ~n38567 ) ;
  assign n38569 = ( n3579 & ~n10817 ) | ( n3579 & n15799 ) | ( ~n10817 & n15799 ) ;
  assign n38570 = ( n3854 & n33787 ) | ( n3854 & ~n34040 ) | ( n33787 & ~n34040 ) ;
  assign n38571 = ~n38569 & n38570 ;
  assign n38574 = n27866 ^ n25589 ^ n20946 ;
  assign n38572 = ( ~n3966 & n8356 ) | ( ~n3966 & n28101 ) | ( n8356 & n28101 ) ;
  assign n38573 = ~n26791 & n38572 ;
  assign n38575 = n38574 ^ n38573 ^ 1'b0 ;
  assign n38576 = n3511 & n7290 ;
  assign n38577 = n38576 ^ n25712 ^ 1'b0 ;
  assign n38578 = n38577 ^ n9910 ^ n7857 ;
  assign n38582 = ( ~x80 & n336 ) | ( ~x80 & n17933 ) | ( n336 & n17933 ) ;
  assign n38579 = n8039 & ~n15086 ;
  assign n38580 = n38579 ^ n33912 ^ 1'b0 ;
  assign n38581 = n38580 ^ n5237 ^ n3725 ;
  assign n38583 = n38582 ^ n38581 ^ n22306 ;
  assign n38584 = ( n1738 & n4168 ) | ( n1738 & n12739 ) | ( n4168 & n12739 ) ;
  assign n38585 = n21352 ^ n874 ^ 1'b0 ;
  assign n38586 = n38584 | n38585 ;
  assign n38587 = n694 & ~n5142 ;
  assign n38588 = n38587 ^ n3158 ^ 1'b0 ;
  assign n38594 = ~n7795 & n23786 ;
  assign n38595 = ~n7199 & n38594 ;
  assign n38589 = n1027 | n7148 ;
  assign n38590 = n6834 & ~n38589 ;
  assign n38591 = n11079 & ~n38590 ;
  assign n38592 = ~n10314 & n38591 ;
  assign n38593 = ( n14184 & ~n20759 ) | ( n14184 & n38592 ) | ( ~n20759 & n38592 ) ;
  assign n38596 = n38595 ^ n38593 ^ n33038 ;
  assign n38600 = n32089 ^ n10761 ^ 1'b0 ;
  assign n38599 = ( n9644 & ~n16836 ) | ( n9644 & n35953 ) | ( ~n16836 & n35953 ) ;
  assign n38597 = n14453 | n16608 ;
  assign n38598 = n38597 ^ n28206 ^ n1406 ;
  assign n38601 = n38600 ^ n38599 ^ n38598 ;
  assign n38602 = n25483 | n36474 ;
  assign n38603 = n31291 ^ n14992 ^ 1'b0 ;
  assign n38604 = n26169 & n28087 ;
  assign n38605 = ~n20651 & n38604 ;
  assign n38606 = ( ~n5958 & n10206 ) | ( ~n5958 & n38605 ) | ( n10206 & n38605 ) ;
  assign n38607 = n38606 ^ n30710 ^ 1'b0 ;
  assign n38608 = n27971 | n38607 ;
  assign n38609 = n28846 ^ n482 ^ 1'b0 ;
  assign n38610 = n3624 & n38609 ;
  assign n38611 = n16444 ^ n9673 ^ 1'b0 ;
  assign n38612 = ( n12492 & n33636 ) | ( n12492 & n34297 ) | ( n33636 & n34297 ) ;
  assign n38615 = ( ~n1920 & n5181 ) | ( ~n1920 & n6195 ) | ( n5181 & n6195 ) ;
  assign n38613 = n23455 ^ n20462 ^ n6687 ;
  assign n38614 = ( ~n3495 & n7460 ) | ( ~n3495 & n38613 ) | ( n7460 & n38613 ) ;
  assign n38616 = n38615 ^ n38614 ^ n37589 ;
  assign n38617 = ( ~n15248 & n18032 ) | ( ~n15248 & n29029 ) | ( n18032 & n29029 ) ;
  assign n38618 = ~n33425 & n38617 ;
  assign n38619 = n38569 ^ n36806 ^ 1'b0 ;
  assign n38620 = n27288 ^ n25274 ^ 1'b0 ;
  assign n38621 = ( n2074 & n6996 ) | ( n2074 & n30061 ) | ( n6996 & n30061 ) ;
  assign n38622 = ( n9479 & n12010 ) | ( n9479 & n38621 ) | ( n12010 & n38621 ) ;
  assign n38623 = n8674 | n38622 ;
  assign n38624 = n22410 | n38623 ;
  assign n38627 = ( n4641 & ~n19894 ) | ( n4641 & n26887 ) | ( ~n19894 & n26887 ) ;
  assign n38625 = n13423 ^ n3399 ^ 1'b0 ;
  assign n38626 = ( n11897 & n18613 ) | ( n11897 & n38625 ) | ( n18613 & n38625 ) ;
  assign n38628 = n38627 ^ n38626 ^ 1'b0 ;
  assign n38629 = n15116 ^ n2949 ^ 1'b0 ;
  assign n38630 = n2029 & ~n38629 ;
  assign n38633 = n24100 ^ n12560 ^ n9054 ;
  assign n38631 = n25244 ^ n8868 ^ 1'b0 ;
  assign n38632 = n11471 | n38631 ;
  assign n38634 = n38633 ^ n38632 ^ n5269 ;
  assign n38635 = ( n11608 & n38630 ) | ( n11608 & ~n38634 ) | ( n38630 & ~n38634 ) ;
  assign n38636 = n23186 ^ n9877 ^ n5602 ;
  assign n38637 = n38636 ^ n29427 ^ n1014 ;
  assign n38638 = n32059 ^ n22446 ^ n12722 ;
  assign n38639 = n19729 ^ n3162 ^ 1'b0 ;
  assign n38640 = n10780 & ~n38639 ;
  assign n38641 = ( n16422 & n19123 ) | ( n16422 & n26133 ) | ( n19123 & n26133 ) ;
  assign n38642 = n1598 | n29938 ;
  assign n38643 = n38641 | n38642 ;
  assign n38644 = n5719 ^ n1143 ^ 1'b0 ;
  assign n38645 = n13098 & n38644 ;
  assign n38646 = n38645 ^ n4422 ^ n1482 ;
  assign n38647 = n38646 ^ n28564 ^ n24588 ;
  assign n38648 = ( n15228 & n15674 ) | ( n15228 & n38647 ) | ( n15674 & n38647 ) ;
  assign n38649 = n409 | n38648 ;
  assign n38652 = n25594 ^ n23961 ^ n15640 ;
  assign n38650 = n1070 & ~n10282 ;
  assign n38651 = ~n11443 & n38650 ;
  assign n38653 = n38652 ^ n38651 ^ 1'b0 ;
  assign n38654 = n9808 & n22574 ;
  assign n38655 = n38654 ^ n3945 ^ 1'b0 ;
  assign n38656 = n2724 & n18174 ;
  assign n38657 = n38656 ^ n38194 ^ 1'b0 ;
  assign n38658 = ( ~n1365 & n3204 ) | ( ~n1365 & n38657 ) | ( n3204 & n38657 ) ;
  assign n38659 = ( ~n4988 & n16586 ) | ( ~n4988 & n38658 ) | ( n16586 & n38658 ) ;
  assign n38660 = n28941 ^ n14632 ^ 1'b0 ;
  assign n38661 = ( ~n17993 & n33168 ) | ( ~n17993 & n38660 ) | ( n33168 & n38660 ) ;
  assign n38662 = n28507 ^ n23896 ^ 1'b0 ;
  assign n38663 = n38662 ^ n27720 ^ n8448 ;
  assign n38664 = n22714 ^ n10321 ^ n7600 ;
  assign n38665 = n38664 ^ n25916 ^ n7676 ;
  assign n38666 = n16954 ^ n15836 ^ x199 ;
  assign n38667 = ~n2292 & n38666 ;
  assign n38668 = n4120 & n38667 ;
  assign n38669 = n11381 | n30432 ;
  assign n38670 = n25847 | n38669 ;
  assign n38672 = ( n4774 & ~n19139 ) | ( n4774 & n20985 ) | ( ~n19139 & n20985 ) ;
  assign n38673 = ( n5158 & n19552 ) | ( n5158 & ~n38672 ) | ( n19552 & ~n38672 ) ;
  assign n38671 = n33163 ^ n16753 ^ n8337 ;
  assign n38674 = n38673 ^ n38671 ^ n21730 ;
  assign n38677 = ~n6505 & n27434 ;
  assign n38678 = ~n23882 & n38677 ;
  assign n38675 = n5532 & ~n6220 ;
  assign n38676 = n20470 & n38675 ;
  assign n38679 = n38678 ^ n38676 ^ n4188 ;
  assign n38680 = n7572 | n11322 ;
  assign n38681 = n38680 ^ n17838 ^ 1'b0 ;
  assign n38682 = n38681 ^ n17897 ^ n14460 ;
  assign n38683 = n11032 | n31438 ;
  assign n38684 = ( ~n5958 & n16118 ) | ( ~n5958 & n38683 ) | ( n16118 & n38683 ) ;
  assign n38685 = n38684 ^ n11710 ^ 1'b0 ;
  assign n38686 = ~n27512 & n38685 ;
  assign n38687 = n22365 & n38686 ;
  assign n38688 = n38687 ^ n14251 ^ 1'b0 ;
  assign n38689 = n36412 & n38688 ;
  assign n38690 = n28141 & n38689 ;
  assign n38691 = ( n8767 & n9303 ) | ( n8767 & ~n20355 ) | ( n9303 & ~n20355 ) ;
  assign n38692 = ( n8246 & n20855 ) | ( n8246 & n38691 ) | ( n20855 & n38691 ) ;
  assign n38693 = ( n5488 & ~n24199 ) | ( n5488 & n33680 ) | ( ~n24199 & n33680 ) ;
  assign n38694 = n16869 ^ n8874 ^ n593 ;
  assign n38695 = n801 & ~n8454 ;
  assign n38696 = ~n28218 & n38695 ;
  assign n38698 = n2142 & ~n8547 ;
  assign n38699 = n15498 & n38698 ;
  assign n38697 = n5985 | n9478 ;
  assign n38700 = n38699 ^ n38697 ^ 1'b0 ;
  assign n38701 = ~n4004 & n4448 ;
  assign n38702 = ( n7277 & ~n14449 ) | ( n7277 & n21829 ) | ( ~n14449 & n21829 ) ;
  assign n38703 = n38702 ^ n19452 ^ 1'b0 ;
  assign n38704 = ( n13681 & n38701 ) | ( n13681 & n38703 ) | ( n38701 & n38703 ) ;
  assign n38705 = ( n706 & n2538 ) | ( n706 & n38704 ) | ( n2538 & n38704 ) ;
  assign n38706 = n5500 & ~n38219 ;
  assign n38707 = ~n5179 & n38706 ;
  assign n38708 = ( n26349 & n30957 ) | ( n26349 & ~n36780 ) | ( n30957 & ~n36780 ) ;
  assign n38709 = n24219 ^ n17186 ^ n4499 ;
  assign n38710 = n30531 ^ n22003 ^ 1'b0 ;
  assign n38711 = n26348 | n38710 ;
  assign n38712 = n34853 ^ n2288 ^ 1'b0 ;
  assign n38713 = n15435 | n38712 ;
  assign n38714 = n27272 ^ n13948 ^ n12020 ;
  assign n38715 = ( n5257 & ~n14515 ) | ( n5257 & n38714 ) | ( ~n14515 & n38714 ) ;
  assign n38716 = ( n21058 & ~n38713 ) | ( n21058 & n38715 ) | ( ~n38713 & n38715 ) ;
  assign n38717 = ( ~n15941 & n30904 ) | ( ~n15941 & n31193 ) | ( n30904 & n31193 ) ;
  assign n38724 = ( n8781 & ~n9064 ) | ( n8781 & n25586 ) | ( ~n9064 & n25586 ) ;
  assign n38721 = n1375 ^ n547 ^ 1'b0 ;
  assign n38722 = n23221 | n38721 ;
  assign n38718 = n26429 ^ n17174 ^ n4339 ;
  assign n38719 = n38718 ^ n21106 ^ 1'b0 ;
  assign n38720 = n28239 & n38719 ;
  assign n38723 = n38722 ^ n38720 ^ n10541 ;
  assign n38725 = n38724 ^ n38723 ^ 1'b0 ;
  assign n38726 = ~n35580 & n38725 ;
  assign n38727 = n24658 ^ n18086 ^ 1'b0 ;
  assign n38728 = n3668 & ~n38727 ;
  assign n38729 = ( ~n3547 & n38726 ) | ( ~n3547 & n38728 ) | ( n38726 & n38728 ) ;
  assign n38730 = n19531 ^ n13999 ^ 1'b0 ;
  assign n38731 = n38730 ^ n34563 ^ n19224 ;
  assign n38732 = ( n6076 & n12372 ) | ( n6076 & n22489 ) | ( n12372 & n22489 ) ;
  assign n38733 = n25025 & n37362 ;
  assign n38734 = ~n28713 & n38733 ;
  assign n38735 = n38005 ^ n21040 ^ 1'b0 ;
  assign n38736 = n33926 | n38735 ;
  assign n38737 = n38736 ^ n17553 ^ n5269 ;
  assign n38738 = n34434 ^ n3006 ^ n2357 ;
  assign n38739 = n36559 ^ n350 ^ 1'b0 ;
  assign n38740 = n38739 ^ n2629 ^ 1'b0 ;
  assign n38741 = ( ~n4995 & n9679 ) | ( ~n4995 & n19015 ) | ( n9679 & n19015 ) ;
  assign n38742 = ( n14047 & n18967 ) | ( n14047 & n38741 ) | ( n18967 & n38741 ) ;
  assign n38743 = ( ~n10346 & n27333 ) | ( ~n10346 & n38742 ) | ( n27333 & n38742 ) ;
  assign n38744 = n18834 ^ n18260 ^ n13209 ;
  assign n38745 = n20049 & ~n38744 ;
  assign n38746 = n8928 & n38745 ;
  assign n38747 = ~n5093 & n17758 ;
  assign n38748 = n38747 ^ n5253 ^ 1'b0 ;
  assign n38749 = ~n38746 & n38748 ;
  assign n38751 = n17427 & ~n20766 ;
  assign n38750 = n4383 & ~n15162 ;
  assign n38752 = n38751 ^ n38750 ^ n1634 ;
  assign n38753 = n19904 ^ n3925 ^ x229 ;
  assign n38754 = n38753 ^ n18898 ^ 1'b0 ;
  assign n38755 = n24142 ^ n19227 ^ n9073 ;
  assign n38756 = x78 & n2794 ;
  assign n38757 = n38756 ^ n23208 ^ 1'b0 ;
  assign n38758 = ( n6077 & n9345 ) | ( n6077 & ~n38757 ) | ( n9345 & ~n38757 ) ;
  assign n38759 = ~n13533 & n33534 ;
  assign n38760 = ~n13545 & n38759 ;
  assign n38761 = n32883 ^ n16815 ^ n9046 ;
  assign n38762 = n26803 ^ n23349 ^ x28 ;
  assign n38763 = n16642 ^ n16471 ^ 1'b0 ;
  assign n38764 = ( ~n20917 & n38762 ) | ( ~n20917 & n38763 ) | ( n38762 & n38763 ) ;
  assign n38765 = ( n7717 & n14199 ) | ( n7717 & n21345 ) | ( n14199 & n21345 ) ;
  assign n38766 = n38765 ^ n20996 ^ n2357 ;
  assign n38767 = n16128 | n38766 ;
  assign n38768 = n18134 & n38767 ;
  assign n38769 = n38768 ^ n37770 ^ n2931 ;
  assign n38770 = n36863 ^ n17743 ^ n1070 ;
  assign n38771 = n5930 ^ n1727 ^ 1'b0 ;
  assign n38772 = ~n11348 & n38771 ;
  assign n38773 = ( ~n13232 & n27057 ) | ( ~n13232 & n35510 ) | ( n27057 & n35510 ) ;
  assign n38774 = ( n12542 & n38772 ) | ( n12542 & ~n38773 ) | ( n38772 & ~n38773 ) ;
  assign n38775 = n20891 | n38774 ;
  assign n38776 = ( n1063 & ~n14014 ) | ( n1063 & n37961 ) | ( ~n14014 & n37961 ) ;
  assign n38777 = n38776 ^ n21494 ^ n343 ;
  assign n38778 = n17933 ^ n8106 ^ 1'b0 ;
  assign n38779 = n3073 | n38778 ;
  assign n38780 = n25583 | n38779 ;
  assign n38781 = n17288 | n38780 ;
  assign n38782 = ~n7211 & n38781 ;
  assign n38783 = n38782 ^ n20736 ^ 1'b0 ;
  assign n38784 = n38783 ^ n1476 ^ 1'b0 ;
  assign n38785 = n3900 | n13109 ;
  assign n38786 = n8690 & ~n38785 ;
  assign n38787 = n38786 ^ n31043 ^ 1'b0 ;
  assign n38788 = n18990 ^ n16111 ^ n7335 ;
  assign n38789 = n11442 ^ n11345 ^ 1'b0 ;
  assign n38790 = n4413 | n6813 ;
  assign n38791 = n38789 & ~n38790 ;
  assign n38792 = ~n8538 & n21634 ;
  assign n38793 = n19143 & n38792 ;
  assign n38794 = n12289 ^ n6963 ^ n1408 ;
  assign n38795 = n28730 & n38794 ;
  assign n38796 = n38795 ^ n8234 ^ 1'b0 ;
  assign n38797 = n37258 ^ n13878 ^ 1'b0 ;
  assign n38798 = n38524 ^ n27619 ^ n11616 ;
  assign n38799 = n38798 ^ n38651 ^ n16530 ;
  assign n38800 = n31400 ^ n30408 ^ n17631 ;
  assign n38801 = ( n15563 & n22501 ) | ( n15563 & ~n38800 ) | ( n22501 & ~n38800 ) ;
  assign n38804 = ( ~n8148 & n8728 ) | ( ~n8148 & n20844 ) | ( n8728 & n20844 ) ;
  assign n38805 = n38804 ^ n35914 ^ n24006 ;
  assign n38802 = n18905 & n22243 ;
  assign n38803 = n10559 & ~n38802 ;
  assign n38806 = n38805 ^ n38803 ^ 1'b0 ;
  assign n38807 = n16515 ^ n16094 ^ 1'b0 ;
  assign n38808 = ~n20362 & n38807 ;
  assign n38809 = ( n431 & n8674 ) | ( n431 & ~n28395 ) | ( n8674 & ~n28395 ) ;
  assign n38810 = ~n13657 & n19842 ;
  assign n38811 = n38809 & n38810 ;
  assign n38812 = n27448 ^ n20623 ^ n14595 ;
  assign n38813 = ~n13663 & n23704 ;
  assign n38814 = n38813 ^ n32993 ^ 1'b0 ;
  assign n38815 = n38814 ^ n10327 ^ 1'b0 ;
  assign n38816 = ( n4138 & n5732 ) | ( n4138 & ~n26165 ) | ( n5732 & ~n26165 ) ;
  assign n38817 = n15805 | n35396 ;
  assign n38818 = ( n5261 & n26691 ) | ( n5261 & n28325 ) | ( n26691 & n28325 ) ;
  assign n38819 = ( n17498 & ~n19574 ) | ( n17498 & n30656 ) | ( ~n19574 & n30656 ) ;
  assign n38820 = n30828 ^ n10973 ^ 1'b0 ;
  assign n38821 = x81 & n38820 ;
  assign n38822 = ~n10206 & n12114 ;
  assign n38823 = n20784 & n38822 ;
  assign n38824 = ( ~n3539 & n38821 ) | ( ~n3539 & n38823 ) | ( n38821 & n38823 ) ;
  assign n38825 = n5348 | n5836 ;
  assign n38826 = n38825 ^ n32128 ^ 1'b0 ;
  assign n38827 = ( n1341 & n30959 ) | ( n1341 & n38826 ) | ( n30959 & n38826 ) ;
  assign n38828 = n13567 & ~n19068 ;
  assign n38829 = n38827 & n38828 ;
  assign n38830 = n36977 ^ n11893 ^ 1'b0 ;
  assign n38831 = ( n6161 & ~n14021 ) | ( n6161 & n38830 ) | ( ~n14021 & n38830 ) ;
  assign n38832 = ~n26019 & n33120 ;
  assign n38833 = n38832 ^ n14777 ^ 1'b0 ;
  assign n38834 = n38831 & ~n38833 ;
  assign n38835 = n38834 ^ n10079 ^ 1'b0 ;
  assign n38836 = n22785 ^ n20833 ^ n17378 ;
  assign n38837 = n4876 & ~n21545 ;
  assign n38839 = n27583 ^ n21194 ^ n18217 ;
  assign n38840 = n14098 & ~n38839 ;
  assign n38838 = n16493 | n32031 ;
  assign n38841 = n38840 ^ n38838 ^ n20940 ;
  assign n38842 = n38321 ^ n20641 ^ n1409 ;
  assign n38843 = n29826 ^ n11242 ^ n1611 ;
  assign n38844 = n6138 & ~n21615 ;
  assign n38845 = n7850 & n38844 ;
  assign n38846 = ( ~n38842 & n38843 ) | ( ~n38842 & n38845 ) | ( n38843 & n38845 ) ;
  assign n38851 = n19766 ^ n7369 ^ n2784 ;
  assign n38852 = n33844 ^ n23419 ^ 1'b0 ;
  assign n38853 = n38851 & n38852 ;
  assign n38848 = n16146 & n19473 ;
  assign n38849 = n38848 ^ n3787 ^ 1'b0 ;
  assign n38847 = ( ~n4373 & n8022 ) | ( ~n4373 & n29283 ) | ( n8022 & n29283 ) ;
  assign n38850 = n38849 ^ n38847 ^ n20369 ;
  assign n38854 = n38853 ^ n38850 ^ 1'b0 ;
  assign n38855 = n37052 & n38854 ;
  assign n38856 = n35249 ^ n4439 ^ 1'b0 ;
  assign n38857 = n22979 & ~n38856 ;
  assign n38858 = n11601 | n27726 ;
  assign n38859 = n38858 ^ n18405 ^ 1'b0 ;
  assign n38861 = n6809 ^ n6085 ^ 1'b0 ;
  assign n38862 = ~n5619 & n38861 ;
  assign n38863 = ( n15689 & ~n18709 ) | ( n15689 & n38862 ) | ( ~n18709 & n38862 ) ;
  assign n38860 = n28423 & ~n34515 ;
  assign n38864 = n38863 ^ n38860 ^ 1'b0 ;
  assign n38865 = n13296 ^ n12927 ^ n7144 ;
  assign n38866 = ( x46 & n38864 ) | ( x46 & n38865 ) | ( n38864 & n38865 ) ;
  assign n38867 = n10360 | n15583 ;
  assign n38868 = n38867 ^ n10171 ^ 1'b0 ;
  assign n38869 = ( n2609 & ~n15992 ) | ( n2609 & n38868 ) | ( ~n15992 & n38868 ) ;
  assign n38870 = n35737 ^ n4875 ^ 1'b0 ;
  assign n38871 = n9393 & ~n38870 ;
  assign n38872 = n38871 ^ n10587 ^ n8724 ;
  assign n38873 = n11689 ^ n5332 ^ 1'b0 ;
  assign n38874 = ( n1090 & n4959 ) | ( n1090 & n38849 ) | ( n4959 & n38849 ) ;
  assign n38875 = n38873 & n38874 ;
  assign n38876 = n19437 | n36579 ;
  assign n38877 = n36414 & n36713 ;
  assign n38878 = ~n5612 & n38877 ;
  assign n38879 = ( n14626 & n23541 ) | ( n14626 & ~n38878 ) | ( n23541 & ~n38878 ) ;
  assign n38880 = n27458 ^ n20657 ^ n10654 ;
  assign n38881 = ( n2440 & n15608 ) | ( n2440 & ~n36545 ) | ( n15608 & ~n36545 ) ;
  assign n38882 = n38881 ^ n30420 ^ n13689 ;
  assign n38885 = n1200 & n9318 ;
  assign n38886 = n38885 ^ n15224 ^ 1'b0 ;
  assign n38887 = n38886 ^ n22859 ^ 1'b0 ;
  assign n38883 = ~n19637 & n26593 ;
  assign n38884 = n29827 & n38883 ;
  assign n38888 = n38887 ^ n38884 ^ n20970 ;
  assign n38889 = n29864 ^ n25665 ^ n15370 ;
  assign n38890 = ( n23419 & n28101 ) | ( n23419 & n38889 ) | ( n28101 & n38889 ) ;
  assign n38891 = ( n18163 & n38888 ) | ( n18163 & n38890 ) | ( n38888 & n38890 ) ;
  assign n38895 = ( n17213 & n28400 ) | ( n17213 & ~n34690 ) | ( n28400 & ~n34690 ) ;
  assign n38892 = n21667 ^ n2022 ^ n1642 ;
  assign n38893 = n3635 & n38892 ;
  assign n38894 = n38893 ^ n38762 ^ n17346 ;
  assign n38896 = n38895 ^ n38894 ^ n15510 ;
  assign n38897 = n19038 ^ n13513 ^ 1'b0 ;
  assign n38898 = ( n688 & ~n22498 ) | ( n688 & n24151 ) | ( ~n22498 & n24151 ) ;
  assign n38899 = ( n10790 & ~n27088 ) | ( n10790 & n34198 ) | ( ~n27088 & n34198 ) ;
  assign n38900 = n38899 ^ n23030 ^ 1'b0 ;
  assign n38901 = n21482 | n38900 ;
  assign n38902 = ( ~n14232 & n20378 ) | ( ~n14232 & n21917 ) | ( n20378 & n21917 ) ;
  assign n38903 = ( n7253 & n24024 ) | ( n7253 & ~n38902 ) | ( n24024 & ~n38902 ) ;
  assign n38904 = n13759 | n15354 ;
  assign n38905 = ( n1248 & ~n35104 ) | ( n1248 & n38904 ) | ( ~n35104 & n38904 ) ;
  assign n38906 = n31460 ^ n17757 ^ n7574 ;
  assign n38907 = n38906 ^ n26511 ^ n20528 ;
  assign n38908 = n4852 & n8023 ;
  assign n38909 = n38908 ^ n16245 ^ n8037 ;
  assign n38910 = ~n38907 & n38909 ;
  assign n38911 = n13560 & ~n29870 ;
  assign n38912 = ( n38905 & n38910 ) | ( n38905 & ~n38911 ) | ( n38910 & ~n38911 ) ;
  assign n38915 = ( n850 & n17312 ) | ( n850 & ~n31455 ) | ( n17312 & ~n31455 ) ;
  assign n38913 = n7826 ^ n4494 ^ 1'b0 ;
  assign n38914 = n3908 & n38913 ;
  assign n38916 = n38915 ^ n38914 ^ n16157 ;
  assign n38917 = n15241 | n18776 ;
  assign n38918 = n33584 | n38917 ;
  assign n38919 = n32627 ^ n1476 ^ 1'b0 ;
  assign n38920 = n11935 & n38919 ;
  assign n38926 = n16635 ^ n12281 ^ n2221 ;
  assign n38927 = n36027 & ~n38926 ;
  assign n38922 = n9442 & n11306 ;
  assign n38923 = ~n3770 & n38922 ;
  assign n38921 = n37096 ^ n25284 ^ n20916 ;
  assign n38924 = n38923 ^ n38921 ^ n9959 ;
  assign n38925 = n38924 ^ n27478 ^ 1'b0 ;
  assign n38928 = n38927 ^ n38925 ^ 1'b0 ;
  assign n38929 = n31723 & n38928 ;
  assign n38933 = n18614 & n30922 ;
  assign n38930 = n12642 ^ n3779 ^ n263 ;
  assign n38931 = n38930 ^ n14412 ^ 1'b0 ;
  assign n38932 = n24278 & n38931 ;
  assign n38934 = n38933 ^ n38932 ^ 1'b0 ;
  assign n38935 = n11750 | n24474 ;
  assign n38936 = ~n36233 & n38935 ;
  assign n38937 = n6668 & n24941 ;
  assign n38938 = n38937 ^ n11825 ^ 1'b0 ;
  assign n38939 = n11919 ^ n9283 ^ n5110 ;
  assign n38940 = ( n19395 & n35428 ) | ( n19395 & ~n38939 ) | ( n35428 & ~n38939 ) ;
  assign n38941 = n4944 & ~n18913 ;
  assign n38942 = ~n23893 & n38941 ;
  assign n38943 = ( n993 & ~n2459 ) | ( n993 & n38942 ) | ( ~n2459 & n38942 ) ;
  assign n38944 = ( ~n27924 & n32879 ) | ( ~n27924 & n38943 ) | ( n32879 & n38943 ) ;
  assign n38945 = n14283 ^ n13555 ^ 1'b0 ;
  assign n38946 = n38945 ^ n14939 ^ 1'b0 ;
  assign n38947 = n27590 ^ n6827 ^ n1842 ;
  assign n38948 = n28317 & n38947 ;
  assign n38949 = n38948 ^ n1279 ^ 1'b0 ;
  assign n38950 = ~n2016 & n7781 ;
  assign n38951 = n38950 ^ n5203 ^ 1'b0 ;
  assign n38952 = n34118 ^ n26274 ^ n23974 ;
  assign n38953 = n3826 | n38952 ;
  assign n38954 = n38951 | n38953 ;
  assign n38955 = n38949 & n38954 ;
  assign n38956 = n11230 ^ n4113 ^ 1'b0 ;
  assign n38957 = n8582 | n38956 ;
  assign n38958 = ~n2782 & n38957 ;
  assign n38959 = ~n11236 & n25116 ;
  assign n38960 = n38959 ^ n1298 ^ 1'b0 ;
  assign n38961 = n24500 ^ n14895 ^ 1'b0 ;
  assign n38962 = n38960 & n38961 ;
  assign n38963 = n21472 & ~n31792 ;
  assign n38964 = n38963 ^ n5662 ^ 1'b0 ;
  assign n38965 = ( ~n3334 & n13639 ) | ( ~n3334 & n35696 ) | ( n13639 & n35696 ) ;
  assign n38966 = n32304 ^ n5684 ^ 1'b0 ;
  assign n38967 = ~n26338 & n38966 ;
  assign n38968 = ( n6546 & n38636 ) | ( n6546 & n38967 ) | ( n38636 & n38967 ) ;
  assign n38969 = n38400 | n38968 ;
  assign n38970 = n7319 ^ n3072 ^ n2408 ;
  assign n38971 = n2910 & ~n20309 ;
  assign n38972 = ( n945 & n3290 ) | ( n945 & ~n18172 ) | ( n3290 & ~n18172 ) ;
  assign n38973 = ( n12471 & ~n38971 ) | ( n12471 & n38972 ) | ( ~n38971 & n38972 ) ;
  assign n38974 = ( n7786 & n38970 ) | ( n7786 & n38973 ) | ( n38970 & n38973 ) ;
  assign n38975 = ( n2059 & ~n3555 ) | ( n2059 & n29086 ) | ( ~n3555 & n29086 ) ;
  assign n38976 = n13458 & ~n38975 ;
  assign n38977 = n23174 ^ n19394 ^ n16542 ;
  assign n38978 = ( ~n19346 & n20038 ) | ( ~n19346 & n35293 ) | ( n20038 & n35293 ) ;
  assign n38979 = ( ~n11158 & n15840 ) | ( ~n11158 & n27369 ) | ( n15840 & n27369 ) ;
  assign n38980 = n6593 | n24868 ;
  assign n38981 = n11423 & ~n38980 ;
  assign n38982 = n21836 ^ n7696 ^ n2273 ;
  assign n38983 = n5054 & n38982 ;
  assign n38984 = ~n9601 & n38983 ;
  assign n38985 = n32581 ^ n10783 ^ n8095 ;
  assign n38986 = ( ~n12095 & n38984 ) | ( ~n12095 & n38985 ) | ( n38984 & n38985 ) ;
  assign n38987 = ( n9686 & ~n23721 ) | ( n9686 & n30192 ) | ( ~n23721 & n30192 ) ;
  assign n38988 = ( n8038 & n27956 ) | ( n8038 & n38987 ) | ( n27956 & n38987 ) ;
  assign n38989 = ( n3097 & n15146 ) | ( n3097 & ~n30587 ) | ( n15146 & ~n30587 ) ;
  assign n38991 = n38306 ^ n14687 ^ n3053 ;
  assign n38990 = n34229 ^ n30311 ^ n6029 ;
  assign n38992 = n38991 ^ n38990 ^ n21834 ;
  assign n38993 = n30297 ^ n16558 ^ 1'b0 ;
  assign n38994 = n8964 & n38993 ;
  assign n38995 = ( n8772 & n23183 ) | ( n8772 & n25034 ) | ( n23183 & n25034 ) ;
  assign n38996 = ( n7462 & n11667 ) | ( n7462 & n23620 ) | ( n11667 & n23620 ) ;
  assign n38997 = ( n25367 & ~n33880 ) | ( n25367 & n38996 ) | ( ~n33880 & n38996 ) ;
  assign n38998 = n38997 ^ n21570 ^ 1'b0 ;
  assign n38999 = n38995 | n38998 ;
  assign n39000 = ( n7558 & ~n7761 ) | ( n7558 & n30385 ) | ( ~n7761 & n30385 ) ;
  assign n39002 = ( ~n3115 & n5202 ) | ( ~n3115 & n13688 ) | ( n5202 & n13688 ) ;
  assign n39003 = n15542 ^ n7817 ^ 1'b0 ;
  assign n39004 = x240 & ~n39003 ;
  assign n39005 = ( n7242 & ~n39002 ) | ( n7242 & n39004 ) | ( ~n39002 & n39004 ) ;
  assign n39001 = n17014 ^ n15497 ^ 1'b0 ;
  assign n39006 = n39005 ^ n39001 ^ n28148 ;
  assign n39009 = n3768 ^ n2800 ^ 1'b0 ;
  assign n39007 = n9618 ^ n6099 ^ n5909 ;
  assign n39008 = ( n1968 & n12834 ) | ( n1968 & n39007 ) | ( n12834 & n39007 ) ;
  assign n39010 = n39009 ^ n39008 ^ n32926 ;
  assign n39011 = n15896 ^ n7678 ^ n6794 ;
  assign n39012 = ~n26010 & n39011 ;
  assign n39013 = n39012 ^ n17140 ^ 1'b0 ;
  assign n39015 = n26924 ^ n24652 ^ n7273 ;
  assign n39014 = ~n9643 & n28403 ;
  assign n39016 = n39015 ^ n39014 ^ 1'b0 ;
  assign n39017 = ( n5463 & ~n18518 ) | ( n5463 & n27232 ) | ( ~n18518 & n27232 ) ;
  assign n39018 = n31587 | n39017 ;
  assign n39019 = n2418 & ~n26615 ;
  assign n39020 = ~n15664 & n39019 ;
  assign n39021 = n39020 ^ n33634 ^ 1'b0 ;
  assign n39022 = ~n30089 & n32005 ;
  assign n39023 = n39022 ^ n37595 ^ 1'b0 ;
  assign n39024 = ( n11447 & n18789 ) | ( n11447 & ~n39023 ) | ( n18789 & ~n39023 ) ;
  assign n39025 = n33203 ^ n18037 ^ 1'b0 ;
  assign n39026 = ( n3211 & n13773 ) | ( n3211 & n17365 ) | ( n13773 & n17365 ) ;
  assign n39027 = ~n5661 & n39026 ;
  assign n39028 = ( n13883 & n23170 ) | ( n13883 & ~n29998 ) | ( n23170 & ~n29998 ) ;
  assign n39029 = n31037 & ~n32726 ;
  assign n39030 = ~n854 & n39029 ;
  assign n39031 = n18018 | n33105 ;
  assign n39032 = ~n22108 & n33613 ;
  assign n39033 = n33950 & n39032 ;
  assign n39034 = n39033 ^ n31698 ^ n21395 ;
  assign n39035 = ( n3690 & n12236 ) | ( n3690 & ~n17613 ) | ( n12236 & ~n17613 ) ;
  assign n39036 = ( n5961 & n20510 ) | ( n5961 & ~n39035 ) | ( n20510 & ~n39035 ) ;
  assign n39037 = ( ~n13645 & n17392 ) | ( ~n13645 & n39036 ) | ( n17392 & n39036 ) ;
  assign n39038 = n5387 | n5722 ;
  assign n39039 = n28861 & ~n39038 ;
  assign n39040 = n38878 ^ n5701 ^ n384 ;
  assign n39041 = n14243 | n20589 ;
  assign n39042 = n3025 & n16999 ;
  assign n39043 = n39042 ^ n11527 ^ 1'b0 ;
  assign n39044 = ( n14931 & ~n25637 ) | ( n14931 & n39043 ) | ( ~n25637 & n39043 ) ;
  assign n39045 = n39044 ^ n24927 ^ 1'b0 ;
  assign n39046 = n32078 ^ n25336 ^ n24395 ;
  assign n39049 = n7537 ^ n3217 ^ n837 ;
  assign n39047 = n12948 ^ n9506 ^ n3331 ;
  assign n39048 = n39047 ^ n34242 ^ n8268 ;
  assign n39050 = n39049 ^ n39048 ^ n24083 ;
  assign n39051 = ( n28001 & n39046 ) | ( n28001 & ~n39050 ) | ( n39046 & ~n39050 ) ;
  assign n39052 = n7379 & n10448 ;
  assign n39053 = n39052 ^ n19844 ^ n1101 ;
  assign n39054 = n13291 | n39053 ;
  assign n39055 = n39054 ^ n20715 ^ 1'b0 ;
  assign n39056 = n39055 ^ n14582 ^ 1'b0 ;
  assign n39057 = n39051 | n39056 ;
  assign n39058 = n2617 & n7403 ;
  assign n39059 = n28242 & n39058 ;
  assign n39060 = n21661 ^ n19548 ^ n1080 ;
  assign n39061 = n13576 ^ n4935 ^ 1'b0 ;
  assign n39062 = n39060 & ~n39061 ;
  assign n39063 = ~n20693 & n39062 ;
  assign n39064 = n39063 ^ n11031 ^ 1'b0 ;
  assign n39065 = n39064 ^ n25227 ^ n9616 ;
  assign n39066 = ( ~n9778 & n13061 ) | ( ~n9778 & n17492 ) | ( n13061 & n17492 ) ;
  assign n39067 = ( n17203 & n21055 ) | ( n17203 & ~n39066 ) | ( n21055 & ~n39066 ) ;
  assign n39068 = n39067 ^ n17508 ^ 1'b0 ;
  assign n39069 = n19038 ^ n15881 ^ 1'b0 ;
  assign n39070 = n39069 ^ n17626 ^ n17056 ;
  assign n39071 = ( ~n6564 & n18541 ) | ( ~n6564 & n22555 ) | ( n18541 & n22555 ) ;
  assign n39072 = n11697 ^ n9908 ^ n922 ;
  assign n39073 = n39072 ^ n33708 ^ n23634 ;
  assign n39074 = ( ~x5 & n13849 ) | ( ~x5 & n31762 ) | ( n13849 & n31762 ) ;
  assign n39075 = n11291 ^ n3430 ^ 1'b0 ;
  assign n39076 = n39074 & ~n39075 ;
  assign n39077 = n1438 & ~n8532 ;
  assign n39079 = n19352 ^ n9877 ^ n7295 ;
  assign n39078 = n18253 ^ n8918 ^ n4582 ;
  assign n39080 = n39079 ^ n39078 ^ n33766 ;
  assign n39081 = n25109 ^ n19101 ^ n2506 ;
  assign n39082 = n20747 | n39081 ;
  assign n39083 = ~n8014 & n36414 ;
  assign n39084 = n39083 ^ n4122 ^ 1'b0 ;
  assign n39085 = n39084 ^ n16770 ^ n11754 ;
  assign n39086 = n32361 ^ n31485 ^ n25694 ;
  assign n39087 = n39086 ^ n35910 ^ n21419 ;
  assign n39088 = ( n11330 & n39085 ) | ( n11330 & n39087 ) | ( n39085 & n39087 ) ;
  assign n39089 = n3646 & ~n13957 ;
  assign n39090 = n39089 ^ n37262 ^ n4792 ;
  assign n39091 = ( n805 & n1668 ) | ( n805 & n8337 ) | ( n1668 & n8337 ) ;
  assign n39094 = n23522 ^ n15637 ^ 1'b0 ;
  assign n39092 = n9298 ^ n6340 ^ 1'b0 ;
  assign n39093 = ( n2962 & n22490 ) | ( n2962 & ~n39092 ) | ( n22490 & ~n39092 ) ;
  assign n39095 = n39094 ^ n39093 ^ n9232 ;
  assign n39096 = ( n26495 & n39091 ) | ( n26495 & ~n39095 ) | ( n39091 & ~n39095 ) ;
  assign n39098 = n13244 ^ n3264 ^ 1'b0 ;
  assign n39099 = ~n10010 & n39098 ;
  assign n39097 = ~n16731 & n17473 ;
  assign n39100 = n39099 ^ n39097 ^ 1'b0 ;
  assign n39101 = n3707 & ~n11493 ;
  assign n39102 = ( n19088 & ~n25131 ) | ( n19088 & n27199 ) | ( ~n25131 & n27199 ) ;
  assign n39103 = ( n10912 & n13634 ) | ( n10912 & n14907 ) | ( n13634 & n14907 ) ;
  assign n39104 = n15572 ^ n2326 ^ 1'b0 ;
  assign n39105 = n39103 | n39104 ;
  assign n39106 = n39105 ^ n17398 ^ 1'b0 ;
  assign n39107 = n26190 ^ n18518 ^ 1'b0 ;
  assign n39108 = ~n2863 & n39107 ;
  assign n39109 = n28854 ^ n24910 ^ n13866 ;
  assign n39110 = n39109 ^ n25505 ^ n24737 ;
  assign n39111 = ( ~n404 & n12727 ) | ( ~n404 & n16474 ) | ( n12727 & n16474 ) ;
  assign n39112 = n13758 ^ n10369 ^ n3888 ;
  assign n39113 = n21503 ^ n4675 ^ 1'b0 ;
  assign n39114 = ( n39111 & ~n39112 ) | ( n39111 & n39113 ) | ( ~n39112 & n39113 ) ;
  assign n39115 = n26176 ^ n6587 ^ n1553 ;
  assign n39116 = n39115 ^ n38464 ^ x120 ;
  assign n39117 = ( n3170 & n12909 ) | ( n3170 & ~n39116 ) | ( n12909 & ~n39116 ) ;
  assign n39118 = n22286 ^ n19893 ^ n16161 ;
  assign n39119 = n15744 ^ n546 ^ 1'b0 ;
  assign n39120 = n39118 | n39119 ;
  assign n39121 = n39120 ^ n28744 ^ n4151 ;
  assign n39122 = ( n6507 & n34723 ) | ( n6507 & n39121 ) | ( n34723 & n39121 ) ;
  assign n39123 = n16006 ^ n7856 ^ n2441 ;
  assign n39124 = n14675 & ~n17450 ;
  assign n39125 = n28684 ^ n27996 ^ 1'b0 ;
  assign n39126 = ~n9729 & n12992 ;
  assign n39127 = n37556 & n39126 ;
  assign n39128 = n23646 & ~n39127 ;
  assign n39129 = n11862 & n39128 ;
  assign n39130 = n6766 | n14411 ;
  assign n39131 = n30942 ^ n19867 ^ 1'b0 ;
  assign n39132 = ( n12357 & n13597 ) | ( n12357 & ~n39131 ) | ( n13597 & ~n39131 ) ;
  assign n39133 = n32428 ^ n12062 ^ n6251 ;
  assign n39134 = ( n19469 & n34438 ) | ( n19469 & ~n39133 ) | ( n34438 & ~n39133 ) ;
  assign n39135 = ( ~n3139 & n16343 ) | ( ~n3139 & n28471 ) | ( n16343 & n28471 ) ;
  assign n39136 = n10529 & ~n21842 ;
  assign n39137 = n34563 & n39136 ;
  assign n39138 = n28025 & ~n39137 ;
  assign n39139 = ~n13251 & n39138 ;
  assign n39140 = ( ~n32752 & n39135 ) | ( ~n32752 & n39139 ) | ( n39135 & n39139 ) ;
  assign n39141 = n16006 & ~n36215 ;
  assign n39142 = n39141 ^ n23821 ^ 1'b0 ;
  assign n39143 = n26399 ^ n17224 ^ n13233 ;
  assign n39144 = n15728 ^ n4743 ^ n2810 ;
  assign n39145 = ( ~n6612 & n28715 ) | ( ~n6612 & n39144 ) | ( n28715 & n39144 ) ;
  assign n39147 = n37963 ^ n3014 ^ n2844 ;
  assign n39146 = n20090 ^ n19228 ^ n1113 ;
  assign n39148 = n39147 ^ n39146 ^ 1'b0 ;
  assign n39149 = ( n522 & ~n5113 ) | ( n522 & n14471 ) | ( ~n5113 & n14471 ) ;
  assign n39150 = n11968 ^ n1352 ^ 1'b0 ;
  assign n39151 = ~n39149 & n39150 ;
  assign n39155 = ( n9885 & n11221 ) | ( n9885 & ~n24586 ) | ( n11221 & ~n24586 ) ;
  assign n39153 = n6433 ^ n1007 ^ n352 ;
  assign n39152 = ~n17348 & n17509 ;
  assign n39154 = n39153 ^ n39152 ^ 1'b0 ;
  assign n39156 = n39155 ^ n39154 ^ n25719 ;
  assign n39158 = ( n4212 & ~n5624 ) | ( n4212 & n7885 ) | ( ~n5624 & n7885 ) ;
  assign n39157 = n13118 & ~n19250 ;
  assign n39159 = n39158 ^ n39157 ^ 1'b0 ;
  assign n39160 = ( ~n3797 & n7883 ) | ( ~n3797 & n10994 ) | ( n7883 & n10994 ) ;
  assign n39161 = n31291 ^ n23499 ^ n13050 ;
  assign n39162 = ( n14502 & n30980 ) | ( n14502 & ~n39161 ) | ( n30980 & ~n39161 ) ;
  assign n39163 = ( n39159 & n39160 ) | ( n39159 & n39162 ) | ( n39160 & n39162 ) ;
  assign n39164 = n21832 ^ n18615 ^ 1'b0 ;
  assign n39165 = n455 | n39164 ;
  assign n39166 = ( ~n7699 & n29889 ) | ( ~n7699 & n39165 ) | ( n29889 & n39165 ) ;
  assign n39167 = n39166 ^ n4433 ^ 1'b0 ;
  assign n39168 = n15361 ^ n10753 ^ n264 ;
  assign n39169 = n9964 & ~n17983 ;
  assign n39170 = ~n39168 & n39169 ;
  assign n39171 = n33412 ^ n27334 ^ n20585 ;
  assign n39172 = n32796 ^ n13012 ^ n11261 ;
  assign n39173 = ( n9289 & n29288 ) | ( n9289 & ~n39172 ) | ( n29288 & ~n39172 ) ;
  assign n39174 = ( ~n1456 & n21355 ) | ( ~n1456 & n21426 ) | ( n21355 & n21426 ) ;
  assign n39175 = ( n16201 & n21140 ) | ( n16201 & ~n39174 ) | ( n21140 & ~n39174 ) ;
  assign n39176 = n39175 ^ n12559 ^ n1896 ;
  assign n39177 = n34599 ^ n1042 ^ 1'b0 ;
  assign n39178 = ~n11408 & n18823 ;
  assign n39179 = n5037 | n26478 ;
  assign n39180 = n2003 & ~n39179 ;
  assign n39181 = n5341 & n16477 ;
  assign n39182 = n39181 ^ n13740 ^ n4288 ;
  assign n39183 = n22890 ^ n10428 ^ 1'b0 ;
  assign n39184 = n20532 & n39183 ;
  assign n39185 = n39184 ^ n11011 ^ n10943 ;
  assign n39186 = n38129 ^ n12203 ^ 1'b0 ;
  assign n39187 = n39186 ^ n37094 ^ 1'b0 ;
  assign n39188 = ( ~n16769 & n17098 ) | ( ~n16769 & n21232 ) | ( n17098 & n21232 ) ;
  assign n39189 = n9363 | n19395 ;
  assign n39190 = n11913 ^ n11828 ^ 1'b0 ;
  assign n39191 = n12912 & ~n39190 ;
  assign n39192 = n39191 ^ n2137 ^ 1'b0 ;
  assign n39193 = ~n30558 & n39192 ;
  assign n39194 = n39193 ^ n8387 ^ 1'b0 ;
  assign n39195 = ~n39189 & n39194 ;
  assign n39196 = n14583 ^ n13683 ^ n8283 ;
  assign n39197 = n2476 | n39196 ;
  assign n39198 = ( n19804 & n31232 ) | ( n19804 & ~n39197 ) | ( n31232 & ~n39197 ) ;
  assign n39199 = ~n11373 & n15845 ;
  assign n39200 = ~n9848 & n39199 ;
  assign n39201 = n12903 & n39200 ;
  assign n39202 = n39201 ^ n33949 ^ 1'b0 ;
  assign n39203 = n39198 & ~n39202 ;
  assign n39205 = n6591 ^ n918 ^ 1'b0 ;
  assign n39204 = n5687 & n37760 ;
  assign n39206 = n39205 ^ n39204 ^ n28330 ;
  assign n39207 = n30361 & ~n39206 ;
  assign n39208 = n39207 ^ n1745 ^ 1'b0 ;
  assign n39209 = n9963 & ~n27053 ;
  assign n39210 = n39208 & n39209 ;
  assign n39213 = n12097 ^ n3731 ^ n2956 ;
  assign n39214 = n39213 ^ n7252 ^ 1'b0 ;
  assign n39215 = n3553 & ~n39214 ;
  assign n39211 = ( n11124 & n14838 ) | ( n11124 & ~n16814 ) | ( n14838 & ~n16814 ) ;
  assign n39212 = n39211 ^ n11347 ^ n3837 ;
  assign n39216 = n39215 ^ n39212 ^ n35398 ;
  assign n39217 = n26571 ^ n6705 ^ 1'b0 ;
  assign n39218 = n29854 & ~n39217 ;
  assign n39219 = n39218 ^ n9972 ^ n4544 ;
  assign n39220 = n32769 ^ n7642 ^ n2278 ;
  assign n39228 = n21216 ^ n11985 ^ n6663 ;
  assign n39222 = n6329 ^ n5896 ^ 1'b0 ;
  assign n39221 = n8740 & n17762 ;
  assign n39223 = n39222 ^ n39221 ^ 1'b0 ;
  assign n39224 = n39223 ^ n8490 ^ 1'b0 ;
  assign n39225 = n13137 & ~n39224 ;
  assign n39226 = ( n14179 & n21252 ) | ( n14179 & n37073 ) | ( n21252 & n37073 ) ;
  assign n39227 = ( n1185 & ~n39225 ) | ( n1185 & n39226 ) | ( ~n39225 & n39226 ) ;
  assign n39229 = n39228 ^ n39227 ^ n28561 ;
  assign n39230 = n10425 & n39229 ;
  assign n39231 = n39230 ^ n12151 ^ 1'b0 ;
  assign n39232 = n35477 ^ n31893 ^ n12483 ;
  assign n39233 = ( ~n658 & n15029 ) | ( ~n658 & n23281 ) | ( n15029 & n23281 ) ;
  assign n39234 = n39233 ^ n38762 ^ n3532 ;
  assign n39237 = ( ~n351 & n9598 ) | ( ~n351 & n34857 ) | ( n9598 & n34857 ) ;
  assign n39235 = n6960 & ~n23881 ;
  assign n39236 = n18938 & n39235 ;
  assign n39238 = n39237 ^ n39236 ^ 1'b0 ;
  assign n39239 = n37657 ^ n19020 ^ 1'b0 ;
  assign n39240 = n15033 ^ n4291 ^ n2147 ;
  assign n39241 = ( ~n15029 & n15287 ) | ( ~n15029 & n39240 ) | ( n15287 & n39240 ) ;
  assign n39242 = ~n23217 & n23470 ;
  assign n39243 = ~n5311 & n39242 ;
  assign n39244 = ( x35 & ~n39241 ) | ( x35 & n39243 ) | ( ~n39241 & n39243 ) ;
  assign n39245 = n39244 ^ n38436 ^ n4831 ;
  assign n39246 = n27999 ^ n22933 ^ 1'b0 ;
  assign n39247 = n29373 & ~n39246 ;
  assign n39248 = n39247 ^ n12521 ^ 1'b0 ;
  assign n39249 = ( n29299 & ~n38326 ) | ( n29299 & n38786 ) | ( ~n38326 & n38786 ) ;
  assign n39250 = ( n18331 & ~n36073 ) | ( n18331 & n39249 ) | ( ~n36073 & n39249 ) ;
  assign n39251 = n39250 ^ n8669 ^ 1'b0 ;
  assign n39255 = ( n9917 & ~n12070 ) | ( n9917 & n35644 ) | ( ~n12070 & n35644 ) ;
  assign n39256 = n39255 ^ n6336 ^ n5065 ;
  assign n39252 = ~x99 & n2719 ;
  assign n39253 = n39252 ^ n32919 ^ 1'b0 ;
  assign n39254 = n39253 ^ n34452 ^ n28647 ;
  assign n39257 = n39256 ^ n39254 ^ n22202 ;
  assign n39258 = ~n3019 & n12003 ;
  assign n39259 = n38681 ^ n31830 ^ n25140 ;
  assign n39260 = ( ~n29187 & n39258 ) | ( ~n29187 & n39259 ) | ( n39258 & n39259 ) ;
  assign n39261 = n39260 ^ n22136 ^ 1'b0 ;
  assign n39262 = ~n8657 & n36325 ;
  assign n39263 = n39262 ^ n4506 ^ 1'b0 ;
  assign n39264 = n24351 ^ n21715 ^ 1'b0 ;
  assign n39265 = n21119 | n39264 ;
  assign n39266 = n28093 ^ n14487 ^ 1'b0 ;
  assign n39267 = n30161 & ~n35728 ;
  assign n39268 = ~n39266 & n39267 ;
  assign n39269 = n30844 ^ n22802 ^ n4269 ;
  assign n39270 = n39269 ^ n35783 ^ 1'b0 ;
  assign n39271 = n27390 ^ n15435 ^ n14757 ;
  assign n39274 = ( n6706 & ~n9603 ) | ( n6706 & n16683 ) | ( ~n9603 & n16683 ) ;
  assign n39272 = n4398 | n7944 ;
  assign n39273 = n39272 ^ n27023 ^ n1307 ;
  assign n39275 = n39274 ^ n39273 ^ n35971 ;
  assign n39276 = n2622 & ~n24435 ;
  assign n39277 = n39276 ^ n1695 ^ 1'b0 ;
  assign n39278 = n2435 & ~n34599 ;
  assign n39279 = ~n1024 & n39278 ;
  assign n39280 = n28174 & ~n39279 ;
  assign n39281 = ~n25036 & n39280 ;
  assign n39283 = n1769 & ~n3653 ;
  assign n39282 = n14799 ^ n9775 ^ n8617 ;
  assign n39284 = n39283 ^ n39282 ^ n12230 ;
  assign n39285 = ( n18243 & n18260 ) | ( n18243 & ~n20635 ) | ( n18260 & ~n20635 ) ;
  assign n39286 = ( ~n23216 & n30911 ) | ( ~n23216 & n39285 ) | ( n30911 & n39285 ) ;
  assign n39287 = n17752 ^ x184 ^ 1'b0 ;
  assign n39288 = n24093 & ~n39287 ;
  assign n39289 = n8578 ^ n5628 ^ 1'b0 ;
  assign n39290 = n34660 ^ n9637 ^ 1'b0 ;
  assign n39291 = n29682 ^ n18335 ^ n3853 ;
  assign n39292 = n4252 & n39291 ;
  assign n39293 = n10175 | n15343 ;
  assign n39294 = n29240 & ~n39293 ;
  assign n39295 = n8004 | n16880 ;
  assign n39296 = n19590 & ~n39295 ;
  assign n39297 = n29759 ^ n15054 ^ n1962 ;
  assign n39298 = n27604 ^ n22071 ^ 1'b0 ;
  assign n39299 = n39297 & ~n39298 ;
  assign n39300 = ( n7957 & ~n23163 ) | ( n7957 & n27431 ) | ( ~n23163 & n27431 ) ;
  assign n39303 = ( n4815 & n4993 ) | ( n4815 & n7181 ) | ( n4993 & n7181 ) ;
  assign n39302 = n33880 ^ n9141 ^ n486 ;
  assign n39304 = n39303 ^ n39302 ^ n8398 ;
  assign n39305 = n39304 ^ n15411 ^ n11269 ;
  assign n39301 = ~n4256 & n18781 ;
  assign n39306 = n39305 ^ n39301 ^ n26444 ;
  assign n39307 = ( n4116 & n12902 ) | ( n4116 & n22982 ) | ( n12902 & n22982 ) ;
  assign n39311 = n21099 ^ n5991 ^ n2198 ;
  assign n39309 = ( n12143 & n15592 ) | ( n12143 & n17465 ) | ( n15592 & n17465 ) ;
  assign n39308 = n27358 ^ n13026 ^ n5469 ;
  assign n39310 = n39309 ^ n39308 ^ n14137 ;
  assign n39312 = n39311 ^ n39310 ^ n28162 ;
  assign n39313 = x152 & ~n24466 ;
  assign n39314 = ~n7910 & n39313 ;
  assign n39315 = ~n15619 & n39314 ;
  assign n39316 = ( n24318 & n26608 ) | ( n24318 & ~n39315 ) | ( n26608 & ~n39315 ) ;
  assign n39317 = ~n19855 & n21212 ;
  assign n39318 = n13335 | n29359 ;
  assign n39319 = n39318 ^ n9179 ^ 1'b0 ;
  assign n39320 = n16551 & ~n34022 ;
  assign n39321 = ( x109 & n18221 ) | ( x109 & ~n26131 ) | ( n18221 & ~n26131 ) ;
  assign n39322 = n31477 ^ n16741 ^ n2926 ;
  assign n39323 = ( ~n5465 & n17188 ) | ( ~n5465 & n37612 ) | ( n17188 & n37612 ) ;
  assign n39324 = ( ~n37635 & n39322 ) | ( ~n37635 & n39323 ) | ( n39322 & n39323 ) ;
  assign n39325 = ( n28300 & n36420 ) | ( n28300 & n39324 ) | ( n36420 & n39324 ) ;
  assign n39326 = n15866 ^ n9949 ^ n5017 ;
  assign n39327 = n23164 | n39326 ;
  assign n39328 = ( ~n6650 & n11155 ) | ( ~n6650 & n34807 ) | ( n11155 & n34807 ) ;
  assign n39329 = ( ~n8090 & n22779 ) | ( ~n8090 & n39328 ) | ( n22779 & n39328 ) ;
  assign n39330 = ~n3828 & n15552 ;
  assign n39331 = n39330 ^ n32123 ^ 1'b0 ;
  assign n39332 = ~n6236 & n21992 ;
  assign n39333 = n31170 ^ n17423 ^ n6277 ;
  assign n39334 = ( x202 & n39332 ) | ( x202 & ~n39333 ) | ( n39332 & ~n39333 ) ;
  assign n39335 = n39334 ^ n29472 ^ n2691 ;
  assign n39336 = n2103 | n35934 ;
  assign n39337 = n39336 ^ n5296 ^ 1'b0 ;
  assign n39339 = n6973 ^ n6317 ^ n3701 ;
  assign n39338 = n15600 ^ n2640 ^ 1'b0 ;
  assign n39340 = n39339 ^ n39338 ^ n28664 ;
  assign n39341 = n39340 ^ n11636 ^ n5698 ;
  assign n39342 = ( ~n10422 & n13007 ) | ( ~n10422 & n32214 ) | ( n13007 & n32214 ) ;
  assign n39343 = n27832 | n39342 ;
  assign n39344 = n39343 ^ n15281 ^ 1'b0 ;
  assign n39345 = ( n11716 & n31948 ) | ( n11716 & n39344 ) | ( n31948 & n39344 ) ;
  assign n39346 = n29740 ^ n23949 ^ n11546 ;
  assign n39347 = n25704 ^ n9482 ^ n3178 ;
  assign n39348 = n37657 ^ n21537 ^ n1583 ;
  assign n39349 = ( ~n13675 & n16618 ) | ( ~n13675 & n39348 ) | ( n16618 & n39348 ) ;
  assign n39350 = n28014 ^ n21199 ^ n9965 ;
  assign n39351 = n28511 ^ n948 ^ 1'b0 ;
  assign n39352 = n39350 | n39351 ;
  assign n39353 = n2414 | n36828 ;
  assign n39354 = n39353 ^ n10318 ^ 1'b0 ;
  assign n39355 = n39352 & n39354 ;
  assign n39356 = n27094 ^ n24863 ^ n4804 ;
  assign n39357 = n10111 & ~n39356 ;
  assign n39359 = ( n1869 & ~n6054 ) | ( n1869 & n17604 ) | ( ~n6054 & n17604 ) ;
  assign n39358 = ( n2490 & n3410 ) | ( n2490 & ~n18321 ) | ( n3410 & ~n18321 ) ;
  assign n39360 = n39359 ^ n39358 ^ 1'b0 ;
  assign n39361 = ( n4859 & n13063 ) | ( n4859 & ~n39360 ) | ( n13063 & ~n39360 ) ;
  assign n39362 = n35860 & n39361 ;
  assign n39363 = n39362 ^ n32342 ^ 1'b0 ;
  assign n39364 = ( n5577 & ~n28908 ) | ( n5577 & n32599 ) | ( ~n28908 & n32599 ) ;
  assign n39365 = ( n14192 & n26831 ) | ( n14192 & ~n30477 ) | ( n26831 & ~n30477 ) ;
  assign n39366 = n30444 ^ n5786 ^ 1'b0 ;
  assign n39367 = n23871 ^ n21119 ^ n18377 ;
  assign n39368 = n39367 ^ n25728 ^ n14110 ;
  assign n39369 = ( ~n29734 & n39366 ) | ( ~n29734 & n39368 ) | ( n39366 & n39368 ) ;
  assign n39374 = ( n6937 & n7979 ) | ( n6937 & ~n8941 ) | ( n7979 & ~n8941 ) ;
  assign n39371 = n4319 | n6079 ;
  assign n39372 = x99 | n39371 ;
  assign n39373 = ( n14090 & ~n25383 ) | ( n14090 & n39372 ) | ( ~n25383 & n39372 ) ;
  assign n39370 = n22494 ^ n5267 ^ n3969 ;
  assign n39375 = n39374 ^ n39373 ^ n39370 ;
  assign n39376 = ( x200 & ~n1823 ) | ( x200 & n11291 ) | ( ~n1823 & n11291 ) ;
  assign n39377 = n39376 ^ n4654 ^ 1'b0 ;
  assign n39378 = n39377 ^ n20370 ^ 1'b0 ;
  assign n39379 = ( n279 & n8035 ) | ( n279 & ~n13425 ) | ( n8035 & ~n13425 ) ;
  assign n39380 = n2195 & n39379 ;
  assign n39381 = n21629 ^ n20554 ^ n5078 ;
  assign n39382 = n27017 & ~n27179 ;
  assign n39383 = n39382 ^ n6173 ^ 1'b0 ;
  assign n39384 = n39381 | n39383 ;
  assign n39385 = ~n11373 & n21788 ;
  assign n39386 = ~n9554 & n39385 ;
  assign n39387 = ( n1002 & n19047 ) | ( n1002 & n39386 ) | ( n19047 & n39386 ) ;
  assign n39388 = n16287 ^ n15148 ^ n1720 ;
  assign n39389 = ( n1315 & n1902 ) | ( n1315 & n1915 ) | ( n1902 & n1915 ) ;
  assign n39390 = n39389 ^ n26820 ^ n13613 ;
  assign n39392 = n28001 ^ n599 ^ 1'b0 ;
  assign n39391 = n8223 ^ n7155 ^ 1'b0 ;
  assign n39393 = n39392 ^ n39391 ^ n24440 ;
  assign n39394 = ( n8143 & ~n12850 ) | ( n8143 & n29847 ) | ( ~n12850 & n29847 ) ;
  assign n39395 = n39394 ^ n6724 ^ n4108 ;
  assign n39396 = n23419 ^ n11537 ^ 1'b0 ;
  assign n39397 = n2533 & n39396 ;
  assign n39398 = n1771 ^ n1016 ^ 1'b0 ;
  assign n39399 = ( n27444 & n39397 ) | ( n27444 & ~n39398 ) | ( n39397 & ~n39398 ) ;
  assign n39400 = n27192 ^ n2995 ^ n655 ;
  assign n39401 = n9948 & n20520 ;
  assign n39402 = n39401 ^ n4000 ^ 1'b0 ;
  assign n39403 = ( n6831 & ~n10331 ) | ( n6831 & n20580 ) | ( ~n10331 & n20580 ) ;
  assign n39404 = n39403 ^ n12318 ^ n7160 ;
  assign n39405 = n6926 ^ n2930 ^ n1214 ;
  assign n39406 = ~n14883 & n35316 ;
  assign n39407 = ~n39405 & n39406 ;
  assign n39408 = n11048 & n39407 ;
  assign n39409 = n16181 ^ n12680 ^ n4673 ;
  assign n39410 = n6243 | n28243 ;
  assign n39411 = n11393 | n39410 ;
  assign n39412 = n9114 ^ n6613 ^ n5311 ;
  assign n39413 = ( ~n16146 & n39411 ) | ( ~n16146 & n39412 ) | ( n39411 & n39412 ) ;
  assign n39414 = ( n9113 & n9895 ) | ( n9113 & n23993 ) | ( n9895 & n23993 ) ;
  assign n39415 = n10548 & ~n39414 ;
  assign n39416 = ~n39413 & n39415 ;
  assign n39417 = n15503 ^ n15030 ^ 1'b0 ;
  assign n39418 = n4527 & ~n39417 ;
  assign n39419 = n11971 | n39418 ;
  assign n39420 = n5071 ^ n2697 ^ 1'b0 ;
  assign n39421 = n2105 | n39420 ;
  assign n39422 = ( n5813 & n16154 ) | ( n5813 & ~n39421 ) | ( n16154 & ~n39421 ) ;
  assign n39423 = n24768 ^ n17678 ^ 1'b0 ;
  assign n39424 = ( n1714 & n27438 ) | ( n1714 & n39423 ) | ( n27438 & n39423 ) ;
  assign n39425 = n36087 ^ n17333 ^ n6859 ;
  assign n39426 = ~n11274 & n20702 ;
  assign n39427 = n39426 ^ n3291 ^ 1'b0 ;
  assign n39428 = n33315 & n39427 ;
  assign n39429 = n28521 ^ n17448 ^ n15446 ;
  assign n39430 = n2177 & n6690 ;
  assign n39431 = n1822 & n39430 ;
  assign n39432 = n39431 ^ n14662 ^ n11630 ;
  assign n39433 = n39432 ^ n3601 ^ x139 ;
  assign n39434 = x183 & ~n5939 ;
  assign n39435 = n39434 ^ n38722 ^ n9318 ;
  assign n39436 = ( n8881 & n12842 ) | ( n8881 & n23712 ) | ( n12842 & n23712 ) ;
  assign n39437 = n1449 ^ n1070 ^ 1'b0 ;
  assign n39438 = n5400 & n39437 ;
  assign n39439 = ( n8673 & n15023 ) | ( n8673 & n39438 ) | ( n15023 & n39438 ) ;
  assign n39440 = ( n23791 & n39359 ) | ( n23791 & ~n39439 ) | ( n39359 & ~n39439 ) ;
  assign n39441 = n28487 ^ n9012 ^ 1'b0 ;
  assign n39442 = n39441 ^ n7594 ^ n5445 ;
  assign n39443 = ( n16057 & ~n31832 ) | ( n16057 & n39442 ) | ( ~n31832 & n39442 ) ;
  assign n39444 = n5232 ^ n2668 ^ 1'b0 ;
  assign n39445 = n11824 & ~n39444 ;
  assign n39446 = n39445 ^ n21169 ^ n3117 ;
  assign n39447 = n39446 ^ n2169 ^ n2125 ;
  assign n39448 = n1269 | n6214 ;
  assign n39449 = n39448 ^ n24971 ^ 1'b0 ;
  assign n39450 = n14144 | n39449 ;
  assign n39451 = n39450 ^ n36722 ^ n23363 ;
  assign n39452 = n19412 | n37458 ;
  assign n39453 = n38511 ^ n15548 ^ 1'b0 ;
  assign n39454 = ( n39366 & n39452 ) | ( n39366 & ~n39453 ) | ( n39452 & ~n39453 ) ;
  assign n39458 = n23502 ^ n2437 ^ 1'b0 ;
  assign n39459 = n39458 ^ n10595 ^ 1'b0 ;
  assign n39460 = ( ~n20170 & n35577 ) | ( ~n20170 & n39459 ) | ( n35577 & n39459 ) ;
  assign n39455 = n28586 ^ n5194 ^ n1452 ;
  assign n39456 = ( n7525 & n8124 ) | ( n7525 & n39455 ) | ( n8124 & n39455 ) ;
  assign n39457 = ~n10231 & n39456 ;
  assign n39461 = n39460 ^ n39457 ^ 1'b0 ;
  assign n39462 = n2433 & n11859 ;
  assign n39463 = n23420 | n28719 ;
  assign n39464 = n3306 & ~n39463 ;
  assign n39465 = n10529 ^ n10164 ^ n6010 ;
  assign n39466 = n39465 ^ n14934 ^ 1'b0 ;
  assign n39467 = ( ~n3489 & n32453 ) | ( ~n3489 & n39466 ) | ( n32453 & n39466 ) ;
  assign n39468 = n39467 ^ n11603 ^ n4209 ;
  assign n39469 = ( ~n39462 & n39464 ) | ( ~n39462 & n39468 ) | ( n39464 & n39468 ) ;
  assign n39470 = n9452 & n21650 ;
  assign n39471 = n29120 ^ n7191 ^ 1'b0 ;
  assign n39472 = n29655 & ~n35167 ;
  assign n39473 = n17517 | n39472 ;
  assign n39474 = n34155 & ~n39473 ;
  assign n39475 = ( n4324 & n4997 ) | ( n4324 & ~n7143 ) | ( n4997 & ~n7143 ) ;
  assign n39476 = n6985 & ~n16532 ;
  assign n39477 = n2934 ^ n1628 ^ 1'b0 ;
  assign n39478 = n11385 & n39477 ;
  assign n39479 = ( n39475 & n39476 ) | ( n39475 & ~n39478 ) | ( n39476 & ~n39478 ) ;
  assign n39480 = n4066 & ~n35866 ;
  assign n39481 = n9570 & n39480 ;
  assign n39482 = ( ~n12859 & n13969 ) | ( ~n12859 & n21710 ) | ( n13969 & n21710 ) ;
  assign n39483 = ~n12786 & n22005 ;
  assign n39484 = n39483 ^ n16706 ^ 1'b0 ;
  assign n39485 = ( n39109 & n39482 ) | ( n39109 & n39484 ) | ( n39482 & n39484 ) ;
  assign n39486 = n16514 ^ n3626 ^ 1'b0 ;
  assign n39487 = ~n11789 & n39486 ;
  assign n39488 = ( n15541 & ~n33575 ) | ( n15541 & n39487 ) | ( ~n33575 & n39487 ) ;
  assign n39489 = ( n8726 & n22227 ) | ( n8726 & ~n33303 ) | ( n22227 & ~n33303 ) ;
  assign n39490 = n36224 ^ n29980 ^ n24236 ;
  assign n39491 = ( n15884 & ~n27705 ) | ( n15884 & n39259 ) | ( ~n27705 & n39259 ) ;
  assign n39492 = n1429 & ~n3826 ;
  assign n39493 = n1258 & n39492 ;
  assign n39494 = ( ~x18 & n4288 ) | ( ~x18 & n7476 ) | ( n4288 & n7476 ) ;
  assign n39495 = n39494 ^ n11304 ^ n2745 ;
  assign n39496 = n18274 & ~n39495 ;
  assign n39497 = n39496 ^ n21529 ^ 1'b0 ;
  assign n39498 = ( n2707 & n39493 ) | ( n2707 & n39497 ) | ( n39493 & n39497 ) ;
  assign n39499 = n39498 ^ n32081 ^ n1930 ;
  assign n39500 = n21075 ^ n14225 ^ n10743 ;
  assign n39501 = n39499 | n39500 ;
  assign n39502 = n5247 ^ x133 ^ 1'b0 ;
  assign n39503 = n20451 | n39502 ;
  assign n39504 = ( n4827 & n8273 ) | ( n4827 & n17082 ) | ( n8273 & n17082 ) ;
  assign n39505 = ~n15029 & n39504 ;
  assign n39506 = n39505 ^ n31484 ^ 1'b0 ;
  assign n39507 = n10862 ^ n6377 ^ 1'b0 ;
  assign n39508 = ~n9289 & n11146 ;
  assign n39509 = n39508 ^ n18636 ^ 1'b0 ;
  assign n39510 = ~n39507 & n39509 ;
  assign n39511 = n30498 ^ n6464 ^ n3492 ;
  assign n39512 = n39511 ^ n29857 ^ n4158 ;
  assign n39514 = n2546 & n22402 ;
  assign n39515 = n39514 ^ n8501 ^ 1'b0 ;
  assign n39513 = n19785 & ~n24604 ;
  assign n39516 = n39515 ^ n39513 ^ n33761 ;
  assign n39517 = n31698 & n39516 ;
  assign n39518 = n15947 & n39517 ;
  assign n39519 = ~n25870 & n39313 ;
  assign n39521 = n17352 ^ n9131 ^ n2342 ;
  assign n39520 = n20885 ^ n860 ^ n552 ;
  assign n39522 = n39521 ^ n39520 ^ n23472 ;
  assign n39523 = n27574 ^ n23483 ^ 1'b0 ;
  assign n39524 = n4502 ^ n2509 ^ 1'b0 ;
  assign n39525 = ~n3593 & n5354 ;
  assign n39526 = ~n36130 & n39525 ;
  assign n39527 = n39526 ^ n24337 ^ n11406 ;
  assign n39528 = ~n4498 & n39527 ;
  assign n39529 = ( n9986 & ~n12920 ) | ( n9986 & n39528 ) | ( ~n12920 & n39528 ) ;
  assign n39530 = ( n19785 & n21277 ) | ( n19785 & n31549 ) | ( n21277 & n31549 ) ;
  assign n39531 = n12986 ^ n6283 ^ n4198 ;
  assign n39532 = n21238 ^ n8887 ^ n8077 ;
  assign n39533 = n23780 & ~n31421 ;
  assign n39534 = ~n39532 & n39533 ;
  assign n39535 = n39531 & n39534 ;
  assign n39536 = ( n4311 & n30838 ) | ( n4311 & ~n39535 ) | ( n30838 & ~n39535 ) ;
  assign n39537 = ( n13205 & n39530 ) | ( n13205 & ~n39536 ) | ( n39530 & ~n39536 ) ;
  assign n39538 = n23989 & n39537 ;
  assign n39539 = n2589 ^ n1435 ^ x173 ;
  assign n39540 = n15839 & ~n39539 ;
  assign n39541 = ( n19477 & n29116 ) | ( n19477 & ~n36711 ) | ( n29116 & ~n36711 ) ;
  assign n39542 = n34563 ^ n27740 ^ 1'b0 ;
  assign n39543 = n11563 ^ n1293 ^ x42 ;
  assign n39544 = ( n4212 & ~n24477 ) | ( n4212 & n29271 ) | ( ~n24477 & n29271 ) ;
  assign n39545 = ( n14865 & n32986 ) | ( n14865 & ~n39544 ) | ( n32986 & ~n39544 ) ;
  assign n39546 = n21320 | n23188 ;
  assign n39547 = n519 & ~n39546 ;
  assign n39548 = n39547 ^ n12859 ^ n3372 ;
  assign n39549 = ( n2272 & n37367 ) | ( n2272 & n39548 ) | ( n37367 & n39548 ) ;
  assign n39550 = n21656 ^ n9383 ^ n9174 ;
  assign n39551 = n33739 ^ n19275 ^ n4017 ;
  assign n39552 = n39550 & n39551 ;
  assign n39553 = n35057 ^ n3169 ^ 1'b0 ;
  assign n39554 = ( n4397 & n17798 ) | ( n4397 & ~n23451 ) | ( n17798 & ~n23451 ) ;
  assign n39555 = n39554 ^ n34662 ^ 1'b0 ;
  assign n39556 = ~n29013 & n39555 ;
  assign n39557 = n6433 & n6911 ;
  assign n39558 = ~n39556 & n39557 ;
  assign n39559 = n7556 | n35761 ;
  assign n39560 = n39559 ^ n37124 ^ 1'b0 ;
  assign n39561 = n21657 ^ n12576 ^ n4010 ;
  assign n39562 = n8953 ^ n327 ^ 1'b0 ;
  assign n39563 = ( n16846 & ~n39561 ) | ( n16846 & n39562 ) | ( ~n39561 & n39562 ) ;
  assign n39565 = n12714 ^ n11527 ^ n2290 ;
  assign n39564 = ( ~n6759 & n8469 ) | ( ~n6759 & n28383 ) | ( n8469 & n28383 ) ;
  assign n39566 = n39565 ^ n39564 ^ n35483 ;
  assign n39567 = n12578 ^ n7153 ^ n3340 ;
  assign n39568 = n39567 ^ n4610 ^ n4228 ;
  assign n39575 = ~n11529 & n16603 ;
  assign n39576 = ( n16016 & ~n19064 ) | ( n16016 & n39575 ) | ( ~n19064 & n39575 ) ;
  assign n39569 = ( ~n630 & n4568 ) | ( ~n630 & n21104 ) | ( n4568 & n21104 ) ;
  assign n39571 = n10730 | n14938 ;
  assign n39572 = n39571 ^ n12914 ^ 1'b0 ;
  assign n39570 = n32438 ^ n22117 ^ n2837 ;
  assign n39573 = n39572 ^ n39570 ^ 1'b0 ;
  assign n39574 = ~n39569 & n39573 ;
  assign n39577 = n39576 ^ n39574 ^ n31052 ;
  assign n39578 = n39577 ^ n27444 ^ n17726 ;
  assign n39579 = x208 & n29151 ;
  assign n39580 = n17205 ^ n16671 ^ n12764 ;
  assign n39581 = ( n14914 & n29629 ) | ( n14914 & ~n39580 ) | ( n29629 & ~n39580 ) ;
  assign n39582 = n12980 & n38270 ;
  assign n39583 = ( n11228 & n39581 ) | ( n11228 & ~n39582 ) | ( n39581 & ~n39582 ) ;
  assign n39584 = n25550 ^ n7869 ^ n2151 ;
  assign n39585 = ( n10651 & n13260 ) | ( n10651 & ~n15041 ) | ( n13260 & ~n15041 ) ;
  assign n39586 = n39585 ^ n15089 ^ n14765 ;
  assign n39587 = n39586 ^ n28584 ^ 1'b0 ;
  assign n39588 = ~n9102 & n39587 ;
  assign n39589 = ( ~n15947 & n39584 ) | ( ~n15947 & n39588 ) | ( n39584 & n39588 ) ;
  assign n39590 = n5697 & n6817 ;
  assign n39591 = n39590 ^ n14381 ^ 1'b0 ;
  assign n39592 = n24971 ^ n10023 ^ 1'b0 ;
  assign n39593 = n39591 & ~n39592 ;
  assign n39594 = ( n10012 & n13959 ) | ( n10012 & ~n14621 ) | ( n13959 & ~n14621 ) ;
  assign n39595 = n39594 ^ n25673 ^ n5464 ;
  assign n39596 = n21696 ^ n8262 ^ 1'b0 ;
  assign n39597 = ~n39595 & n39596 ;
  assign n39598 = n27348 ^ n20950 ^ n6169 ;
  assign n39599 = n39598 ^ n12057 ^ 1'b0 ;
  assign n39600 = n22819 | n33844 ;
  assign n39601 = ( n19509 & ~n39599 ) | ( n19509 & n39600 ) | ( ~n39599 & n39600 ) ;
  assign n39603 = n31076 ^ n9869 ^ 1'b0 ;
  assign n39602 = ( ~n10625 & n12231 ) | ( ~n10625 & n27112 ) | ( n12231 & n27112 ) ;
  assign n39604 = n39603 ^ n39602 ^ n13935 ;
  assign n39605 = ~n3486 & n7177 ;
  assign n39606 = n39605 ^ n3280 ^ 1'b0 ;
  assign n39607 = n29140 ^ n20579 ^ n18883 ;
  assign n39608 = ( n1464 & n2350 ) | ( n1464 & ~n7828 ) | ( n2350 & ~n7828 ) ;
  assign n39609 = n12095 & ~n39608 ;
  assign n39610 = n18050 ^ n11965 ^ 1'b0 ;
  assign n39611 = ~n9592 & n39610 ;
  assign n39612 = n7122 | n21471 ;
  assign n39613 = n39612 ^ n35786 ^ 1'b0 ;
  assign n39614 = n32501 ^ n21797 ^ 1'b0 ;
  assign n39615 = n2992 & n39614 ;
  assign n39616 = n36542 ^ n35124 ^ n30509 ;
  assign n39617 = n11895 ^ n11037 ^ 1'b0 ;
  assign n39618 = n39617 ^ n17561 ^ n6974 ;
  assign n39619 = n33543 ^ n13055 ^ n10921 ;
  assign n39620 = n39619 ^ n8944 ^ x227 ;
  assign n39621 = ( n1243 & n3800 ) | ( n1243 & ~n11617 ) | ( n3800 & ~n11617 ) ;
  assign n39622 = ( ~n2949 & n18738 ) | ( ~n2949 & n32937 ) | ( n18738 & n32937 ) ;
  assign n39623 = ( n35099 & ~n39621 ) | ( n35099 & n39622 ) | ( ~n39621 & n39622 ) ;
  assign n39624 = ( n8651 & n13645 ) | ( n8651 & ~n31912 ) | ( n13645 & ~n31912 ) ;
  assign n39625 = n15978 ^ n8891 ^ 1'b0 ;
  assign n39626 = n35511 ^ n28248 ^ n27226 ;
  assign n39627 = n15902 ^ n955 ^ 1'b0 ;
  assign n39628 = n39626 | n39627 ;
  assign n39629 = ( n5529 & ~n6607 ) | ( n5529 & n12999 ) | ( ~n6607 & n12999 ) ;
  assign n39630 = ( n20433 & n25450 ) | ( n20433 & n39629 ) | ( n25450 & n39629 ) ;
  assign n39631 = n1928 & ~n18954 ;
  assign n39633 = ( n4203 & n5136 ) | ( n4203 & ~n7749 ) | ( n5136 & ~n7749 ) ;
  assign n39632 = n20844 | n29326 ;
  assign n39634 = n39633 ^ n39632 ^ 1'b0 ;
  assign n39635 = n39634 ^ n38068 ^ n2737 ;
  assign n39636 = ( n9117 & n15459 ) | ( n9117 & n16745 ) | ( n15459 & n16745 ) ;
  assign n39637 = ( n18134 & ~n29842 ) | ( n18134 & n39636 ) | ( ~n29842 & n39636 ) ;
  assign n39638 = n39637 ^ n37692 ^ n8919 ;
  assign n39639 = n33425 ^ n22228 ^ n11876 ;
  assign n39640 = n39639 ^ n31332 ^ n13954 ;
  assign n39641 = ( n2803 & ~n31290 ) | ( n2803 & n38053 ) | ( ~n31290 & n38053 ) ;
  assign n39642 = n39641 ^ n23660 ^ n23372 ;
  assign n39643 = ( n4072 & ~n11267 ) | ( n4072 & n39642 ) | ( ~n11267 & n39642 ) ;
  assign n39644 = n20748 ^ n11792 ^ 1'b0 ;
  assign n39645 = n39643 | n39644 ;
  assign n39646 = n6189 & n31499 ;
  assign n39648 = n20246 ^ n8122 ^ n7180 ;
  assign n39650 = n7419 ^ n429 ^ x11 ;
  assign n39649 = n22335 ^ n6723 ^ x44 ;
  assign n39651 = n39650 ^ n39649 ^ n7659 ;
  assign n39652 = ( ~n10398 & n39648 ) | ( ~n10398 & n39651 ) | ( n39648 & n39651 ) ;
  assign n39647 = n19903 ^ n18191 ^ n15562 ;
  assign n39653 = n39652 ^ n39647 ^ n27466 ;
  assign n39654 = n23626 ^ n21181 ^ n18268 ;
  assign n39656 = ( n1930 & n2370 ) | ( n1930 & n4922 ) | ( n2370 & n4922 ) ;
  assign n39655 = ( n12629 & n26399 ) | ( n12629 & ~n31202 ) | ( n26399 & ~n31202 ) ;
  assign n39657 = n39656 ^ n39655 ^ n24321 ;
  assign n39658 = ~n18084 & n26055 ;
  assign n39659 = n39658 ^ n29902 ^ 1'b0 ;
  assign n39660 = n39659 ^ n18516 ^ 1'b0 ;
  assign n39661 = n24703 & n39660 ;
  assign n39662 = ( x169 & n20277 ) | ( x169 & n39661 ) | ( n20277 & n39661 ) ;
  assign n39663 = n11775 ^ n6025 ^ n2849 ;
  assign n39664 = n39663 ^ n3816 ^ 1'b0 ;
  assign n39665 = n34940 ^ n29503 ^ n22787 ;
  assign n39666 = ( n3647 & ~n32438 ) | ( n3647 & n39665 ) | ( ~n32438 & n39665 ) ;
  assign n39667 = n21640 ^ n13551 ^ n13083 ;
  assign n39668 = n39667 ^ n30967 ^ n9062 ;
  assign n39669 = ( n2508 & n13583 ) | ( n2508 & ~n27739 ) | ( n13583 & ~n27739 ) ;
  assign n39670 = n39669 ^ n25660 ^ n11920 ;
  assign n39671 = n13587 ^ n11201 ^ n9510 ;
  assign n39672 = ( ~n5293 & n39670 ) | ( ~n5293 & n39671 ) | ( n39670 & n39671 ) ;
  assign n39673 = n9772 ^ n9170 ^ n5106 ;
  assign n39674 = ( n1819 & ~n35040 ) | ( n1819 & n39673 ) | ( ~n35040 & n39673 ) ;
  assign n39675 = n17757 ^ n9349 ^ 1'b0 ;
  assign n39676 = n27793 ^ n9533 ^ 1'b0 ;
  assign n39677 = n12639 ^ n5357 ^ n2232 ;
  assign n39678 = ( n681 & n28706 ) | ( n681 & n39677 ) | ( n28706 & n39677 ) ;
  assign n39679 = n39678 ^ n30839 ^ n19068 ;
  assign n39680 = n21571 ^ n17745 ^ n684 ;
  assign n39681 = n39680 ^ n31936 ^ n11916 ;
  assign n39682 = n16542 ^ n14040 ^ n10654 ;
  assign n39683 = n36990 ^ n18972 ^ n17754 ;
  assign n39684 = n17760 | n21049 ;
  assign n39685 = n3690 & n18107 ;
  assign n39686 = ~n34101 & n39685 ;
  assign n39687 = n8090 | n39686 ;
  assign n39688 = n39687 ^ n36649 ^ 1'b0 ;
  assign n39689 = n7279 ^ n3362 ^ 1'b0 ;
  assign n39690 = n39688 | n39689 ;
  assign n39691 = n22308 & n39690 ;
  assign n39692 = n16467 ^ n3200 ^ 1'b0 ;
  assign n39693 = n27089 ^ n24841 ^ 1'b0 ;
  assign n39694 = ( n4293 & n6959 ) | ( n4293 & ~n39693 ) | ( n6959 & ~n39693 ) ;
  assign n39695 = n18304 & n34184 ;
  assign n39696 = n34149 ^ n33784 ^ 1'b0 ;
  assign n39697 = n39695 & ~n39696 ;
  assign n39698 = n7330 & n31401 ;
  assign n39699 = n39698 ^ n7094 ^ 1'b0 ;
  assign n39700 = n25589 ^ n21535 ^ n4834 ;
  assign n39701 = ( n24307 & ~n26803 ) | ( n24307 & n39700 ) | ( ~n26803 & n39700 ) ;
  assign n39702 = ( ~n9758 & n14083 ) | ( ~n9758 & n28882 ) | ( n14083 & n28882 ) ;
  assign n39703 = ~n12295 & n19965 ;
  assign n39704 = ( n39418 & n39702 ) | ( n39418 & n39703 ) | ( n39702 & n39703 ) ;
  assign n39705 = n19704 & ~n24053 ;
  assign n39706 = ( n5873 & n8557 ) | ( n5873 & ~n39705 ) | ( n8557 & ~n39705 ) ;
  assign n39707 = n39706 ^ n24548 ^ n5107 ;
  assign n39708 = n20731 & n38577 ;
  assign n39709 = ( n2367 & n27732 ) | ( n2367 & n34028 ) | ( n27732 & n34028 ) ;
  assign n39710 = n15734 ^ n11891 ^ n7618 ;
  assign n39711 = n11547 | n39710 ;
  assign n39712 = x227 | n39711 ;
  assign n39713 = n28186 ^ n28102 ^ 1'b0 ;
  assign n39714 = n27205 ^ n21289 ^ 1'b0 ;
  assign n39715 = n39714 ^ n11918 ^ x238 ;
  assign n39716 = n33901 ^ n32086 ^ n21031 ;
  assign n39717 = n39716 ^ n18097 ^ n1352 ;
  assign n39718 = n39717 ^ n10545 ^ n6465 ;
  assign n39719 = n36513 ^ n13471 ^ n6877 ;
  assign n39724 = n19271 ^ n13674 ^ n6864 ;
  assign n39723 = n1476 & n6341 ;
  assign n39725 = n39724 ^ n39723 ^ 1'b0 ;
  assign n39720 = ( n3360 & ~n8549 ) | ( n3360 & n21532 ) | ( ~n8549 & n21532 ) ;
  assign n39721 = n4878 ^ n913 ^ 1'b0 ;
  assign n39722 = n39720 | n39721 ;
  assign n39726 = n39725 ^ n39722 ^ n8798 ;
  assign n39727 = ~n2631 & n4213 ;
  assign n39728 = ~n27343 & n39727 ;
  assign n39729 = n23720 & ~n32534 ;
  assign n39730 = ~n27045 & n39729 ;
  assign n39731 = n19076 ^ n1111 ^ 1'b0 ;
  assign n39732 = n39731 ^ n9098 ^ 1'b0 ;
  assign n39733 = ( n8644 & n36054 ) | ( n8644 & ~n39732 ) | ( n36054 & ~n39732 ) ;
  assign n39734 = n21777 ^ n18806 ^ n11972 ;
  assign n39735 = n32158 ^ n27434 ^ n10665 ;
  assign n39736 = n19444 & ~n19802 ;
  assign n39737 = n39736 ^ n34563 ^ 1'b0 ;
  assign n39738 = n34995 ^ n24292 ^ 1'b0 ;
  assign n39739 = ( n21165 & n39737 ) | ( n21165 & ~n39738 ) | ( n39737 & ~n39738 ) ;
  assign n39740 = ~n2780 & n10246 ;
  assign n39741 = n39740 ^ n10781 ^ 1'b0 ;
  assign n39742 = n18325 ^ n3990 ^ 1'b0 ;
  assign n39743 = n23594 ^ n15913 ^ 1'b0 ;
  assign n39744 = n35938 | n39743 ;
  assign n39745 = n39742 | n39744 ;
  assign n39746 = ( n11553 & ~n37487 ) | ( n11553 & n39745 ) | ( ~n37487 & n39745 ) ;
  assign n39750 = n36736 ^ n13641 ^ 1'b0 ;
  assign n39748 = n1071 & ~n24148 ;
  assign n39749 = n39748 ^ n16011 ^ 1'b0 ;
  assign n39747 = n10062 ^ n8378 ^ n6978 ;
  assign n39751 = n39750 ^ n39749 ^ n39747 ;
  assign n39752 = n5703 | n7691 ;
  assign n39753 = ~n672 & n17388 ;
  assign n39754 = n35090 ^ n11979 ^ n1236 ;
  assign n39755 = n22503 | n39754 ;
  assign n39756 = n3770 | n39755 ;
  assign n39760 = n21989 & ~n29584 ;
  assign n39761 = n39760 ^ n14532 ^ 1'b0 ;
  assign n39757 = ( n907 & n3310 ) | ( n907 & ~n16158 ) | ( n3310 & ~n16158 ) ;
  assign n39758 = ( n906 & n23979 ) | ( n906 & n39757 ) | ( n23979 & n39757 ) ;
  assign n39759 = n39758 ^ n18388 ^ n7169 ;
  assign n39762 = n39761 ^ n39759 ^ n31255 ;
  assign n39763 = n39762 ^ n360 ^ 1'b0 ;
  assign n39764 = n25925 & n39763 ;
  assign n39765 = ( n2156 & n7035 ) | ( n2156 & ~n18651 ) | ( n7035 & ~n18651 ) ;
  assign n39766 = ( n2785 & n7111 ) | ( n2785 & ~n30340 ) | ( n7111 & ~n30340 ) ;
  assign n39767 = n39766 ^ n25128 ^ n19890 ;
  assign n39768 = n6065 & ~n14917 ;
  assign n39769 = ( n14545 & n34331 ) | ( n14545 & n39768 ) | ( n34331 & n39768 ) ;
  assign n39770 = ( n3659 & n12806 ) | ( n3659 & ~n32555 ) | ( n12806 & ~n32555 ) ;
  assign n39771 = ( n9994 & n39769 ) | ( n9994 & ~n39770 ) | ( n39769 & ~n39770 ) ;
  assign n39772 = n19745 & n20207 ;
  assign n39773 = ( ~n5276 & n7326 ) | ( ~n5276 & n16148 ) | ( n7326 & n16148 ) ;
  assign n39774 = n16055 ^ n14834 ^ n8059 ;
  assign n39775 = ( n20784 & n39773 ) | ( n20784 & n39774 ) | ( n39773 & n39774 ) ;
  assign n39776 = ( ~n22785 & n39772 ) | ( ~n22785 & n39775 ) | ( n39772 & n39775 ) ;
  assign n39778 = n6952 | n27167 ;
  assign n39777 = n5560 & n21399 ;
  assign n39779 = n39778 ^ n39777 ^ n11103 ;
  assign n39780 = n4353 & ~n5247 ;
  assign n39781 = ~n9771 & n39780 ;
  assign n39782 = n39781 ^ n16309 ^ n15526 ;
  assign n39783 = ( ~n27522 & n37858 ) | ( ~n27522 & n39782 ) | ( n37858 & n39782 ) ;
  assign n39784 = n25319 ^ n5220 ^ 1'b0 ;
  assign n39785 = n5996 | n34975 ;
  assign n39786 = n39548 ^ n10908 ^ 1'b0 ;
  assign n39787 = n33490 & ~n39786 ;
  assign n39788 = ( ~n5444 & n32889 ) | ( ~n5444 & n33986 ) | ( n32889 & n33986 ) ;
  assign n39789 = n27624 ^ n21994 ^ 1'b0 ;
  assign n39790 = n39788 | n39789 ;
  assign n39792 = n17784 | n34669 ;
  assign n39793 = n1972 & ~n39792 ;
  assign n39791 = n5003 & n33134 ;
  assign n39794 = n39793 ^ n39791 ^ n16862 ;
  assign n39795 = ( n7653 & n9621 ) | ( n7653 & ~n39794 ) | ( n9621 & ~n39794 ) ;
  assign n39796 = n5649 & n19315 ;
  assign n39797 = ~n16874 & n39796 ;
  assign n39798 = n39797 ^ n31237 ^ x143 ;
  assign n39800 = ( n5454 & n9395 ) | ( n5454 & ~n15162 ) | ( n9395 & ~n15162 ) ;
  assign n39799 = n38702 ^ n17406 ^ n10792 ;
  assign n39801 = n39800 ^ n39799 ^ x27 ;
  assign n39802 = ( n8293 & n8644 ) | ( n8293 & ~n10752 ) | ( n8644 & ~n10752 ) ;
  assign n39803 = ( n642 & n8402 ) | ( n642 & ~n39802 ) | ( n8402 & ~n39802 ) ;
  assign n39804 = n39803 ^ n25709 ^ n12307 ;
  assign n39805 = n16258 & n19939 ;
  assign n39806 = ~n39411 & n39805 ;
  assign n39807 = ( n13465 & n30877 ) | ( n13465 & n39806 ) | ( n30877 & n39806 ) ;
  assign n39808 = n2948 ^ n2826 ^ 1'b0 ;
  assign n39809 = ( n10426 & n15232 ) | ( n10426 & ~n39808 ) | ( n15232 & ~n39808 ) ;
  assign n39810 = n27922 ^ n10117 ^ n9321 ;
  assign n39811 = ( n2429 & ~n22410 ) | ( n2429 & n39810 ) | ( ~n22410 & n39810 ) ;
  assign n39812 = n39811 ^ n36587 ^ n21262 ;
  assign n39813 = ~n697 & n3471 ;
  assign n39814 = n39812 & n39813 ;
  assign n39815 = n16982 ^ n12068 ^ 1'b0 ;
  assign n39816 = n5282 | n39815 ;
  assign n39817 = n987 | n39816 ;
  assign n39818 = ~n12658 & n24268 ;
  assign n39819 = n18601 & n39818 ;
  assign n39820 = ( n5290 & ~n7721 ) | ( n5290 & n17196 ) | ( ~n7721 & n17196 ) ;
  assign n39821 = ~n10111 & n39820 ;
  assign n39822 = n33637 ^ n28330 ^ n1016 ;
  assign n39823 = n22931 & ~n23204 ;
  assign n39824 = n39823 ^ n15822 ^ n1726 ;
  assign n39825 = ( n1044 & n32999 ) | ( n1044 & ~n39824 ) | ( n32999 & ~n39824 ) ;
  assign n39826 = n7250 ^ n2389 ^ 1'b0 ;
  assign n39827 = ~n1950 & n39826 ;
  assign n39828 = n39827 ^ n39196 ^ n38358 ;
  assign n39829 = n11745 ^ n11609 ^ n10723 ;
  assign n39830 = ~n6693 & n39829 ;
  assign n39831 = n28907 ^ n20041 ^ 1'b0 ;
  assign n39832 = ( ~n29512 & n39830 ) | ( ~n29512 & n39831 ) | ( n39830 & n39831 ) ;
  assign n39833 = n34327 ^ n31562 ^ 1'b0 ;
  assign n39834 = n38926 ^ n8671 ^ 1'b0 ;
  assign n39835 = n18973 & ~n39834 ;
  assign n39836 = n24771 ^ n16312 ^ n15473 ;
  assign n39837 = n39836 ^ n16385 ^ n12350 ;
  assign n39838 = n39837 ^ n20826 ^ n12402 ;
  assign n39839 = n39838 ^ n3822 ^ 1'b0 ;
  assign n39840 = n2292 | n27887 ;
  assign n39841 = n6719 & n14657 ;
  assign n39842 = ( n5737 & n14410 ) | ( n5737 & n39841 ) | ( n14410 & n39841 ) ;
  assign n39843 = ~n6703 & n39842 ;
  assign n39844 = n15783 ^ n12009 ^ n7086 ;
  assign n39845 = n37725 ^ n12563 ^ n12476 ;
  assign n39846 = n22467 ^ n11061 ^ n4474 ;
  assign n39847 = ( ~n5794 & n10746 ) | ( ~n5794 & n33549 ) | ( n10746 & n33549 ) ;
  assign n39848 = ( n5911 & ~n14769 ) | ( n5911 & n39847 ) | ( ~n14769 & n39847 ) ;
  assign n39849 = n39848 ^ n29049 ^ n15363 ;
  assign n39850 = n15506 & ~n29631 ;
  assign n39851 = ( n1029 & n13854 ) | ( n1029 & ~n16993 ) | ( n13854 & ~n16993 ) ;
  assign n39852 = n17944 ^ n17075 ^ n2094 ;
  assign n39853 = ( n17683 & n39851 ) | ( n17683 & n39852 ) | ( n39851 & n39852 ) ;
  assign n39854 = n39853 ^ n7545 ^ 1'b0 ;
  assign n39855 = ~n1236 & n29159 ;
  assign n39856 = n39855 ^ n13092 ^ n4529 ;
  assign n39857 = n30321 ^ n16611 ^ 1'b0 ;
  assign n39858 = ~n39603 & n39857 ;
  assign n39859 = n39858 ^ n37530 ^ n10859 ;
  assign n39860 = n9589 ^ n1793 ^ n775 ;
  assign n39861 = n39860 ^ n33426 ^ n27991 ;
  assign n39862 = n30925 ^ n19491 ^ 1'b0 ;
  assign n39863 = n13460 & ~n14358 ;
  assign n39864 = ~n16164 & n39863 ;
  assign n39865 = ~n12250 & n18175 ;
  assign n39866 = n39865 ^ n21777 ^ 1'b0 ;
  assign n39869 = n23144 ^ n3724 ^ 1'b0 ;
  assign n39870 = n39869 ^ n29797 ^ 1'b0 ;
  assign n39867 = n22182 ^ n4818 ^ n598 ;
  assign n39868 = ~n6578 & n39867 ;
  assign n39871 = n39870 ^ n39868 ^ n653 ;
  assign n39872 = n2803 | n4671 ;
  assign n39873 = n39872 ^ n22111 ^ 1'b0 ;
  assign n39874 = ( n8694 & n32755 ) | ( n8694 & ~n35520 ) | ( n32755 & ~n35520 ) ;
  assign n39875 = ( ~n7351 & n39873 ) | ( ~n7351 & n39874 ) | ( n39873 & n39874 ) ;
  assign n39876 = n14383 ^ n7113 ^ n4590 ;
  assign n39877 = ( n14678 & n17161 ) | ( n14678 & ~n39876 ) | ( n17161 & ~n39876 ) ;
  assign n39878 = n39464 ^ n31801 ^ n15925 ;
  assign n39883 = n17514 ^ n16456 ^ n10903 ;
  assign n39879 = ~n23807 & n28332 ;
  assign n39880 = n39879 ^ n33490 ^ 1'b0 ;
  assign n39881 = ( n20596 & ~n20697 ) | ( n20596 & n39880 ) | ( ~n20697 & n39880 ) ;
  assign n39882 = ( n30529 & ~n35701 ) | ( n30529 & n39881 ) | ( ~n35701 & n39881 ) ;
  assign n39884 = n39883 ^ n39882 ^ n21451 ;
  assign n39886 = n39658 ^ n39120 ^ n21604 ;
  assign n39885 = n4442 & n7358 ;
  assign n39887 = n39886 ^ n39885 ^ 1'b0 ;
  assign n39888 = ~n26547 & n39887 ;
  assign n39889 = n35636 ^ n13603 ^ 1'b0 ;
  assign n39890 = n23479 | n39889 ;
  assign n39891 = ~n33268 & n39890 ;
  assign n39892 = n2047 & ~n26121 ;
  assign n39893 = ~n34102 & n39892 ;
  assign n39894 = n13772 ^ n1256 ^ 1'b0 ;
  assign n39895 = n39893 | n39894 ;
  assign n39896 = n1709 & n32728 ;
  assign n39897 = n12135 ^ n4764 ^ 1'b0 ;
  assign n39898 = n39897 ^ n10595 ^ n3097 ;
  assign n39899 = n12455 & n39898 ;
  assign n39900 = n39896 & n39899 ;
  assign n39901 = n22052 ^ n3657 ^ 1'b0 ;
  assign n39902 = ( n9888 & n14189 ) | ( n9888 & n21278 ) | ( n14189 & n21278 ) ;
  assign n39903 = ( ~n24670 & n39901 ) | ( ~n24670 & n39902 ) | ( n39901 & n39902 ) ;
  assign n39904 = n22901 ^ n3164 ^ n711 ;
  assign n39905 = ~n31076 & n34165 ;
  assign n39906 = ( ~n15265 & n39904 ) | ( ~n15265 & n39905 ) | ( n39904 & n39905 ) ;
  assign n39907 = n34243 ^ n22012 ^ n4346 ;
  assign n39908 = n14795 ^ n6396 ^ 1'b0 ;
  assign n39909 = n18932 ^ n14874 ^ 1'b0 ;
  assign n39910 = n7039 | n7878 ;
  assign n39911 = n39910 ^ n10415 ^ n705 ;
  assign n39912 = n13903 & n39911 ;
  assign n39913 = n39912 ^ n28050 ^ 1'b0 ;
  assign n39914 = n30830 ^ n21577 ^ n13536 ;
  assign n39915 = n39914 ^ n37776 ^ n9080 ;
  assign n39916 = n39915 ^ n35550 ^ n1688 ;
  assign n39917 = n28102 ^ n1299 ^ 1'b0 ;
  assign n39918 = n39917 ^ n27120 ^ n3606 ;
  assign n39919 = n23325 ^ n8294 ^ 1'b0 ;
  assign n39920 = ( n1399 & n5812 ) | ( n1399 & ~n32539 ) | ( n5812 & ~n32539 ) ;
  assign n39921 = ( n2617 & n25123 ) | ( n2617 & ~n39920 ) | ( n25123 & ~n39920 ) ;
  assign n39922 = n28214 ^ n20478 ^ n3824 ;
  assign n39923 = ( n4247 & ~n39777 ) | ( n4247 & n39922 ) | ( ~n39777 & n39922 ) ;
  assign n39924 = ( ~n6669 & n22619 ) | ( ~n6669 & n39923 ) | ( n22619 & n39923 ) ;
  assign n39925 = n29155 ^ n1124 ^ 1'b0 ;
  assign n39926 = n6546 | n39925 ;
  assign n39927 = n5203 ^ n563 ^ 1'b0 ;
  assign n39928 = ~n39926 & n39927 ;
  assign n39929 = n34449 ^ n25539 ^ n6651 ;
  assign n39938 = n31290 ^ n25853 ^ n24822 ;
  assign n39939 = n10215 & n39938 ;
  assign n39932 = n7774 ^ n6903 ^ 1'b0 ;
  assign n39933 = ~n18141 & n39932 ;
  assign n39934 = n39933 ^ n13013 ^ n5087 ;
  assign n39930 = ( ~n2453 & n11156 ) | ( ~n2453 & n17584 ) | ( n11156 & n17584 ) ;
  assign n39931 = ~n3715 & n39930 ;
  assign n39935 = n39934 ^ n39931 ^ n16513 ;
  assign n39936 = n37325 ^ n17861 ^ 1'b0 ;
  assign n39937 = n39935 & ~n39936 ;
  assign n39940 = n39939 ^ n39937 ^ n11989 ;
  assign n39941 = ( x108 & n19655 ) | ( x108 & n33070 ) | ( n19655 & n33070 ) ;
  assign n39942 = n39940 | n39941 ;
  assign n39943 = ( n7869 & n31396 ) | ( n7869 & ~n34095 ) | ( n31396 & ~n34095 ) ;
  assign n39944 = n17378 & n39943 ;
  assign n39945 = n39944 ^ n6892 ^ n2714 ;
  assign n39946 = n28597 ^ n10473 ^ n3210 ;
  assign n39947 = ( n649 & n6330 ) | ( n649 & n11201 ) | ( n6330 & n11201 ) ;
  assign n39948 = n10095 & ~n22399 ;
  assign n39949 = ( n16254 & ~n39947 ) | ( n16254 & n39948 ) | ( ~n39947 & n39948 ) ;
  assign n39950 = n39949 ^ n2539 ^ 1'b0 ;
  assign n39951 = ( n4392 & n24486 ) | ( n4392 & n28707 ) | ( n24486 & n28707 ) ;
  assign n39952 = n39951 ^ n12882 ^ 1'b0 ;
  assign n39953 = ( n4438 & n7437 ) | ( n4438 & n13117 ) | ( n7437 & n13117 ) ;
  assign n39954 = ( n17060 & n39952 ) | ( n17060 & ~n39953 ) | ( n39952 & ~n39953 ) ;
  assign n39955 = ~n8305 & n18775 ;
  assign n39956 = n13063 & n39955 ;
  assign n39957 = ~n18115 & n18124 ;
  assign n39958 = n39957 ^ n16515 ^ 1'b0 ;
  assign n39959 = n8535 | n9707 ;
  assign n39960 = n9866 & ~n39959 ;
  assign n39961 = n6442 ^ n3208 ^ n358 ;
  assign n39962 = ( n15121 & ~n39960 ) | ( n15121 & n39961 ) | ( ~n39960 & n39961 ) ;
  assign n39963 = ~n19364 & n20913 ;
  assign n39964 = n37952 ^ n31808 ^ n31330 ;
  assign n39965 = n33002 & n39304 ;
  assign n39967 = ( n3371 & n7304 ) | ( n3371 & n19359 ) | ( n7304 & n19359 ) ;
  assign n39968 = ~n13724 & n39967 ;
  assign n39969 = n39968 ^ n4702 ^ 1'b0 ;
  assign n39970 = ( n4694 & ~n10012 ) | ( n4694 & n39969 ) | ( ~n10012 & n39969 ) ;
  assign n39971 = n9596 | n39970 ;
  assign n39972 = n22087 & ~n39971 ;
  assign n39966 = n21003 ^ n13351 ^ n7990 ;
  assign n39973 = n39972 ^ n39966 ^ n9521 ;
  assign n39974 = n4143 | n15696 ;
  assign n39975 = ( n1886 & ~n2568 ) | ( n1886 & n28199 ) | ( ~n2568 & n28199 ) ;
  assign n39976 = ( n6370 & ~n21274 ) | ( n6370 & n39975 ) | ( ~n21274 & n39975 ) ;
  assign n39977 = ( n6775 & n9379 ) | ( n6775 & ~n39976 ) | ( n9379 & ~n39976 ) ;
  assign n39978 = ( n1380 & ~n11205 ) | ( n1380 & n16628 ) | ( ~n11205 & n16628 ) ;
  assign n39979 = n39978 ^ n22178 ^ n9098 ;
  assign n39980 = n39979 ^ n30375 ^ n17945 ;
  assign n39981 = n39980 ^ n33843 ^ 1'b0 ;
  assign n39986 = ~n10028 & n12689 ;
  assign n39987 = n39986 ^ n3649 ^ 1'b0 ;
  assign n39985 = n6488 ^ n5719 ^ 1'b0 ;
  assign n39982 = n8915 ^ n6015 ^ n5804 ;
  assign n39983 = n14649 | n39982 ;
  assign n39984 = n2966 | n39983 ;
  assign n39988 = n39987 ^ n39985 ^ n39984 ;
  assign n39989 = n5503 | n23102 ;
  assign n39990 = n39772 ^ n30520 ^ n310 ;
  assign n39991 = n38570 ^ n26440 ^ 1'b0 ;
  assign n39992 = ( n1722 & ~n3330 ) | ( n1722 & n25025 ) | ( ~n3330 & n25025 ) ;
  assign n39993 = n35237 ^ n16444 ^ n1862 ;
  assign n39994 = ( ~n14492 & n39547 ) | ( ~n14492 & n39993 ) | ( n39547 & n39993 ) ;
  assign n39995 = ( ~n6324 & n13497 ) | ( ~n6324 & n19399 ) | ( n13497 & n19399 ) ;
  assign n39996 = n29088 ^ n20377 ^ n10694 ;
  assign n39997 = ( n7160 & ~n11772 ) | ( n7160 & n27036 ) | ( ~n11772 & n27036 ) ;
  assign n39998 = ( n14383 & n20238 ) | ( n14383 & n39997 ) | ( n20238 & n39997 ) ;
  assign n39999 = n23912 | n39998 ;
  assign n40000 = n39999 ^ n27791 ^ 1'b0 ;
  assign n40001 = n3009 & ~n13666 ;
  assign n40002 = n40001 ^ n12810 ^ 1'b0 ;
  assign n40003 = n1967 & ~n40002 ;
  assign n40004 = ~n9830 & n40003 ;
  assign n40005 = n4456 & ~n11172 ;
  assign n40006 = n39799 & n40005 ;
  assign n40007 = ( x160 & n40004 ) | ( x160 & n40006 ) | ( n40004 & n40006 ) ;
  assign n40008 = n35269 ^ n22762 ^ n14237 ;
  assign n40009 = n12891 & ~n40008 ;
  assign n40010 = n40007 & n40009 ;
  assign n40011 = ( n3126 & n8556 ) | ( n3126 & ~n26307 ) | ( n8556 & ~n26307 ) ;
  assign n40012 = n38332 ^ n14878 ^ n9704 ;
  assign n40013 = n3636 & ~n11985 ;
  assign n40014 = ~n2527 & n21884 ;
  assign n40015 = n22209 ^ n882 ^ x20 ;
  assign n40016 = n40015 ^ n22343 ^ 1'b0 ;
  assign n40017 = ~n8160 & n9930 ;
  assign n40018 = ~n9274 & n40017 ;
  assign n40019 = n822 | n40018 ;
  assign n40020 = n23517 | n40019 ;
  assign n40021 = ( x99 & ~n10347 ) | ( x99 & n10928 ) | ( ~n10347 & n10928 ) ;
  assign n40022 = ( ~n353 & n935 ) | ( ~n353 & n40021 ) | ( n935 & n40021 ) ;
  assign n40023 = n40022 ^ n24723 ^ n9181 ;
  assign n40024 = n40020 & ~n40023 ;
  assign n40025 = n23379 ^ n6106 ^ 1'b0 ;
  assign n40026 = n34663 ^ n21878 ^ 1'b0 ;
  assign n40027 = n40025 & n40026 ;
  assign n40028 = n33318 | n38298 ;
  assign n40029 = n40028 ^ n2794 ^ 1'b0 ;
  assign n40030 = n31359 ^ n30615 ^ n8845 ;
  assign n40031 = n33788 ^ n8302 ^ n3960 ;
  assign n40032 = n30665 ^ n7318 ^ 1'b0 ;
  assign n40033 = n10169 ^ n5389 ^ n4911 ;
  assign n40034 = ( ~n8738 & n19329 ) | ( ~n8738 & n40033 ) | ( n19329 & n40033 ) ;
  assign n40035 = n6985 ^ n3340 ^ n1130 ;
  assign n40036 = ( n1505 & n5871 ) | ( n1505 & n13354 ) | ( n5871 & n13354 ) ;
  assign n40037 = n23148 ^ n8691 ^ 1'b0 ;
  assign n40038 = n40036 & ~n40037 ;
  assign n40039 = n40035 & n40038 ;
  assign n40040 = n39509 ^ n3664 ^ 1'b0 ;
  assign n40041 = n26071 ^ n6345 ^ 1'b0 ;
  assign n40042 = n15459 & ~n40041 ;
  assign n40043 = ( n26104 & n26734 ) | ( n26104 & n35624 ) | ( n26734 & n35624 ) ;
  assign n40045 = ~n9602 & n16132 ;
  assign n40046 = n40045 ^ n5964 ^ 1'b0 ;
  assign n40044 = n23844 & n25131 ;
  assign n40047 = n40046 ^ n40044 ^ 1'b0 ;
  assign n40048 = n40047 ^ n24756 ^ 1'b0 ;
  assign n40049 = n14060 ^ n7673 ^ 1'b0 ;
  assign n40050 = n13210 | n40049 ;
  assign n40051 = n40050 ^ n16150 ^ n7779 ;
  assign n40052 = n40051 ^ n12156 ^ n10106 ;
  assign n40053 = ( n25824 & n27678 ) | ( n25824 & n30722 ) | ( n27678 & n30722 ) ;
  assign n40054 = n449 | n4258 ;
  assign n40059 = n8063 ^ n1702 ^ x230 ;
  assign n40055 = n4957 | n9339 ;
  assign n40056 = n40055 ^ n3900 ^ 1'b0 ;
  assign n40057 = n3944 | n15175 ;
  assign n40058 = ( n14388 & n40056 ) | ( n14388 & n40057 ) | ( n40056 & n40057 ) ;
  assign n40060 = n40059 ^ n40058 ^ n36784 ;
  assign n40061 = ( n1269 & ~n28269 ) | ( n1269 & n33592 ) | ( ~n28269 & n33592 ) ;
  assign n40062 = n40061 ^ n27717 ^ 1'b0 ;
  assign n40063 = n35901 & n40062 ;
  assign n40064 = n22017 ^ n14127 ^ n10330 ;
  assign n40065 = ( ~n21236 & n32058 ) | ( ~n21236 & n40064 ) | ( n32058 & n40064 ) ;
  assign n40066 = ( n7573 & ~n22163 ) | ( n7573 & n25639 ) | ( ~n22163 & n25639 ) ;
  assign n40067 = n40066 ^ n1279 ^ 1'b0 ;
  assign n40068 = n40065 | n40067 ;
  assign n40069 = ( n7560 & ~n23182 ) | ( n7560 & n24145 ) | ( ~n23182 & n24145 ) ;
  assign n40070 = n15841 ^ n11791 ^ 1'b0 ;
  assign n40071 = n14399 & n40070 ;
  assign n40072 = ( n12626 & n37612 ) | ( n12626 & n40071 ) | ( n37612 & n40071 ) ;
  assign n40075 = n5955 ^ n2933 ^ n959 ;
  assign n40076 = n15067 & n40075 ;
  assign n40073 = n39979 ^ n33845 ^ 1'b0 ;
  assign n40074 = n19861 & ~n40073 ;
  assign n40077 = n40076 ^ n40074 ^ n35694 ;
  assign n40078 = n16568 ^ n11791 ^ 1'b0 ;
  assign n40079 = n15506 & n40078 ;
  assign n40084 = n7078 ^ n4176 ^ n2466 ;
  assign n40085 = n40084 ^ n8250 ^ n1460 ;
  assign n40080 = n5929 & ~n9668 ;
  assign n40081 = ~n13016 & n40080 ;
  assign n40082 = ( n18860 & n24584 ) | ( n18860 & ~n40081 ) | ( n24584 & ~n40081 ) ;
  assign n40083 = n13137 & ~n40082 ;
  assign n40086 = n40085 ^ n40083 ^ 1'b0 ;
  assign n40087 = n40079 & n40086 ;
  assign n40088 = ( ~n327 & n8083 ) | ( ~n327 & n28566 ) | ( n8083 & n28566 ) ;
  assign n40089 = ( n11669 & n23763 ) | ( n11669 & n40088 ) | ( n23763 & n40088 ) ;
  assign n40090 = n1956 & n24010 ;
  assign n40091 = n40090 ^ n23145 ^ 1'b0 ;
  assign n40092 = n9064 & n40091 ;
  assign n40093 = n31406 ^ n22781 ^ n8194 ;
  assign n40094 = n22971 ^ n14771 ^ 1'b0 ;
  assign n40095 = ( ~n10980 & n12131 ) | ( ~n10980 & n22164 ) | ( n12131 & n22164 ) ;
  assign n40096 = ( n606 & n1650 ) | ( n606 & ~n16726 ) | ( n1650 & ~n16726 ) ;
  assign n40097 = ( n18242 & ~n40095 ) | ( n18242 & n40096 ) | ( ~n40095 & n40096 ) ;
  assign n40098 = n11893 ^ n4141 ^ 1'b0 ;
  assign n40099 = n13315 ^ n2189 ^ 1'b0 ;
  assign n40101 = n1095 | n1590 ;
  assign n40102 = n24880 | n40101 ;
  assign n40100 = n7142 | n33263 ;
  assign n40103 = n40102 ^ n40100 ^ 1'b0 ;
  assign n40104 = ( n497 & n12801 ) | ( n497 & n19398 ) | ( n12801 & n19398 ) ;
  assign n40105 = n30605 | n40104 ;
  assign n40106 = n40105 ^ n4574 ^ 1'b0 ;
  assign n40107 = n22677 | n24910 ;
  assign n40108 = n40107 ^ n23128 ^ 1'b0 ;
  assign n40109 = n19052 & n40108 ;
  assign n40110 = n35753 ^ n23507 ^ 1'b0 ;
  assign n40111 = n40109 & ~n40110 ;
  assign n40112 = n18910 ^ n17446 ^ n2867 ;
  assign n40113 = ( ~n11625 & n23627 ) | ( ~n11625 & n26944 ) | ( n23627 & n26944 ) ;
  assign n40114 = n3708 | n40113 ;
  assign n40115 = n40114 ^ n30290 ^ n19284 ;
  assign n40117 = n6101 & n14122 ;
  assign n40118 = n40117 ^ n35649 ^ 1'b0 ;
  assign n40116 = n3326 & ~n37351 ;
  assign n40119 = n40118 ^ n40116 ^ 1'b0 ;
  assign n40120 = ( ~n4426 & n26951 ) | ( ~n4426 & n40119 ) | ( n26951 & n40119 ) ;
  assign n40121 = n37788 ^ n19159 ^ n5533 ;
  assign n40122 = ( n8784 & n23479 ) | ( n8784 & n24626 ) | ( n23479 & n24626 ) ;
  assign n40123 = n19136 ^ n9929 ^ 1'b0 ;
  assign n40124 = ( ~n17944 & n40122 ) | ( ~n17944 & n40123 ) | ( n40122 & n40123 ) ;
  assign n40125 = n4004 & ~n32388 ;
  assign n40126 = n40125 ^ n33002 ^ 1'b0 ;
  assign n40127 = ( n5717 & n7004 ) | ( n5717 & ~n13149 ) | ( n7004 & ~n13149 ) ;
  assign n40128 = n40127 ^ n10920 ^ 1'b0 ;
  assign n40129 = ~n1712 & n40128 ;
  assign n40130 = ~n12084 & n13683 ;
  assign n40131 = n11895 ^ n3240 ^ n2308 ;
  assign n40132 = ~n24376 & n40131 ;
  assign n40133 = ~n16885 & n32173 ;
  assign n40134 = n39562 ^ n20016 ^ 1'b0 ;
  assign n40135 = ( n24015 & ~n40133 ) | ( n24015 & n40134 ) | ( ~n40133 & n40134 ) ;
  assign n40140 = n9772 | n31223 ;
  assign n40141 = n40140 ^ n9872 ^ 1'b0 ;
  assign n40137 = n19707 ^ n15959 ^ 1'b0 ;
  assign n40138 = ~n16480 & n40137 ;
  assign n40139 = x74 & ~n40138 ;
  assign n40136 = n21360 ^ n15298 ^ n1125 ;
  assign n40142 = n40141 ^ n40139 ^ n40136 ;
  assign n40143 = n31955 ^ n24943 ^ 1'b0 ;
  assign n40144 = n8135 & ~n40143 ;
  assign n40145 = n40144 ^ n22599 ^ 1'b0 ;
  assign n40146 = ( n2685 & ~n2795 ) | ( n2685 & n11530 ) | ( ~n2795 & n11530 ) ;
  assign n40147 = n36583 ^ n35593 ^ n22887 ;
  assign n40148 = n29155 ^ n16695 ^ n3596 ;
  assign n40149 = n40148 ^ n13793 ^ 1'b0 ;
  assign n40150 = ( n40146 & ~n40147 ) | ( n40146 & n40149 ) | ( ~n40147 & n40149 ) ;
  assign n40152 = ( n5143 & n18813 ) | ( n5143 & n37259 ) | ( n18813 & n37259 ) ;
  assign n40151 = n25497 | n33686 ;
  assign n40153 = n40152 ^ n40151 ^ 1'b0 ;
  assign n40154 = n16083 ^ n4060 ^ 1'b0 ;
  assign n40155 = n13134 | n40154 ;
  assign n40156 = ( x29 & n17611 ) | ( x29 & ~n37176 ) | ( n17611 & ~n37176 ) ;
  assign n40157 = n23854 ^ n6465 ^ n5861 ;
  assign n40158 = ( n7529 & ~n11311 ) | ( n7529 & n40157 ) | ( ~n11311 & n40157 ) ;
  assign n40159 = n24370 ^ n14391 ^ 1'b0 ;
  assign n40160 = n27612 & n40159 ;
  assign n40161 = ( n28512 & n40158 ) | ( n28512 & ~n40160 ) | ( n40158 & ~n40160 ) ;
  assign n40162 = n19789 ^ n5201 ^ 1'b0 ;
  assign n40163 = n13771 ^ n13477 ^ 1'b0 ;
  assign n40164 = n40163 ^ n36316 ^ n9398 ;
  assign n40165 = n22710 ^ n15315 ^ 1'b0 ;
  assign n40166 = ( n16925 & ~n16959 ) | ( n16925 & n34849 ) | ( ~n16959 & n34849 ) ;
  assign n40167 = ( ~n16880 & n40165 ) | ( ~n16880 & n40166 ) | ( n40165 & n40166 ) ;
  assign n40168 = n2951 & n40167 ;
  assign n40169 = n40168 ^ n17822 ^ 1'b0 ;
  assign n40172 = n15979 ^ n9050 ^ n7577 ;
  assign n40170 = n39650 ^ n6130 ^ n438 ;
  assign n40171 = n7091 & ~n40170 ;
  assign n40173 = n40172 ^ n40171 ^ 1'b0 ;
  assign n40174 = ( n12331 & ~n15438 ) | ( n12331 & n16773 ) | ( ~n15438 & n16773 ) ;
  assign n40175 = ( ~n4128 & n11039 ) | ( ~n4128 & n16411 ) | ( n11039 & n16411 ) ;
  assign n40176 = ( ~n6388 & n6463 ) | ( ~n6388 & n40175 ) | ( n6463 & n40175 ) ;
  assign n40177 = n40176 ^ n32477 ^ n29861 ;
  assign n40178 = n9884 ^ n4841 ^ n854 ;
  assign n40179 = n40178 ^ n29204 ^ n27876 ;
  assign n40180 = n40179 ^ n8578 ^ 1'b0 ;
  assign n40181 = ( n6193 & n19588 ) | ( n6193 & n40180 ) | ( n19588 & n40180 ) ;
  assign n40182 = n23914 ^ n11847 ^ 1'b0 ;
  assign n40183 = n16683 & n40182 ;
  assign n40184 = n40183 ^ n37254 ^ n11245 ;
  assign n40186 = n13689 ^ n1871 ^ 1'b0 ;
  assign n40185 = ~n5948 & n13214 ;
  assign n40187 = n40186 ^ n40185 ^ n24139 ;
  assign n40188 = ( n1482 & ~n10095 ) | ( n1482 & n40187 ) | ( ~n10095 & n40187 ) ;
  assign n40189 = n36109 ^ n10259 ^ n7582 ;
  assign n40190 = n15634 & n40189 ;
  assign n40191 = n13773 ^ n13078 ^ 1'b0 ;
  assign n40192 = n25400 ^ n25305 ^ n17175 ;
  assign n40195 = n27443 ^ n8887 ^ n5617 ;
  assign n40193 = n33539 | n36079 ;
  assign n40194 = n40193 ^ n11626 ^ 1'b0 ;
  assign n40196 = n40195 ^ n40194 ^ n21691 ;
  assign n40197 = ( n10840 & n32746 ) | ( n10840 & n33438 ) | ( n32746 & n33438 ) ;
  assign n40198 = n38090 ^ n1461 ^ 1'b0 ;
  assign n40199 = n5948 & n40198 ;
  assign n40200 = n38552 & n40199 ;
  assign n40201 = n40197 & n40200 ;
  assign n40202 = ( ~n24665 & n30852 ) | ( ~n24665 & n35148 ) | ( n30852 & n35148 ) ;
  assign n40203 = n2657 & ~n40202 ;
  assign n40204 = n8794 | n12332 ;
  assign n40205 = n40204 ^ n21081 ^ 1'b0 ;
  assign n40206 = n40205 ^ n12320 ^ 1'b0 ;
  assign n40207 = n15034 | n15296 ;
  assign n40208 = n25075 ^ n18252 ^ n12853 ;
  assign n40209 = n6444 ^ n5247 ^ n1061 ;
  assign n40210 = ~n23460 & n37406 ;
  assign n40211 = n40209 & n40210 ;
  assign n40212 = n29711 & ~n31710 ;
  assign n40213 = ( ~n24092 & n36542 ) | ( ~n24092 & n38984 ) | ( n36542 & n38984 ) ;
  assign n40214 = ( n986 & n1062 ) | ( n986 & n16517 ) | ( n1062 & n16517 ) ;
  assign n40215 = n40214 ^ n13513 ^ n1708 ;
  assign n40216 = ( ~n18597 & n21456 ) | ( ~n18597 & n40215 ) | ( n21456 & n40215 ) ;
  assign n40217 = n20894 ^ n14960 ^ n4357 ;
  assign n40218 = n40217 ^ n6628 ^ 1'b0 ;
  assign n40219 = ~n13130 & n25376 ;
  assign n40220 = ( n5808 & n20974 ) | ( n5808 & ~n32513 ) | ( n20974 & ~n32513 ) ;
  assign n40221 = n16175 | n18103 ;
  assign n40222 = n11238 | n40221 ;
  assign n40223 = n20379 ^ n6592 ^ 1'b0 ;
  assign n40225 = n32971 ^ n16809 ^ 1'b0 ;
  assign n40226 = n5341 & n40225 ;
  assign n40224 = n1402 | n16175 ;
  assign n40227 = n40226 ^ n40224 ^ 1'b0 ;
  assign n40228 = ( ~n3271 & n23871 ) | ( ~n3271 & n28438 ) | ( n23871 & n28438 ) ;
  assign n40229 = n40228 ^ n19994 ^ n12321 ;
  assign n40230 = n40229 ^ n14242 ^ 1'b0 ;
  assign n40231 = ( n1476 & ~n5978 ) | ( n1476 & n20343 ) | ( ~n5978 & n20343 ) ;
  assign n40232 = n27176 & ~n37511 ;
  assign n40233 = ( n31646 & n40231 ) | ( n31646 & ~n40232 ) | ( n40231 & ~n40232 ) ;
  assign n40234 = ( n17627 & n22376 ) | ( n17627 & ~n40233 ) | ( n22376 & ~n40233 ) ;
  assign n40236 = n7265 ^ n5684 ^ n4457 ;
  assign n40237 = ( n6609 & n13922 ) | ( n6609 & n40236 ) | ( n13922 & n40236 ) ;
  assign n40238 = n19626 ^ n6987 ^ n4330 ;
  assign n40239 = ( n9288 & n40237 ) | ( n9288 & ~n40238 ) | ( n40237 & ~n40238 ) ;
  assign n40235 = ( n2527 & ~n18946 ) | ( n2527 & n32937 ) | ( ~n18946 & n32937 ) ;
  assign n40240 = n40239 ^ n40235 ^ n31620 ;
  assign n40241 = n6992 ^ n4901 ^ 1'b0 ;
  assign n40242 = n30588 ^ n29550 ^ 1'b0 ;
  assign n40243 = ~n12206 & n40242 ;
  assign n40244 = n40243 ^ x16 ^ 1'b0 ;
  assign n40245 = n11989 | n23387 ;
  assign n40246 = ( n40241 & n40244 ) | ( n40241 & ~n40245 ) | ( n40244 & ~n40245 ) ;
  assign n40247 = n22235 ^ n11808 ^ 1'b0 ;
  assign n40248 = n21232 & n40247 ;
  assign n40249 = n3562 ^ n287 ^ 1'b0 ;
  assign n40250 = ( n12519 & n27271 ) | ( n12519 & ~n40249 ) | ( n27271 & ~n40249 ) ;
  assign n40251 = n9956 ^ n6268 ^ n5617 ;
  assign n40252 = ( ~n11893 & n21348 ) | ( ~n11893 & n40251 ) | ( n21348 & n40251 ) ;
  assign n40253 = n40252 ^ n402 ^ x5 ;
  assign n40254 = n6592 & n7127 ;
  assign n40255 = n21888 ^ n2659 ^ n257 ;
  assign n40256 = n2150 & ~n28295 ;
  assign n40257 = n12699 ^ n3505 ^ 1'b0 ;
  assign n40258 = ( ~n20446 & n24525 ) | ( ~n20446 & n25738 ) | ( n24525 & n25738 ) ;
  assign n40259 = n12421 & ~n40258 ;
  assign n40260 = n10442 & ~n40259 ;
  assign n40261 = n40257 & n40260 ;
  assign n40262 = n40256 | n40261 ;
  assign n40263 = n23669 & ~n40262 ;
  assign n40264 = ( n40254 & n40255 ) | ( n40254 & n40263 ) | ( n40255 & n40263 ) ;
  assign n40265 = n38407 ^ n28882 ^ 1'b0 ;
  assign n40266 = n2086 & n40265 ;
  assign n40267 = n40266 ^ n12666 ^ n496 ;
  assign n40268 = n21859 & n33572 ;
  assign n40269 = n40268 ^ n6214 ^ 1'b0 ;
  assign n40270 = n9074 | n18581 ;
  assign n40271 = n40270 ^ n4116 ^ 1'b0 ;
  assign n40272 = n40269 & ~n40271 ;
  assign n40273 = n5561 & ~n39788 ;
  assign n40274 = n40273 ^ n34050 ^ 1'b0 ;
  assign n40275 = ( n3328 & n32540 ) | ( n3328 & n40274 ) | ( n32540 & n40274 ) ;
  assign n40276 = n15836 ^ n12001 ^ n3806 ;
  assign n40277 = ( n4108 & n17109 ) | ( n4108 & n40276 ) | ( n17109 & n40276 ) ;
  assign n40278 = n6476 & n40277 ;
  assign n40279 = n40278 ^ n9654 ^ 1'b0 ;
  assign n40280 = ( n9233 & n40079 ) | ( n9233 & n40279 ) | ( n40079 & n40279 ) ;
  assign n40281 = n6458 & n24374 ;
  assign n40282 = n40281 ^ n12470 ^ 1'b0 ;
  assign n40283 = n40282 ^ n9577 ^ 1'b0 ;
  assign n40284 = ( n21271 & ~n24840 ) | ( n21271 & n32937 ) | ( ~n24840 & n32937 ) ;
  assign n40285 = n40284 ^ n33754 ^ n21552 ;
  assign n40286 = ~n7562 & n18295 ;
  assign n40287 = n22245 ^ n9758 ^ 1'b0 ;
  assign n40289 = n17909 & ~n26301 ;
  assign n40288 = n11707 & n27144 ;
  assign n40290 = n40289 ^ n40288 ^ 1'b0 ;
  assign n40291 = n15415 | n26793 ;
  assign n40292 = n27368 & n40291 ;
  assign n40293 = ~n16685 & n40292 ;
  assign n40294 = ~n6524 & n7168 ;
  assign n40295 = n14207 ^ n2699 ^ 1'b0 ;
  assign n40296 = n798 & n40295 ;
  assign n40297 = n8840 & n40296 ;
  assign n40298 = ~n40294 & n40297 ;
  assign n40299 = ~n5668 & n40298 ;
  assign n40300 = n22524 | n25104 ;
  assign n40301 = n40300 ^ n6558 ^ 1'b0 ;
  assign n40302 = n25873 ^ n18598 ^ n6717 ;
  assign n40303 = n4155 | n4341 ;
  assign n40304 = n40303 ^ x76 ^ 1'b0 ;
  assign n40305 = n40304 ^ n33889 ^ 1'b0 ;
  assign n40306 = n9507 & ~n32503 ;
  assign n40307 = n10660 & n40306 ;
  assign n40308 = n39827 ^ n9274 ^ n8137 ;
  assign n40309 = ( n37144 & n40307 ) | ( n37144 & ~n40308 ) | ( n40307 & ~n40308 ) ;
  assign n40310 = ( n28304 & n40305 ) | ( n28304 & n40309 ) | ( n40305 & n40309 ) ;
  assign n40311 = n40310 ^ n19813 ^ n3144 ;
  assign n40312 = ( n21781 & n29116 ) | ( n21781 & n40311 ) | ( n29116 & n40311 ) ;
  assign n40313 = ( n931 & n21290 ) | ( n931 & ~n30116 ) | ( n21290 & ~n30116 ) ;
  assign n40322 = ( n16339 & ~n27626 ) | ( n16339 & n32361 ) | ( ~n27626 & n32361 ) ;
  assign n40323 = ( ~n4420 & n10925 ) | ( ~n4420 & n40322 ) | ( n10925 & n40322 ) ;
  assign n40314 = n22858 ^ n17381 ^ n6496 ;
  assign n40315 = ( n1898 & n12836 ) | ( n1898 & n15660 ) | ( n12836 & n15660 ) ;
  assign n40316 = n4448 | n40315 ;
  assign n40317 = n40316 ^ n30340 ^ n8195 ;
  assign n40318 = ( n10454 & n23948 ) | ( n10454 & ~n40317 ) | ( n23948 & ~n40317 ) ;
  assign n40319 = ~n10761 & n40318 ;
  assign n40320 = ~n1058 & n40319 ;
  assign n40321 = n40314 & ~n40320 ;
  assign n40324 = n40323 ^ n40321 ^ n22310 ;
  assign n40325 = ~n412 & n40324 ;
  assign n40326 = n22726 ^ x180 ^ 1'b0 ;
  assign n40327 = ( ~n1893 & n12000 ) | ( ~n1893 & n14105 ) | ( n12000 & n14105 ) ;
  assign n40328 = n40327 ^ n39388 ^ 1'b0 ;
  assign n40329 = n6947 & ~n40328 ;
  assign n40330 = n20333 | n24317 ;
  assign n40331 = n3389 | n40330 ;
  assign n40332 = n381 & n40331 ;
  assign n40333 = ~n15950 & n40332 ;
  assign n40334 = ~n1780 & n19500 ;
  assign n40335 = n33563 ^ n16806 ^ n6333 ;
  assign n40340 = n12270 & ~n14255 ;
  assign n40338 = n9905 ^ n8252 ^ n781 ;
  assign n40339 = n40338 ^ n23166 ^ n18258 ;
  assign n40336 = ( n959 & n1189 ) | ( n959 & n2081 ) | ( n1189 & n2081 ) ;
  assign n40337 = n6789 | n40336 ;
  assign n40341 = n40340 ^ n40339 ^ n40337 ;
  assign n40342 = ( n3609 & n13226 ) | ( n3609 & ~n40341 ) | ( n13226 & ~n40341 ) ;
  assign n40343 = n26254 ^ n4549 ^ 1'b0 ;
  assign n40344 = ( ~n13765 & n27839 ) | ( ~n13765 & n40343 ) | ( n27839 & n40343 ) ;
  assign n40345 = n733 & ~n8873 ;
  assign n40346 = n30817 ^ n29119 ^ 1'b0 ;
  assign n40347 = n12210 & ~n40346 ;
  assign n40348 = ( n8318 & n40345 ) | ( n8318 & ~n40347 ) | ( n40345 & ~n40347 ) ;
  assign n40349 = ( n26769 & n32872 ) | ( n26769 & ~n40348 ) | ( n32872 & ~n40348 ) ;
  assign n40350 = n2232 & n7085 ;
  assign n40351 = n40350 ^ n11251 ^ n5225 ;
  assign n40352 = n21134 ^ n14948 ^ n7101 ;
  assign n40353 = ( n3641 & ~n5789 ) | ( n3641 & n40352 ) | ( ~n5789 & n40352 ) ;
  assign n40354 = ( ~n23186 & n40351 ) | ( ~n23186 & n40353 ) | ( n40351 & n40353 ) ;
  assign n40355 = n23363 ^ n17838 ^ n9618 ;
  assign n40356 = n23803 & ~n40355 ;
  assign n40357 = n14227 ^ n12240 ^ n7830 ;
  assign n40358 = n12302 & n40357 ;
  assign n40359 = n30971 ^ n5844 ^ n2536 ;
  assign n40360 = n5328 | n7362 ;
  assign n40361 = n40360 ^ n23674 ^ 1'b0 ;
  assign n40362 = ( ~n5247 & n40359 ) | ( ~n5247 & n40361 ) | ( n40359 & n40361 ) ;
  assign n40363 = n17345 | n34476 ;
  assign n40364 = ( n16893 & n36520 ) | ( n16893 & n40363 ) | ( n36520 & n40363 ) ;
  assign n40365 = ( n9586 & ~n16718 ) | ( n9586 & n31971 ) | ( ~n16718 & n31971 ) ;
  assign n40366 = ( n5928 & ~n19746 ) | ( n5928 & n32698 ) | ( ~n19746 & n32698 ) ;
  assign n40367 = n40366 ^ n28343 ^ n2953 ;
  assign n40368 = n40367 ^ n38446 ^ n35501 ;
  assign n40373 = n20222 ^ n7794 ^ n1014 ;
  assign n40369 = n18246 ^ n14629 ^ 1'b0 ;
  assign n40370 = n16212 & n40369 ;
  assign n40371 = n21945 ^ n7329 ^ 1'b0 ;
  assign n40372 = ( n10394 & n40370 ) | ( n10394 & ~n40371 ) | ( n40370 & ~n40371 ) ;
  assign n40374 = n40373 ^ n40372 ^ n39350 ;
  assign n40375 = n37096 ^ n5925 ^ 1'b0 ;
  assign n40376 = n2668 | n40375 ;
  assign n40377 = ( n5843 & n40374 ) | ( n5843 & ~n40376 ) | ( n40374 & ~n40376 ) ;
  assign n40379 = ( ~n602 & n3685 ) | ( ~n602 & n32304 ) | ( n3685 & n32304 ) ;
  assign n40378 = n35845 ^ n7062 ^ 1'b0 ;
  assign n40380 = n40379 ^ n40378 ^ x6 ;
  assign n40383 = n12239 ^ n3058 ^ x170 ;
  assign n40381 = n3267 & n6314 ;
  assign n40382 = n40381 ^ n11779 ^ n4906 ;
  assign n40384 = n40383 ^ n40382 ^ n9842 ;
  assign n40385 = n40384 ^ n22935 ^ n4562 ;
  assign n40386 = n40385 ^ n16885 ^ 1'b0 ;
  assign n40387 = n15903 & n40386 ;
  assign n40388 = n8061 | n17450 ;
  assign n40389 = n482 | n40388 ;
  assign n40390 = n40389 ^ n3054 ^ 1'b0 ;
  assign n40391 = n17509 ^ n6398 ^ n1242 ;
  assign n40392 = n13120 & ~n32982 ;
  assign n40393 = ~n40391 & n40392 ;
  assign n40394 = ( ~n20503 & n33337 ) | ( ~n20503 & n35701 ) | ( n33337 & n35701 ) ;
  assign n40395 = n10047 ^ n5411 ^ n4431 ;
  assign n40396 = ( n5147 & n10209 ) | ( n5147 & ~n28947 ) | ( n10209 & ~n28947 ) ;
  assign n40397 = n2909 ^ n1039 ^ 1'b0 ;
  assign n40398 = ( n938 & n3061 ) | ( n938 & ~n40397 ) | ( n3061 & ~n40397 ) ;
  assign n40399 = ( x11 & ~n8360 ) | ( x11 & n40398 ) | ( ~n8360 & n40398 ) ;
  assign n40400 = n31045 ^ n10523 ^ n1146 ;
  assign n40401 = n40400 ^ n32093 ^ 1'b0 ;
  assign n40402 = n7467 | n38652 ;
  assign n40403 = n22830 | n40402 ;
  assign n40404 = ( n5502 & n25827 ) | ( n5502 & ~n40403 ) | ( n25827 & ~n40403 ) ;
  assign n40409 = ( n2245 & ~n6088 ) | ( n2245 & n6105 ) | ( ~n6088 & n6105 ) ;
  assign n40405 = n26115 ^ n6343 ^ 1'b0 ;
  assign n40406 = n4371 & ~n40405 ;
  assign n40407 = ( x65 & n21091 ) | ( x65 & ~n28602 ) | ( n21091 & ~n28602 ) ;
  assign n40408 = n40406 & ~n40407 ;
  assign n40410 = n40409 ^ n40408 ^ 1'b0 ;
  assign n40411 = ( n3588 & n10217 ) | ( n3588 & n16087 ) | ( n10217 & n16087 ) ;
  assign n40412 = n40411 ^ n5014 ^ 1'b0 ;
  assign n40413 = n15531 & n40412 ;
  assign n40414 = n652 & n11986 ;
  assign n40415 = n19203 & n40414 ;
  assign n40416 = n40415 ^ n7120 ^ 1'b0 ;
  assign n40417 = n40413 & n40416 ;
  assign n40418 = ( ~n10072 & n16802 ) | ( ~n10072 & n37326 ) | ( n16802 & n37326 ) ;
  assign n40419 = n13336 ^ n9330 ^ n4354 ;
  assign n40420 = ( n22351 & ~n25299 ) | ( n22351 & n35512 ) | ( ~n25299 & n35512 ) ;
  assign n40421 = n7070 | n38739 ;
  assign n40422 = n22448 ^ n12988 ^ n3998 ;
  assign n40423 = ( n8941 & n40421 ) | ( n8941 & n40422 ) | ( n40421 & n40422 ) ;
  assign n40424 = ~n19126 & n32558 ;
  assign n40425 = n40424 ^ n27931 ^ 1'b0 ;
  assign n40426 = n6255 & n25398 ;
  assign n40427 = n14890 & ~n33467 ;
  assign n40428 = n40426 & n40427 ;
  assign n40429 = ( ~n20525 & n35176 ) | ( ~n20525 & n35277 ) | ( n35176 & n35277 ) ;
  assign n40430 = n36512 ^ n9829 ^ n3417 ;
  assign n40431 = n40430 ^ n28876 ^ n23222 ;
  assign n40432 = n20081 ^ n9994 ^ 1'b0 ;
  assign n40433 = n40432 ^ n32618 ^ n11680 ;
  assign n40434 = n12825 & n19444 ;
  assign n40435 = ~n6896 & n7700 ;
  assign n40436 = n6466 & ~n40435 ;
  assign n40437 = n11240 | n15477 ;
  assign n40438 = n461 | n40437 ;
  assign n40439 = ( n17081 & n40307 ) | ( n17081 & ~n40438 ) | ( n40307 & ~n40438 ) ;
  assign n40440 = n17004 & n34787 ;
  assign n40441 = ( n14939 & n40439 ) | ( n14939 & ~n40440 ) | ( n40439 & ~n40440 ) ;
  assign n40442 = n40441 ^ n38437 ^ 1'b0 ;
  assign n40443 = n6362 ^ n5588 ^ 1'b0 ;
  assign n40444 = n1169 & n40443 ;
  assign n40445 = ( n3060 & ~n26675 ) | ( n3060 & n40444 ) | ( ~n26675 & n40444 ) ;
  assign n40446 = ( n2540 & n9608 ) | ( n2540 & ~n15153 ) | ( n9608 & ~n15153 ) ;
  assign n40447 = n39091 ^ n1007 ^ 1'b0 ;
  assign n40448 = n23914 ^ n18581 ^ 1'b0 ;
  assign n40449 = n40447 & n40448 ;
  assign n40450 = n40449 ^ n22345 ^ 1'b0 ;
  assign n40451 = n40446 | n40450 ;
  assign n40452 = n20693 ^ n11641 ^ 1'b0 ;
  assign n40453 = ( n5205 & n15458 ) | ( n5205 & ~n37839 ) | ( n15458 & ~n37839 ) ;
  assign n40454 = ( n19055 & n40452 ) | ( n19055 & n40453 ) | ( n40452 & n40453 ) ;
  assign n40455 = n6296 & ~n12564 ;
  assign n40456 = n40455 ^ n37042 ^ 1'b0 ;
  assign n40457 = n40456 ^ n35507 ^ 1'b0 ;
  assign n40458 = n40454 & ~n40457 ;
  assign n40459 = n28204 ^ n26658 ^ n17224 ;
  assign n40460 = ( ~n785 & n10240 ) | ( ~n785 & n28132 ) | ( n10240 & n28132 ) ;
  assign n40461 = n40460 ^ n21046 ^ n8638 ;
  assign n40462 = n38414 ^ n22509 ^ n21274 ;
  assign n40463 = n23070 ^ n10569 ^ 1'b0 ;
  assign n40464 = ( n7479 & ~n8026 ) | ( n7479 & n40463 ) | ( ~n8026 & n40463 ) ;
  assign n40465 = n40464 ^ n38975 ^ 1'b0 ;
  assign n40466 = n38293 ^ n16615 ^ n298 ;
  assign n40467 = n13233 | n25468 ;
  assign n40468 = n26940 & n35060 ;
  assign n40469 = n37723 ^ n28257 ^ n4761 ;
  assign n40470 = n40469 ^ n27109 ^ 1'b0 ;
  assign n40471 = n40468 | n40470 ;
  assign n40473 = n20273 ^ n18086 ^ n3757 ;
  assign n40472 = ~n4464 & n31029 ;
  assign n40474 = n40473 ^ n40472 ^ 1'b0 ;
  assign n40475 = n40474 ^ n31207 ^ n19257 ;
  assign n40476 = ( n978 & n13481 ) | ( n978 & n33437 ) | ( n13481 & n33437 ) ;
  assign n40477 = ( n17977 & ~n29436 ) | ( n17977 & n40476 ) | ( ~n29436 & n40476 ) ;
  assign n40480 = n16581 ^ n16157 ^ n10381 ;
  assign n40478 = n4945 | n6673 ;
  assign n40479 = n36514 & n40478 ;
  assign n40481 = n40480 ^ n40479 ^ n22178 ;
  assign n40482 = ( ~n933 & n19030 ) | ( ~n933 & n20903 ) | ( n19030 & n20903 ) ;
  assign n40483 = ~n271 & n29676 ;
  assign n40484 = n14047 ^ n7270 ^ 1'b0 ;
  assign n40485 = ~n17914 & n40484 ;
  assign n40486 = n40485 ^ n3564 ^ 1'b0 ;
  assign n40487 = n9293 & ~n40486 ;
  assign n40488 = n8308 & n20107 ;
  assign n40489 = x37 & n40488 ;
  assign n40490 = n40489 ^ n15891 ^ 1'b0 ;
  assign n40491 = ( ~n21143 & n30446 ) | ( ~n21143 & n40490 ) | ( n30446 & n40490 ) ;
  assign n40492 = ( n15194 & ~n22337 ) | ( n15194 & n22879 ) | ( ~n22337 & n22879 ) ;
  assign n40493 = n40492 ^ n40473 ^ n23712 ;
  assign n40494 = ~n16544 & n34847 ;
  assign n40495 = n5398 | n40494 ;
  assign n40496 = n3423 | n40495 ;
  assign n40497 = ( ~n2708 & n16704 ) | ( ~n2708 & n40496 ) | ( n16704 & n40496 ) ;
  assign n40498 = n17671 & n34521 ;
  assign n40499 = ( n17507 & ~n19550 ) | ( n17507 & n40498 ) | ( ~n19550 & n40498 ) ;
  assign n40500 = n11676 ^ n4957 ^ 1'b0 ;
  assign n40501 = ( x8 & n3593 ) | ( x8 & n10896 ) | ( n3593 & n10896 ) ;
  assign n40502 = n40501 ^ n16354 ^ n12917 ;
  assign n40503 = n40502 ^ n20871 ^ 1'b0 ;
  assign n40504 = ~n2098 & n40503 ;
  assign n40505 = n40504 ^ n33138 ^ n20793 ;
  assign n40506 = n7703 & n20285 ;
  assign n40507 = n40506 ^ n5694 ^ 1'b0 ;
  assign n40508 = ( n11686 & ~n14575 ) | ( n11686 & n40507 ) | ( ~n14575 & n40507 ) ;
  assign n40509 = ( n40500 & n40505 ) | ( n40500 & n40508 ) | ( n40505 & n40508 ) ;
  assign n40510 = n26010 ^ n11183 ^ 1'b0 ;
  assign n40511 = n14414 & n40510 ;
  assign n40512 = n40511 ^ n8926 ^ n922 ;
  assign n40516 = n21756 ^ n6632 ^ n733 ;
  assign n40517 = ( ~n19432 & n28510 ) | ( ~n19432 & n40516 ) | ( n28510 & n40516 ) ;
  assign n40514 = n30772 ^ n4247 ^ 1'b0 ;
  assign n40515 = ~n2355 & n40514 ;
  assign n40513 = n25522 ^ n23254 ^ n9496 ;
  assign n40518 = n40517 ^ n40515 ^ n40513 ;
  assign n40519 = n35183 ^ n21219 ^ n1797 ;
  assign n40520 = ( ~n16175 & n27810 ) | ( ~n16175 & n40519 ) | ( n27810 & n40519 ) ;
  assign n40521 = n34250 ^ n9333 ^ 1'b0 ;
  assign n40522 = ( n5065 & n23856 ) | ( n5065 & ~n40521 ) | ( n23856 & ~n40521 ) ;
  assign n40523 = ( ~n40518 & n40520 ) | ( ~n40518 & n40522 ) | ( n40520 & n40522 ) ;
  assign n40524 = ( n2508 & ~n4710 ) | ( n2508 & n9932 ) | ( ~n4710 & n9932 ) ;
  assign n40525 = n16598 & ~n20592 ;
  assign n40526 = n40524 & n40525 ;
  assign n40527 = ( n3739 & n5015 ) | ( n3739 & ~n18540 ) | ( n5015 & ~n18540 ) ;
  assign n40528 = n40527 ^ n36889 ^ n21223 ;
  assign n40529 = n8745 | n18687 ;
  assign n40530 = ( n8422 & n15853 ) | ( n8422 & n40529 ) | ( n15853 & n40529 ) ;
  assign n40531 = n40530 ^ n33686 ^ n15496 ;
  assign n40534 = ( n10434 & ~n25882 ) | ( n10434 & n26121 ) | ( ~n25882 & n26121 ) ;
  assign n40532 = ( n1905 & ~n5598 ) | ( n1905 & n7825 ) | ( ~n5598 & n7825 ) ;
  assign n40533 = n14702 & ~n40532 ;
  assign n40535 = n40534 ^ n40533 ^ n21859 ;
  assign n40536 = n18584 & ~n21096 ;
  assign n40537 = n40536 ^ n29319 ^ 1'b0 ;
  assign n40538 = n6890 ^ n6340 ^ n1037 ;
  assign n40539 = n40538 ^ x87 ^ 1'b0 ;
  assign n40540 = n3983 & n40539 ;
  assign n40541 = n6706 | n38990 ;
  assign n40542 = n40540 | n40541 ;
  assign n40543 = n16260 ^ n13647 ^ 1'b0 ;
  assign n40544 = n40543 ^ n7021 ^ 1'b0 ;
  assign n40545 = n14927 & ~n40544 ;
  assign n40548 = n15377 ^ n14485 ^ n4235 ;
  assign n40549 = ( n6887 & n23066 ) | ( n6887 & n40548 ) | ( n23066 & n40548 ) ;
  assign n40547 = n271 & ~n5062 ;
  assign n40546 = n18544 ^ n11480 ^ n2383 ;
  assign n40550 = n40549 ^ n40547 ^ n40546 ;
  assign n40551 = n28221 ^ n4743 ^ n4128 ;
  assign n40552 = ~n37304 & n40551 ;
  assign n40553 = ( n13955 & n16513 ) | ( n13955 & n40552 ) | ( n16513 & n40552 ) ;
  assign n40554 = ~n14603 & n18428 ;
  assign n40555 = n12566 ^ n8605 ^ 1'b0 ;
  assign n40556 = n40555 ^ n7764 ^ 1'b0 ;
  assign n40557 = n40554 | n40556 ;
  assign n40558 = n40557 ^ n7029 ^ n5139 ;
  assign n40559 = ( n40550 & n40553 ) | ( n40550 & ~n40558 ) | ( n40553 & ~n40558 ) ;
  assign n40560 = ( ~n3934 & n18179 ) | ( ~n3934 & n26121 ) | ( n18179 & n26121 ) ;
  assign n40561 = n40560 ^ n31844 ^ n17233 ;
  assign n40562 = ( n26422 & ~n29246 ) | ( n26422 & n40561 ) | ( ~n29246 & n40561 ) ;
  assign n40563 = n40562 ^ n29992 ^ n21532 ;
  assign n40564 = n7694 & ~n16455 ;
  assign n40565 = n40564 ^ n29031 ^ n18865 ;
  assign n40566 = n12199 & n40565 ;
  assign n40567 = n40566 ^ n32551 ^ 1'b0 ;
  assign n40568 = ~n24223 & n33998 ;
  assign n40569 = ( n9254 & n30156 ) | ( n9254 & n30665 ) | ( n30156 & n30665 ) ;
  assign n40570 = ~n6772 & n23748 ;
  assign n40571 = n40570 ^ n18280 ^ 1'b0 ;
  assign n40572 = ( n16611 & ~n40569 ) | ( n16611 & n40571 ) | ( ~n40569 & n40571 ) ;
  assign n40573 = ( n5765 & n8504 ) | ( n5765 & ~n40572 ) | ( n8504 & ~n40572 ) ;
  assign n40574 = n25452 ^ n19141 ^ n14948 ;
  assign n40575 = n25816 ^ n17124 ^ 1'b0 ;
  assign n40576 = ( ~n22132 & n28816 ) | ( ~n22132 & n40575 ) | ( n28816 & n40575 ) ;
  assign n40577 = n1202 | n6017 ;
  assign n40578 = n35575 ^ n15321 ^ n8770 ;
  assign n40579 = ( n7360 & n40577 ) | ( n7360 & ~n40578 ) | ( n40577 & ~n40578 ) ;
  assign n40580 = n14078 ^ n11955 ^ 1'b0 ;
  assign n40581 = n17172 & ~n26589 ;
  assign n40582 = n40580 & ~n40581 ;
  assign n40583 = n35633 ^ n33770 ^ n33437 ;
  assign n40584 = ~n14645 & n40583 ;
  assign n40585 = ( ~n6380 & n23876 ) | ( ~n6380 & n30148 ) | ( n23876 & n30148 ) ;
  assign n40586 = n520 | n40585 ;
  assign n40587 = n2031 | n40586 ;
  assign n40588 = n11536 ^ n11506 ^ 1'b0 ;
  assign n40589 = n18836 ^ n15303 ^ 1'b0 ;
  assign n40590 = ( ~n6618 & n13443 ) | ( ~n6618 & n28600 ) | ( n13443 & n28600 ) ;
  assign n40591 = ( ~n11614 & n40589 ) | ( ~n11614 & n40590 ) | ( n40589 & n40590 ) ;
  assign n40592 = ( n8534 & ~n14635 ) | ( n8534 & n17772 ) | ( ~n14635 & n17772 ) ;
  assign n40599 = n19255 | n24724 ;
  assign n40600 = n12336 & ~n40599 ;
  assign n40597 = n11720 ^ n11682 ^ 1'b0 ;
  assign n40593 = n29529 ^ n2296 ^ 1'b0 ;
  assign n40594 = n4301 & n40593 ;
  assign n40595 = n40594 ^ n25514 ^ n21801 ;
  assign n40596 = n20381 & n40595 ;
  assign n40598 = n40597 ^ n40596 ^ 1'b0 ;
  assign n40601 = n40600 ^ n40598 ^ n36474 ;
  assign n40602 = n27119 ^ n19382 ^ 1'b0 ;
  assign n40603 = n40602 ^ n21862 ^ n298 ;
  assign n40604 = ~n11520 & n19047 ;
  assign n40605 = ~n29855 & n40604 ;
  assign n40606 = n3036 | n40605 ;
  assign n40607 = n40606 ^ n21711 ^ 1'b0 ;
  assign n40608 = n25785 ^ n5765 ^ 1'b0 ;
  assign n40609 = ~n35924 & n40608 ;
  assign n40610 = ~n12595 & n16749 ;
  assign n40611 = ( ~n14367 & n14793 ) | ( ~n14367 & n40610 ) | ( n14793 & n40610 ) ;
  assign n40612 = n1248 & ~n33129 ;
  assign n40613 = ( n13314 & n40611 ) | ( n13314 & n40612 ) | ( n40611 & n40612 ) ;
  assign n40614 = n13731 ^ n2584 ^ 1'b0 ;
  assign n40615 = n13127 & ~n40614 ;
  assign n40616 = n40615 ^ n6261 ^ 1'b0 ;
  assign n40617 = ( n7227 & ~n14877 ) | ( n7227 & n40616 ) | ( ~n14877 & n40616 ) ;
  assign n40618 = n9000 | n11025 ;
  assign n40619 = n40618 ^ n39743 ^ 1'b0 ;
  assign n40620 = n40619 ^ n21675 ^ 1'b0 ;
  assign n40621 = n6869 & n9922 ;
  assign n40622 = n9176 & n40621 ;
  assign n40623 = n40622 ^ n35817 ^ n32926 ;
  assign n40624 = n20069 ^ n9032 ^ 1'b0 ;
  assign n40625 = n30720 | n40624 ;
  assign n40626 = n37789 & ~n40625 ;
  assign n40627 = n40626 ^ n9223 ^ 1'b0 ;
  assign n40628 = n30547 ^ n30330 ^ 1'b0 ;
  assign n40629 = n34444 & n40628 ;
  assign n40630 = ( n5212 & n21982 ) | ( n5212 & ~n28052 ) | ( n21982 & ~n28052 ) ;
  assign n40631 = n40630 ^ n30898 ^ n20169 ;
  assign n40632 = n40631 ^ n494 ^ 1'b0 ;
  assign n40633 = ( n341 & ~n6290 ) | ( n341 & n36049 ) | ( ~n6290 & n36049 ) ;
  assign n40634 = n4383 & n8554 ;
  assign n40635 = ( n12087 & n39310 ) | ( n12087 & ~n40634 ) | ( n39310 & ~n40634 ) ;
  assign n40640 = n25554 ^ n21172 ^ n13199 ;
  assign n40636 = n17191 ^ n3914 ^ 1'b0 ;
  assign n40637 = n38540 | n40636 ;
  assign n40638 = n40637 ^ n23988 ^ n23749 ;
  assign n40639 = ( n8501 & n18979 ) | ( n8501 & n40638 ) | ( n18979 & n40638 ) ;
  assign n40641 = n40640 ^ n40639 ^ n22935 ;
  assign n40642 = ( n1319 & ~n40294 ) | ( n1319 & n40641 ) | ( ~n40294 & n40641 ) ;
  assign n40643 = ( n6342 & ~n39446 ) | ( n6342 & n40642 ) | ( ~n39446 & n40642 ) ;
  assign n40644 = n31382 ^ n27527 ^ n15889 ;
  assign n40645 = n40644 ^ n22208 ^ n21782 ;
  assign n40646 = n9179 & n24357 ;
  assign n40647 = n40646 ^ n29911 ^ n1538 ;
  assign n40648 = ( n951 & ~n7775 ) | ( n951 & n28238 ) | ( ~n7775 & n28238 ) ;
  assign n40649 = n22481 | n32637 ;
  assign n40650 = n40648 & ~n40649 ;
  assign n40651 = n13143 & ~n40650 ;
  assign n40652 = ~n40647 & n40651 ;
  assign n40653 = n4567 | n6139 ;
  assign n40654 = n40653 ^ n23830 ^ 1'b0 ;
  assign n40655 = n40654 ^ n13657 ^ 1'b0 ;
  assign n40656 = ( n7389 & ~n14625 ) | ( n7389 & n27918 ) | ( ~n14625 & n27918 ) ;
  assign n40657 = n40655 | n40656 ;
  assign n40658 = ( ~n1757 & n4034 ) | ( ~n1757 & n12936 ) | ( n4034 & n12936 ) ;
  assign n40659 = ( ~n10349 & n29345 ) | ( ~n10349 & n31415 ) | ( n29345 & n31415 ) ;
  assign n40660 = ( n9251 & n20519 ) | ( n9251 & ~n40659 ) | ( n20519 & ~n40659 ) ;
  assign n40661 = ( n8611 & n23533 ) | ( n8611 & ~n40660 ) | ( n23533 & ~n40660 ) ;
  assign n40662 = n1849 & n2392 ;
  assign n40663 = ( ~n7126 & n25206 ) | ( ~n7126 & n40662 ) | ( n25206 & n40662 ) ;
  assign n40664 = n5107 & n28600 ;
  assign n40665 = n40664 ^ n32010 ^ n4583 ;
  assign n40666 = ( ~n28575 & n40663 ) | ( ~n28575 & n40665 ) | ( n40663 & n40665 ) ;
  assign n40667 = ~n12745 & n16093 ;
  assign n40668 = n40667 ^ n1855 ^ 1'b0 ;
  assign n40669 = n12216 & n40668 ;
  assign n40670 = ( n5421 & n37667 ) | ( n5421 & ~n40669 ) | ( n37667 & ~n40669 ) ;
  assign n40671 = ( n7327 & ~n8588 ) | ( n7327 & n38138 ) | ( ~n8588 & n38138 ) ;
  assign n40676 = n735 & ~n14021 ;
  assign n40672 = ( ~n20883 & n27171 ) | ( ~n20883 & n28858 ) | ( n27171 & n28858 ) ;
  assign n40673 = n21936 | n23755 ;
  assign n40674 = n33953 & ~n40673 ;
  assign n40675 = n40672 | n40674 ;
  assign n40677 = n40676 ^ n40675 ^ 1'b0 ;
  assign n40678 = n19497 ^ n6557 ^ 1'b0 ;
  assign n40679 = n4965 ^ n4615 ^ 1'b0 ;
  assign n40680 = n1880 & n40679 ;
  assign n40681 = ( n3720 & n15748 ) | ( n3720 & ~n40680 ) | ( n15748 & ~n40680 ) ;
  assign n40682 = n40681 ^ n16278 ^ 1'b0 ;
  assign n40683 = n27543 & n40682 ;
  assign n40684 = n40683 ^ n34462 ^ n5599 ;
  assign n40685 = n29950 ^ n13594 ^ n7819 ;
  assign n40686 = n39876 ^ n7981 ^ 1'b0 ;
  assign n40687 = n16689 & ~n40686 ;
  assign n40688 = ( n20338 & ~n22222 ) | ( n20338 & n40687 ) | ( ~n22222 & n40687 ) ;
  assign n40689 = n1046 ^ n772 ^ 1'b0 ;
  assign n40690 = n40689 ^ n24701 ^ n20052 ;
  assign n40691 = n31066 ^ n15932 ^ 1'b0 ;
  assign n40692 = n37704 ^ n22506 ^ 1'b0 ;
  assign n40693 = n23865 ^ n21069 ^ 1'b0 ;
  assign n40694 = n40692 | n40693 ;
  assign n40698 = n15252 ^ n10949 ^ n513 ;
  assign n40695 = ~n2903 & n13941 ;
  assign n40696 = n40695 ^ n591 ^ 1'b0 ;
  assign n40697 = ( n5663 & ~n31180 ) | ( n5663 & n40696 ) | ( ~n31180 & n40696 ) ;
  assign n40699 = n40698 ^ n40697 ^ n32971 ;
  assign n40700 = n18381 ^ n14215 ^ n9985 ;
  assign n40701 = n40700 ^ n18407 ^ n8079 ;
  assign n40702 = ( n13163 & ~n16278 ) | ( n13163 & n40701 ) | ( ~n16278 & n40701 ) ;
  assign n40703 = n16010 ^ n4896 ^ n3067 ;
  assign n40704 = n33648 ^ n13719 ^ n7649 ;
  assign n40705 = ( n34852 & n40703 ) | ( n34852 & n40704 ) | ( n40703 & n40704 ) ;
  assign n40706 = n39982 ^ n39737 ^ n12205 ;
  assign n40707 = n40706 ^ n22959 ^ n17639 ;
  assign n40710 = n12442 & n13922 ;
  assign n40708 = n31935 ^ n10873 ^ n7810 ;
  assign n40709 = n16267 & n40708 ;
  assign n40711 = n40710 ^ n40709 ^ 1'b0 ;
  assign n40712 = n24731 ^ n5078 ^ 1'b0 ;
  assign n40713 = ( ~n1152 & n7403 ) | ( ~n1152 & n17142 ) | ( n7403 & n17142 ) ;
  assign n40714 = n40713 ^ n11055 ^ n903 ;
  assign n40715 = n15345 ^ n4609 ^ n4017 ;
  assign n40716 = n16510 & ~n40715 ;
  assign n40717 = ( n16954 & n18402 ) | ( n16954 & ~n38907 ) | ( n18402 & ~n38907 ) ;
  assign n40718 = ( n502 & n7054 ) | ( n502 & n7761 ) | ( n7054 & n7761 ) ;
  assign n40719 = n11821 ^ n2017 ^ 1'b0 ;
  assign n40720 = ~n40718 & n40719 ;
  assign n40721 = ~n20088 & n40720 ;
  assign n40722 = n7152 & n40721 ;
  assign n40723 = ( ~n20993 & n21365 ) | ( ~n20993 & n22273 ) | ( n21365 & n22273 ) ;
  assign n40724 = n34336 ^ n13592 ^ n8122 ;
  assign n40729 = n39297 ^ n36023 ^ 1'b0 ;
  assign n40725 = n34816 ^ n11710 ^ n9239 ;
  assign n40726 = n40725 ^ n19499 ^ n5319 ;
  assign n40727 = n5627 | n40726 ;
  assign n40728 = n40727 ^ n15269 ^ 1'b0 ;
  assign n40730 = n40729 ^ n40728 ^ n23877 ;
  assign n40731 = ( n10307 & ~n16004 ) | ( n10307 & n24424 ) | ( ~n16004 & n24424 ) ;
  assign n40732 = n40731 ^ n6062 ^ 1'b0 ;
  assign n40733 = n24317 ^ n21787 ^ n1936 ;
  assign n40734 = n40733 ^ n10476 ^ 1'b0 ;
  assign n40735 = ( n4757 & n17906 ) | ( n4757 & n40734 ) | ( n17906 & n40734 ) ;
  assign n40736 = n11292 ^ n2111 ^ n365 ;
  assign n40737 = n40736 ^ n8237 ^ 1'b0 ;
  assign n40738 = ~n13462 & n40737 ;
  assign n40739 = n40738 ^ n19585 ^ 1'b0 ;
  assign n40740 = n40739 ^ n10958 ^ n7909 ;
  assign n40741 = n40740 ^ n12366 ^ n5534 ;
  assign n40742 = n38223 ^ n7018 ^ 1'b0 ;
  assign n40743 = ~n40741 & n40742 ;
  assign n40744 = ( ~n8391 & n10676 ) | ( ~n8391 & n16630 ) | ( n10676 & n16630 ) ;
  assign n40745 = ( ~n6204 & n25833 ) | ( ~n6204 & n40744 ) | ( n25833 & n40744 ) ;
  assign n40746 = ( n14896 & ~n18198 ) | ( n14896 & n21812 ) | ( ~n18198 & n21812 ) ;
  assign n40747 = ( n1665 & ~n6370 ) | ( n1665 & n21002 ) | ( ~n6370 & n21002 ) ;
  assign n40748 = n11797 ^ n7662 ^ 1'b0 ;
  assign n40749 = ~n38718 & n40748 ;
  assign n40750 = ~n10490 & n13506 ;
  assign n40751 = n40750 ^ n13759 ^ 1'b0 ;
  assign n40752 = ( n6407 & ~n29143 ) | ( n6407 & n40751 ) | ( ~n29143 & n40751 ) ;
  assign n40753 = n40752 ^ n2528 ^ 1'b0 ;
  assign n40754 = n39372 & ~n40753 ;
  assign n40755 = ( n28032 & ~n40749 ) | ( n28032 & n40754 ) | ( ~n40749 & n40754 ) ;
  assign n40756 = n4161 & n22343 ;
  assign n40757 = ( n809 & n18963 ) | ( n809 & n40756 ) | ( n18963 & n40756 ) ;
  assign n40758 = ( n2846 & n4663 ) | ( n2846 & n33844 ) | ( n4663 & n33844 ) ;
  assign n40759 = n11577 ^ x84 ^ 1'b0 ;
  assign n40760 = n40759 ^ n13849 ^ 1'b0 ;
  assign n40761 = n7141 & ~n40760 ;
  assign n40762 = n40758 & n40761 ;
  assign n40763 = n26087 ^ n24162 ^ n20109 ;
  assign n40764 = n40763 ^ n12840 ^ 1'b0 ;
  assign n40765 = ~n20958 & n40764 ;
  assign n40766 = n2846 ^ n2741 ^ 1'b0 ;
  assign n40767 = n40765 & n40766 ;
  assign n40768 = n14209 & n40767 ;
  assign n40769 = n28482 ^ n16066 ^ 1'b0 ;
  assign n40770 = n4916 & n31452 ;
  assign n40771 = ( n10523 & n14434 ) | ( n10523 & n40770 ) | ( n14434 & n40770 ) ;
  assign n40772 = ( n9864 & n13817 ) | ( n9864 & n30305 ) | ( n13817 & n30305 ) ;
  assign n40773 = n21309 ^ n17116 ^ 1'b0 ;
  assign n40774 = n922 & n40773 ;
  assign n40775 = n40772 & n40774 ;
  assign n40776 = ( n674 & n24203 ) | ( n674 & n40775 ) | ( n24203 & n40775 ) ;
  assign n40777 = n16784 ^ n8963 ^ n6515 ;
  assign n40778 = n40777 ^ n30711 ^ n18804 ;
  assign n40779 = ( ~n23127 & n27216 ) | ( ~n23127 & n40778 ) | ( n27216 & n40778 ) ;
  assign n40780 = ( n10808 & ~n27984 ) | ( n10808 & n40779 ) | ( ~n27984 & n40779 ) ;
  assign n40781 = ( ~n27830 & n33961 ) | ( ~n27830 & n35132 ) | ( n33961 & n35132 ) ;
  assign n40782 = ( ~n2186 & n17183 ) | ( ~n2186 & n36319 ) | ( n17183 & n36319 ) ;
  assign n40783 = n17204 ^ n12209 ^ n6169 ;
  assign n40784 = n4312 ^ n3990 ^ 1'b0 ;
  assign n40785 = ~n6464 & n40784 ;
  assign n40786 = n3071 & n40785 ;
  assign n40787 = ( n24422 & ~n40783 ) | ( n24422 & n40786 ) | ( ~n40783 & n40786 ) ;
  assign n40788 = ~n13775 & n22539 ;
  assign n40791 = ( n820 & ~n1243 ) | ( n820 & n5042 ) | ( ~n1243 & n5042 ) ;
  assign n40792 = ( ~n4645 & n5429 ) | ( ~n4645 & n26773 ) | ( n5429 & n26773 ) ;
  assign n40793 = ( n32593 & n40791 ) | ( n32593 & ~n40792 ) | ( n40791 & ~n40792 ) ;
  assign n40789 = n31665 ^ n11578 ^ n6450 ;
  assign n40790 = n40789 ^ n9464 ^ 1'b0 ;
  assign n40794 = n40793 ^ n40790 ^ n27503 ;
  assign n40795 = n6029 & n19493 ;
  assign n40796 = ( n478 & ~n5911 ) | ( n478 & n19793 ) | ( ~n5911 & n19793 ) ;
  assign n40797 = n40796 ^ n12652 ^ 1'b0 ;
  assign n40798 = ( n30668 & n32536 ) | ( n30668 & n40585 ) | ( n32536 & n40585 ) ;
  assign n40799 = ~n1646 & n2175 ;
  assign n40800 = n40799 ^ n31733 ^ n11308 ;
  assign n40801 = ( n18982 & n20503 ) | ( n18982 & n40800 ) | ( n20503 & n40800 ) ;
  assign n40802 = n9516 & n40801 ;
  assign n40803 = ( n4579 & n10530 ) | ( n4579 & n30277 ) | ( n10530 & n30277 ) ;
  assign n40804 = n21522 ^ n14658 ^ 1'b0 ;
  assign n40805 = ~n34954 & n40804 ;
  assign n40806 = n270 | n8585 ;
  assign n40807 = n2943 | n40806 ;
  assign n40808 = ( n779 & n2964 ) | ( n779 & n3212 ) | ( n2964 & n3212 ) ;
  assign n40809 = n8163 ^ n5312 ^ 1'b0 ;
  assign n40810 = ( ~n19729 & n40808 ) | ( ~n19729 & n40809 ) | ( n40808 & n40809 ) ;
  assign n40811 = n8707 ^ n6537 ^ 1'b0 ;
  assign n40812 = n5332 | n40811 ;
  assign n40813 = n3239 & ~n40812 ;
  assign n40814 = ~n40810 & n40813 ;
  assign n40815 = n40580 ^ n10207 ^ n6730 ;
  assign n40816 = ( ~n6621 & n19349 ) | ( ~n6621 & n40815 ) | ( n19349 & n40815 ) ;
  assign n40817 = ( n17232 & n25378 ) | ( n17232 & n38744 ) | ( n25378 & n38744 ) ;
  assign n40818 = n17335 ^ n4328 ^ 1'b0 ;
  assign n40822 = n4633 & n11748 ;
  assign n40823 = ~n11748 & n40822 ;
  assign n40824 = n9896 & ~n40823 ;
  assign n40825 = ~n9896 & n40824 ;
  assign n40819 = n16925 & n19342 ;
  assign n40820 = n40819 ^ n4097 ^ 1'b0 ;
  assign n40821 = n18318 | n40820 ;
  assign n40826 = n40825 ^ n40821 ^ 1'b0 ;
  assign n40827 = n40826 ^ n39711 ^ n23236 ;
  assign n40829 = ( n14407 & ~n16013 ) | ( n14407 & n27632 ) | ( ~n16013 & n27632 ) ;
  assign n40828 = ~n2828 & n20025 ;
  assign n40830 = n40829 ^ n40828 ^ 1'b0 ;
  assign n40831 = n6982 & n40830 ;
  assign n40832 = ~n11195 & n17516 ;
  assign n40833 = n40832 ^ n33692 ^ 1'b0 ;
  assign n40834 = ( n14602 & n19549 ) | ( n14602 & ~n25956 ) | ( n19549 & ~n25956 ) ;
  assign n40835 = ~n19239 & n23849 ;
  assign n40836 = n40835 ^ n37326 ^ 1'b0 ;
  assign n40837 = n2015 | n11625 ;
  assign n40838 = n38985 ^ n24514 ^ 1'b0 ;
  assign n40839 = n9536 ^ n8856 ^ n5440 ;
  assign n40840 = n17407 ^ n13181 ^ n1635 ;
  assign n40841 = n33681 & n40840 ;
  assign n40842 = n40841 ^ n22344 ^ 1'b0 ;
  assign n40843 = ( ~n6972 & n18096 ) | ( ~n6972 & n40842 ) | ( n18096 & n40842 ) ;
  assign n40844 = n23576 ^ n13071 ^ n5216 ;
  assign n40845 = n22486 ^ n11760 ^ 1'b0 ;
  assign n40846 = ( n26332 & ~n30917 ) | ( n26332 & n31874 ) | ( ~n30917 & n31874 ) ;
  assign n40847 = n40846 ^ n13652 ^ 1'b0 ;
  assign n40854 = ( ~n11634 & n23095 ) | ( ~n11634 & n28186 ) | ( n23095 & n28186 ) ;
  assign n40855 = n40854 ^ n9252 ^ 1'b0 ;
  assign n40856 = n16689 & n40855 ;
  assign n40850 = n9674 ^ n6669 ^ n3309 ;
  assign n40851 = n40850 ^ n2884 ^ 1'b0 ;
  assign n40849 = ( n1933 & n2626 ) | ( n1933 & ~n11793 ) | ( n2626 & ~n11793 ) ;
  assign n40848 = n23399 ^ n10311 ^ n257 ;
  assign n40852 = n40851 ^ n40849 ^ n40848 ;
  assign n40853 = n40852 ^ n15853 ^ n15205 ;
  assign n40857 = n40856 ^ n40853 ^ n4092 ;
  assign n40858 = n25549 ^ n11740 ^ n8986 ;
  assign n40859 = n2504 & n16125 ;
  assign n40860 = ( n22880 & ~n40858 ) | ( n22880 & n40859 ) | ( ~n40858 & n40859 ) ;
  assign n40861 = n10766 & ~n34021 ;
  assign n40862 = ~n19089 & n40861 ;
  assign n40863 = n12165 | n40862 ;
  assign n40864 = ( n18369 & n18952 ) | ( n18369 & n40863 ) | ( n18952 & n40863 ) ;
  assign n40865 = n17547 ^ n3068 ^ 1'b0 ;
  assign n40866 = n21798 ^ n7940 ^ n706 ;
  assign n40867 = ( n11505 & n40865 ) | ( n11505 & n40866 ) | ( n40865 & n40866 ) ;
  assign n40868 = ( n4342 & n13166 ) | ( n4342 & ~n25882 ) | ( n13166 & ~n25882 ) ;
  assign n40869 = n4934 | n18820 ;
  assign n40870 = n10735 & ~n40869 ;
  assign n40871 = n9210 & ~n40870 ;
  assign n40872 = n40871 ^ n21101 ^ 1'b0 ;
  assign n40873 = n22565 & ~n40872 ;
  assign n40874 = n40873 ^ n37112 ^ 1'b0 ;
  assign n40875 = ( n33495 & n40868 ) | ( n33495 & n40874 ) | ( n40868 & n40874 ) ;
  assign n40876 = ~n3356 & n32951 ;
  assign n40877 = n40876 ^ n24518 ^ 1'b0 ;
  assign n40878 = n19671 ^ n6166 ^ n5240 ;
  assign n40879 = n18663 | n24253 ;
  assign n40880 = n40878 & ~n40879 ;
  assign n40881 = ~n33237 & n35133 ;
  assign n40882 = ~n16947 & n20429 ;
  assign n40883 = n40882 ^ n1637 ^ 1'b0 ;
  assign n40884 = n40883 ^ n38746 ^ n25681 ;
  assign n40885 = n2113 | n4155 ;
  assign n40886 = n21927 | n40885 ;
  assign n40887 = ( n15674 & n30463 ) | ( n15674 & n40886 ) | ( n30463 & n40886 ) ;
  assign n40888 = n3134 & n40887 ;
  assign n40889 = n33529 ^ n21200 ^ 1'b0 ;
  assign n40892 = n9071 ^ n3259 ^ 1'b0 ;
  assign n40893 = n25610 | n40892 ;
  assign n40890 = n32714 ^ n25869 ^ n16321 ;
  assign n40891 = n8647 & ~n40890 ;
  assign n40894 = n40893 ^ n40891 ^ 1'b0 ;
  assign n40895 = n38939 ^ n38189 ^ n3097 ;
  assign n40896 = n40895 ^ n34715 ^ 1'b0 ;
  assign n40897 = n33591 ^ n2890 ^ x36 ;
  assign n40898 = n15925 & n40897 ;
  assign n40899 = n40898 ^ n19918 ^ 1'b0 ;
  assign n40900 = n36086 ^ n26701 ^ 1'b0 ;
  assign n40901 = n1619 | n5261 ;
  assign n40902 = ( n2011 & n32544 ) | ( n2011 & n40901 ) | ( n32544 & n40901 ) ;
  assign n40903 = ( n27373 & n39269 ) | ( n27373 & n40902 ) | ( n39269 & n40902 ) ;
  assign n40904 = n27080 ^ n17591 ^ n9653 ;
  assign n40905 = ( x212 & n25049 ) | ( x212 & ~n30577 ) | ( n25049 & ~n30577 ) ;
  assign n40906 = n40905 ^ n4181 ^ 1'b0 ;
  assign n40907 = ( ~n8116 & n25080 ) | ( ~n8116 & n40906 ) | ( n25080 & n40906 ) ;
  assign n40908 = n32186 ^ n29529 ^ n21875 ;
  assign n40909 = ( ~n22393 & n28592 ) | ( ~n22393 & n40908 ) | ( n28592 & n40908 ) ;
  assign n40910 = ( n15459 & n24702 ) | ( n15459 & n40909 ) | ( n24702 & n40909 ) ;
  assign n40911 = ( n1126 & n33823 ) | ( n1126 & ~n40910 ) | ( n33823 & ~n40910 ) ;
  assign n40912 = n20054 ^ n11036 ^ 1'b0 ;
  assign n40913 = n3769 & ~n40912 ;
  assign n40914 = n40913 ^ n14498 ^ n3766 ;
  assign n40915 = n40914 ^ n2516 ^ 1'b0 ;
  assign n40916 = ( n25712 & n40911 ) | ( n25712 & ~n40915 ) | ( n40911 & ~n40915 ) ;
  assign n40917 = ( n4527 & n17731 ) | ( n4527 & ~n33523 ) | ( n17731 & ~n33523 ) ;
  assign n40918 = ~n6387 & n22981 ;
  assign n40919 = n526 & n23225 ;
  assign n40920 = n40919 ^ n7889 ^ 1'b0 ;
  assign n40923 = n10913 & n14116 ;
  assign n40924 = n40923 ^ n9748 ^ 1'b0 ;
  assign n40925 = n40924 ^ n28953 ^ n13823 ;
  assign n40921 = n35052 ^ n16431 ^ n3691 ;
  assign n40922 = n20465 | n40921 ;
  assign n40926 = n40925 ^ n40922 ^ 1'b0 ;
  assign n40927 = n25383 ^ n16086 ^ n2736 ;
  assign n40928 = n40927 ^ n22188 ^ n11617 ;
  assign n40929 = n32475 ^ n13957 ^ n2603 ;
  assign n40930 = ( n7254 & ~n24474 ) | ( n7254 & n37137 ) | ( ~n24474 & n37137 ) ;
  assign n40931 = n40930 ^ n24963 ^ 1'b0 ;
  assign n40932 = n15383 & ~n28665 ;
  assign n40933 = n9144 ^ n4366 ^ n1101 ;
  assign n40934 = n40933 ^ n16657 ^ n15677 ;
  assign n40935 = n40934 ^ n13846 ^ 1'b0 ;
  assign n40936 = ~n20104 & n40935 ;
  assign n40937 = ( n33916 & ~n40932 ) | ( n33916 & n40936 ) | ( ~n40932 & n40936 ) ;
  assign n40938 = n383 & ~n33815 ;
  assign n40940 = n24871 ^ n8413 ^ n8034 ;
  assign n40939 = n11871 ^ n2092 ^ 1'b0 ;
  assign n40941 = n40940 ^ n40939 ^ n11209 ;
  assign n40942 = ~n8190 & n9463 ;
  assign n40943 = n14594 ^ n4339 ^ 1'b0 ;
  assign n40944 = n30173 & ~n40943 ;
  assign n40945 = n19068 ^ n14749 ^ 1'b0 ;
  assign n40946 = n5020 & ~n11137 ;
  assign n40947 = n40946 ^ n2850 ^ 1'b0 ;
  assign n40948 = ( n17186 & n23612 ) | ( n17186 & ~n40947 ) | ( n23612 & ~n40947 ) ;
  assign n40949 = ( n1560 & ~n28424 ) | ( n1560 & n40948 ) | ( ~n28424 & n40948 ) ;
  assign n40950 = n35846 ^ n13970 ^ 1'b0 ;
  assign n40951 = n29162 ^ n12884 ^ n4689 ;
  assign n40952 = n40951 ^ n22519 ^ 1'b0 ;
  assign n40953 = ( ~n317 & n7290 ) | ( ~n317 & n40952 ) | ( n7290 & n40952 ) ;
  assign n40954 = n29801 ^ n26566 ^ 1'b0 ;
  assign n40955 = n27732 & n40954 ;
  assign n40956 = n14745 ^ n10753 ^ 1'b0 ;
  assign n40957 = n40956 ^ n33973 ^ n7679 ;
  assign n40958 = ~n8026 & n35053 ;
  assign n40959 = ( n40955 & n40957 ) | ( n40955 & ~n40958 ) | ( n40957 & ~n40958 ) ;
  assign n40960 = n29241 ^ n5847 ^ n2797 ;
  assign n40961 = ( ~n19834 & n26412 ) | ( ~n19834 & n40960 ) | ( n26412 & n40960 ) ;
  assign n40962 = n22308 ^ n2963 ^ 1'b0 ;
  assign n40966 = n16882 ^ n8212 ^ n1787 ;
  assign n40963 = n33830 ^ n3225 ^ n906 ;
  assign n40964 = n532 & n40963 ;
  assign n40965 = n7991 & ~n40964 ;
  assign n40967 = n40966 ^ n40965 ^ 1'b0 ;
  assign n40968 = n16423 & ~n38592 ;
  assign n40969 = ~n4960 & n40968 ;
  assign n40970 = ( n22111 & n28666 ) | ( n22111 & ~n35825 ) | ( n28666 & ~n35825 ) ;
  assign n40971 = n20358 ^ n18536 ^ n11590 ;
  assign n40972 = n5762 ^ n4606 ^ n4172 ;
  assign n40973 = ( ~n14705 & n32265 ) | ( ~n14705 & n40972 ) | ( n32265 & n40972 ) ;
  assign n40974 = n4680 | n40973 ;
  assign n40975 = n40974 ^ n28769 ^ 1'b0 ;
  assign n40976 = ( n16429 & ~n40971 ) | ( n16429 & n40975 ) | ( ~n40971 & n40975 ) ;
  assign n40977 = ( n6275 & n16860 ) | ( n6275 & ~n28005 ) | ( n16860 & ~n28005 ) ;
  assign n40978 = n40977 ^ n5146 ^ n2527 ;
  assign n40981 = ( n3600 & n9514 ) | ( n3600 & ~n14173 ) | ( n9514 & ~n14173 ) ;
  assign n40982 = ~n13544 & n40981 ;
  assign n40983 = n40982 ^ n2200 ^ 1'b0 ;
  assign n40979 = n10995 & n35457 ;
  assign n40980 = n40979 ^ n16128 ^ 1'b0 ;
  assign n40984 = n40983 ^ n40980 ^ n34840 ;
  assign n40985 = ~n6166 & n11907 ;
  assign n40986 = n40985 ^ n1785 ^ 1'b0 ;
  assign n40987 = n17400 ^ n2725 ^ n2186 ;
  assign n40988 = n40987 ^ n33441 ^ n18869 ;
  assign n40989 = n10455 & ~n39427 ;
  assign n40990 = ~n4446 & n35930 ;
  assign n40991 = n12013 ^ n10919 ^ 1'b0 ;
  assign n40992 = n40990 & ~n40991 ;
  assign n40993 = n40992 ^ n36624 ^ n4320 ;
  assign n40995 = n33200 ^ n9465 ^ n3143 ;
  assign n40994 = ( ~n17953 & n37975 ) | ( ~n17953 & n39824 ) | ( n37975 & n39824 ) ;
  assign n40996 = n40995 ^ n40994 ^ n35746 ;
  assign n40997 = n22755 ^ n7556 ^ 1'b0 ;
  assign n40998 = n22743 | n40997 ;
  assign n40999 = n40998 ^ n18794 ^ n3672 ;
  assign n41000 = n23508 ^ n4817 ^ 1'b0 ;
  assign n41001 = ~n40999 & n41000 ;
  assign n41002 = n41001 ^ n20504 ^ n4842 ;
  assign n41005 = ( n4174 & n21644 ) | ( n4174 & ~n22092 ) | ( n21644 & ~n22092 ) ;
  assign n41003 = n10513 ^ n7204 ^ 1'b0 ;
  assign n41004 = ~n33119 & n41003 ;
  assign n41006 = n41005 ^ n41004 ^ n34526 ;
  assign n41007 = n38577 ^ n32978 ^ n29802 ;
  assign n41008 = n3675 | n27585 ;
  assign n41009 = n16481 | n41008 ;
  assign n41010 = ( ~n643 & n3162 ) | ( ~n643 & n19257 ) | ( n3162 & n19257 ) ;
  assign n41011 = n41010 ^ n10841 ^ n7345 ;
  assign n41012 = n7080 & ~n33056 ;
  assign n41013 = n41012 ^ n21969 ^ 1'b0 ;
  assign n41014 = ( n3575 & ~n6668 ) | ( n3575 & n15589 ) | ( ~n6668 & n15589 ) ;
  assign n41015 = ( n496 & n41013 ) | ( n496 & n41014 ) | ( n41013 & n41014 ) ;
  assign n41016 = n39933 ^ n13992 ^ x78 ;
  assign n41017 = n31341 ^ n12143 ^ 1'b0 ;
  assign n41018 = ( n36931 & ~n41016 ) | ( n36931 & n41017 ) | ( ~n41016 & n41017 ) ;
  assign n41019 = n10328 | n10638 ;
  assign n41020 = n21747 & ~n41019 ;
  assign n41021 = n41020 ^ n19429 ^ n10734 ;
  assign n41022 = n36447 ^ n13268 ^ n7830 ;
  assign n41023 = n452 | n30607 ;
  assign n41024 = n41023 ^ n25056 ^ 1'b0 ;
  assign n41025 = ( n21474 & n22297 ) | ( n21474 & n36668 ) | ( n22297 & n36668 ) ;
  assign n41026 = n7987 ^ n2186 ^ 1'b0 ;
  assign n41027 = ~n1405 & n41026 ;
  assign n41028 = n41027 ^ n22608 ^ 1'b0 ;
  assign n41029 = n41025 & ~n41028 ;
  assign n41030 = n4132 | n16692 ;
  assign n41031 = n35812 & ~n41030 ;
  assign n41032 = n26088 & ~n41031 ;
  assign n41033 = ~n7393 & n41032 ;
  assign n41034 = ~n4181 & n7101 ;
  assign n41035 = n747 & n41034 ;
  assign n41037 = ( n30322 & n33357 ) | ( n30322 & ~n34169 ) | ( n33357 & ~n34169 ) ;
  assign n41036 = ( n1759 & ~n8647 ) | ( n1759 & n36480 ) | ( ~n8647 & n36480 ) ;
  assign n41038 = n41037 ^ n41036 ^ n30294 ;
  assign n41039 = n6021 & n12664 ;
  assign n41040 = n41039 ^ n10557 ^ 1'b0 ;
  assign n41041 = ( n2688 & n29498 ) | ( n2688 & ~n41040 ) | ( n29498 & ~n41040 ) ;
  assign n41042 = ( n7235 & n9418 ) | ( n7235 & ~n29509 ) | ( n9418 & ~n29509 ) ;
  assign n41043 = n41042 ^ n21398 ^ 1'b0 ;
  assign n41044 = n24544 ^ n6990 ^ 1'b0 ;
  assign n41045 = n18769 ^ n10943 ^ n4272 ;
  assign n41046 = n12661 & ~n41045 ;
  assign n41047 = n21155 & ~n41046 ;
  assign n41048 = ~n18461 & n41047 ;
  assign n41049 = n28063 ^ n1032 ^ 1'b0 ;
  assign n41050 = n24885 & ~n41049 ;
  assign n41051 = n33926 ^ n6339 ^ x243 ;
  assign n41052 = n41051 ^ n22293 ^ 1'b0 ;
  assign n41053 = ( n10600 & ~n15950 ) | ( n10600 & n17064 ) | ( ~n15950 & n17064 ) ;
  assign n41055 = n28791 ^ n22925 ^ n8432 ;
  assign n41056 = ( n6650 & n9085 ) | ( n6650 & n24288 ) | ( n9085 & n24288 ) ;
  assign n41057 = n41056 ^ n5344 ^ n3822 ;
  assign n41058 = n10037 & ~n41057 ;
  assign n41059 = n2648 & n41058 ;
  assign n41060 = ~n36583 & n41059 ;
  assign n41061 = ( n2209 & n41055 ) | ( n2209 & ~n41060 ) | ( n41055 & ~n41060 ) ;
  assign n41054 = n7294 | n16937 ;
  assign n41062 = n41061 ^ n41054 ^ 1'b0 ;
  assign n41063 = n33705 ^ n19646 ^ n19207 ;
  assign n41064 = n27664 ^ n9836 ^ 1'b0 ;
  assign n41065 = n41063 & ~n41064 ;
  assign n41066 = n733 & ~n2486 ;
  assign n41067 = n41066 ^ n31591 ^ n3847 ;
  assign n41068 = n29518 & n41067 ;
  assign n41069 = n39533 ^ n29797 ^ n13733 ;
  assign n41070 = ( n3813 & ~n6598 ) | ( n3813 & n25837 ) | ( ~n6598 & n25837 ) ;
  assign n41071 = n41070 ^ n29175 ^ n23715 ;
  assign n41073 = ~n570 & n29838 ;
  assign n41074 = ~n5739 & n41073 ;
  assign n41072 = n5980 & n13470 ;
  assign n41075 = n41074 ^ n41072 ^ n25150 ;
  assign n41076 = ( n4611 & n5107 ) | ( n4611 & n17496 ) | ( n5107 & n17496 ) ;
  assign n41077 = ( n5808 & n22891 ) | ( n5808 & n41076 ) | ( n22891 & n41076 ) ;
  assign n41078 = n3574 & n7862 ;
  assign n41079 = n41078 ^ n39637 ^ 1'b0 ;
  assign n41081 = n22330 ^ n17172 ^ n14560 ;
  assign n41080 = x177 & ~n22069 ;
  assign n41082 = n41081 ^ n41080 ^ 1'b0 ;
  assign n41083 = n2550 & n13578 ;
  assign n41084 = n41083 ^ n16633 ^ 1'b0 ;
  assign n41085 = n29630 ^ n17333 ^ n3859 ;
  assign n41086 = n41085 ^ n36545 ^ n30203 ;
  assign n41087 = n4735 | n26525 ;
  assign n41088 = ( ~n1569 & n13983 ) | ( ~n1569 & n41087 ) | ( n13983 & n41087 ) ;
  assign n41089 = ( n5082 & n9111 ) | ( n5082 & n15232 ) | ( n9111 & n15232 ) ;
  assign n41090 = n41089 ^ n30106 ^ n16181 ;
  assign n41091 = n296 & ~n9279 ;
  assign n41092 = n35544 ^ n7603 ^ 1'b0 ;
  assign n41094 = ( n5151 & n10735 ) | ( n5151 & n17406 ) | ( n10735 & n17406 ) ;
  assign n41093 = ~n21878 & n38836 ;
  assign n41095 = n41094 ^ n41093 ^ 1'b0 ;
  assign n41096 = n14813 & n27769 ;
  assign n41097 = n31707 ^ n31648 ^ n4216 ;
  assign n41104 = n13776 ^ n10730 ^ 1'b0 ;
  assign n41105 = n12067 & ~n41104 ;
  assign n41103 = n16329 ^ n7939 ^ 1'b0 ;
  assign n41099 = ( n7242 & n8206 ) | ( n7242 & ~n12136 ) | ( n8206 & ~n12136 ) ;
  assign n41098 = n3398 & n17520 ;
  assign n41100 = n41099 ^ n41098 ^ 1'b0 ;
  assign n41101 = ( n5186 & n17147 ) | ( n5186 & n41100 ) | ( n17147 & n41100 ) ;
  assign n41102 = n1368 | n41101 ;
  assign n41106 = n41105 ^ n41103 ^ n41102 ;
  assign n41107 = n24169 ^ n14256 ^ n10465 ;
  assign n41108 = n13763 | n38135 ;
  assign n41109 = ( n4352 & ~n28440 ) | ( n4352 & n41108 ) | ( ~n28440 & n41108 ) ;
  assign n41110 = ( n6429 & n9346 ) | ( n6429 & n35060 ) | ( n9346 & n35060 ) ;
  assign n41111 = n26124 ^ n18257 ^ 1'b0 ;
  assign n41112 = x108 & n41111 ;
  assign n41114 = ( n5291 & ~n30335 ) | ( n5291 & n33810 ) | ( ~n30335 & n33810 ) ;
  assign n41113 = n15715 | n17096 ;
  assign n41115 = n41114 ^ n41113 ^ 1'b0 ;
  assign n41116 = n13687 ^ n4616 ^ 1'b0 ;
  assign n41117 = n22017 | n41116 ;
  assign n41118 = n15184 & n36457 ;
  assign n41119 = n41118 ^ n12160 ^ n7673 ;
  assign n41120 = n41117 & n41119 ;
  assign n41121 = ~n478 & n16389 ;
  assign n41122 = n41121 ^ n22526 ^ 1'b0 ;
  assign n41123 = n6924 & ~n41122 ;
  assign n41124 = n41123 ^ n17157 ^ 1'b0 ;
  assign n41125 = ( n19856 & n41120 ) | ( n19856 & n41124 ) | ( n41120 & n41124 ) ;
  assign n41126 = ( x162 & ~n8166 ) | ( x162 & n9254 ) | ( ~n8166 & n9254 ) ;
  assign n41127 = n41126 ^ n36503 ^ n12507 ;
  assign n41128 = n35281 ^ n31790 ^ n2397 ;
  assign n41129 = n346 & n30345 ;
  assign n41130 = n41129 ^ n31800 ^ 1'b0 ;
  assign n41132 = n8267 ^ n5938 ^ n5691 ;
  assign n41131 = n37155 ^ n28854 ^ n15436 ;
  assign n41133 = n41132 ^ n41131 ^ n21687 ;
  assign n41134 = n13324 ^ x219 ^ 1'b0 ;
  assign n41135 = ~n7364 & n41134 ;
  assign n41136 = ~n15144 & n41135 ;
  assign n41137 = n11388 ^ n9773 ^ n6933 ;
  assign n41138 = n41137 ^ n6940 ^ 1'b0 ;
  assign n41139 = ~n41136 & n41138 ;
  assign n41140 = n41139 ^ n39330 ^ n32591 ;
  assign n41141 = ~n1256 & n40763 ;
  assign n41142 = n33467 ^ n29567 ^ n15537 ;
  assign n41143 = n41142 ^ n33339 ^ n28055 ;
  assign n41144 = n29989 ^ n15114 ^ n5487 ;
  assign n41145 = ( n8892 & n22955 ) | ( n8892 & n38968 ) | ( n22955 & n38968 ) ;
  assign n41146 = ( n24546 & n25556 ) | ( n24546 & n41145 ) | ( n25556 & n41145 ) ;
  assign n41147 = ( ~n14996 & n15988 ) | ( ~n14996 & n23748 ) | ( n15988 & n23748 ) ;
  assign n41150 = ~n7994 & n24190 ;
  assign n41151 = n28691 | n41150 ;
  assign n41148 = n308 & n19660 ;
  assign n41149 = n6664 | n41148 ;
  assign n41152 = n41151 ^ n41149 ^ 1'b0 ;
  assign n41153 = n33287 ^ n19005 ^ n12000 ;
  assign n41154 = n41153 ^ n38597 ^ 1'b0 ;
  assign n41155 = ( n10880 & ~n12760 ) | ( n10880 & n20824 ) | ( ~n12760 & n20824 ) ;
  assign n41156 = n41155 ^ n39475 ^ n3166 ;
  assign n41157 = n23162 ^ n14926 ^ n4531 ;
  assign n41158 = n7914 & n22861 ;
  assign n41159 = ( n3592 & n25614 ) | ( n3592 & n41158 ) | ( n25614 & n41158 ) ;
  assign n41160 = n30277 ^ n4444 ^ 1'b0 ;
  assign n41163 = n632 | n13082 ;
  assign n41164 = n41163 ^ n19014 ^ 1'b0 ;
  assign n41165 = n41164 ^ n31869 ^ n12405 ;
  assign n41161 = ( ~n4232 & n9130 ) | ( ~n4232 & n12121 ) | ( n9130 & n12121 ) ;
  assign n41162 = n5304 & ~n41161 ;
  assign n41166 = n41165 ^ n41162 ^ 1'b0 ;
  assign n41167 = n38043 & n41166 ;
  assign n41168 = n41167 ^ n26427 ^ 1'b0 ;
  assign n41169 = ( n3155 & ~n31649 ) | ( n3155 & n41168 ) | ( ~n31649 & n41168 ) ;
  assign n41170 = ~n25788 & n35878 ;
  assign n41171 = ( n6377 & n14818 ) | ( n6377 & ~n41170 ) | ( n14818 & ~n41170 ) ;
  assign n41172 = ( ~n5907 & n8172 ) | ( ~n5907 & n34120 ) | ( n8172 & n34120 ) ;
  assign n41173 = n24196 ^ n7447 ^ 1'b0 ;
  assign n41174 = n6906 & n41173 ;
  assign n41175 = n41174 ^ n21238 ^ n18388 ;
  assign n41176 = n28847 ^ n17749 ^ n8758 ;
  assign n41177 = n41176 ^ n17867 ^ n15119 ;
  assign n41178 = n32706 ^ n21457 ^ 1'b0 ;
  assign n41179 = n4764 ^ x90 ^ 1'b0 ;
  assign n41180 = n18626 ^ n14745 ^ n1668 ;
  assign n41181 = ( n16290 & n17075 ) | ( n16290 & n41180 ) | ( n17075 & n41180 ) ;
  assign n41182 = ( n4795 & ~n41179 ) | ( n4795 & n41181 ) | ( ~n41179 & n41181 ) ;
  assign n41183 = ( n16114 & n17424 ) | ( n16114 & n41182 ) | ( n17424 & n41182 ) ;
  assign n41184 = ~n15912 & n29423 ;
  assign n41185 = n17267 & n41184 ;
  assign n41186 = n15376 | n17006 ;
  assign n41187 = n41186 ^ n1599 ^ 1'b0 ;
  assign n41188 = n959 & ~n1625 ;
  assign n41189 = n41188 ^ n2091 ^ 1'b0 ;
  assign n41190 = n22325 ^ n16527 ^ n3439 ;
  assign n41191 = n39060 ^ n1121 ^ n1079 ;
  assign n41192 = n18347 ^ n2801 ^ 1'b0 ;
  assign n41193 = n20189 ^ n15856 ^ 1'b0 ;
  assign n41194 = n20894 ^ n12335 ^ 1'b0 ;
  assign n41195 = ~n3991 & n41194 ;
  assign n41196 = ( n13964 & ~n15481 ) | ( n13964 & n41195 ) | ( ~n15481 & n41195 ) ;
  assign n41197 = n39867 ^ n27043 ^ n1141 ;
  assign n41198 = ( ~n16608 & n17787 ) | ( ~n16608 & n29140 ) | ( n17787 & n29140 ) ;
  assign n41199 = n4698 & ~n41198 ;
  assign n41200 = n7747 ^ n3488 ^ n2711 ;
  assign n41201 = n9243 & ~n41200 ;
  assign n41202 = n7928 | n41201 ;
  assign n41203 = n41199 & ~n41202 ;
  assign n41204 = ( n7486 & n31039 ) | ( n7486 & ~n41203 ) | ( n31039 & ~n41203 ) ;
  assign n41205 = n22640 ^ n16148 ^ 1'b0 ;
  assign n41206 = ~n7666 & n14051 ;
  assign n41207 = ~n6207 & n33267 ;
  assign n41208 = n24781 ^ n20931 ^ n15110 ;
  assign n41209 = ( ~x109 & n19957 ) | ( ~x109 & n24198 ) | ( n19957 & n24198 ) ;
  assign n41210 = n41208 | n41209 ;
  assign n41211 = ~n9739 & n22979 ;
  assign n41212 = n5773 & ~n19835 ;
  assign n41213 = ( ~n405 & n16338 ) | ( ~n405 & n41212 ) | ( n16338 & n41212 ) ;
  assign n41214 = n41213 ^ n21055 ^ n606 ;
  assign n41215 = n17107 & n36560 ;
  assign n41216 = ( ~n2674 & n19920 ) | ( ~n2674 & n26134 ) | ( n19920 & n26134 ) ;
  assign n41217 = n9098 & ~n34258 ;
  assign n41218 = ~n41216 & n41217 ;
  assign n41219 = n4135 & ~n17752 ;
  assign n41220 = n41219 ^ n12105 ^ 1'b0 ;
  assign n41221 = n31315 ^ n5465 ^ 1'b0 ;
  assign n41222 = ~n14627 & n41221 ;
  assign n41223 = n41220 & n41222 ;
  assign n41224 = n3751 ^ n400 ^ 1'b0 ;
  assign n41225 = ( n9426 & n19483 ) | ( n9426 & n19695 ) | ( n19483 & n19695 ) ;
  assign n41226 = n11480 | n41225 ;
  assign n41227 = n41224 | n41226 ;
  assign n41231 = n23151 | n27229 ;
  assign n41232 = n41231 ^ n7723 ^ 1'b0 ;
  assign n41228 = n11811 & n23539 ;
  assign n41229 = n38794 & n41228 ;
  assign n41230 = ( n30630 & ~n31485 ) | ( n30630 & n41229 ) | ( ~n31485 & n41229 ) ;
  assign n41233 = n41232 ^ n41230 ^ n5385 ;
  assign n41234 = n16942 ^ n15397 ^ n7537 ;
  assign n41235 = n35582 ^ n14699 ^ n5766 ;
  assign n41236 = n41235 ^ n16263 ^ 1'b0 ;
  assign n41237 = n11453 ^ n4910 ^ 1'b0 ;
  assign n41238 = ~n6525 & n13111 ;
  assign n41239 = n41238 ^ n23931 ^ 1'b0 ;
  assign n41240 = n41239 ^ n30577 ^ n14127 ;
  assign n41241 = n2417 & n30938 ;
  assign n41242 = n13768 & n25139 ;
  assign n41243 = ( n1338 & n20411 ) | ( n1338 & n39600 ) | ( n20411 & n39600 ) ;
  assign n41244 = n1023 & n7747 ;
  assign n41245 = ( n10280 & n31925 ) | ( n10280 & ~n41244 ) | ( n31925 & ~n41244 ) ;
  assign n41246 = n41245 ^ n2960 ^ 1'b0 ;
  assign n41247 = n41243 & n41246 ;
  assign n41248 = n4789 & ~n22455 ;
  assign n41249 = n41248 ^ n4303 ^ 1'b0 ;
  assign n41250 = n20875 ^ n10434 ^ 1'b0 ;
  assign n41251 = n13438 ^ n1799 ^ n1012 ;
  assign n41252 = ( n15290 & n32937 ) | ( n15290 & ~n37566 ) | ( n32937 & ~n37566 ) ;
  assign n41253 = n40924 ^ n17123 ^ 1'b0 ;
  assign n41254 = ( x201 & n38702 ) | ( x201 & ~n41253 ) | ( n38702 & ~n41253 ) ;
  assign n41255 = n20945 ^ n3445 ^ x112 ;
  assign n41256 = n20824 ^ n5162 ^ 1'b0 ;
  assign n41257 = ~n30975 & n41256 ;
  assign n41258 = n25506 ^ n5367 ^ n903 ;
  assign n41259 = ( ~n20858 & n26786 ) | ( ~n20858 & n41258 ) | ( n26786 & n41258 ) ;
  assign n41262 = ( n14957 & ~n18602 ) | ( n14957 & n24613 ) | ( ~n18602 & n24613 ) ;
  assign n41260 = ( n4147 & n17349 ) | ( n4147 & n32187 ) | ( n17349 & n32187 ) ;
  assign n41261 = n41260 ^ n39504 ^ n25475 ;
  assign n41263 = n41262 ^ n41261 ^ n16027 ;
  assign n41264 = n9482 ^ n6555 ^ n1436 ;
  assign n41265 = ( n4238 & n20071 ) | ( n4238 & ~n35497 ) | ( n20071 & ~n35497 ) ;
  assign n41266 = ( n35150 & n39353 ) | ( n35150 & n41265 ) | ( n39353 & n41265 ) ;
  assign n41267 = n32317 & n41266 ;
  assign n41268 = n38080 ^ n13897 ^ n447 ;
  assign n41269 = n3082 | n24443 ;
  assign n41270 = n4774 | n41269 ;
  assign n41271 = n41270 ^ n21217 ^ n16600 ;
  assign n41272 = n1231 & ~n29071 ;
  assign n41274 = n4485 ^ n4189 ^ n2403 ;
  assign n41275 = n6495 ^ n5671 ^ 1'b0 ;
  assign n41276 = ~n41274 & n41275 ;
  assign n41273 = n2733 & n40592 ;
  assign n41277 = n41276 ^ n41273 ^ 1'b0 ;
  assign n41280 = n22228 ^ n10433 ^ 1'b0 ;
  assign n41281 = n35313 & n41280 ;
  assign n41282 = n27080 & n41281 ;
  assign n41278 = n5576 | n33393 ;
  assign n41279 = n41278 ^ n7316 ^ 1'b0 ;
  assign n41283 = n41282 ^ n41279 ^ 1'b0 ;
  assign n41284 = n35555 & n41283 ;
  assign n41285 = n41284 ^ n6411 ^ 1'b0 ;
  assign n41287 = n31566 ^ n20581 ^ 1'b0 ;
  assign n41288 = n41287 ^ n17232 ^ 1'b0 ;
  assign n41286 = n32530 ^ n27505 ^ n7159 ;
  assign n41289 = n41288 ^ n41286 ^ n10917 ;
  assign n41293 = n3479 | n16156 ;
  assign n41294 = n6395 & ~n41293 ;
  assign n41290 = n17071 | n18237 ;
  assign n41291 = n41290 ^ n20207 ^ 1'b0 ;
  assign n41292 = n41291 ^ n13118 ^ 1'b0 ;
  assign n41295 = n41294 ^ n41292 ^ n36890 ;
  assign n41296 = n40079 ^ n34093 ^ 1'b0 ;
  assign n41297 = n6717 ^ n2433 ^ 1'b0 ;
  assign n41298 = n41297 ^ n1713 ^ 1'b0 ;
  assign n41299 = ( n8153 & ~n29132 ) | ( n8153 & n41298 ) | ( ~n29132 & n41298 ) ;
  assign n41300 = ~n11035 & n20126 ;
  assign n41301 = ~n13914 & n41300 ;
  assign n41302 = n991 & ~n41301 ;
  assign n41303 = n41302 ^ n16036 ^ 1'b0 ;
  assign n41304 = n29990 ^ n7227 ^ 1'b0 ;
  assign n41305 = n25837 & ~n41304 ;
  assign n41306 = ~n37140 & n41305 ;
  assign n41307 = n22142 ^ n13932 ^ 1'b0 ;
  assign n41308 = ( n5259 & n22128 ) | ( n5259 & n30383 ) | ( n22128 & n30383 ) ;
  assign n41309 = n41308 ^ n22745 ^ n22202 ;
  assign n41310 = n25963 ^ n25368 ^ n7107 ;
  assign n41311 = n14740 | n41310 ;
  assign n41312 = n5613 ^ n3977 ^ n2631 ;
  assign n41313 = ( n903 & ~n9344 ) | ( n903 & n41312 ) | ( ~n9344 & n41312 ) ;
  assign n41314 = n41313 ^ n38274 ^ n9769 ;
  assign n41315 = n41314 ^ n13366 ^ n6926 ;
  assign n41316 = n13839 ^ n9030 ^ n4906 ;
  assign n41318 = n10943 ^ n2566 ^ 1'b0 ;
  assign n41317 = n29087 & n29422 ;
  assign n41319 = n41318 ^ n41317 ^ 1'b0 ;
  assign n41320 = ~n1956 & n41319 ;
  assign n41322 = n26531 ^ n8513 ^ 1'b0 ;
  assign n41323 = n3508 & ~n41322 ;
  assign n41324 = ( n11513 & ~n34054 ) | ( n11513 & n41323 ) | ( ~n34054 & n41323 ) ;
  assign n41321 = n21757 ^ n12235 ^ 1'b0 ;
  assign n41325 = n41324 ^ n41321 ^ n7387 ;
  assign n41326 = n26340 & ~n41325 ;
  assign n41327 = n41320 & n41326 ;
  assign n41328 = n30317 ^ n10893 ^ 1'b0 ;
  assign n41329 = n4130 & ~n41328 ;
  assign n41330 = n34279 | n36318 ;
  assign n41331 = n41330 ^ n37521 ^ n10767 ;
  assign n41332 = ( n3800 & n6639 ) | ( n3800 & ~n13285 ) | ( n6639 & ~n13285 ) ;
  assign n41333 = n585 & n17427 ;
  assign n41335 = n19394 ^ n14292 ^ 1'b0 ;
  assign n41334 = n18270 ^ n6572 ^ n3759 ;
  assign n41336 = n41335 ^ n41334 ^ n30297 ;
  assign n41337 = n30570 ^ n3812 ^ 1'b0 ;
  assign n41338 = n41337 ^ n26457 ^ n3609 ;
  assign n41339 = n41338 ^ n26531 ^ 1'b0 ;
  assign n41340 = n11457 & ~n41339 ;
  assign n41341 = ~n10032 & n41340 ;
  assign n41342 = n20094 ^ n7125 ^ n6242 ;
  assign n41343 = n41342 ^ n28972 ^ n1413 ;
  assign n41344 = n41343 ^ n28614 ^ n5833 ;
  assign n41345 = ( n7483 & ~n22423 ) | ( n7483 & n41344 ) | ( ~n22423 & n41344 ) ;
  assign n41346 = ~n3492 & n41345 ;
  assign n41347 = n6466 & n41346 ;
  assign n41348 = ( ~n11572 & n19614 ) | ( ~n11572 & n26999 ) | ( n19614 & n26999 ) ;
  assign n41349 = n19099 ^ n8409 ^ 1'b0 ;
  assign n41350 = ( n14194 & n40088 ) | ( n14194 & ~n41349 ) | ( n40088 & ~n41349 ) ;
  assign n41351 = ( n28379 & n36840 ) | ( n28379 & ~n38239 ) | ( n36840 & ~n38239 ) ;
  assign n41352 = n41351 ^ n16060 ^ 1'b0 ;
  assign n41353 = n41350 & ~n41352 ;
  assign n41354 = ~n41348 & n41353 ;
  assign n41355 = ~n29676 & n41354 ;
  assign n41356 = n39745 ^ n20104 ^ n17462 ;
  assign n41357 = n16432 | n41356 ;
  assign n41358 = n34236 ^ n24025 ^ n8429 ;
  assign n41359 = ( n22323 & n31002 ) | ( n22323 & n41358 ) | ( n31002 & n41358 ) ;
  assign n41360 = n41359 ^ n32573 ^ n19412 ;
  assign n41361 = n24497 ^ n4779 ^ 1'b0 ;
  assign n41362 = ( ~n18322 & n27343 ) | ( ~n18322 & n31222 ) | ( n27343 & n31222 ) ;
  assign n41363 = ( n9514 & n16752 ) | ( n9514 & n23718 ) | ( n16752 & n23718 ) ;
  assign n41364 = n41363 ^ n19626 ^ n17900 ;
  assign n41365 = n21817 ^ n4709 ^ 1'b0 ;
  assign n41366 = ~n41364 & n41365 ;
  assign n41367 = n41366 ^ n29288 ^ n3906 ;
  assign n41368 = ( n24859 & ~n25405 ) | ( n24859 & n41367 ) | ( ~n25405 & n41367 ) ;
  assign n41369 = n10599 | n16175 ;
  assign n41370 = n41369 ^ n34507 ^ 1'b0 ;
  assign n41371 = n17182 & ~n41370 ;
  assign n41372 = n503 & ~n9097 ;
  assign n41373 = n38945 & n41372 ;
  assign n41374 = ~n14602 & n33478 ;
  assign n41375 = ~n2923 & n41374 ;
  assign n41376 = n35512 ^ n18906 ^ n15851 ;
  assign n41377 = ( ~n3629 & n18210 ) | ( ~n3629 & n22448 ) | ( n18210 & n22448 ) ;
  assign n41378 = ~n3249 & n18702 ;
  assign n41379 = n41378 ^ n8652 ^ x66 ;
  assign n41380 = n39495 ^ n26203 ^ n25150 ;
  assign n41381 = n6302 & n34000 ;
  assign n41382 = n41381 ^ n9707 ^ 1'b0 ;
  assign n41383 = n30584 ^ n9092 ^ n3313 ;
  assign n41384 = ( n9330 & ~n13339 ) | ( n9330 & n17732 ) | ( ~n13339 & n17732 ) ;
  assign n41385 = ( x55 & ~n271 ) | ( x55 & n17312 ) | ( ~n271 & n17312 ) ;
  assign n41386 = n41385 ^ n24224 ^ n16416 ;
  assign n41387 = n19478 & n20613 ;
  assign n41388 = n16936 & ~n25453 ;
  assign n41389 = n24253 ^ n1020 ^ 1'b0 ;
  assign n41390 = ( n25329 & ~n29927 ) | ( n25329 & n41389 ) | ( ~n29927 & n41389 ) ;
  assign n41391 = n29333 & ~n41390 ;
  assign n41392 = n23969 ^ n17816 ^ 1'b0 ;
  assign n41393 = n19662 ^ n6585 ^ n3767 ;
  assign n41394 = n29681 ^ n20752 ^ n2334 ;
  assign n41395 = n41394 ^ n33038 ^ n18116 ;
  assign n41396 = n41395 ^ n26896 ^ n10314 ;
  assign n41397 = ( ~n2627 & n35775 ) | ( ~n2627 & n41396 ) | ( n35775 & n41396 ) ;
  assign n41398 = ( n2540 & n2603 ) | ( n2540 & ~n41397 ) | ( n2603 & ~n41397 ) ;
  assign n41400 = n14596 ^ n7490 ^ n4960 ;
  assign n41399 = ~n19241 & n37080 ;
  assign n41401 = n41400 ^ n41399 ^ 1'b0 ;
  assign n41402 = ( n25855 & ~n35963 ) | ( n25855 & n41401 ) | ( ~n35963 & n41401 ) ;
  assign n41403 = n41402 ^ n23734 ^ 1'b0 ;
  assign n41404 = n41403 ^ n21966 ^ 1'b0 ;
  assign n41405 = n40759 ^ n9492 ^ 1'b0 ;
  assign n41406 = n41405 ^ n16596 ^ n6515 ;
  assign n41407 = n7568 & n41406 ;
  assign n41408 = ~n32639 & n41407 ;
  assign n41409 = n41408 ^ n26404 ^ n22622 ;
  assign n41410 = n10702 ^ n9736 ^ n997 ;
  assign n41411 = n27264 & ~n28592 ;
  assign n41412 = n21624 & ~n24320 ;
  assign n41413 = n41412 ^ n1039 ^ 1'b0 ;
  assign n41414 = ~n34826 & n41413 ;
  assign n41415 = n31099 ^ n28050 ^ n1734 ;
  assign n41416 = n35334 ^ n2251 ^ n1406 ;
  assign n41417 = n32692 ^ n16818 ^ 1'b0 ;
  assign n41422 = ~n11968 & n27714 ;
  assign n41420 = n34471 ^ n13936 ^ n4482 ;
  assign n41418 = n4431 & n40548 ;
  assign n41419 = ( n7732 & ~n28377 ) | ( n7732 & n41418 ) | ( ~n28377 & n41418 ) ;
  assign n41421 = n41420 ^ n41419 ^ n37039 ;
  assign n41423 = n41422 ^ n41421 ^ n28139 ;
  assign n41426 = ( n13858 & n33118 ) | ( n13858 & n35646 ) | ( n33118 & n35646 ) ;
  assign n41424 = n11153 ^ n10196 ^ n5440 ;
  assign n41425 = n12339 & ~n41424 ;
  assign n41427 = n41426 ^ n41425 ^ n7375 ;
  assign n41428 = ~n10130 & n41427 ;
  assign n41429 = n37138 & n41428 ;
  assign n41430 = ( ~n10022 & n14002 ) | ( ~n10022 & n23631 ) | ( n14002 & n23631 ) ;
  assign n41431 = n41430 ^ n32834 ^ n4657 ;
  assign n41432 = n41431 ^ n16314 ^ n3059 ;
  assign n41433 = n7247 & n34509 ;
  assign n41435 = ( ~n3528 & n6359 ) | ( ~n3528 & n12901 ) | ( n6359 & n12901 ) ;
  assign n41434 = n11144 ^ n6352 ^ n1386 ;
  assign n41436 = n41435 ^ n41434 ^ n13264 ;
  assign n41437 = ( ~n3916 & n11184 ) | ( ~n3916 & n29262 ) | ( n11184 & n29262 ) ;
  assign n41438 = n25594 & ~n41437 ;
  assign n41439 = ( n19827 & n41436 ) | ( n19827 & ~n41438 ) | ( n41436 & ~n41438 ) ;
  assign n41440 = ( ~n7105 & n11063 ) | ( ~n7105 & n41439 ) | ( n11063 & n41439 ) ;
  assign n41441 = n7100 ^ n2816 ^ x56 ;
  assign n41442 = n41441 ^ n37579 ^ 1'b0 ;
  assign n41443 = n12374 ^ n12114 ^ n3949 ;
  assign n41444 = ( x126 & n4664 ) | ( x126 & n9762 ) | ( n4664 & n9762 ) ;
  assign n41445 = ~n41312 & n41444 ;
  assign n41446 = ~n24699 & n41445 ;
  assign n41447 = ~n15931 & n39377 ;
  assign n41448 = n41447 ^ n7326 ^ 1'b0 ;
  assign n41449 = n41448 ^ n20570 ^ 1'b0 ;
  assign n41450 = n41446 | n41449 ;
  assign n41451 = n26764 & ~n29433 ;
  assign n41452 = n24412 ^ n21810 ^ n16284 ;
  assign n41453 = n22012 ^ n19766 ^ n2863 ;
  assign n41454 = n41453 ^ n18477 ^ n10986 ;
  assign n41455 = ( n28453 & ~n36988 ) | ( n28453 & n41454 ) | ( ~n36988 & n41454 ) ;
  assign n41456 = n41455 ^ n20396 ^ 1'b0 ;
  assign n41457 = n41452 & ~n41456 ;
  assign n41460 = n6172 ^ n1909 ^ 1'b0 ;
  assign n41458 = n29842 ^ n8517 ^ n7286 ;
  assign n41459 = n41458 ^ n40698 ^ n27918 ;
  assign n41461 = n41460 ^ n41459 ^ n34877 ;
  assign n41462 = ( n406 & ~n1836 ) | ( n406 & n9123 ) | ( ~n1836 & n9123 ) ;
  assign n41463 = ( n6414 & n40214 ) | ( n6414 & n41462 ) | ( n40214 & n41462 ) ;
  assign n41466 = n22863 & ~n24266 ;
  assign n41467 = ~n41056 & n41466 ;
  assign n41468 = n41467 ^ n31724 ^ n12681 ;
  assign n41464 = n26441 ^ n23957 ^ n11545 ;
  assign n41465 = ( ~n18233 & n35204 ) | ( ~n18233 & n41464 ) | ( n35204 & n41464 ) ;
  assign n41469 = n41468 ^ n41465 ^ 1'b0 ;
  assign n41470 = n37556 ^ n4024 ^ n452 ;
  assign n41471 = n20335 | n41470 ;
  assign n41472 = n41471 ^ n19677 ^ 1'b0 ;
  assign n41473 = ( n422 & n8475 ) | ( n422 & ~n15199 ) | ( n8475 & ~n15199 ) ;
  assign n41474 = n930 & n20553 ;
  assign n41475 = ( ~n1598 & n3811 ) | ( ~n1598 & n37570 ) | ( n3811 & n37570 ) ;
  assign n41476 = ( n5201 & n41474 ) | ( n5201 & n41475 ) | ( n41474 & n41475 ) ;
  assign n41477 = n41476 ^ n1329 ^ 1'b0 ;
  assign n41478 = n41473 & n41477 ;
  assign n41479 = ~n9755 & n28194 ;
  assign n41483 = ( n10545 & ~n14413 ) | ( n10545 & n16522 ) | ( ~n14413 & n16522 ) ;
  assign n41484 = n22453 ^ n10144 ^ 1'b0 ;
  assign n41485 = n41483 | n41484 ;
  assign n41481 = n13940 ^ n6377 ^ 1'b0 ;
  assign n41480 = ( n15673 & n18889 ) | ( n15673 & n22056 ) | ( n18889 & n22056 ) ;
  assign n41482 = n41481 ^ n41480 ^ 1'b0 ;
  assign n41486 = n41485 ^ n41482 ^ n14020 ;
  assign n41487 = n8062 ^ n267 ^ 1'b0 ;
  assign n41488 = n34072 ^ n14861 ^ n3868 ;
  assign n41489 = ~n38907 & n41488 ;
  assign n41490 = n12844 ^ n7085 ^ n815 ;
  assign n41491 = ~n3258 & n28830 ;
  assign n41492 = ( ~n4161 & n28722 ) | ( ~n4161 & n32660 ) | ( n28722 & n32660 ) ;
  assign n41493 = ( n8891 & n12068 ) | ( n8891 & ~n20747 ) | ( n12068 & ~n20747 ) ;
  assign n41494 = n4697 | n41493 ;
  assign n41495 = n41494 ^ n8456 ^ n6505 ;
  assign n41496 = n5888 | n25226 ;
  assign n41497 = n41495 | n41496 ;
  assign n41498 = ( ~n12951 & n34341 ) | ( ~n12951 & n34648 ) | ( n34341 & n34648 ) ;
  assign n41499 = ( n28226 & ~n37747 ) | ( n28226 & n41498 ) | ( ~n37747 & n41498 ) ;
  assign n41500 = n21232 & n31076 ;
  assign n41501 = n19021 & n41500 ;
  assign n41502 = n8681 & ~n41501 ;
  assign n41503 = n36793 ^ n18922 ^ n587 ;
  assign n41504 = n16788 ^ n10692 ^ n2726 ;
  assign n41505 = ( n395 & n35824 ) | ( n395 & n41504 ) | ( n35824 & n41504 ) ;
  assign n41506 = n26096 ^ n25594 ^ n852 ;
  assign n41507 = n41506 ^ n21443 ^ n2736 ;
  assign n41508 = n41507 ^ n13545 ^ n13125 ;
  assign n41511 = n8885 & ~n15203 ;
  assign n41509 = ( n2646 & n20822 ) | ( n2646 & n28075 ) | ( n20822 & n28075 ) ;
  assign n41510 = ( n4109 & n7478 ) | ( n4109 & ~n41509 ) | ( n7478 & ~n41509 ) ;
  assign n41512 = n41511 ^ n41510 ^ n6111 ;
  assign n41515 = n38042 ^ n416 ^ 1'b0 ;
  assign n41516 = ( n13666 & ~n33112 ) | ( n13666 & n41515 ) | ( ~n33112 & n41515 ) ;
  assign n41513 = n13053 ^ n2176 ^ 1'b0 ;
  assign n41514 = ~n12336 & n41513 ;
  assign n41517 = n41516 ^ n41514 ^ n6898 ;
  assign n41518 = ~n35520 & n38317 ;
  assign n41519 = n41518 ^ n15928 ^ 1'b0 ;
  assign n41520 = n21801 ^ n10996 ^ n10870 ;
  assign n41521 = ( n14284 & n21110 ) | ( n14284 & n41520 ) | ( n21110 & n41520 ) ;
  assign n41522 = ~n2187 & n5233 ;
  assign n41523 = ~n41521 & n41522 ;
  assign n41524 = n40178 ^ n7525 ^ n3294 ;
  assign n41525 = n41524 ^ n13771 ^ n542 ;
  assign n41526 = n14523 | n15912 ;
  assign n41527 = n2645 & ~n41526 ;
  assign n41528 = ~n41525 & n41527 ;
  assign n41529 = n29964 ^ n5086 ^ 1'b0 ;
  assign n41530 = ~n1009 & n20875 ;
  assign n41531 = ~n1944 & n41530 ;
  assign n41532 = ( n7385 & ~n14477 ) | ( n7385 & n41531 ) | ( ~n14477 & n41531 ) ;
  assign n41533 = ( n21729 & ~n41529 ) | ( n21729 & n41532 ) | ( ~n41529 & n41532 ) ;
  assign n41535 = n30686 ^ n14339 ^ 1'b0 ;
  assign n41534 = n15563 & ~n36828 ;
  assign n41536 = n41535 ^ n41534 ^ 1'b0 ;
  assign n41537 = n33848 ^ n27289 ^ n22548 ;
  assign n41538 = ~n41536 & n41537 ;
  assign n41540 = n32948 ^ n17770 ^ 1'b0 ;
  assign n41541 = n41137 & ~n41540 ;
  assign n41542 = ( ~n5130 & n20817 ) | ( ~n5130 & n41541 ) | ( n20817 & n41541 ) ;
  assign n41539 = n1756 & n35518 ;
  assign n41543 = n41542 ^ n41539 ^ 1'b0 ;
  assign n41544 = ~n13075 & n22727 ;
  assign n41545 = n28667 ^ n17841 ^ n10495 ;
  assign n41546 = ( n15983 & n38580 ) | ( n15983 & n41545 ) | ( n38580 & n41545 ) ;
  assign n41547 = n20389 ^ n2501 ^ n1433 ;
  assign n41548 = n33109 ^ n20040 ^ n2161 ;
  assign n41549 = n41548 ^ n25147 ^ n10319 ;
  assign n41550 = n41549 ^ n34066 ^ 1'b0 ;
  assign n41554 = n17373 ^ n12558 ^ 1'b0 ;
  assign n41555 = x16 & ~n41554 ;
  assign n41552 = ~n5913 & n27096 ;
  assign n41553 = n22736 | n41552 ;
  assign n41556 = n41555 ^ n41553 ^ 1'b0 ;
  assign n41551 = n14436 & n24550 ;
  assign n41557 = n41556 ^ n41551 ^ n4048 ;
  assign n41558 = n5990 ^ n3866 ^ 1'b0 ;
  assign n41559 = n12697 & ~n41558 ;
  assign n41560 = n3372 & ~n20681 ;
  assign n41561 = n41560 ^ n36134 ^ 1'b0 ;
  assign n41562 = ( n764 & ~n2397 ) | ( n764 & n12889 ) | ( ~n2397 & n12889 ) ;
  assign n41563 = n13351 ^ n8236 ^ n7125 ;
  assign n41564 = ( n17861 & n41562 ) | ( n17861 & n41563 ) | ( n41562 & n41563 ) ;
  assign n41565 = n41564 ^ n13106 ^ n10899 ;
  assign n41566 = ~n8140 & n36503 ;
  assign n41567 = ( n7000 & n9018 ) | ( n7000 & ~n25451 ) | ( n9018 & ~n25451 ) ;
  assign n41568 = ~n1350 & n6356 ;
  assign n41569 = ( n20454 & n37575 ) | ( n20454 & ~n41568 ) | ( n37575 & ~n41568 ) ;
  assign n41570 = n22195 & ~n38517 ;
  assign n41571 = n41570 ^ n30254 ^ 1'b0 ;
  assign n41572 = n3673 | n32462 ;
  assign n41573 = n39619 & ~n41572 ;
  assign n41574 = n26191 ^ n1875 ^ x35 ;
  assign n41575 = n41574 ^ n33133 ^ n24535 ;
  assign n41576 = ( n587 & n26572 ) | ( n587 & ~n41575 ) | ( n26572 & ~n41575 ) ;
  assign n41577 = ( n2486 & n26242 ) | ( n2486 & n32009 ) | ( n26242 & n32009 ) ;
  assign n41578 = n41577 ^ n29060 ^ 1'b0 ;
  assign n41579 = n41576 & n41578 ;
  assign n41580 = n35021 ^ n7904 ^ 1'b0 ;
  assign n41581 = n9344 & ~n41580 ;
  assign n41582 = n38906 ^ n8277 ^ n4478 ;
  assign n41583 = n11266 ^ n9836 ^ 1'b0 ;
  assign n41584 = ( n30710 & n33268 ) | ( n30710 & n41583 ) | ( n33268 & n41583 ) ;
  assign n41585 = n2581 & ~n23466 ;
  assign n41586 = n2105 & n41585 ;
  assign n41587 = ( n8069 & n8209 ) | ( n8069 & ~n41586 ) | ( n8209 & ~n41586 ) ;
  assign n41588 = n26941 ^ n17757 ^ n10351 ;
  assign n41589 = n41587 & ~n41588 ;
  assign n41590 = n9996 & n21032 ;
  assign n41591 = n41590 ^ n27637 ^ 1'b0 ;
  assign n41592 = n12703 ^ x248 ^ 1'b0 ;
  assign n41593 = n10780 & ~n41592 ;
  assign n41594 = ( n25078 & ~n41591 ) | ( n25078 & n41593 ) | ( ~n41591 & n41593 ) ;
  assign n41595 = ~n7091 & n23370 ;
  assign n41596 = ( ~n4046 & n5542 ) | ( ~n4046 & n9449 ) | ( n5542 & n9449 ) ;
  assign n41597 = n38664 ^ n573 ^ 1'b0 ;
  assign n41598 = n41596 & n41597 ;
  assign n41599 = ( ~n25822 & n41595 ) | ( ~n25822 & n41598 ) | ( n41595 & n41598 ) ;
  assign n41600 = n41599 ^ n18751 ^ n10690 ;
  assign n41601 = ( n9611 & n11857 ) | ( n9611 & ~n36181 ) | ( n11857 & ~n36181 ) ;
  assign n41602 = ( ~n795 & n1906 ) | ( ~n795 & n41601 ) | ( n1906 & n41601 ) ;
  assign n41603 = n12624 & ~n40032 ;
  assign n41604 = n41603 ^ n14172 ^ 1'b0 ;
  assign n41605 = ( n4358 & n24511 ) | ( n4358 & n26985 ) | ( n24511 & n26985 ) ;
  assign n41606 = n41605 ^ n23203 ^ 1'b0 ;
  assign n41607 = n2806 | n41606 ;
  assign n41608 = n24123 ^ n4601 ^ n4239 ;
  assign n41609 = n16076 | n41608 ;
  assign n41610 = n26032 | n41609 ;
  assign n41611 = n1031 & ~n6841 ;
  assign n41612 = n41611 ^ n3242 ^ 1'b0 ;
  assign n41613 = n41612 ^ n11743 ^ 1'b0 ;
  assign n41614 = n3864 & ~n41613 ;
  assign n41615 = ( n10786 & n15256 ) | ( n10786 & n41614 ) | ( n15256 & n41614 ) ;
  assign n41616 = ( n23490 & ~n32389 ) | ( n23490 & n41615 ) | ( ~n32389 & n41615 ) ;
  assign n41617 = n2605 ^ n2502 ^ 1'b0 ;
  assign n41618 = n4237 & ~n8625 ;
  assign n41619 = n41618 ^ n7753 ^ 1'b0 ;
  assign n41620 = n41619 ^ n21167 ^ n19957 ;
  assign n41621 = n28615 ^ n4181 ^ 1'b0 ;
  assign n41622 = n4525 & ~n41621 ;
  assign n41623 = n41622 ^ n30908 ^ 1'b0 ;
  assign n41624 = n41623 ^ n30605 ^ 1'b0 ;
  assign n41625 = n13460 | n41624 ;
  assign n41626 = ~n12688 & n16634 ;
  assign n41627 = n41626 ^ n7756 ^ 1'b0 ;
  assign n41628 = ~n37879 & n41627 ;
  assign n41629 = n36878 ^ n14256 ^ n7743 ;
  assign n41630 = n23081 ^ n17805 ^ 1'b0 ;
  assign n41631 = n38204 | n41630 ;
  assign n41632 = ( n12930 & n15099 ) | ( n12930 & ~n27714 ) | ( n15099 & ~n27714 ) ;
  assign n41633 = ( n34569 & n41631 ) | ( n34569 & n41632 ) | ( n41631 & n41632 ) ;
  assign n41634 = n41633 ^ n29801 ^ n22397 ;
  assign n41635 = n37839 ^ n37038 ^ n12430 ;
  assign n41636 = n41635 ^ n24787 ^ n5479 ;
  assign n41637 = n12521 ^ n4102 ^ n2373 ;
  assign n41638 = n39961 ^ n24705 ^ n14725 ;
  assign n41639 = n39322 ^ n31948 ^ n3303 ;
  assign n41640 = ( ~n10176 & n41638 ) | ( ~n10176 & n41639 ) | ( n41638 & n41639 ) ;
  assign n41641 = n32045 ^ n14492 ^ 1'b0 ;
  assign n41642 = ~n26218 & n41641 ;
  assign n41643 = n2241 | n25019 ;
  assign n41644 = n20221 & ~n41643 ;
  assign n41645 = n9755 ^ n6836 ^ n4442 ;
  assign n41646 = ( n4441 & n8705 ) | ( n4441 & ~n20663 ) | ( n8705 & ~n20663 ) ;
  assign n41647 = n41646 ^ n10654 ^ 1'b0 ;
  assign n41648 = ~n41645 & n41647 ;
  assign n41649 = ( n11871 & n13194 ) | ( n11871 & ~n41648 ) | ( n13194 & ~n41648 ) ;
  assign n41650 = ~n10592 & n11072 ;
  assign n41651 = n41649 & n41650 ;
  assign n41652 = n14647 ^ n4985 ^ 1'b0 ;
  assign n41653 = ( n5129 & n10086 ) | ( n5129 & n41652 ) | ( n10086 & n41652 ) ;
  assign n41654 = n41653 ^ n38304 ^ n26388 ;
  assign n41655 = n22372 ^ n3573 ^ 1'b0 ;
  assign n41656 = n34864 ^ n10363 ^ 1'b0 ;
  assign n41657 = ( ~n27221 & n32469 ) | ( ~n27221 & n41656 ) | ( n32469 & n41656 ) ;
  assign n41658 = ~n8804 & n19363 ;
  assign n41659 = ( n3088 & ~n4894 ) | ( n3088 & n23518 ) | ( ~n4894 & n23518 ) ;
  assign n41660 = n41659 ^ n16448 ^ 1'b0 ;
  assign n41661 = n8679 | n36828 ;
  assign n41662 = n9999 | n41661 ;
  assign n41663 = ( n14899 & n41660 ) | ( n14899 & ~n41662 ) | ( n41660 & ~n41662 ) ;
  assign n41664 = ( n10426 & n24950 ) | ( n10426 & n41663 ) | ( n24950 & n41663 ) ;
  assign n41665 = n19706 ^ n3278 ^ 1'b0 ;
  assign n41666 = n7054 | n41665 ;
  assign n41667 = n19839 | n28198 ;
  assign n41668 = n41667 ^ n4496 ^ 1'b0 ;
  assign n41669 = n39923 ^ n22413 ^ n4950 ;
  assign n41670 = ( ~n11019 & n13750 ) | ( ~n11019 & n27618 ) | ( n13750 & n27618 ) ;
  assign n41671 = n41670 ^ n31260 ^ n21787 ;
  assign n41672 = n14606 ^ n11144 ^ n10415 ;
  assign n41673 = n41672 ^ n27974 ^ n9217 ;
  assign n41674 = ( x28 & ~n20899 ) | ( x28 & n41673 ) | ( ~n20899 & n41673 ) ;
  assign n41675 = n22046 ^ n18839 ^ n12341 ;
  assign n41676 = ~n11244 & n11271 ;
  assign n41677 = n41676 ^ n34787 ^ 1'b0 ;
  assign n41678 = n33765 ^ n17067 ^ n7283 ;
  assign n41679 = ( ~n41675 & n41677 ) | ( ~n41675 & n41678 ) | ( n41677 & n41678 ) ;
  assign n41680 = n12121 ^ n5804 ^ n2334 ;
  assign n41681 = n10017 | n19891 ;
  assign n41682 = n41681 ^ n12388 ^ 1'b0 ;
  assign n41683 = n28857 ^ n2995 ^ 1'b0 ;
  assign n41684 = n41682 | n41683 ;
  assign n41685 = n461 & n29418 ;
  assign n41686 = n16118 ^ n6908 ^ 1'b0 ;
  assign n41687 = ~n1258 & n41686 ;
  assign n41688 = x69 & n32948 ;
  assign n41689 = ( ~n5726 & n13179 ) | ( ~n5726 & n25095 ) | ( n13179 & n25095 ) ;
  assign n41690 = n36725 ^ n32047 ^ 1'b0 ;
  assign n41691 = n5556 ^ n2516 ^ n1655 ;
  assign n41692 = n7121 & ~n13131 ;
  assign n41693 = n41692 ^ n10270 ^ 1'b0 ;
  assign n41694 = ( n4212 & n6771 ) | ( n4212 & n24054 ) | ( n6771 & n24054 ) ;
  assign n41695 = ( ~n817 & n13371 ) | ( ~n817 & n13950 ) | ( n13371 & n13950 ) ;
  assign n41696 = n41695 ^ n20481 ^ 1'b0 ;
  assign n41697 = n41694 | n41696 ;
  assign n41698 = ( ~n17386 & n41693 ) | ( ~n17386 & n41697 ) | ( n41693 & n41697 ) ;
  assign n41699 = ( ~n7149 & n16764 ) | ( ~n7149 & n20851 ) | ( n16764 & n20851 ) ;
  assign n41700 = ( n5991 & ~n7845 ) | ( n5991 & n41699 ) | ( ~n7845 & n41699 ) ;
  assign n41701 = n41700 ^ n33804 ^ n18798 ;
  assign n41702 = n20970 & ~n41701 ;
  assign n41703 = ~n7957 & n36734 ;
  assign n41704 = n36928 ^ n11694 ^ n8163 ;
  assign n41707 = n25752 ^ n5109 ^ n355 ;
  assign n41705 = n26138 ^ n14744 ^ 1'b0 ;
  assign n41706 = n41705 ^ n37595 ^ n17251 ;
  assign n41708 = n41707 ^ n41706 ^ n27734 ;
  assign n41709 = n41708 ^ n18665 ^ n7688 ;
  assign n41710 = n32865 ^ n13162 ^ 1'b0 ;
  assign n41711 = n7566 & n24573 ;
  assign n41712 = n41465 ^ n19431 ^ n9525 ;
  assign n41713 = n18352 ^ n693 ^ 1'b0 ;
  assign n41714 = n1927 | n41713 ;
  assign n41715 = ~n19858 & n23613 ;
  assign n41720 = n34136 ^ n18595 ^ 1'b0 ;
  assign n41716 = n4803 & n20943 ;
  assign n41717 = ( n8014 & n13096 ) | ( n8014 & ~n41716 ) | ( n13096 & ~n41716 ) ;
  assign n41718 = n14346 ^ n8470 ^ n4987 ;
  assign n41719 = ( n11860 & ~n41717 ) | ( n11860 & n41718 ) | ( ~n41717 & n41718 ) ;
  assign n41721 = n41720 ^ n41719 ^ n34454 ;
  assign n41722 = n15073 | n24470 ;
  assign n41723 = n9277 | n41722 ;
  assign n41724 = ( n1034 & n5219 ) | ( n1034 & n41723 ) | ( n5219 & n41723 ) ;
  assign n41725 = n35071 ^ n34003 ^ n21495 ;
  assign n41728 = n8814 ^ n3207 ^ n1806 ;
  assign n41726 = n21436 ^ n15273 ^ 1'b0 ;
  assign n41727 = n27595 | n41726 ;
  assign n41729 = n41728 ^ n41727 ^ n25114 ;
  assign n41730 = ( n9999 & ~n17357 ) | ( n9999 & n41729 ) | ( ~n17357 & n41729 ) ;
  assign n41731 = n39873 ^ n38200 ^ n13808 ;
  assign n41732 = ( n8223 & n32612 ) | ( n8223 & n36038 ) | ( n32612 & n36038 ) ;
  assign n41733 = n2347 & ~n11680 ;
  assign n41734 = n18786 ^ n9922 ^ n5983 ;
  assign n41735 = ( n5994 & n39099 ) | ( n5994 & ~n41734 ) | ( n39099 & ~n41734 ) ;
  assign n41736 = ( n9142 & n41733 ) | ( n9142 & n41735 ) | ( n41733 & n41735 ) ;
  assign n41737 = n41736 ^ n21787 ^ n19321 ;
  assign n41738 = ( n8841 & n15785 ) | ( n8841 & ~n41737 ) | ( n15785 & ~n41737 ) ;
  assign n41739 = n41738 ^ n35330 ^ 1'b0 ;
  assign n41740 = ( n942 & n18397 ) | ( n942 & ~n38826 ) | ( n18397 & ~n38826 ) ;
  assign n41741 = n41740 ^ n22398 ^ 1'b0 ;
  assign n41742 = n10106 & n41741 ;
  assign n41743 = n10848 | n28808 ;
  assign n41746 = n32044 ^ n22097 ^ n1090 ;
  assign n41744 = n34929 ^ n15699 ^ n10132 ;
  assign n41745 = n41744 ^ n37080 ^ n4132 ;
  assign n41747 = n41746 ^ n41745 ^ n27999 ;
  assign n41751 = n7956 ^ n405 ^ 1'b0 ;
  assign n41752 = ( n4263 & n12387 ) | ( n4263 & n41751 ) | ( n12387 & n41751 ) ;
  assign n41753 = ( n11601 & n17183 ) | ( n11601 & n41752 ) | ( n17183 & n41752 ) ;
  assign n41750 = ( n14094 & n20658 ) | ( n14094 & ~n27269 ) | ( n20658 & ~n27269 ) ;
  assign n41748 = n13599 | n25466 ;
  assign n41749 = n41748 ^ n31438 ^ 1'b0 ;
  assign n41754 = n41753 ^ n41750 ^ n41749 ;
  assign n41755 = n27186 ^ n928 ^ n858 ;
  assign n41756 = n9603 ^ n5594 ^ n4054 ;
  assign n41757 = n41756 ^ n29989 ^ n14674 ;
  assign n41758 = ( ~n8323 & n41755 ) | ( ~n8323 & n41757 ) | ( n41755 & n41757 ) ;
  assign n41759 = ( ~n13226 & n13257 ) | ( ~n13226 & n41758 ) | ( n13257 & n41758 ) ;
  assign n41760 = n36236 ^ n28265 ^ n1246 ;
  assign n41761 = ( n3399 & n4168 ) | ( n3399 & n41760 ) | ( n4168 & n41760 ) ;
  assign n41763 = n1600 | n19394 ;
  assign n41764 = n41763 ^ n38722 ^ n11790 ;
  assign n41762 = ( n3108 & n22629 ) | ( n3108 & ~n35657 ) | ( n22629 & ~n35657 ) ;
  assign n41765 = n41764 ^ n41762 ^ n33545 ;
  assign n41766 = ~n2597 & n18228 ;
  assign n41767 = ~n7074 & n41766 ;
  assign n41768 = ~n3944 & n6508 ;
  assign n41769 = ( n7781 & ~n41767 ) | ( n7781 & n41768 ) | ( ~n41767 & n41768 ) ;
  assign n41770 = ~n14563 & n27006 ;
  assign n41771 = n41770 ^ n2913 ^ 1'b0 ;
  assign n41772 = n3006 & n30967 ;
  assign n41773 = n41771 & n41772 ;
  assign n41774 = n15606 ^ n9670 ^ 1'b0 ;
  assign n41775 = n13920 | n41774 ;
  assign n41776 = n34259 ^ n26337 ^ 1'b0 ;
  assign n41777 = ( ~x221 & n18397 ) | ( ~x221 & n41776 ) | ( n18397 & n41776 ) ;
  assign n41778 = ( n20058 & n28135 ) | ( n20058 & n31549 ) | ( n28135 & n31549 ) ;
  assign n41779 = n17756 ^ n4590 ^ 1'b0 ;
  assign n41780 = n41778 & ~n41779 ;
  assign n41781 = n26942 ^ n12789 ^ 1'b0 ;
  assign n41782 = ( n2003 & n41780 ) | ( n2003 & ~n41781 ) | ( n41780 & ~n41781 ) ;
  assign n41783 = ~n4177 & n15756 ;
  assign n41784 = n28861 ^ n2926 ^ 1'b0 ;
  assign n41785 = ( n16557 & n20552 ) | ( n16557 & n26349 ) | ( n20552 & n26349 ) ;
  assign n41787 = n19412 ^ n15448 ^ n1538 ;
  assign n41786 = x67 | n3526 ;
  assign n41788 = n41787 ^ n41786 ^ 1'b0 ;
  assign n41789 = ( n6707 & n41785 ) | ( n6707 & n41788 ) | ( n41785 & n41788 ) ;
  assign n41790 = n8150 ^ n7522 ^ 1'b0 ;
  assign n41791 = n23772 & ~n41790 ;
  assign n41793 = ( n4935 & n7365 ) | ( n4935 & n21452 ) | ( n7365 & n21452 ) ;
  assign n41794 = ( ~n15813 & n22244 ) | ( ~n15813 & n41793 ) | ( n22244 & n41793 ) ;
  assign n41792 = n28597 & n31529 ;
  assign n41795 = n41794 ^ n41792 ^ 1'b0 ;
  assign n41797 = ( n306 & n3449 ) | ( n306 & ~n38715 ) | ( n3449 & ~n38715 ) ;
  assign n41796 = n19924 | n30400 ;
  assign n41798 = n41797 ^ n41796 ^ 1'b0 ;
  assign n41799 = n10814 & ~n21906 ;
  assign n41800 = ~n15288 & n41799 ;
  assign n41801 = ( ~n19869 & n41480 ) | ( ~n19869 & n41800 ) | ( n41480 & n41800 ) ;
  assign n41802 = ( n1151 & ~n35441 ) | ( n1151 & n36115 ) | ( ~n35441 & n36115 ) ;
  assign n41803 = ~n3929 & n10216 ;
  assign n41804 = n41803 ^ n33216 ^ 1'b0 ;
  assign n41805 = ( ~n17022 & n22209 ) | ( ~n17022 & n41804 ) | ( n22209 & n41804 ) ;
  assign n41806 = ~n17705 & n30193 ;
  assign n41807 = n41806 ^ n2572 ^ 1'b0 ;
  assign n41808 = n8654 ^ n2186 ^ 1'b0 ;
  assign n41809 = n15574 ^ n3881 ^ n3747 ;
  assign n41810 = ~n9552 & n41809 ;
  assign n41811 = ( ~n28571 & n40023 ) | ( ~n28571 & n41810 ) | ( n40023 & n41810 ) ;
  assign n41812 = n36546 ^ n13268 ^ 1'b0 ;
  assign n41813 = n21884 ^ n21485 ^ n15502 ;
  assign n41814 = ~n2271 & n34009 ;
  assign n41815 = ~n41813 & n41814 ;
  assign n41816 = n40569 ^ n399 ^ 1'b0 ;
  assign n41817 = n32219 ^ n19889 ^ 1'b0 ;
  assign n41818 = ( n14208 & ~n22173 ) | ( n14208 & n35521 ) | ( ~n22173 & n35521 ) ;
  assign n41819 = n1476 & n21326 ;
  assign n41820 = n41819 ^ n710 ^ 1'b0 ;
  assign n41823 = n18801 ^ n16770 ^ n10031 ;
  assign n41824 = n41823 ^ n16418 ^ n5667 ;
  assign n41825 = n41824 ^ n24770 ^ 1'b0 ;
  assign n41826 = n7642 ^ n1651 ^ 1'b0 ;
  assign n41827 = n41825 | n41826 ;
  assign n41821 = n14303 ^ n13923 ^ n13140 ;
  assign n41822 = n15297 & ~n41821 ;
  assign n41828 = n41827 ^ n41822 ^ 1'b0 ;
  assign n41829 = n18845 & ~n19248 ;
  assign n41830 = ~n22245 & n41829 ;
  assign n41831 = ( n5897 & ~n24060 ) | ( n5897 & n30142 ) | ( ~n24060 & n30142 ) ;
  assign n41832 = ( ~n4665 & n7736 ) | ( ~n4665 & n9944 ) | ( n7736 & n9944 ) ;
  assign n41833 = n41832 ^ n32446 ^ n7782 ;
  assign n41835 = ( n419 & n6223 ) | ( n419 & n17907 ) | ( n6223 & n17907 ) ;
  assign n41834 = n7878 | n19058 ;
  assign n41836 = n41835 ^ n41834 ^ 1'b0 ;
  assign n41837 = n41836 ^ n41243 ^ n22557 ;
  assign n41838 = ( n10209 & n35556 ) | ( n10209 & ~n41837 ) | ( n35556 & ~n41837 ) ;
  assign n41839 = n13042 & ~n13629 ;
  assign n41840 = ( n10245 & n20306 ) | ( n10245 & ~n22336 ) | ( n20306 & ~n22336 ) ;
  assign n41841 = ( ~n1395 & n19712 ) | ( ~n1395 & n22579 ) | ( n19712 & n22579 ) ;
  assign n41842 = n34634 ^ n7749 ^ n7037 ;
  assign n41843 = n41842 ^ n30630 ^ n2667 ;
  assign n41844 = ~n3083 & n17446 ;
  assign n41845 = ~n36849 & n41844 ;
  assign n41846 = n31028 & n41845 ;
  assign n41847 = n41846 ^ n1357 ^ 1'b0 ;
  assign n41848 = n24179 & ~n41847 ;
  assign n41849 = ( n797 & n18539 ) | ( n797 & n25542 ) | ( n18539 & n25542 ) ;
  assign n41850 = n8892 & ~n11262 ;
  assign n41851 = n41850 ^ n6058 ^ 1'b0 ;
  assign n41852 = n18718 | n33108 ;
  assign n41853 = n14693 & ~n41852 ;
  assign n41854 = n41853 ^ n933 ^ 1'b0 ;
  assign n41855 = n38935 ^ n20916 ^ n4306 ;
  assign n41858 = x211 & n1129 ;
  assign n41859 = n25665 & n41858 ;
  assign n41856 = ( ~n912 & n1612 ) | ( ~n912 & n7043 ) | ( n1612 & n7043 ) ;
  assign n41857 = ~n18971 & n41856 ;
  assign n41860 = n41859 ^ n41857 ^ n16762 ;
  assign n41861 = ( ~n9168 & n18850 ) | ( ~n9168 & n27703 ) | ( n18850 & n27703 ) ;
  assign n41865 = n31748 ^ n29092 ^ n15139 ;
  assign n41866 = ~n28161 & n41865 ;
  assign n41867 = n41866 ^ n15090 ^ 1'b0 ;
  assign n41862 = n16438 & n25673 ;
  assign n41863 = n41862 ^ n5085 ^ 1'b0 ;
  assign n41864 = ~n3735 & n41863 ;
  assign n41868 = n41867 ^ n41864 ^ 1'b0 ;
  assign n41869 = ( ~n37590 & n41861 ) | ( ~n37590 & n41868 ) | ( n41861 & n41868 ) ;
  assign n41872 = n20244 ^ n15919 ^ n6071 ;
  assign n41871 = n11176 | n17687 ;
  assign n41873 = n41872 ^ n41871 ^ 1'b0 ;
  assign n41870 = ~n15718 & n21969 ;
  assign n41874 = n41873 ^ n41870 ^ 1'b0 ;
  assign n41875 = n12134 ^ n8541 ^ 1'b0 ;
  assign n41876 = n10488 & n41875 ;
  assign n41877 = n3595 & n41876 ;
  assign n41878 = n41877 ^ n14035 ^ 1'b0 ;
  assign n41879 = n18760 ^ n17540 ^ n15657 ;
  assign n41880 = n25485 & n41879 ;
  assign n41881 = n41878 & n41880 ;
  assign n41885 = ( n19723 & n26767 ) | ( n19723 & ~n29537 ) | ( n26767 & ~n29537 ) ;
  assign n41882 = ~n15278 & n27037 ;
  assign n41883 = ~n22376 & n41882 ;
  assign n41884 = n930 | n41883 ;
  assign n41886 = n41885 ^ n41884 ^ 1'b0 ;
  assign n41887 = ( n5233 & n9707 ) | ( n5233 & ~n18163 ) | ( n9707 & ~n18163 ) ;
  assign n41888 = n16423 & ~n37315 ;
  assign n41889 = n41888 ^ n39584 ^ 1'b0 ;
  assign n41890 = ( n27931 & n41887 ) | ( n27931 & n41889 ) | ( n41887 & n41889 ) ;
  assign n41891 = n37259 ^ x27 ^ 1'b0 ;
  assign n41892 = ( n3130 & n30494 ) | ( n3130 & ~n41891 ) | ( n30494 & ~n41891 ) ;
  assign n41893 = ( n36334 & n41890 ) | ( n36334 & ~n41892 ) | ( n41890 & ~n41892 ) ;
  assign n41894 = n33957 ^ n13000 ^ n5402 ;
  assign n41895 = n6327 & n17821 ;
  assign n41896 = n41895 ^ n21768 ^ 1'b0 ;
  assign n41897 = ( n8585 & ~n21316 ) | ( n8585 & n41879 ) | ( ~n21316 & n41879 ) ;
  assign n41898 = ( n15023 & n41896 ) | ( n15023 & n41897 ) | ( n41896 & n41897 ) ;
  assign n41899 = n34291 ^ n19244 ^ n17502 ;
  assign n41900 = n20710 ^ n18866 ^ 1'b0 ;
  assign n41901 = ( n4359 & n20934 ) | ( n4359 & n24756 ) | ( n20934 & n24756 ) ;
  assign n41902 = n41901 ^ n12638 ^ 1'b0 ;
  assign n41903 = ~n41900 & n41902 ;
  assign n41907 = n36519 ^ n25837 ^ n20076 ;
  assign n41904 = n23027 ^ n12089 ^ 1'b0 ;
  assign n41905 = ~n5253 & n41904 ;
  assign n41906 = n17982 & n41905 ;
  assign n41908 = n41907 ^ n41906 ^ 1'b0 ;
  assign n41909 = n31271 | n34631 ;
  assign n41910 = n39516 ^ n11404 ^ n8085 ;
  assign n41913 = n40654 ^ n16711 ^ n12810 ;
  assign n41911 = n4136 | n6750 ;
  assign n41912 = n41911 ^ n34451 ^ n10775 ;
  assign n41914 = n41913 ^ n41912 ^ n36621 ;
  assign n41915 = n30884 ^ n15493 ^ n9727 ;
  assign n41916 = n21801 ^ n5240 ^ 1'b0 ;
  assign n41917 = ( n4366 & n9178 ) | ( n4366 & n41340 ) | ( n9178 & n41340 ) ;
  assign n41918 = n41917 ^ n39100 ^ n4297 ;
  assign n41919 = n1991 | n12291 ;
  assign n41920 = ( ~n418 & n3636 ) | ( ~n418 & n3772 ) | ( n3636 & n3772 ) ;
  assign n41921 = n12837 & ~n41920 ;
  assign n41922 = ~n7231 & n41921 ;
  assign n41923 = n6599 ^ n5144 ^ 1'b0 ;
  assign n41924 = n13634 | n41923 ;
  assign n41925 = ~n19427 & n28908 ;
  assign n41926 = n41924 & n41925 ;
  assign n41927 = ~n9583 & n21305 ;
  assign n41928 = n41927 ^ n26883 ^ 1'b0 ;
  assign n41929 = n1327 & ~n41928 ;
  assign n41930 = n36807 ^ n22453 ^ 1'b0 ;
  assign n41931 = ~n10651 & n41930 ;
  assign n41932 = n41931 ^ n38094 ^ n10212 ;
  assign n41933 = n32874 ^ n16489 ^ 1'b0 ;
  assign n41934 = n37691 ^ n8119 ^ n5587 ;
  assign n41935 = ( n416 & n15585 ) | ( n416 & ~n24687 ) | ( n15585 & ~n24687 ) ;
  assign n41936 = ( n14131 & ~n41934 ) | ( n14131 & n41935 ) | ( ~n41934 & n41935 ) ;
  assign n41937 = n4576 & n23069 ;
  assign n41938 = n32748 & n41937 ;
  assign n41939 = ( n26255 & n28486 ) | ( n26255 & n41938 ) | ( n28486 & n41938 ) ;
  assign n41940 = n29329 ^ n19150 ^ 1'b0 ;
  assign n41941 = n19258 | n41940 ;
  assign n41942 = n15091 & n41941 ;
  assign n41943 = n41942 ^ n27044 ^ 1'b0 ;
  assign n41944 = n25218 ^ n19983 ^ n8190 ;
  assign n41945 = n2278 & ~n41944 ;
  assign n41946 = ( n6333 & n11421 ) | ( n6333 & ~n41945 ) | ( n11421 & ~n41945 ) ;
  assign n41947 = ( n5758 & n16638 ) | ( n5758 & n32790 ) | ( n16638 & n32790 ) ;
  assign n41948 = n41947 ^ n25801 ^ n12013 ;
  assign n41949 = ( n18702 & n22942 ) | ( n18702 & n40081 ) | ( n22942 & n40081 ) ;
  assign n41950 = n41949 ^ n27458 ^ n25810 ;
  assign n41951 = n16300 & ~n34061 ;
  assign n41952 = ~n15729 & n41951 ;
  assign n41953 = n41952 ^ n17213 ^ n1312 ;
  assign n41954 = n39548 ^ n25244 ^ n4277 ;
  assign n41955 = ( ~n6971 & n22249 ) | ( ~n6971 & n41954 ) | ( n22249 & n41954 ) ;
  assign n41956 = n41718 ^ n35592 ^ 1'b0 ;
  assign n41957 = n5871 & n41956 ;
  assign n41958 = n24236 & n31864 ;
  assign n41959 = n26441 & ~n35154 ;
  assign n41960 = n39530 ^ n35563 ^ x157 ;
  assign n41961 = n14992 ^ n6626 ^ n5780 ;
  assign n41962 = ( n10573 & ~n21902 ) | ( n10573 & n40485 ) | ( ~n21902 & n40485 ) ;
  assign n41963 = n24680 ^ n11199 ^ 1'b0 ;
  assign n41964 = n41963 ^ x202 ^ 1'b0 ;
  assign n41966 = n37140 ^ n5763 ^ n1725 ;
  assign n41965 = ~n28633 & n37789 ;
  assign n41967 = n41966 ^ n41965 ^ 1'b0 ;
  assign n41969 = ( n473 & n4181 ) | ( n473 & ~n20856 ) | ( n4181 & ~n20856 ) ;
  assign n41968 = ( n3110 & n16200 ) | ( n3110 & ~n21802 ) | ( n16200 & ~n21802 ) ;
  assign n41970 = n41969 ^ n41968 ^ 1'b0 ;
  assign n41971 = n920 & ~n13394 ;
  assign n41972 = n41971 ^ n14038 ^ n6974 ;
  assign n41973 = n26803 ^ n16846 ^ n6967 ;
  assign n41974 = n9553 ^ n4026 ^ 1'b0 ;
  assign n41975 = n6611 & n41974 ;
  assign n41976 = ( n299 & ~n20932 ) | ( n299 & n41975 ) | ( ~n20932 & n41975 ) ;
  assign n41977 = n18708 ^ n9998 ^ n4336 ;
  assign n41978 = n26020 | n41977 ;
  assign n41979 = n24513 ^ n7060 ^ 1'b0 ;
  assign n41980 = n38681 ^ n13683 ^ 1'b0 ;
  assign n41981 = ~n22705 & n41980 ;
  assign n41982 = n22879 ^ n6069 ^ n2878 ;
  assign n41983 = ( n41979 & n41981 ) | ( n41979 & n41982 ) | ( n41981 & n41982 ) ;
  assign n41984 = ( n8714 & n41978 ) | ( n8714 & n41983 ) | ( n41978 & n41983 ) ;
  assign n41985 = n29773 ^ n11577 ^ 1'b0 ;
  assign n41986 = n2341 & ~n41985 ;
  assign n41987 = n6211 & ~n19426 ;
  assign n41988 = n3523 & ~n41987 ;
  assign n41989 = n41986 & n41988 ;
  assign n41997 = ( n2353 & n8445 ) | ( n2353 & ~n10783 ) | ( n8445 & ~n10783 ) ;
  assign n41998 = n41997 ^ n9221 ^ 1'b0 ;
  assign n41999 = n4566 & ~n41998 ;
  assign n41990 = ~n14054 & n16036 ;
  assign n41991 = ~n2041 & n41990 ;
  assign n41992 = n20910 | n41991 ;
  assign n41993 = n41992 ^ n23493 ^ 1'b0 ;
  assign n41994 = n20758 ^ n20481 ^ n16978 ;
  assign n41995 = n41994 ^ n6610 ^ 1'b0 ;
  assign n41996 = n41993 | n41995 ;
  assign n42000 = n41999 ^ n41996 ^ n19067 ;
  assign n42001 = ( ~n13787 & n19353 ) | ( ~n13787 & n37727 ) | ( n19353 & n37727 ) ;
  assign n42002 = ( n2218 & n34818 ) | ( n2218 & ~n42001 ) | ( n34818 & ~n42001 ) ;
  assign n42003 = n33253 ^ n16457 ^ n1738 ;
  assign n42004 = ( n5464 & n10781 ) | ( n5464 & ~n16373 ) | ( n10781 & ~n16373 ) ;
  assign n42005 = n42004 ^ n16371 ^ n5731 ;
  assign n42006 = n28801 ^ n19378 ^ 1'b0 ;
  assign n42007 = n26925 | n42006 ;
  assign n42008 = ~n19938 & n23861 ;
  assign n42009 = ( n39656 & n42007 ) | ( n39656 & ~n42008 ) | ( n42007 & ~n42008 ) ;
  assign n42010 = n27079 & n30563 ;
  assign n42011 = n5693 | n42010 ;
  assign n42012 = n30696 | n42011 ;
  assign n42013 = n41577 ^ n21125 ^ 1'b0 ;
  assign n42014 = n14255 | n42013 ;
  assign n42015 = n3107 & n9740 ;
  assign n42016 = n42015 ^ n10050 ^ 1'b0 ;
  assign n42026 = n16039 & ~n28042 ;
  assign n42024 = n9771 & ~n10241 ;
  assign n42025 = n42024 ^ n3535 ^ 1'b0 ;
  assign n42017 = n9134 & ~n11688 ;
  assign n42018 = n4011 & n42017 ;
  assign n42019 = n3326 & ~n14215 ;
  assign n42020 = n15868 & n42019 ;
  assign n42021 = n16568 ^ n14016 ^ 1'b0 ;
  assign n42022 = n42020 | n42021 ;
  assign n42023 = ( ~n27030 & n42018 ) | ( ~n27030 & n42022 ) | ( n42018 & n42022 ) ;
  assign n42027 = n42026 ^ n42025 ^ n42023 ;
  assign n42028 = ( ~x115 & n15583 ) | ( ~x115 & n33014 ) | ( n15583 & n33014 ) ;
  assign n42029 = n12346 ^ n2247 ^ n2044 ;
  assign n42030 = n42029 ^ n13724 ^ n4221 ;
  assign n42032 = ( n4388 & n9754 ) | ( n4388 & n13879 ) | ( n9754 & n13879 ) ;
  assign n42033 = ( n861 & ~n36186 ) | ( n861 & n42032 ) | ( ~n36186 & n42032 ) ;
  assign n42034 = ( n26279 & n29408 ) | ( n26279 & ~n42033 ) | ( n29408 & ~n42033 ) ;
  assign n42031 = n36447 ^ n27706 ^ n7586 ;
  assign n42035 = n42034 ^ n42031 ^ n22991 ;
  assign n42036 = n23526 ^ n1599 ^ 1'b0 ;
  assign n42037 = n34175 ^ n31722 ^ 1'b0 ;
  assign n42038 = n42036 & ~n42037 ;
  assign n42039 = n42038 ^ n32651 ^ n7676 ;
  assign n42040 = n42039 ^ n31801 ^ n21742 ;
  assign n42041 = ~n19099 & n36661 ;
  assign n42042 = ~n15074 & n42041 ;
  assign n42043 = n20300 ^ n12930 ^ 1'b0 ;
  assign n42044 = n30431 ^ n3065 ^ n2536 ;
  assign n42045 = n12248 & ~n42044 ;
  assign n42046 = n42043 & n42045 ;
  assign n42047 = n27928 ^ n14804 ^ 1'b0 ;
  assign n42048 = n42046 | n42047 ;
  assign n42049 = n38595 ^ n24452 ^ n17039 ;
  assign n42050 = n39007 ^ n20449 ^ n20398 ;
  assign n42051 = ( n2868 & ~n25813 ) | ( n2868 & n42050 ) | ( ~n25813 & n42050 ) ;
  assign n42052 = n42049 | n42051 ;
  assign n42053 = n42052 ^ n1570 ^ 1'b0 ;
  assign n42054 = ~n13245 & n26918 ;
  assign n42055 = ( n13880 & n15902 ) | ( n13880 & ~n21957 ) | ( n15902 & ~n21957 ) ;
  assign n42056 = n42055 ^ n41928 ^ 1'b0 ;
  assign n42062 = ( ~n3299 & n6459 ) | ( ~n3299 & n26871 ) | ( n6459 & n26871 ) ;
  assign n42057 = n2525 & n6694 ;
  assign n42058 = n42057 ^ n21253 ^ 1'b0 ;
  assign n42059 = n23891 ^ n14308 ^ 1'b0 ;
  assign n42060 = ~n17281 & n42059 ;
  assign n42061 = ( n9447 & n42058 ) | ( n9447 & n42060 ) | ( n42058 & n42060 ) ;
  assign n42063 = n42062 ^ n42061 ^ 1'b0 ;
  assign n42064 = ( n13924 & n28754 ) | ( n13924 & ~n37597 ) | ( n28754 & ~n37597 ) ;
  assign n42065 = n17773 ^ n7492 ^ n3266 ;
  assign n42066 = n26716 ^ n11730 ^ 1'b0 ;
  assign n42067 = ( n2247 & ~n5296 ) | ( n2247 & n12850 ) | ( ~n5296 & n12850 ) ;
  assign n42068 = n42067 ^ n29638 ^ n5323 ;
  assign n42069 = ( n7348 & n19439 ) | ( n7348 & ~n27330 ) | ( n19439 & ~n27330 ) ;
  assign n42070 = ( n558 & ~n42068 ) | ( n558 & n42069 ) | ( ~n42068 & n42069 ) ;
  assign n42071 = ( n11421 & n42066 ) | ( n11421 & ~n42070 ) | ( n42066 & ~n42070 ) ;
  assign n42072 = ( n13689 & n16349 ) | ( n13689 & ~n18773 ) | ( n16349 & ~n18773 ) ;
  assign n42073 = n42072 ^ n34690 ^ n915 ;
  assign n42074 = n12153 ^ n2510 ^ 1'b0 ;
  assign n42075 = n5994 & ~n42074 ;
  assign n42076 = ( n8970 & ~n26622 ) | ( n8970 & n42075 ) | ( ~n26622 & n42075 ) ;
  assign n42078 = n14498 ^ n1851 ^ n1292 ;
  assign n42079 = n23304 & ~n42078 ;
  assign n42080 = ~n8873 & n42079 ;
  assign n42077 = n30975 ^ n19883 ^ n11426 ;
  assign n42081 = n42080 ^ n42077 ^ n21653 ;
  assign n42082 = n30678 ^ n30486 ^ 1'b0 ;
  assign n42083 = n16590 & ~n42082 ;
  assign n42084 = n4406 | n10942 ;
  assign n42085 = ( n1409 & ~n15089 ) | ( n1409 & n42084 ) | ( ~n15089 & n42084 ) ;
  assign n42086 = n42085 ^ n33390 ^ n31836 ;
  assign n42087 = ~n11291 & n36452 ;
  assign n42088 = n29759 ^ n17170 ^ n17166 ;
  assign n42089 = n20800 & n42088 ;
  assign n42090 = n19712 ^ x234 ^ 1'b0 ;
  assign n42091 = n39778 ^ n26377 ^ n11577 ;
  assign n42092 = n42091 ^ n39851 ^ n33033 ;
  assign n42093 = n25332 ^ n1573 ^ 1'b0 ;
  assign n42094 = ~n27520 & n42093 ;
  assign n42095 = ( n31049 & n32973 ) | ( n31049 & n42094 ) | ( n32973 & n42094 ) ;
  assign n42096 = n12944 ^ n9258 ^ n4043 ;
  assign n42097 = ~n31877 & n42096 ;
  assign n42098 = n33738 & n42097 ;
  assign n42099 = n34352 | n42098 ;
  assign n42100 = n5134 & ~n42099 ;
  assign n42101 = ~n28573 & n42100 ;
  assign n42103 = n5526 & ~n20283 ;
  assign n42102 = n24354 ^ n24236 ^ n3092 ;
  assign n42104 = n42103 ^ n42102 ^ n19250 ;
  assign n42105 = ( n18517 & n34782 ) | ( n18517 & n42104 ) | ( n34782 & n42104 ) ;
  assign n42106 = n15976 ^ n9361 ^ n8235 ;
  assign n42107 = ( n6495 & n9866 ) | ( n6495 & n42106 ) | ( n9866 & n42106 ) ;
  assign n42108 = n42107 ^ n32341 ^ n431 ;
  assign n42109 = n40504 ^ n22139 ^ n3733 ;
  assign n42112 = n2133 | n13478 ;
  assign n42110 = n21674 & ~n40492 ;
  assign n42111 = ~n340 & n42110 ;
  assign n42113 = n42112 ^ n42111 ^ n3991 ;
  assign n42114 = n15829 ^ n8422 ^ 1'b0 ;
  assign n42115 = n18992 | n42114 ;
  assign n42116 = n42115 ^ n3773 ^ 1'b0 ;
  assign n42117 = n28109 ^ n19822 ^ n15964 ;
  assign n42118 = n42117 ^ n28246 ^ 1'b0 ;
  assign n42119 = n5766 & n13315 ;
  assign n42120 = n41883 & n42119 ;
  assign n42122 = ( ~n1652 & n3934 ) | ( ~n1652 & n27421 ) | ( n3934 & n27421 ) ;
  assign n42121 = n2306 & n11934 ;
  assign n42123 = n42122 ^ n42121 ^ 1'b0 ;
  assign n42124 = ( n3952 & n13217 ) | ( n3952 & n29348 ) | ( n13217 & n29348 ) ;
  assign n42125 = n42124 ^ n25655 ^ 1'b0 ;
  assign n42126 = ~n22372 & n42125 ;
  assign n42127 = ~n10054 & n10121 ;
  assign n42128 = n42127 ^ n7865 ^ 1'b0 ;
  assign n42129 = n9270 & n42128 ;
  assign n42130 = n42129 ^ n20656 ^ 1'b0 ;
  assign n42131 = ( n6685 & n10347 ) | ( n6685 & n42130 ) | ( n10347 & n42130 ) ;
  assign n42132 = n22974 & ~n42131 ;
  assign n42133 = ( n6723 & n11911 ) | ( n6723 & n42132 ) | ( n11911 & n42132 ) ;
  assign n42134 = n31440 ^ n17802 ^ n11143 ;
  assign n42135 = ( n21710 & n39663 ) | ( n21710 & ~n42134 ) | ( n39663 & ~n42134 ) ;
  assign n42136 = ( n2939 & n15553 ) | ( n2939 & ~n25380 ) | ( n15553 & ~n25380 ) ;
  assign n42137 = ( ~n4909 & n13013 ) | ( ~n4909 & n24854 ) | ( n13013 & n24854 ) ;
  assign n42138 = n42137 ^ n3452 ^ n334 ;
  assign n42139 = ( ~n25008 & n34476 ) | ( ~n25008 & n42138 ) | ( n34476 & n42138 ) ;
  assign n42140 = ( ~n14094 & n42136 ) | ( ~n14094 & n42139 ) | ( n42136 & n42139 ) ;
  assign n42141 = n3307 ^ n1529 ^ 1'b0 ;
  assign n42142 = n1384 & ~n42141 ;
  assign n42143 = n22109 ^ n12066 ^ n1668 ;
  assign n42144 = ( n15155 & n42142 ) | ( n15155 & n42143 ) | ( n42142 & n42143 ) ;
  assign n42145 = ( n2935 & ~n29024 ) | ( n2935 & n40792 ) | ( ~n29024 & n40792 ) ;
  assign n42146 = n42145 ^ n35298 ^ n33064 ;
  assign n42147 = ( n5459 & ~n8397 ) | ( n5459 & n18533 ) | ( ~n8397 & n18533 ) ;
  assign n42148 = ( n26742 & n34657 ) | ( n26742 & n42147 ) | ( n34657 & n42147 ) ;
  assign n42149 = n26175 & ~n35342 ;
  assign n42153 = ( ~n4820 & n6701 ) | ( ~n4820 & n28730 ) | ( n6701 & n28730 ) ;
  assign n42150 = n13839 ^ n4621 ^ n2394 ;
  assign n42151 = n34717 ^ n9722 ^ 1'b0 ;
  assign n42152 = n42150 | n42151 ;
  assign n42154 = n42153 ^ n42152 ^ 1'b0 ;
  assign n42155 = n15850 ^ x252 ^ 1'b0 ;
  assign n42156 = n4092 & ~n42155 ;
  assign n42157 = ~n3956 & n20856 ;
  assign n42158 = n10742 ^ n7901 ^ n4751 ;
  assign n42159 = n42158 ^ n7473 ^ 1'b0 ;
  assign n42160 = n16644 ^ n12648 ^ 1'b0 ;
  assign n42161 = n3137 & ~n42160 ;
  assign n42162 = n28876 ^ n7153 ^ n4347 ;
  assign n42163 = n42162 ^ n17604 ^ 1'b0 ;
  assign n42164 = ( n42159 & n42161 ) | ( n42159 & n42163 ) | ( n42161 & n42163 ) ;
  assign n42165 = ( ~n42156 & n42157 ) | ( ~n42156 & n42164 ) | ( n42157 & n42164 ) ;
  assign n42166 = n29136 ^ n2562 ^ 1'b0 ;
  assign n42167 = n29228 ^ n16869 ^ n1813 ;
  assign n42168 = ~n11983 & n34446 ;
  assign n42169 = ( n24620 & n42167 ) | ( n24620 & ~n42168 ) | ( n42167 & ~n42168 ) ;
  assign n42170 = n41025 ^ n9175 ^ 1'b0 ;
  assign n42171 = n35257 | n42170 ;
  assign n42172 = n26919 ^ n12910 ^ n1386 ;
  assign n42173 = n42172 ^ n25198 ^ n3356 ;
  assign n42174 = n42173 ^ n23885 ^ 1'b0 ;
  assign n42175 = n11055 & ~n42174 ;
  assign n42176 = n39616 ^ n30348 ^ 1'b0 ;
  assign n42177 = n7498 ^ n5260 ^ n4629 ;
  assign n42178 = ~n13573 & n42177 ;
  assign n42179 = ( n17159 & n24126 ) | ( n17159 & ~n38224 ) | ( n24126 & ~n38224 ) ;
  assign n42180 = n8961 | n24076 ;
  assign n42181 = ( n39940 & n42179 ) | ( n39940 & ~n42180 ) | ( n42179 & ~n42180 ) ;
  assign n42182 = n26502 ^ n18135 ^ 1'b0 ;
  assign n42183 = n10550 ^ x31 ^ 1'b0 ;
  assign n42184 = ~n20931 & n42183 ;
  assign n42185 = n18097 & n42184 ;
  assign n42186 = n34417 ^ n20082 ^ n15481 ;
  assign n42187 = n42186 ^ n24254 ^ n16013 ;
  assign n42188 = n25022 ^ n24443 ^ n2241 ;
  assign n42190 = ( n2501 & n4273 ) | ( n2501 & ~n16729 ) | ( n4273 & ~n16729 ) ;
  assign n42189 = ( ~n8779 & n23164 ) | ( ~n8779 & n24508 ) | ( n23164 & n24508 ) ;
  assign n42191 = n42190 ^ n42189 ^ n16532 ;
  assign n42192 = n42188 | n42191 ;
  assign n42193 = n10869 ^ n9146 ^ n2528 ;
  assign n42194 = ~n36938 & n42193 ;
  assign n42195 = n27844 ^ n528 ^ 1'b0 ;
  assign n42196 = n25560 & ~n42195 ;
  assign n42197 = n32264 ^ n17002 ^ n1703 ;
  assign n42198 = n42197 ^ n4262 ^ 1'b0 ;
  assign n42199 = n26734 & ~n42198 ;
  assign n42200 = ( ~n5056 & n7920 ) | ( ~n5056 & n42050 ) | ( n7920 & n42050 ) ;
  assign n42201 = ( ~n23341 & n29878 ) | ( ~n23341 & n38023 ) | ( n29878 & n38023 ) ;
  assign n42202 = ( n8090 & ~n29196 ) | ( n8090 & n37176 ) | ( ~n29196 & n37176 ) ;
  assign n42203 = ( ~x31 & x82 ) | ( ~x31 & n33645 ) | ( x82 & n33645 ) ;
  assign n42204 = n38517 ^ n4524 ^ 1'b0 ;
  assign n42205 = ~n42203 & n42204 ;
  assign n42206 = n32807 ^ n13685 ^ 1'b0 ;
  assign n42207 = n27758 ^ n18797 ^ n15371 ;
  assign n42208 = ( n21223 & ~n25368 ) | ( n21223 & n25778 ) | ( ~n25368 & n25778 ) ;
  assign n42209 = n36196 ^ n26512 ^ 1'b0 ;
  assign n42210 = n32398 ^ n12337 ^ n4196 ;
  assign n42211 = n33210 ^ n4728 ^ n4469 ;
  assign n42212 = ~n8966 & n42211 ;
  assign n42213 = n22376 | n34773 ;
  assign n42214 = n38152 ^ n1227 ^ 1'b0 ;
  assign n42215 = n42213 & ~n42214 ;
  assign n42216 = n37183 ^ n25179 ^ n7094 ;
  assign n42218 = ( n683 & ~n34102 ) | ( n683 & n38739 ) | ( ~n34102 & n38739 ) ;
  assign n42217 = n12446 & ~n23757 ;
  assign n42219 = n42218 ^ n42217 ^ 1'b0 ;
  assign n42220 = n10976 ^ n7060 ^ x130 ;
  assign n42221 = ~n6624 & n42220 ;
  assign n42222 = n42221 ^ n36110 ^ n29721 ;
  assign n42223 = n26187 ^ n18511 ^ n13009 ;
  assign n42224 = n22517 & n42223 ;
  assign n42225 = n34412 ^ n16332 ^ n4645 ;
  assign n42227 = ( n14291 & ~n17294 ) | ( n14291 & n22611 ) | ( ~n17294 & n22611 ) ;
  assign n42226 = n3073 | n26829 ;
  assign n42228 = n42227 ^ n42226 ^ 1'b0 ;
  assign n42229 = ( n5241 & n8321 ) | ( n5241 & n32642 ) | ( n8321 & n32642 ) ;
  assign n42230 = ~n8301 & n24092 ;
  assign n42231 = n42230 ^ n25428 ^ n15215 ;
  assign n42232 = ~n42229 & n42231 ;
  assign n42233 = ( ~n3510 & n30191 ) | ( ~n3510 & n41037 ) | ( n30191 & n41037 ) ;
  assign n42234 = n21533 ^ n18466 ^ n1647 ;
  assign n42236 = n4520 | n14206 ;
  assign n42237 = n42236 ^ n22288 ^ 1'b0 ;
  assign n42238 = n42237 ^ n32649 ^ n5044 ;
  assign n42239 = n42238 ^ n12579 ^ x123 ;
  assign n42240 = ~n18020 & n42239 ;
  assign n42235 = n12077 ^ n8463 ^ n3947 ;
  assign n42241 = n42240 ^ n42235 ^ n9160 ;
  assign n42242 = n42241 ^ n12920 ^ 1'b0 ;
  assign n42244 = n2530 | n25767 ;
  assign n42245 = ( n3327 & n5544 ) | ( n3327 & n35316 ) | ( n5544 & n35316 ) ;
  assign n42246 = ( ~n14478 & n42244 ) | ( ~n14478 & n42245 ) | ( n42244 & n42245 ) ;
  assign n42243 = n37521 ^ n11285 ^ 1'b0 ;
  assign n42247 = n42246 ^ n42243 ^ n31214 ;
  assign n42248 = n42242 | n42247 ;
  assign n42249 = n11384 ^ n8315 ^ n989 ;
  assign n42250 = n13729 ^ n3937 ^ 1'b0 ;
  assign n42251 = ( ~n14162 & n40655 ) | ( ~n14162 & n42250 ) | ( n40655 & n42250 ) ;
  assign n42252 = n32654 ^ n23872 ^ n967 ;
  assign n42253 = ( n42249 & n42251 ) | ( n42249 & n42252 ) | ( n42251 & n42252 ) ;
  assign n42254 = n16933 ^ n12004 ^ n2630 ;
  assign n42255 = ~n1544 & n28368 ;
  assign n42256 = n42255 ^ n34945 ^ 1'b0 ;
  assign n42257 = n4884 & ~n42256 ;
  assign n42258 = ( n12120 & n42254 ) | ( n12120 & ~n42257 ) | ( n42254 & ~n42257 ) ;
  assign n42260 = ( n3059 & n17964 ) | ( n3059 & ~n39987 ) | ( n17964 & ~n39987 ) ;
  assign n42259 = n13190 & ~n19490 ;
  assign n42261 = n42260 ^ n42259 ^ 1'b0 ;
  assign n42262 = n18892 | n31486 ;
  assign n42263 = n42261 & ~n42262 ;
  assign n42264 = ( ~n7133 & n14240 ) | ( ~n7133 & n18670 ) | ( n14240 & n18670 ) ;
  assign n42265 = n42264 ^ n37866 ^ n4606 ;
  assign n42266 = n19762 ^ n361 ^ 1'b0 ;
  assign n42269 = ~n9306 & n11448 ;
  assign n42267 = n15583 | n20221 ;
  assign n42268 = n26704 & ~n42267 ;
  assign n42270 = n42269 ^ n42268 ^ n22667 ;
  assign n42271 = n42270 ^ n15020 ^ n14618 ;
  assign n42272 = n9597 | n30556 ;
  assign n42273 = n10739 | n42272 ;
  assign n42274 = n11164 & ~n32635 ;
  assign n42275 = ( ~n25632 & n42273 ) | ( ~n25632 & n42274 ) | ( n42273 & n42274 ) ;
  assign n42276 = n5794 ^ n3829 ^ n604 ;
  assign n42277 = n42276 ^ n23746 ^ n6925 ;
  assign n42278 = ( n17484 & n40540 ) | ( n17484 & n42277 ) | ( n40540 & n42277 ) ;
  assign n42279 = ~n30322 & n31717 ;
  assign n42280 = n42278 & n42279 ;
  assign n42281 = ( ~n1191 & n3617 ) | ( ~n1191 & n24513 ) | ( n3617 & n24513 ) ;
  assign n42282 = n29736 ^ n28366 ^ n655 ;
  assign n42284 = x166 & n12834 ;
  assign n42285 = n42284 ^ n1945 ^ 1'b0 ;
  assign n42283 = n29808 ^ n23899 ^ n4563 ;
  assign n42286 = n42285 ^ n42283 ^ n12558 ;
  assign n42287 = n42286 ^ n24476 ^ n15212 ;
  assign n42288 = n42287 ^ n14123 ^ n1560 ;
  assign n42289 = n34202 ^ n28886 ^ n12836 ;
  assign n42290 = n42289 ^ n42026 ^ n2747 ;
  assign n42291 = n42290 ^ n35584 ^ n8200 ;
  assign n42292 = n22763 ^ n3951 ^ 1'b0 ;
  assign n42293 = n40700 ^ n4255 ^ n2863 ;
  assign n42294 = n42293 ^ n23628 ^ 1'b0 ;
  assign n42295 = ( ~n10084 & n20389 ) | ( ~n10084 & n42294 ) | ( n20389 & n42294 ) ;
  assign n42296 = n9444 & ~n12147 ;
  assign n42297 = n21949 & n42296 ;
  assign n42298 = n42297 ^ n36357 ^ n28039 ;
  assign n42300 = ~n6312 & n9344 ;
  assign n42301 = n42300 ^ n6232 ^ 1'b0 ;
  assign n42299 = n28137 ^ n8541 ^ 1'b0 ;
  assign n42302 = n42301 ^ n42299 ^ n16481 ;
  assign n42303 = n7949 & ~n18520 ;
  assign n42304 = n42303 ^ x33 ^ 1'b0 ;
  assign n42305 = n20008 | n22408 ;
  assign n42306 = n42304 | n42305 ;
  assign n42307 = n42098 | n42306 ;
  assign n42308 = n41568 ^ n39155 ^ n12683 ;
  assign n42309 = ~n1631 & n21572 ;
  assign n42310 = n42309 ^ n14436 ^ n2886 ;
  assign n42311 = ~n18575 & n33843 ;
  assign n42312 = n16790 ^ n6151 ^ 1'b0 ;
  assign n42313 = n42311 & ~n42312 ;
  assign n42314 = n32907 ^ n16870 ^ 1'b0 ;
  assign n42315 = n18832 ^ n5576 ^ 1'b0 ;
  assign n42316 = ( n6050 & n25548 ) | ( n6050 & n40178 ) | ( n25548 & n40178 ) ;
  assign n42317 = ( n14243 & ~n36525 ) | ( n14243 & n42316 ) | ( ~n36525 & n42316 ) ;
  assign n42318 = n12607 ^ n3597 ^ 1'b0 ;
  assign n42319 = ( n19248 & n36063 ) | ( n19248 & ~n42318 ) | ( n36063 & ~n42318 ) ;
  assign n42327 = n8584 & ~n11527 ;
  assign n42328 = n42327 ^ n508 ^ 1'b0 ;
  assign n42321 = n21186 ^ n6880 ^ n992 ;
  assign n42322 = n11889 ^ n7505 ^ 1'b0 ;
  assign n42323 = n42321 & ~n42322 ;
  assign n42324 = ( n20711 & n37999 ) | ( n20711 & ~n42323 ) | ( n37999 & ~n42323 ) ;
  assign n42325 = n4776 & ~n42324 ;
  assign n42326 = n25210 & n42325 ;
  assign n42329 = n42328 ^ n42326 ^ n18967 ;
  assign n42330 = n42329 ^ n29084 ^ n28380 ;
  assign n42320 = ~n6069 & n24046 ;
  assign n42331 = n42330 ^ n42320 ^ n38593 ;
  assign n42332 = n33714 ^ n24186 ^ n2302 ;
  assign n42333 = n37872 ^ n25080 ^ n9586 ;
  assign n42334 = n25799 ^ n11560 ^ 1'b0 ;
  assign n42335 = n15986 & n42334 ;
  assign n42336 = ~n1329 & n37747 ;
  assign n42337 = ( n2580 & ~n5456 ) | ( n2580 & n41635 ) | ( ~n5456 & n41635 ) ;
  assign n42338 = n42337 ^ n24727 ^ n17693 ;
  assign n42339 = n36867 ^ n21419 ^ n10933 ;
  assign n42340 = n20765 ^ n14050 ^ n3852 ;
  assign n42341 = ~n7101 & n42340 ;
  assign n42344 = ( n17008 & n20271 ) | ( n17008 & n41832 ) | ( n20271 & n41832 ) ;
  assign n42342 = ~n19437 & n30470 ;
  assign n42343 = n42342 ^ n10395 ^ 1'b0 ;
  assign n42345 = n42344 ^ n42343 ^ 1'b0 ;
  assign n42347 = n3278 & n27083 ;
  assign n42346 = ( ~n11871 & n27761 ) | ( ~n11871 & n39462 ) | ( n27761 & n39462 ) ;
  assign n42348 = n42347 ^ n42346 ^ n26012 ;
  assign n42349 = ( n22915 & ~n42345 ) | ( n22915 & n42348 ) | ( ~n42345 & n42348 ) ;
  assign n42350 = n15829 ^ n7780 ^ n6017 ;
  assign n42351 = n42350 ^ n24560 ^ n23233 ;
  assign n42352 = ( n3113 & n22111 ) | ( n3113 & n36425 ) | ( n22111 & n36425 ) ;
  assign n42353 = ( n23289 & n42351 ) | ( n23289 & n42352 ) | ( n42351 & n42352 ) ;
  assign n42354 = n34920 ^ n34189 ^ n27689 ;
  assign n42355 = ( n3799 & n8189 ) | ( n3799 & n17775 ) | ( n8189 & n17775 ) ;
  assign n42356 = n3107 & ~n8578 ;
  assign n42357 = ~n42355 & n42356 ;
  assign n42358 = n4984 | n37543 ;
  assign n42359 = n40064 ^ n39935 ^ n5006 ;
  assign n42360 = ~n5010 & n25267 ;
  assign n42361 = ~n42359 & n42360 ;
  assign n42362 = ~n527 & n24500 ;
  assign n42363 = n4171 & n42362 ;
  assign n42364 = ( n21179 & ~n32392 ) | ( n21179 & n42363 ) | ( ~n32392 & n42363 ) ;
  assign n42365 = n36583 ^ n11505 ^ n11106 ;
  assign n42366 = n42365 ^ n598 ^ 1'b0 ;
  assign n42367 = ~n7272 & n14988 ;
  assign n42368 = ~n8669 & n42367 ;
  assign n42369 = n42368 ^ n20864 ^ n11948 ;
  assign n42370 = ( ~x52 & n6053 ) | ( ~x52 & n8220 ) | ( n6053 & n8220 ) ;
  assign n42371 = n17278 | n42370 ;
  assign n42376 = ( n6286 & n11432 ) | ( n6286 & ~n31553 ) | ( n11432 & ~n31553 ) ;
  assign n42372 = n19785 ^ n7544 ^ n389 ;
  assign n42373 = n42372 ^ n30337 ^ 1'b0 ;
  assign n42374 = ~n23680 & n42373 ;
  assign n42375 = ~n24953 & n42374 ;
  assign n42377 = n42376 ^ n42375 ^ 1'b0 ;
  assign n42378 = n34693 ^ n9896 ^ 1'b0 ;
  assign n42379 = n26174 & ~n42378 ;
  assign n42380 = ~n23439 & n35136 ;
  assign n42381 = n20524 ^ n18484 ^ 1'b0 ;
  assign n42382 = n42381 ^ n25095 ^ n17790 ;
  assign n42383 = ( n39550 & ~n42380 ) | ( n39550 & n42382 ) | ( ~n42380 & n42382 ) ;
  assign n42384 = ( n21742 & ~n42379 ) | ( n21742 & n42383 ) | ( ~n42379 & n42383 ) ;
  assign n42385 = ~n9369 & n17414 ;
  assign n42386 = n30330 | n42385 ;
  assign n42387 = ~n15661 & n20001 ;
  assign n42388 = n42387 ^ n14231 ^ 1'b0 ;
  assign n42389 = n42388 ^ n26771 ^ n14262 ;
  assign n42390 = ( n1871 & n2382 ) | ( n1871 & ~n11037 ) | ( n2382 & ~n11037 ) ;
  assign n42391 = ( n7629 & n23149 ) | ( n7629 & n42390 ) | ( n23149 & n42390 ) ;
  assign n42392 = n38703 ^ n24863 ^ n8701 ;
  assign n42393 = n42227 ^ n41304 ^ 1'b0 ;
  assign n42394 = ( x119 & ~n16608 ) | ( x119 & n28408 ) | ( ~n16608 & n28408 ) ;
  assign n42395 = n42394 ^ n27562 ^ 1'b0 ;
  assign n42396 = ~n32740 & n42395 ;
  assign n42397 = n32019 ^ n8730 ^ n487 ;
  assign n42398 = n42397 ^ n40830 ^ n1141 ;
  assign n42400 = ( n2863 & n12938 ) | ( n2863 & ~n26108 ) | ( n12938 & ~n26108 ) ;
  assign n42399 = n28882 ^ n12395 ^ 1'b0 ;
  assign n42401 = n42400 ^ n42399 ^ n6351 ;
  assign n42402 = n35948 ^ n27269 ^ 1'b0 ;
  assign n42403 = n17098 ^ n1000 ^ 1'b0 ;
  assign n42404 = n42403 ^ n24600 ^ n15825 ;
  assign n42405 = n18362 ^ n9898 ^ n9680 ;
  assign n42406 = n42405 ^ n41944 ^ n28289 ;
  assign n42407 = ( n37137 & n42404 ) | ( n37137 & n42406 ) | ( n42404 & n42406 ) ;
  assign n42408 = ( ~n27129 & n40799 ) | ( ~n27129 & n42407 ) | ( n40799 & n42407 ) ;
  assign n42409 = n26708 ^ n24772 ^ 1'b0 ;
  assign n42410 = n11710 & n42409 ;
  assign n42411 = ( ~n11372 & n27350 ) | ( ~n11372 & n34215 ) | ( n27350 & n34215 ) ;
  assign n42412 = n23500 ^ n20336 ^ n20298 ;
  assign n42413 = n18466 & n39442 ;
  assign n42414 = n30337 ^ n19718 ^ n3450 ;
  assign n42415 = n37995 ^ n37093 ^ n11497 ;
  assign n42416 = n15364 & ~n39493 ;
  assign n42417 = n42416 ^ n22307 ^ 1'b0 ;
  assign n42418 = n42417 ^ n26466 ^ 1'b0 ;
  assign n42419 = n12488 & ~n42418 ;
  assign n42420 = n26449 & n31731 ;
  assign n42421 = n28359 & n42420 ;
  assign n42422 = n32612 ^ n3980 ^ n3722 ;
  assign n42423 = n11750 ^ n8651 ^ 1'b0 ;
  assign n42424 = ( n25032 & n29258 ) | ( n25032 & n42423 ) | ( n29258 & n42423 ) ;
  assign n42425 = ~n8794 & n40178 ;
  assign n42426 = n42425 ^ n2175 ^ 1'b0 ;
  assign n42427 = n42426 ^ n18092 ^ n13748 ;
  assign n42428 = n42427 ^ n19748 ^ n7331 ;
  assign n42429 = n7155 | n17583 ;
  assign n42430 = n42429 ^ n843 ^ 1'b0 ;
  assign n42431 = n42430 ^ n32826 ^ n8517 ;
  assign n42432 = n34976 & ~n42431 ;
  assign n42433 = n13387 & ~n20685 ;
  assign n42434 = n14508 ^ n8096 ^ 1'b0 ;
  assign n42435 = n5261 & n20826 ;
  assign n42436 = n42435 ^ n2741 ^ 1'b0 ;
  assign n42437 = n2979 | n3691 ;
  assign n42438 = ( n19833 & ~n20649 ) | ( n19833 & n42437 ) | ( ~n20649 & n42437 ) ;
  assign n42439 = ( ~x214 & n8839 ) | ( ~x214 & n42438 ) | ( n8839 & n42438 ) ;
  assign n42440 = n42439 ^ n3601 ^ n747 ;
  assign n42441 = n1498 & n42440 ;
  assign n42442 = n16193 & n42441 ;
  assign n42443 = n5743 ^ n5020 ^ n4768 ;
  assign n42444 = n11824 & ~n17560 ;
  assign n42445 = ( n29109 & n42443 ) | ( n29109 & n42444 ) | ( n42443 & n42444 ) ;
  assign n42450 = ( n8825 & n11553 ) | ( n8825 & n16911 ) | ( n11553 & n16911 ) ;
  assign n42451 = n1209 ^ n1033 ^ x134 ;
  assign n42452 = n42451 ^ n16237 ^ 1'b0 ;
  assign n42453 = n42450 | n42452 ;
  assign n42454 = n42453 ^ n1805 ^ x218 ;
  assign n42447 = n17490 ^ n17047 ^ 1'b0 ;
  assign n42448 = n14731 & n42447 ;
  assign n42446 = n18423 ^ n11348 ^ n1764 ;
  assign n42449 = n42448 ^ n42446 ^ n20358 ;
  assign n42455 = n42454 ^ n42449 ^ n19358 ;
  assign n42456 = n22219 ^ n20336 ^ n9943 ;
  assign n42457 = ( n21661 & n28450 ) | ( n21661 & ~n38437 ) | ( n28450 & ~n38437 ) ;
  assign n42458 = ( n12146 & n42456 ) | ( n12146 & ~n42457 ) | ( n42456 & ~n42457 ) ;
  assign n42459 = n16171 ^ n12313 ^ n4226 ;
  assign n42460 = ( n6796 & ~n14004 ) | ( n6796 & n42459 ) | ( ~n14004 & n42459 ) ;
  assign n42461 = n40655 ^ n32079 ^ n3889 ;
  assign n42462 = n42461 ^ n28659 ^ 1'b0 ;
  assign n42463 = n42460 | n42462 ;
  assign n42464 = n28220 ^ n3506 ^ 1'b0 ;
  assign n42465 = n42463 | n42464 ;
  assign n42466 = n23067 ^ n3107 ^ 1'b0 ;
  assign n42467 = n42301 ^ n30377 ^ n28221 ;
  assign n42468 = n8038 & ~n15469 ;
  assign n42469 = n30565 ^ n20693 ^ n11721 ;
  assign n42470 = ( ~n2904 & n19967 ) | ( ~n2904 & n22374 ) | ( n19967 & n22374 ) ;
  assign n42471 = n16625 & ~n30786 ;
  assign n42472 = n28843 ^ n3045 ^ 1'b0 ;
  assign n42473 = n18527 | n42472 ;
  assign n42474 = n23741 | n24906 ;
  assign n42475 = n42474 ^ n22844 ^ 1'b0 ;
  assign n42476 = n12593 ^ n6389 ^ n4303 ;
  assign n42477 = n42476 ^ n14030 ^ n1949 ;
  assign n42478 = ~n1710 & n34289 ;
  assign n42479 = n26587 ^ n10448 ^ n535 ;
  assign n42480 = ( n15351 & n16121 ) | ( n15351 & ~n42479 ) | ( n16121 & ~n42479 ) ;
  assign n42481 = n37605 ^ n31961 ^ n20572 ;
  assign n42482 = n19253 & n32027 ;
  assign n42483 = n11466 & n42482 ;
  assign n42484 = ( ~n9594 & n42481 ) | ( ~n9594 & n42483 ) | ( n42481 & n42483 ) ;
  assign n42485 = ( n13171 & ~n16733 ) | ( n13171 & n27049 ) | ( ~n16733 & n27049 ) ;
  assign n42488 = n21883 ^ n19483 ^ 1'b0 ;
  assign n42486 = n360 | n12000 ;
  assign n42487 = n42486 ^ n16007 ^ 1'b0 ;
  assign n42489 = n42488 ^ n42487 ^ n39250 ;
  assign n42490 = n31878 ^ n4935 ^ 1'b0 ;
  assign n42491 = n6454 & n42490 ;
  assign n42492 = n30145 ^ n18060 ^ 1'b0 ;
  assign n42493 = n8784 | n38354 ;
  assign n42494 = n42493 ^ n18000 ^ 1'b0 ;
  assign n42495 = n28815 ^ n25813 ^ n3202 ;
  assign n42504 = n786 & n15446 ;
  assign n42496 = n21878 ^ n7983 ^ n4586 ;
  assign n42497 = n20162 ^ n6940 ^ n4014 ;
  assign n42498 = ( n17210 & ~n23393 ) | ( n17210 & n38077 ) | ( ~n23393 & n38077 ) ;
  assign n42499 = ( n20013 & ~n40221 ) | ( n20013 & n42498 ) | ( ~n40221 & n42498 ) ;
  assign n42500 = n24183 ^ n18017 ^ 1'b0 ;
  assign n42501 = n42499 | n42500 ;
  assign n42502 = ( n12351 & ~n42497 ) | ( n12351 & n42501 ) | ( ~n42497 & n42501 ) ;
  assign n42503 = ( n9924 & n42496 ) | ( n9924 & n42502 ) | ( n42496 & n42502 ) ;
  assign n42505 = n42504 ^ n42503 ^ n8882 ;
  assign n42506 = ( n3145 & ~n5713 ) | ( n3145 & n39938 ) | ( ~n5713 & n39938 ) ;
  assign n42507 = n42506 ^ n22434 ^ n13091 ;
  assign n42508 = ( ~n4004 & n14523 ) | ( ~n4004 & n22100 ) | ( n14523 & n22100 ) ;
  assign n42509 = n16233 ^ n3983 ^ 1'b0 ;
  assign n42510 = n42508 | n42509 ;
  assign n42511 = n42510 ^ n6911 ^ 1'b0 ;
  assign n42512 = n12535 ^ n8692 ^ 1'b0 ;
  assign n42513 = ~n23955 & n42512 ;
  assign n42514 = ( n20732 & n41287 ) | ( n20732 & n42513 ) | ( n41287 & n42513 ) ;
  assign n42515 = n42514 ^ n15241 ^ 1'b0 ;
  assign n42516 = n21868 ^ n9383 ^ 1'b0 ;
  assign n42517 = n42515 & n42516 ;
  assign n42518 = ( n7556 & ~n9463 ) | ( n7556 & n27861 ) | ( ~n9463 & n27861 ) ;
  assign n42519 = n13322 & n39778 ;
  assign n42520 = ( x58 & n5495 ) | ( x58 & n14288 ) | ( n5495 & n14288 ) ;
  assign n42521 = n42520 ^ n13190 ^ n2883 ;
  assign n42522 = ( ~n6867 & n17976 ) | ( ~n6867 & n42521 ) | ( n17976 & n42521 ) ;
  assign n42523 = ~n2670 & n24374 ;
  assign n42524 = n8777 & ~n25226 ;
  assign n42525 = ~n12353 & n42524 ;
  assign n42526 = n42525 ^ n14286 ^ n10824 ;
  assign n42527 = n42523 | n42526 ;
  assign n42528 = n38429 ^ n9088 ^ n4834 ;
  assign n42529 = ( ~n15076 & n21429 ) | ( ~n15076 & n22168 ) | ( n21429 & n22168 ) ;
  assign n42531 = ( n9501 & n15875 ) | ( n9501 & n32826 ) | ( n15875 & n32826 ) ;
  assign n42532 = n14860 ^ n12308 ^ 1'b0 ;
  assign n42533 = n42531 & n42532 ;
  assign n42530 = n16862 & ~n24607 ;
  assign n42534 = n42533 ^ n42530 ^ 1'b0 ;
  assign n42535 = n3593 | n42534 ;
  assign n42536 = n42529 | n42535 ;
  assign n42537 = n18354 | n23435 ;
  assign n42538 = n42537 ^ n15683 ^ 1'b0 ;
  assign n42539 = n4880 & n11151 ;
  assign n42540 = n42539 ^ n11985 ^ 1'b0 ;
  assign n42541 = n42540 ^ n35018 ^ n4299 ;
  assign n42542 = n11012 | n36480 ;
  assign n42543 = n8602 & ~n42542 ;
  assign n42544 = n28303 ^ n13370 ^ 1'b0 ;
  assign n42545 = ~n42543 & n42544 ;
  assign n42546 = ~n42541 & n42545 ;
  assign n42547 = n27719 ^ n23601 ^ n4174 ;
  assign n42548 = ( n13961 & ~n18738 ) | ( n13961 & n18819 ) | ( ~n18738 & n18819 ) ;
  assign n42549 = n42548 ^ n19294 ^ n5230 ;
  assign n42550 = n40741 ^ n12066 ^ n7818 ;
  assign n42551 = n34849 ^ n28366 ^ n14789 ;
  assign n42552 = n41058 ^ n8626 ^ 1'b0 ;
  assign n42553 = n34669 ^ n22224 ^ n1040 ;
  assign n42554 = ( n5302 & n39084 ) | ( n5302 & n42553 ) | ( n39084 & n42553 ) ;
  assign n42555 = n42554 ^ n21785 ^ n19358 ;
  assign n42556 = n20218 & n42555 ;
  assign n42557 = n12465 ^ n10700 ^ n10364 ;
  assign n42558 = n40910 ^ n6480 ^ 1'b0 ;
  assign n42559 = ( ~n34820 & n42557 ) | ( ~n34820 & n42558 ) | ( n42557 & n42558 ) ;
  assign n42560 = ( ~n7226 & n30743 ) | ( ~n7226 & n42559 ) | ( n30743 & n42559 ) ;
  assign n42561 = ( n8112 & n22132 ) | ( n8112 & n30997 ) | ( n22132 & n30997 ) ;
  assign n42562 = ( n9679 & n39441 ) | ( n9679 & n40789 ) | ( n39441 & n40789 ) ;
  assign n42563 = ( n9285 & n42561 ) | ( n9285 & n42562 ) | ( n42561 & n42562 ) ;
  assign n42564 = n10343 ^ n9282 ^ 1'b0 ;
  assign n42565 = ~n6318 & n42564 ;
  assign n42566 = n41074 ^ n41060 ^ 1'b0 ;
  assign n42567 = n3386 & n42566 ;
  assign n42568 = n28512 | n35270 ;
  assign n42569 = n42567 | n42568 ;
  assign n42570 = ~n16947 & n32788 ;
  assign n42571 = ~n8694 & n42570 ;
  assign n42572 = n15878 ^ n5947 ^ n3226 ;
  assign n42573 = n5366 & ~n42572 ;
  assign n42574 = n42573 ^ n17777 ^ 1'b0 ;
  assign n42575 = n4431 & n42574 ;
  assign n42576 = n29423 ^ n14291 ^ 1'b0 ;
  assign n42577 = n35817 | n42576 ;
  assign n42578 = ( ~n13105 & n42575 ) | ( ~n13105 & n42577 ) | ( n42575 & n42577 ) ;
  assign n42579 = ( ~n325 & n906 ) | ( ~n325 & n4527 ) | ( n906 & n4527 ) ;
  assign n42580 = n42579 ^ n23056 ^ n3736 ;
  assign n42581 = n15987 ^ n15737 ^ n9352 ;
  assign n42582 = n3411 & ~n11594 ;
  assign n42583 = ~n42581 & n42582 ;
  assign n42584 = n4427 | n10877 ;
  assign n42585 = n42583 & ~n42584 ;
  assign n42586 = n8916 & ~n25454 ;
  assign n42587 = n42586 ^ n20042 ^ 1'b0 ;
  assign n42588 = ( n19271 & n42585 ) | ( n19271 & n42587 ) | ( n42585 & n42587 ) ;
  assign n42593 = n7185 ^ n1582 ^ x235 ;
  assign n42594 = x191 | n24692 ;
  assign n42595 = n13386 | n42594 ;
  assign n42596 = ( x215 & n42593 ) | ( x215 & n42595 ) | ( n42593 & n42595 ) ;
  assign n42589 = ~n811 & n5261 ;
  assign n42590 = n42589 ^ n26052 ^ 1'b0 ;
  assign n42591 = n9866 | n42590 ;
  assign n42592 = ~n8506 & n42591 ;
  assign n42597 = n42596 ^ n42592 ^ 1'b0 ;
  assign n42599 = n27046 ^ n6448 ^ n3469 ;
  assign n42600 = n12905 & n42599 ;
  assign n42601 = n42600 ^ n9081 ^ 1'b0 ;
  assign n42598 = n15035 ^ n14455 ^ n14316 ;
  assign n42602 = n42601 ^ n42598 ^ n36717 ;
  assign n42603 = n20737 | n42602 ;
  assign n42604 = n15949 ^ n11273 ^ 1'b0 ;
  assign n42605 = n1689 | n42604 ;
  assign n42606 = ~n9045 & n42605 ;
  assign n42608 = n23618 ^ n6318 ^ 1'b0 ;
  assign n42609 = ~n15736 & n42608 ;
  assign n42607 = n15939 & ~n35193 ;
  assign n42610 = n42609 ^ n42607 ^ n12467 ;
  assign n42611 = n19579 & ~n24765 ;
  assign n42612 = n12017 & n42611 ;
  assign n42613 = ( n3341 & n15602 ) | ( n3341 & n19693 ) | ( n15602 & n19693 ) ;
  assign n42614 = n10246 & ~n42613 ;
  assign n42615 = n42612 | n42614 ;
  assign n42616 = n28221 ^ n21261 ^ n7912 ;
  assign n42617 = ~n5454 & n14986 ;
  assign n42618 = ( n5920 & ~n42616 ) | ( n5920 & n42617 ) | ( ~n42616 & n42617 ) ;
  assign n42619 = n20103 ^ n9169 ^ n8438 ;
  assign n42620 = n42619 ^ n16482 ^ n5133 ;
  assign n42621 = n26750 ^ n8459 ^ 1'b0 ;
  assign n42622 = ( ~n2175 & n9186 ) | ( ~n2175 & n25925 ) | ( n9186 & n25925 ) ;
  assign n42623 = ( ~n42072 & n42621 ) | ( ~n42072 & n42622 ) | ( n42621 & n42622 ) ;
  assign n42625 = n39497 ^ n23606 ^ 1'b0 ;
  assign n42624 = ( n25270 & n25539 ) | ( n25270 & n30012 ) | ( n25539 & n30012 ) ;
  assign n42626 = n42625 ^ n42624 ^ n31503 ;
  assign n42627 = ( ~n5976 & n10657 ) | ( ~n5976 & n14430 ) | ( n10657 & n14430 ) ;
  assign n42628 = n41297 ^ n22196 ^ n8875 ;
  assign n42629 = ( n30173 & n39617 ) | ( n30173 & ~n42628 ) | ( n39617 & ~n42628 ) ;
  assign n42630 = ( n11609 & n30185 ) | ( n11609 & ~n30500 ) | ( n30185 & ~n30500 ) ;
  assign n42631 = n42630 ^ n32264 ^ x5 ;
  assign n42632 = n5279 | n41262 ;
  assign n42633 = n42632 ^ n19494 ^ n5689 ;
  assign n42634 = n35255 ^ n6135 ^ 1'b0 ;
  assign n42635 = n24659 ^ n9580 ^ 1'b0 ;
  assign n42636 = ~n3130 & n42635 ;
  assign n42637 = ~n4051 & n42636 ;
  assign n42638 = n12510 & n42637 ;
  assign n42639 = n28362 ^ n28218 ^ n17323 ;
  assign n42640 = ( ~n5952 & n8779 ) | ( ~n5952 & n25176 ) | ( n8779 & n25176 ) ;
  assign n42641 = ( n6668 & n30875 ) | ( n6668 & ~n42640 ) | ( n30875 & ~n42640 ) ;
  assign n42642 = n33233 ^ n12436 ^ n11789 ;
  assign n42643 = n42642 ^ n22208 ^ 1'b0 ;
  assign n42644 = n4337 ^ n3484 ^ 1'b0 ;
  assign n42645 = n8981 & ~n42644 ;
  assign n42646 = n8979 & ~n14206 ;
  assign n42647 = n42646 ^ n12867 ^ 1'b0 ;
  assign n42648 = n42647 ^ n15899 ^ 1'b0 ;
  assign n42649 = n42645 & n42648 ;
  assign n42650 = ( n25381 & ~n31556 ) | ( n25381 & n42649 ) | ( ~n31556 & n42649 ) ;
  assign n42651 = n8595 & ~n17026 ;
  assign n42652 = n4524 | n42364 ;
  assign n42653 = n42652 ^ n6281 ^ 1'b0 ;
  assign n42654 = ( n2447 & ~n3535 ) | ( n2447 & n11372 ) | ( ~n3535 & n11372 ) ;
  assign n42655 = n18937 & n42654 ;
  assign n42656 = n41532 & n42655 ;
  assign n42657 = n9034 ^ n7419 ^ 1'b0 ;
  assign n42658 = n4389 & n42657 ;
  assign n42659 = ( n11450 & n19508 ) | ( n11450 & ~n27636 ) | ( n19508 & ~n27636 ) ;
  assign n42660 = ( n1619 & ~n29299 ) | ( n1619 & n42659 ) | ( ~n29299 & n42659 ) ;
  assign n42661 = n35786 ^ n620 ^ 1'b0 ;
  assign n42662 = ~n16588 & n42661 ;
  assign n42663 = n42662 ^ n35059 ^ n4978 ;
  assign n42664 = n16483 ^ n6034 ^ 1'b0 ;
  assign n42665 = ~n12445 & n42664 ;
  assign n42666 = ( x58 & n10841 ) | ( x58 & n42665 ) | ( n10841 & n42665 ) ;
  assign n42667 = n23599 ^ n16322 ^ n4557 ;
  assign n42668 = ( n3811 & ~n36838 ) | ( n3811 & n42667 ) | ( ~n36838 & n42667 ) ;
  assign n42669 = ( n14480 & n42666 ) | ( n14480 & ~n42668 ) | ( n42666 & ~n42668 ) ;
  assign n42670 = ( n15289 & ~n34137 ) | ( n15289 & n42669 ) | ( ~n34137 & n42669 ) ;
  assign n42671 = n9357 & ~n9903 ;
  assign n42672 = n42671 ^ n40256 ^ n35340 ;
  assign n42673 = n42672 ^ n24028 ^ n18152 ;
  assign n42674 = n33200 ^ n25886 ^ n22248 ;
  assign n42675 = ( n21768 & ~n38080 ) | ( n21768 & n42674 ) | ( ~n38080 & n42674 ) ;
  assign n42676 = n23225 & ~n26680 ;
  assign n42677 = n4405 & n11092 ;
  assign n42678 = n42677 ^ n20925 ^ 1'b0 ;
  assign n42679 = n41708 ^ n24109 ^ 1'b0 ;
  assign n42680 = ~n26941 & n42679 ;
  assign n42682 = ( n7198 & n10846 ) | ( n7198 & n33459 ) | ( n10846 & n33459 ) ;
  assign n42681 = ( n500 & ~n33766 ) | ( n500 & n33889 ) | ( ~n33766 & n33889 ) ;
  assign n42683 = n42682 ^ n42681 ^ n21371 ;
  assign n42684 = n37547 ^ n28308 ^ n4876 ;
  assign n42685 = ( n4879 & n11262 ) | ( n4879 & ~n42684 ) | ( n11262 & ~n42684 ) ;
  assign n42686 = n3423 | n3539 ;
  assign n42687 = n42686 ^ n953 ^ 1'b0 ;
  assign n42688 = n42687 ^ n30377 ^ n20529 ;
  assign n42689 = n24074 ^ n19282 ^ n6117 ;
  assign n42690 = n35579 ^ n32241 ^ n25685 ;
  assign n42691 = n41181 ^ n4640 ^ 1'b0 ;
  assign n42692 = ( n5106 & ~n16431 ) | ( n5106 & n22404 ) | ( ~n16431 & n22404 ) ;
  assign n42695 = ( n5986 & n8845 ) | ( n5986 & ~n35492 ) | ( n8845 & ~n35492 ) ;
  assign n42693 = n13124 ^ n12136 ^ n1707 ;
  assign n42694 = ( n11682 & ~n13231 ) | ( n11682 & n42693 ) | ( ~n13231 & n42693 ) ;
  assign n42696 = n42695 ^ n42694 ^ n37705 ;
  assign n42697 = ( n17733 & n42692 ) | ( n17733 & n42696 ) | ( n42692 & n42696 ) ;
  assign n42698 = n5514 & n22908 ;
  assign n42699 = ~n42697 & n42698 ;
  assign n42700 = ~n8356 & n20175 ;
  assign n42701 = ( n23166 & ~n28218 ) | ( n23166 & n39667 ) | ( ~n28218 & n39667 ) ;
  assign n42702 = n29721 ^ n15276 ^ n5574 ;
  assign n42703 = ~n5151 & n19555 ;
  assign n42704 = n20170 & n42703 ;
  assign n42705 = n15891 ^ n15504 ^ n14300 ;
  assign n42706 = ( n36522 & n42704 ) | ( n36522 & n42705 ) | ( n42704 & n42705 ) ;
  assign n42707 = n5673 ^ n3603 ^ 1'b0 ;
  assign n42708 = n5928 & n42707 ;
  assign n42709 = n42708 ^ n31173 ^ n5113 ;
  assign n42710 = ~n5619 & n42709 ;
  assign n42711 = n42710 ^ n27036 ^ 1'b0 ;
  assign n42712 = n22082 | n40493 ;
  assign n42713 = n41203 & ~n42712 ;
  assign n42715 = n30141 ^ n23567 ^ n21807 ;
  assign n42714 = n17646 & n35780 ;
  assign n42716 = n42715 ^ n42714 ^ 1'b0 ;
  assign n42717 = n28314 ^ n4209 ^ n2451 ;
  assign n42718 = ( ~n5312 & n17429 ) | ( ~n5312 & n42717 ) | ( n17429 & n42717 ) ;
  assign n42719 = ~n19233 & n42718 ;
  assign n42720 = ~n327 & n42719 ;
  assign n42721 = n9795 ^ x195 ^ 1'b0 ;
  assign n42722 = n4350 | n42721 ;
  assign n42723 = ( n14631 & n29138 ) | ( n14631 & ~n42722 ) | ( n29138 & ~n42722 ) ;
  assign n42724 = n22284 & n36550 ;
  assign n42725 = n42724 ^ n19556 ^ 1'b0 ;
  assign n42726 = ( n13583 & n20148 ) | ( n13583 & ~n42725 ) | ( n20148 & ~n42725 ) ;
  assign n42727 = n39531 ^ n29333 ^ n11307 ;
  assign n42728 = n8685 ^ n3951 ^ 1'b0 ;
  assign n42729 = n14306 | n42728 ;
  assign n42730 = n42729 ^ n3317 ^ 1'b0 ;
  assign n42731 = n17694 ^ n1680 ^ 1'b0 ;
  assign n42732 = ( n8216 & n19946 ) | ( n8216 & n42731 ) | ( n19946 & n42731 ) ;
  assign n42733 = ( x205 & n18697 ) | ( x205 & ~n20702 ) | ( n18697 & ~n20702 ) ;
  assign n42735 = ~n35552 & n39322 ;
  assign n42736 = n42735 ^ n15471 ^ 1'b0 ;
  assign n42737 = ( n1787 & n39797 ) | ( n1787 & n42736 ) | ( n39797 & n42736 ) ;
  assign n42734 = n26742 & ~n33821 ;
  assign n42738 = n42737 ^ n42734 ^ 1'b0 ;
  assign n42739 = n11131 | n42738 ;
  assign n42740 = n11075 | n42739 ;
  assign n42741 = n25614 ^ n328 ^ 1'b0 ;
  assign n42742 = x163 | n34432 ;
  assign n42743 = n42742 ^ n37335 ^ 1'b0 ;
  assign n42744 = n42743 ^ n42654 ^ 1'b0 ;
  assign n42745 = ~n22278 & n25578 ;
  assign n42746 = n42745 ^ n21565 ^ 1'b0 ;
  assign n42747 = n17454 ^ n5032 ^ n3988 ;
  assign n42748 = n42747 ^ n6646 ^ 1'b0 ;
  assign n42749 = ( n8445 & ~n12564 ) | ( n8445 & n42748 ) | ( ~n12564 & n42748 ) ;
  assign n42753 = n2819 & n16599 ;
  assign n42751 = n25255 ^ n13456 ^ n11455 ;
  assign n42750 = ~n4439 & n14725 ;
  assign n42752 = n42751 ^ n42750 ^ 1'b0 ;
  assign n42754 = n42753 ^ n42752 ^ 1'b0 ;
  assign n42755 = ( n7182 & ~n22589 ) | ( n7182 & n26095 ) | ( ~n22589 & n26095 ) ;
  assign n42756 = ( n15765 & ~n22087 ) | ( n15765 & n35228 ) | ( ~n22087 & n35228 ) ;
  assign n42757 = n42756 ^ n40697 ^ n17479 ;
  assign n42758 = n41395 ^ n7788 ^ n3938 ;
  assign n42759 = ( ~n2798 & n17405 ) | ( ~n2798 & n42758 ) | ( n17405 & n42758 ) ;
  assign n42760 = n40359 & n42759 ;
  assign n42761 = n42760 ^ n5921 ^ n1697 ;
  assign n42762 = ( n12345 & n14038 ) | ( n12345 & n42761 ) | ( n14038 & n42761 ) ;
  assign n42763 = ~n4869 & n15734 ;
  assign n42764 = n42763 ^ n22860 ^ 1'b0 ;
  assign n42765 = n31026 ^ n27619 ^ n6754 ;
  assign n42766 = n5540 & n42765 ;
  assign n42767 = n42764 & n42766 ;
  assign n42769 = ~n26772 & n37461 ;
  assign n42770 = n42769 ^ n539 ^ 1'b0 ;
  assign n42768 = n3742 & ~n40252 ;
  assign n42771 = n42770 ^ n42768 ^ 1'b0 ;
  assign n42772 = n13813 | n24901 ;
  assign n42773 = n42772 ^ n37577 ^ 1'b0 ;
  assign n42774 = ( n17558 & n25082 ) | ( n17558 & n42773 ) | ( n25082 & n42773 ) ;
  assign n42775 = n2057 & n12344 ;
  assign n42776 = ( n28675 & ~n28942 ) | ( n28675 & n42775 ) | ( ~n28942 & n42775 ) ;
  assign n42777 = ~n3779 & n17838 ;
  assign n42778 = n42777 ^ n21303 ^ 1'b0 ;
  assign n42779 = n42778 ^ n18751 ^ n9632 ;
  assign n42780 = ~n35703 & n42779 ;
  assign n42781 = ~n31273 & n42780 ;
  assign n42782 = n42781 ^ n42388 ^ 1'b0 ;
  assign n42789 = ( ~n287 & n13104 ) | ( ~n287 & n33931 ) | ( n13104 & n33931 ) ;
  assign n42785 = n5305 ^ n3254 ^ 1'b0 ;
  assign n42786 = n20624 | n42785 ;
  assign n42787 = n13883 & n18158 ;
  assign n42788 = n42786 & n42787 ;
  assign n42783 = ~n29609 & n36874 ;
  assign n42784 = n42783 ^ n2573 ^ 1'b0 ;
  assign n42790 = n42789 ^ n42788 ^ n42784 ;
  assign n42793 = ( ~n329 & n2451 ) | ( ~n329 & n20594 ) | ( n2451 & n20594 ) ;
  assign n42791 = ( n4480 & ~n16590 ) | ( n4480 & n18270 ) | ( ~n16590 & n18270 ) ;
  assign n42792 = ( n5564 & ~n19522 ) | ( n5564 & n42791 ) | ( ~n19522 & n42791 ) ;
  assign n42794 = n42793 ^ n42792 ^ n17510 ;
  assign n42795 = n24486 ^ n24149 ^ n22310 ;
  assign n42796 = n9484 & n42795 ;
  assign n42797 = n26070 ^ n24818 ^ n8177 ;
  assign n42798 = n12991 ^ n799 ^ 1'b0 ;
  assign n42799 = n20229 & n42798 ;
  assign n42800 = n30576 ^ n26639 ^ n5858 ;
  assign n42801 = n42800 ^ n24818 ^ n5612 ;
  assign n42802 = n42801 ^ n9188 ^ n8209 ;
  assign n42803 = n5110 & n13034 ;
  assign n42804 = ~n42802 & n42803 ;
  assign n42805 = ( n23865 & n26729 ) | ( n23865 & ~n36886 ) | ( n26729 & ~n36886 ) ;
  assign n42806 = n32660 ^ n18604 ^ n10677 ;
  assign n42807 = n42806 ^ n37860 ^ n25369 ;
  assign n42808 = n36892 ^ n2099 ^ 1'b0 ;
  assign n42809 = n20150 | n42808 ;
  assign n42810 = ( n15836 & n42807 ) | ( n15836 & n42809 ) | ( n42807 & n42809 ) ;
  assign n42811 = n22884 ^ n7676 ^ n4012 ;
  assign n42812 = n28805 ^ n4209 ^ 1'b0 ;
  assign n42813 = ( n26176 & n26861 ) | ( n26176 & ~n42812 ) | ( n26861 & ~n42812 ) ;
  assign n42814 = ~n3879 & n12396 ;
  assign n42815 = n42814 ^ n33278 ^ n33250 ;
  assign n42816 = n16011 | n27686 ;
  assign n42817 = n42816 ^ n534 ^ n280 ;
  assign n42818 = n42049 ^ n23875 ^ n15460 ;
  assign n42819 = ( n3553 & n16752 ) | ( n3553 & ~n41975 ) | ( n16752 & ~n41975 ) ;
  assign n42820 = ~n16454 & n42819 ;
  assign n42821 = n11277 & n42820 ;
  assign n42822 = ( ~n8565 & n15144 ) | ( ~n8565 & n15273 ) | ( n15144 & n15273 ) ;
  assign n42823 = n29580 ^ n9318 ^ 1'b0 ;
  assign n42824 = ( n1365 & n2875 ) | ( n1365 & ~n5096 ) | ( n2875 & ~n5096 ) ;
  assign n42825 = ~n14931 & n42824 ;
  assign n42826 = n27395 ^ n973 ^ 1'b0 ;
  assign n42827 = ( n8079 & n23510 ) | ( n8079 & ~n42826 ) | ( n23510 & ~n42826 ) ;
  assign n42828 = n42827 ^ n8728 ^ 1'b0 ;
  assign n42829 = n4161 & n35383 ;
  assign n42830 = n41749 & n42829 ;
  assign n42831 = n2243 & ~n28929 ;
  assign n42832 = n42831 ^ n20801 ^ n19742 ;
  assign n42833 = n499 & ~n9965 ;
  assign n42834 = n42833 ^ n12302 ^ 1'b0 ;
  assign n42835 = n3749 | n12814 ;
  assign n42836 = n42835 ^ x147 ^ 1'b0 ;
  assign n42837 = n42836 ^ n11933 ^ n1369 ;
  assign n42838 = ( ~n5511 & n42834 ) | ( ~n5511 & n42837 ) | ( n42834 & n42837 ) ;
  assign n42839 = ( n9986 & n14889 ) | ( n9986 & n18234 ) | ( n14889 & n18234 ) ;
  assign n42840 = ( n5956 & ~n6177 ) | ( n5956 & n42839 ) | ( ~n6177 & n42839 ) ;
  assign n42841 = ~x219 & n16461 ;
  assign n42843 = n33279 | n34526 ;
  assign n42842 = n21832 ^ n20205 ^ n1429 ;
  assign n42844 = n42843 ^ n42842 ^ n5418 ;
  assign n42845 = n27068 ^ n21388 ^ n8872 ;
  assign n42846 = ( ~n580 & n19560 ) | ( ~n580 & n26349 ) | ( n19560 & n26349 ) ;
  assign n42847 = n7243 & ~n42846 ;
  assign n42848 = n6611 ^ n1596 ^ 1'b0 ;
  assign n42849 = n1155 | n42848 ;
  assign n42850 = n18300 ^ n15294 ^ 1'b0 ;
  assign n42851 = ( ~n21840 & n42849 ) | ( ~n21840 & n42850 ) | ( n42849 & n42850 ) ;
  assign n42852 = n13719 ^ n9030 ^ n2684 ;
  assign n42853 = ( n42847 & n42851 ) | ( n42847 & n42852 ) | ( n42851 & n42852 ) ;
  assign n42854 = n32730 ^ n6377 ^ 1'b0 ;
  assign n42855 = n38558 & ~n42854 ;
  assign n42856 = n2825 & n42855 ;
  assign n42858 = n4230 & ~n15407 ;
  assign n42859 = n42858 ^ n21140 ^ 1'b0 ;
  assign n42857 = n1818 & ~n5109 ;
  assign n42860 = n42859 ^ n42857 ^ 1'b0 ;
  assign n42861 = n5304 ^ x99 ^ 1'b0 ;
  assign n42862 = n42861 ^ n29920 ^ n12276 ;
  assign n42863 = ~n1789 & n42862 ;
  assign n42864 = ~n7024 & n19897 ;
  assign n42865 = n42864 ^ n8598 ^ 1'b0 ;
  assign n42866 = n3245 | n22955 ;
  assign n42867 = ( ~n41763 & n42865 ) | ( ~n41763 & n42866 ) | ( n42865 & n42866 ) ;
  assign n42868 = ( n1960 & n22478 ) | ( n1960 & n24892 ) | ( n22478 & n24892 ) ;
  assign n42869 = ( n12705 & ~n17868 ) | ( n12705 & n40830 ) | ( ~n17868 & n40830 ) ;
  assign n42870 = n6654 & n7312 ;
  assign n42871 = ( n12595 & ~n29810 ) | ( n12595 & n42870 ) | ( ~n29810 & n42870 ) ;
  assign n42872 = ( n5565 & n20490 ) | ( n5565 & ~n32597 ) | ( n20490 & ~n32597 ) ;
  assign n42873 = n857 | n15009 ;
  assign n42874 = n20827 | n42873 ;
  assign n42875 = ~n15147 & n26487 ;
  assign n42876 = n42875 ^ n34203 ^ 1'b0 ;
  assign n42877 = ( ~n42872 & n42874 ) | ( ~n42872 & n42876 ) | ( n42874 & n42876 ) ;
  assign n42878 = n25057 ^ n15452 ^ n9550 ;
  assign n42879 = n414 & n13895 ;
  assign n42880 = n3980 & n22021 ;
  assign n42881 = n42880 ^ n20987 ^ 1'b0 ;
  assign n42882 = n16893 ^ n14804 ^ n9221 ;
  assign n42883 = ( n16071 & n35343 ) | ( n16071 & ~n42882 ) | ( n35343 & ~n42882 ) ;
  assign n42887 = n26380 ^ n10374 ^ n6112 ;
  assign n42884 = n27548 ^ n8722 ^ 1'b0 ;
  assign n42885 = n22358 & ~n42884 ;
  assign n42886 = n42885 ^ n41452 ^ n28267 ;
  assign n42888 = n42887 ^ n42886 ^ n943 ;
  assign n42889 = ( ~n1151 & n5425 ) | ( ~n1151 & n25431 ) | ( n5425 & n25431 ) ;
  assign n42890 = ( n22863 & n29662 ) | ( n22863 & ~n42889 ) | ( n29662 & ~n42889 ) ;
  assign n42891 = ( n2412 & n10212 ) | ( n2412 & n24796 ) | ( n10212 & n24796 ) ;
  assign n42892 = n22645 ^ n9877 ^ 1'b0 ;
  assign n42893 = n4734 & n42892 ;
  assign n42895 = n25428 & n42355 ;
  assign n42894 = n13875 & n14538 ;
  assign n42896 = n42895 ^ n42894 ^ 1'b0 ;
  assign n42897 = n13395 & n24095 ;
  assign n42898 = n42257 ^ n37094 ^ n16812 ;
  assign n42899 = n28947 ^ n5280 ^ 1'b0 ;
  assign n42900 = ~n1735 & n42899 ;
  assign n42901 = n42900 ^ n41982 ^ n17962 ;
  assign n42902 = ( n8428 & n12855 ) | ( n8428 & n25183 ) | ( n12855 & n25183 ) ;
  assign n42904 = n42849 ^ n8213 ^ 1'b0 ;
  assign n42905 = n38225 ^ n23764 ^ 1'b0 ;
  assign n42906 = n42904 | n42905 ;
  assign n42903 = n35852 ^ n10371 ^ n4288 ;
  assign n42907 = n42906 ^ n42903 ^ n8205 ;
  assign n42908 = n9127 | n10642 ;
  assign n42909 = n25458 ^ n23289 ^ 1'b0 ;
  assign n42910 = n7729 ^ n5118 ^ 1'b0 ;
  assign n42911 = n41206 & ~n42910 ;
  assign n42912 = n7859 & ~n8137 ;
  assign n42913 = n42912 ^ n2485 ^ 1'b0 ;
  assign n42914 = n31922 ^ n18532 ^ 1'b0 ;
  assign n42915 = ( n29680 & ~n34370 ) | ( n29680 & n42914 ) | ( ~n34370 & n42914 ) ;
  assign n42916 = n30917 ^ n11899 ^ n7679 ;
  assign n42918 = n9565 ^ n7183 ^ 1'b0 ;
  assign n42919 = ~n34279 & n42918 ;
  assign n42920 = ~n28212 & n42919 ;
  assign n42921 = n42920 ^ n28500 ^ 1'b0 ;
  assign n42917 = n29253 ^ n20060 ^ 1'b0 ;
  assign n42922 = n42921 ^ n42917 ^ n17141 ;
  assign n42923 = n836 | n18258 ;
  assign n42924 = n30199 ^ n17045 ^ n8152 ;
  assign n42928 = ( n5704 & ~n6601 ) | ( n5704 & n11599 ) | ( ~n6601 & n11599 ) ;
  assign n42925 = n17959 ^ n12208 ^ 1'b0 ;
  assign n42926 = n30875 & n42925 ;
  assign n42927 = n8909 & n42926 ;
  assign n42929 = n42928 ^ n42927 ^ 1'b0 ;
  assign n42930 = n28144 ^ n20985 ^ 1'b0 ;
  assign n42931 = n40002 ^ n11443 ^ n3250 ;
  assign n42933 = n15635 & ~n19819 ;
  assign n42934 = n42933 ^ n12609 ^ 1'b0 ;
  assign n42932 = ( n981 & n15146 ) | ( n981 & n17229 ) | ( n15146 & n17229 ) ;
  assign n42935 = n42934 ^ n42932 ^ n29096 ;
  assign n42936 = n13434 ^ n6710 ^ n5336 ;
  assign n42937 = ( n1054 & ~n28285 ) | ( n1054 & n42936 ) | ( ~n28285 & n42936 ) ;
  assign n42938 = n40720 ^ n38261 ^ n33649 ;
  assign n42939 = ~n6584 & n34565 ;
  assign n42940 = ~n29084 & n42939 ;
  assign n42941 = n7013 ^ n6964 ^ 1'b0 ;
  assign n42942 = n20908 | n42941 ;
  assign n42943 = n42942 ^ n40022 ^ n5282 ;
  assign n42946 = n11402 ^ n8520 ^ n6945 ;
  assign n42947 = n42946 ^ n23058 ^ 1'b0 ;
  assign n42948 = n21565 & n42947 ;
  assign n42944 = ( n7735 & n18356 ) | ( n7735 & n32832 ) | ( n18356 & n32832 ) ;
  assign n42945 = n42944 ^ n20069 ^ n14283 ;
  assign n42949 = n42948 ^ n42945 ^ n22526 ;
  assign n42950 = n886 & n6728 ;
  assign n42951 = n42950 ^ n35641 ^ n30096 ;
  assign n42952 = n42951 ^ n16214 ^ 1'b0 ;
  assign n42953 = ( n13972 & n21247 ) | ( n13972 & n41638 ) | ( n21247 & n41638 ) ;
  assign n42954 = ~n5124 & n23815 ;
  assign n42955 = n11612 ^ n6865 ^ n5572 ;
  assign n42956 = ( n24214 & ~n42954 ) | ( n24214 & n42955 ) | ( ~n42954 & n42955 ) ;
  assign n42957 = n24475 ^ n23828 ^ n9591 ;
  assign n42958 = n17034 ^ n11710 ^ 1'b0 ;
  assign n42959 = n29260 ^ n18487 ^ 1'b0 ;
  assign n42960 = n3426 ^ n2926 ^ 1'b0 ;
  assign n42961 = n42959 & n42960 ;
  assign n42962 = n32002 ^ n20542 ^ 1'b0 ;
  assign n42963 = ~n10929 & n42962 ;
  assign n42964 = n42963 ^ n12151 ^ 1'b0 ;
  assign n42965 = ( n3932 & n12950 ) | ( n3932 & ~n42964 ) | ( n12950 & ~n42964 ) ;
  assign n42966 = n34669 ^ n31313 ^ n28635 ;
  assign n42967 = ( ~n1758 & n3385 ) | ( ~n1758 & n13730 ) | ( n3385 & n13730 ) ;
  assign n42968 = ~n8408 & n33070 ;
  assign n42969 = ( n15400 & n19603 ) | ( n15400 & ~n42968 ) | ( n19603 & ~n42968 ) ;
  assign n42970 = n20182 ^ n14094 ^ 1'b0 ;
  assign n42971 = ~n766 & n5344 ;
  assign n42972 = n42971 ^ x5 ^ 1'b0 ;
  assign n42973 = ~n3848 & n15321 ;
  assign n42974 = n42973 ^ n8469 ^ 1'b0 ;
  assign n42975 = n35503 ^ n20292 ^ n19934 ;
  assign n42976 = ( n26971 & n34357 ) | ( n26971 & ~n42975 ) | ( n34357 & ~n42975 ) ;
  assign n42977 = ( ~n12575 & n16372 ) | ( ~n12575 & n21816 ) | ( n16372 & n21816 ) ;
  assign n42978 = n42977 ^ n28037 ^ 1'b0 ;
  assign n42979 = ( ~n2866 & n21525 ) | ( ~n2866 & n33607 ) | ( n21525 & n33607 ) ;
  assign n42980 = n28438 ^ n8293 ^ n3948 ;
  assign n42981 = n42980 ^ n33600 ^ n32244 ;
  assign n42982 = n42981 ^ n33274 ^ n16027 ;
  assign n42983 = n4115 & ~n40914 ;
  assign n42985 = ( ~n2105 & n9003 ) | ( ~n2105 & n9227 ) | ( n9003 & n9227 ) ;
  assign n42984 = n38152 ^ n22287 ^ n8213 ;
  assign n42986 = n42985 ^ n42984 ^ n3504 ;
  assign n42987 = n24910 ^ n24366 ^ n12870 ;
  assign n42988 = n2401 | n41963 ;
  assign n42989 = n39824 ^ n39561 ^ n7641 ;
  assign n42990 = ( ~n2851 & n23934 ) | ( ~n2851 & n31490 ) | ( n23934 & n31490 ) ;
  assign n42991 = ~n8236 & n42990 ;
  assign n42992 = n30810 ^ n26530 ^ n13247 ;
  assign n42993 = ( n26835 & ~n37888 ) | ( n26835 & n42992 ) | ( ~n37888 & n42992 ) ;
  assign n42994 = ( n2244 & ~n33202 ) | ( n2244 & n41787 ) | ( ~n33202 & n41787 ) ;
  assign n42995 = n23748 & ~n42994 ;
  assign n42996 = ~n17548 & n42995 ;
  assign n42997 = n42996 ^ n5327 ^ 1'b0 ;
  assign n42998 = ~n42993 & n42997 ;
  assign n42999 = ~n1336 & n42507 ;
  assign n43000 = n42999 ^ n20746 ^ 1'b0 ;
  assign n43002 = ( n2631 & n15615 ) | ( n2631 & n16280 ) | ( n15615 & n16280 ) ;
  assign n43003 = n43002 ^ n10598 ^ 1'b0 ;
  assign n43004 = ( n8618 & n33538 ) | ( n8618 & n43003 ) | ( n33538 & n43003 ) ;
  assign n43001 = n16999 & n17587 ;
  assign n43005 = n43004 ^ n43001 ^ 1'b0 ;
  assign n43006 = ( n3856 & ~n21355 ) | ( n3856 & n23444 ) | ( ~n21355 & n23444 ) ;
  assign n43007 = ( n12598 & n39241 ) | ( n12598 & n43006 ) | ( n39241 & n43006 ) ;
  assign n43008 = n43007 ^ n17772 ^ n11197 ;
  assign n43009 = ( ~n11406 & n12998 ) | ( ~n11406 & n30616 ) | ( n12998 & n30616 ) ;
  assign n43010 = ~n8582 & n43009 ;
  assign n43011 = ( n1732 & n37324 ) | ( n1732 & ~n42824 ) | ( n37324 & ~n42824 ) ;
  assign n43012 = n25468 ^ n24863 ^ 1'b0 ;
  assign n43013 = n42443 ^ n7539 ^ 1'b0 ;
  assign n43014 = n13420 | n33697 ;
  assign n43015 = n33944 & ~n43014 ;
  assign n43016 = x235 & ~n12212 ;
  assign n43017 = n43016 ^ n10016 ^ 1'b0 ;
  assign n43018 = n43017 ^ n12691 ^ 1'b0 ;
  assign n43019 = n21532 | n41395 ;
  assign n43020 = n43019 ^ n28316 ^ n23197 ;
  assign n43021 = ( ~n17442 & n29329 ) | ( ~n17442 & n34356 ) | ( n29329 & n34356 ) ;
  assign n43022 = ( n24204 & ~n29347 ) | ( n24204 & n43021 ) | ( ~n29347 & n43021 ) ;
  assign n43023 = n43022 ^ n16157 ^ n814 ;
  assign n43024 = n43023 ^ n1404 ^ 1'b0 ;
  assign n43025 = ~n43020 & n43024 ;
  assign n43026 = ( n739 & n4376 ) | ( n739 & n12376 ) | ( n4376 & n12376 ) ;
  assign n43027 = ( ~n1126 & n4841 ) | ( ~n1126 & n41924 ) | ( n4841 & n41924 ) ;
  assign n43028 = ( n18488 & n37703 ) | ( n18488 & n43027 ) | ( n37703 & n43027 ) ;
  assign n43029 = n43028 ^ n26868 ^ 1'b0 ;
  assign n43032 = n8488 & n31400 ;
  assign n43030 = ~n31916 & n41994 ;
  assign n43031 = n43030 ^ n16372 ^ 1'b0 ;
  assign n43033 = n43032 ^ n43031 ^ n40540 ;
  assign n43034 = ( n11049 & ~n14740 ) | ( n11049 & n25579 ) | ( ~n14740 & n25579 ) ;
  assign n43035 = n18517 ^ n14341 ^ n1594 ;
  assign n43036 = n3789 & n43035 ;
  assign n43037 = n18684 ^ n7227 ^ n4609 ;
  assign n43038 = n43037 ^ n12476 ^ 1'b0 ;
  assign n43039 = n43038 ^ n13210 ^ n5104 ;
  assign n43040 = n3865 & n6754 ;
  assign n43041 = ~n27397 & n43040 ;
  assign n43042 = n43041 ^ n17426 ^ 1'b0 ;
  assign n43043 = n20371 & n43042 ;
  assign n43044 = ~n13789 & n37384 ;
  assign n43045 = n43044 ^ n4611 ^ 1'b0 ;
  assign n43046 = n43043 & n43045 ;
  assign n43047 = n5611 & ~n9904 ;
  assign n43048 = n11069 ^ n6028 ^ 1'b0 ;
  assign n43049 = n43047 | n43048 ;
  assign n43055 = n24211 ^ n9083 ^ 1'b0 ;
  assign n43051 = ( n5038 & n6889 ) | ( n5038 & ~n30804 ) | ( n6889 & ~n30804 ) ;
  assign n43052 = n40456 ^ n37556 ^ 1'b0 ;
  assign n43053 = ( n14123 & n43051 ) | ( n14123 & ~n43052 ) | ( n43051 & ~n43052 ) ;
  assign n43050 = n13423 & ~n16033 ;
  assign n43054 = n43053 ^ n43050 ^ 1'b0 ;
  assign n43056 = n43055 ^ n43054 ^ 1'b0 ;
  assign n43057 = n41367 ^ n37458 ^ 1'b0 ;
  assign n43059 = n26675 ^ n7456 ^ 1'b0 ;
  assign n43060 = ~n28001 & n43059 ;
  assign n43058 = ( n5828 & n7197 ) | ( n5828 & n21289 ) | ( n7197 & n21289 ) ;
  assign n43061 = n43060 ^ n43058 ^ n37999 ;
  assign n43062 = n21810 ^ n21262 ^ n18473 ;
  assign n43063 = n19441 ^ n18094 ^ 1'b0 ;
  assign n43064 = n15184 & n43063 ;
  assign n43065 = n24664 ^ n8899 ^ 1'b0 ;
  assign n43066 = n43064 & n43065 ;
  assign n43067 = ~n23395 & n43066 ;
  assign n43068 = n43067 ^ n30128 ^ n23260 ;
  assign n43069 = n5323 & ~n22020 ;
  assign n43070 = ~n23120 & n43069 ;
  assign n43071 = n37417 ^ n32770 ^ 1'b0 ;
  assign n43072 = n42350 ^ n2614 ^ 1'b0 ;
  assign n43073 = n43072 ^ n7361 ^ 1'b0 ;
  assign n43074 = n34614 ^ n12774 ^ n6864 ;
  assign n43075 = n12286 | n38957 ;
  assign n43076 = n43075 ^ n26345 ^ 1'b0 ;
  assign n43077 = ( ~n20462 & n43074 ) | ( ~n20462 & n43076 ) | ( n43074 & n43076 ) ;
  assign n43079 = n15481 ^ n12040 ^ n6141 ;
  assign n43078 = ( n34452 & ~n36223 ) | ( n34452 & n37732 ) | ( ~n36223 & n37732 ) ;
  assign n43080 = n43079 ^ n43078 ^ n16539 ;
  assign n43081 = n9603 | n13635 ;
  assign n43082 = ( n15980 & n21982 ) | ( n15980 & ~n43081 ) | ( n21982 & ~n43081 ) ;
  assign n43083 = n43082 ^ n30073 ^ n8390 ;
  assign n43084 = ( n14621 & n24145 ) | ( n14621 & n39910 ) | ( n24145 & n39910 ) ;
  assign n43085 = ( n22041 & ~n35167 ) | ( n22041 & n43084 ) | ( ~n35167 & n43084 ) ;
  assign n43086 = n28481 ^ n21024 ^ n10592 ;
  assign n43087 = n43086 ^ n30172 ^ n22599 ;
  assign n43088 = n43087 ^ n24502 ^ n23061 ;
  assign n43089 = n18343 & n41174 ;
  assign n43090 = ~n7153 & n13345 ;
  assign n43091 = n43090 ^ n1222 ^ 1'b0 ;
  assign n43092 = n2173 & n43091 ;
  assign n43093 = n14525 & n36249 ;
  assign n43094 = n43093 ^ n12863 ^ 1'b0 ;
  assign n43095 = ( n12705 & n20312 ) | ( n12705 & ~n21262 ) | ( n20312 & ~n21262 ) ;
  assign n43096 = ( ~n4477 & n17150 ) | ( ~n4477 & n43095 ) | ( n17150 & n43095 ) ;
  assign n43097 = n5672 | n24407 ;
  assign n43098 = n43097 ^ n3031 ^ 1'b0 ;
  assign n43099 = n9306 ^ n6752 ^ n3053 ;
  assign n43100 = ( ~n35269 & n43098 ) | ( ~n35269 & n43099 ) | ( n43098 & n43099 ) ;
  assign n43101 = ( n41481 & n43096 ) | ( n41481 & n43100 ) | ( n43096 & n43100 ) ;
  assign n43102 = ( n3737 & n9264 ) | ( n3737 & n42827 ) | ( n9264 & n42827 ) ;
  assign n43103 = n24342 ^ n7202 ^ 1'b0 ;
  assign n43104 = ( n11649 & n22081 ) | ( n11649 & ~n43098 ) | ( n22081 & ~n43098 ) ;
  assign n43105 = ( n2911 & n10967 ) | ( n2911 & n14602 ) | ( n10967 & n14602 ) ;
  assign n43106 = ~n13958 & n14948 ;
  assign n43107 = n40339 | n43106 ;
  assign n43108 = n16697 ^ n7857 ^ 1'b0 ;
  assign n43109 = ~n39617 & n43108 ;
  assign n43110 = n30500 | n43109 ;
  assign n43111 = n32328 ^ n15598 ^ 1'b0 ;
  assign n43112 = n7651 | n43111 ;
  assign n43113 = n13658 & n21835 ;
  assign n43115 = ~n11216 & n26672 ;
  assign n43116 = n5513 & n43115 ;
  assign n43114 = n7842 | n35680 ;
  assign n43117 = n43116 ^ n43114 ^ 1'b0 ;
  assign n43118 = n1057 | n14996 ;
  assign n43119 = n13746 & ~n43118 ;
  assign n43120 = ( n9486 & n28483 ) | ( n9486 & ~n43119 ) | ( n28483 & ~n43119 ) ;
  assign n43121 = n8303 ^ n4057 ^ 1'b0 ;
  assign n43122 = ~n6912 & n31912 ;
  assign n43123 = ( n8917 & n17405 ) | ( n8917 & n43122 ) | ( n17405 & n43122 ) ;
  assign n43124 = n29260 & ~n43123 ;
  assign n43125 = ( n2124 & n43121 ) | ( n2124 & n43124 ) | ( n43121 & n43124 ) ;
  assign n43126 = ( n13243 & n27013 ) | ( n13243 & n29094 ) | ( n27013 & n29094 ) ;
  assign n43127 = ( n32989 & n35011 ) | ( n32989 & n43126 ) | ( n35011 & n43126 ) ;
  assign n43128 = n10137 | n15180 ;
  assign n43129 = n10359 & ~n43128 ;
  assign n43130 = n2273 & ~n43129 ;
  assign n43131 = ( ~n3345 & n8752 ) | ( ~n3345 & n21199 ) | ( n8752 & n21199 ) ;
  assign n43132 = ( n672 & n31341 ) | ( n672 & n31507 ) | ( n31341 & n31507 ) ;
  assign n43133 = n7056 ^ n5134 ^ 1'b0 ;
  assign n43134 = n43133 ^ n19891 ^ n16083 ;
  assign n43135 = ( n14665 & n21842 ) | ( n14665 & n29645 ) | ( n21842 & n29645 ) ;
  assign n43136 = n41991 ^ n8670 ^ 1'b0 ;
  assign n43137 = n5110 & n43136 ;
  assign n43138 = n27653 & n43137 ;
  assign n43139 = n17827 ^ n13370 ^ n12901 ;
  assign n43140 = ~n14677 & n19198 ;
  assign n43141 = n35499 & n43140 ;
  assign n43142 = ~n11151 & n23231 ;
  assign n43143 = ( n1871 & n9867 ) | ( n1871 & n14395 ) | ( n9867 & n14395 ) ;
  assign n43144 = ( ~n917 & n9222 ) | ( ~n917 & n43143 ) | ( n9222 & n43143 ) ;
  assign n43145 = ( n4249 & n8860 ) | ( n4249 & n33285 ) | ( n8860 & n33285 ) ;
  assign n43147 = n29203 ^ n1725 ^ n1472 ;
  assign n43146 = n1338 | n4277 ;
  assign n43148 = n43147 ^ n43146 ^ n28848 ;
  assign n43149 = n14658 & ~n25961 ;
  assign n43150 = n43149 ^ n3358 ^ 1'b0 ;
  assign n43151 = n43150 ^ n13148 ^ 1'b0 ;
  assign n43152 = ( ~n6489 & n26892 ) | ( ~n6489 & n43151 ) | ( n26892 & n43151 ) ;
  assign n43153 = n23619 ^ n17388 ^ n8378 ;
  assign n43154 = n21381 ^ n7488 ^ 1'b0 ;
  assign n43155 = ( x208 & ~n16569 ) | ( x208 & n43154 ) | ( ~n16569 & n43154 ) ;
  assign n43156 = n30476 ^ n12665 ^ n6255 ;
  assign n43157 = ~n4211 & n43156 ;
  assign n43158 = ~n43155 & n43157 ;
  assign n43159 = n19835 ^ n15857 ^ n10222 ;
  assign n43160 = n6136 & n39976 ;
  assign n43161 = ~n43159 & n43160 ;
  assign n43162 = n42866 ^ n30241 ^ 1'b0 ;
  assign n43163 = n12703 | n43162 ;
  assign n43164 = n32820 ^ n20385 ^ n14722 ;
  assign n43165 = n5990 & ~n43164 ;
  assign n43166 = n43165 ^ n26794 ^ 1'b0 ;
  assign n43167 = n5765 | n9084 ;
  assign n43168 = n3285 | n43167 ;
  assign n43169 = ( n28362 & ~n37988 ) | ( n28362 & n43168 ) | ( ~n37988 & n43168 ) ;
  assign n43170 = n6314 ^ n4417 ^ 1'b0 ;
  assign n43171 = n18617 & n43170 ;
  assign n43172 = ( ~n25538 & n33579 ) | ( ~n25538 & n43171 ) | ( n33579 & n43171 ) ;
  assign n43173 = n43172 ^ n8824 ^ n3612 ;
  assign n43175 = n28703 ^ n10267 ^ n6142 ;
  assign n43174 = n23849 ^ n17910 ^ n14880 ;
  assign n43176 = n43175 ^ n43174 ^ n3507 ;
  assign n43177 = n3405 & n27343 ;
  assign n43178 = n43177 ^ n29935 ^ n13060 ;
  assign n43179 = n5643 & ~n43178 ;
  assign n43180 = n43179 ^ n872 ^ 1'b0 ;
  assign n43181 = n33693 ^ n23680 ^ n2830 ;
  assign n43182 = ( ~n10998 & n43180 ) | ( ~n10998 & n43181 ) | ( n43180 & n43181 ) ;
  assign n43183 = n12455 | n33108 ;
  assign n43184 = ~n3015 & n41934 ;
  assign n43185 = ~n20454 & n43184 ;
  assign n43186 = n43185 ^ n29585 ^ n4551 ;
  assign n43187 = n25534 ^ n19324 ^ 1'b0 ;
  assign n43188 = n43187 ^ n16235 ^ 1'b0 ;
  assign n43189 = n16333 | n43188 ;
  assign n43190 = n42585 ^ n3622 ^ 1'b0 ;
  assign n43191 = n17140 ^ n5282 ^ n4570 ;
  assign n43192 = ( n11580 & n13245 ) | ( n11580 & n43191 ) | ( n13245 & n43191 ) ;
  assign n43193 = n43192 ^ n32364 ^ 1'b0 ;
  assign n43194 = ~n4165 & n23062 ;
  assign n43195 = n5328 & ~n25415 ;
  assign n43196 = ( n8806 & ~n9514 ) | ( n8806 & n15141 ) | ( ~n9514 & n15141 ) ;
  assign n43197 = n43196 ^ n24493 ^ 1'b0 ;
  assign n43198 = n8102 ^ n7434 ^ n6996 ;
  assign n43199 = ( n15383 & n43197 ) | ( n15383 & ~n43198 ) | ( n43197 & ~n43198 ) ;
  assign n43200 = ( n4963 & ~n10736 ) | ( n4963 & n42751 ) | ( ~n10736 & n42751 ) ;
  assign n43201 = n43200 ^ n20257 ^ n19941 ;
  assign n43202 = n16309 ^ n10665 ^ n9168 ;
  assign n43203 = n33412 ^ n33021 ^ 1'b0 ;
  assign n43204 = n7672 & n43203 ;
  assign n43205 = n4853 ^ n4589 ^ 1'b0 ;
  assign n43206 = n20334 & ~n43205 ;
  assign n43207 = ( n917 & n18812 ) | ( n917 & ~n20231 ) | ( n18812 & ~n20231 ) ;
  assign n43208 = ( n17101 & ~n24025 ) | ( n17101 & n25554 ) | ( ~n24025 & n25554 ) ;
  assign n43209 = n13107 | n42103 ;
  assign n43210 = n10831 & ~n43209 ;
  assign n43211 = ( n11491 & n43208 ) | ( n11491 & ~n43210 ) | ( n43208 & ~n43210 ) ;
  assign n43212 = n6824 & n23662 ;
  assign n43213 = n43212 ^ n17552 ^ n10108 ;
  assign n43214 = n43213 ^ n18177 ^ 1'b0 ;
  assign n43215 = n21216 | n37263 ;
  assign n43216 = n6010 | n43215 ;
  assign n43217 = n3942 & n7597 ;
  assign n43218 = n27301 & n41994 ;
  assign n43219 = n43218 ^ n16460 ^ 1'b0 ;
  assign n43220 = ( n43216 & n43217 ) | ( n43216 & n43219 ) | ( n43217 & n43219 ) ;
  assign n43221 = n23127 | n32354 ;
  assign n43222 = n43221 ^ n38730 ^ 1'b0 ;
  assign n43223 = ( n17189 & ~n40104 ) | ( n17189 & n43222 ) | ( ~n40104 & n43222 ) ;
  assign n43225 = ~n1015 & n17478 ;
  assign n43226 = n14626 & n43225 ;
  assign n43227 = ( n3669 & n37258 ) | ( n3669 & ~n43226 ) | ( n37258 & ~n43226 ) ;
  assign n43224 = n8233 & ~n32346 ;
  assign n43228 = n43227 ^ n43224 ^ 1'b0 ;
  assign n43229 = n11289 ^ n9287 ^ 1'b0 ;
  assign n43230 = n2450 & ~n43229 ;
  assign n43231 = n43230 ^ n5514 ^ n3619 ;
  assign n43232 = ~n18589 & n43231 ;
  assign n43233 = n34592 ^ n28662 ^ n28572 ;
  assign n43234 = n43233 ^ n28434 ^ 1'b0 ;
  assign n43235 = ( n35457 & ~n36848 ) | ( n35457 & n41040 ) | ( ~n36848 & n41040 ) ;
  assign n43236 = n41535 ^ n12178 ^ n4677 ;
  assign n43237 = n27261 ^ n21445 ^ 1'b0 ;
  assign n43238 = n13850 | n43237 ;
  assign n43239 = ( n33017 & n40852 ) | ( n33017 & ~n43238 ) | ( n40852 & ~n43238 ) ;
  assign n43240 = n7265 | n18921 ;
  assign n43241 = ( x142 & n750 ) | ( x142 & ~n7636 ) | ( n750 & ~n7636 ) ;
  assign n43242 = n43241 ^ n33248 ^ n16649 ;
  assign n43243 = ( ~n11956 & n43240 ) | ( ~n11956 & n43242 ) | ( n43240 & n43242 ) ;
  assign n43244 = ~n25073 & n43243 ;
  assign n43245 = n43244 ^ n17391 ^ 1'b0 ;
  assign n43246 = ( ~n5959 & n17909 ) | ( ~n5959 & n18054 ) | ( n17909 & n18054 ) ;
  assign n43247 = n26511 ^ n16532 ^ n14870 ;
  assign n43248 = n43247 ^ n34248 ^ n7267 ;
  assign n43249 = n43246 & n43248 ;
  assign n43250 = n6173 & n43249 ;
  assign n43251 = n8645 & n43250 ;
  assign n43252 = n25321 ^ n1205 ^ 1'b0 ;
  assign n43253 = n22686 ^ n21157 ^ n10068 ;
  assign n43254 = n22714 ^ n18805 ^ 1'b0 ;
  assign n43255 = n26956 | n43254 ;
  assign n43256 = ( n8549 & n42579 ) | ( n8549 & n43255 ) | ( n42579 & n43255 ) ;
  assign n43257 = n43253 & n43256 ;
  assign n43258 = n43252 & n43257 ;
  assign n43259 = n1475 & n38722 ;
  assign n43260 = n43259 ^ n41785 ^ n26087 ;
  assign n43261 = ( n8766 & n10306 ) | ( n8766 & ~n17277 ) | ( n10306 & ~n17277 ) ;
  assign n43262 = n43261 ^ n38960 ^ n36595 ;
  assign n43263 = ( n2385 & n16704 ) | ( n2385 & ~n22027 ) | ( n16704 & ~n22027 ) ;
  assign n43264 = n13931 ^ n13098 ^ 1'b0 ;
  assign n43265 = ( ~n24377 & n33481 ) | ( ~n24377 & n33529 ) | ( n33481 & n33529 ) ;
  assign n43266 = ( n30309 & n43264 ) | ( n30309 & ~n43265 ) | ( n43264 & ~n43265 ) ;
  assign n43267 = ~n3402 & n18792 ;
  assign n43268 = n22060 & n43267 ;
  assign n43269 = ( n14670 & n19716 ) | ( n14670 & n43268 ) | ( n19716 & n43268 ) ;
  assign n43270 = n43269 ^ n18477 ^ n6460 ;
  assign n43271 = ( ~n3244 & n12922 ) | ( ~n3244 & n13977 ) | ( n12922 & n13977 ) ;
  assign n43272 = n36787 ^ n15428 ^ n7509 ;
  assign n43273 = n21803 & n43272 ;
  assign n43274 = ~n43271 & n43273 ;
  assign n43275 = ( n993 & ~n10100 ) | ( n993 & n13846 ) | ( ~n10100 & n13846 ) ;
  assign n43276 = ( ~n17635 & n41427 ) | ( ~n17635 & n43275 ) | ( n41427 & n43275 ) ;
  assign n43277 = n24294 ^ n14381 ^ n11620 ;
  assign n43278 = ( n491 & n1076 ) | ( n491 & ~n20817 ) | ( n1076 & ~n20817 ) ;
  assign n43279 = ~n7550 & n43278 ;
  assign n43280 = n43279 ^ n14829 ^ 1'b0 ;
  assign n43281 = n43280 ^ n11656 ^ 1'b0 ;
  assign n43282 = ~n35245 & n41304 ;
  assign n43283 = n19528 ^ n9096 ^ 1'b0 ;
  assign n43284 = n34336 & n43283 ;
  assign n43285 = n43284 ^ n26558 ^ n5218 ;
  assign n43286 = n33803 ^ n10125 ^ n9208 ;
  assign n43287 = n33145 & ~n43286 ;
  assign n43288 = n34499 ^ n30887 ^ n21596 ;
  assign n43289 = n43288 ^ n3094 ^ n1205 ;
  assign n43290 = n6179 ^ n6052 ^ 1'b0 ;
  assign n43291 = n43290 ^ n7491 ^ n485 ;
  assign n43292 = ~n39100 & n43291 ;
  assign n43293 = n43292 ^ n15933 ^ 1'b0 ;
  assign n43294 = n15193 & n43293 ;
  assign n43295 = n31430 ^ n21538 ^ n6067 ;
  assign n43297 = n2680 & n7941 ;
  assign n43298 = ~n4078 & n43297 ;
  assign n43296 = n14738 & ~n41244 ;
  assign n43299 = n43298 ^ n43296 ^ n5515 ;
  assign n43300 = n43299 ^ n42355 ^ n41515 ;
  assign n43302 = ( ~n5037 & n17690 ) | ( ~n5037 & n20687 ) | ( n17690 & n20687 ) ;
  assign n43301 = n24175 & n30298 ;
  assign n43303 = n43302 ^ n43301 ^ n4635 ;
  assign n43304 = ( n3437 & n20960 ) | ( n3437 & ~n28588 ) | ( n20960 & ~n28588 ) ;
  assign n43305 = n10096 & n33579 ;
  assign n43306 = n43305 ^ n26104 ^ 1'b0 ;
  assign n43307 = n43304 & ~n43306 ;
  assign n43308 = n2437 & ~n12876 ;
  assign n43309 = n22265 & ~n43308 ;
  assign n43310 = n14562 & n27755 ;
  assign n43311 = n43309 & n43310 ;
  assign n43312 = x40 & ~n12859 ;
  assign n43313 = n43311 & n43312 ;
  assign n43315 = n4369 | n21748 ;
  assign n43316 = n43315 ^ n36532 ^ 1'b0 ;
  assign n43317 = ( n16013 & ~n16513 ) | ( n16013 & n43316 ) | ( ~n16513 & n43316 ) ;
  assign n43314 = ( n11944 & n17686 ) | ( n11944 & n17841 ) | ( n17686 & n17841 ) ;
  assign n43318 = n43317 ^ n43314 ^ n13884 ;
  assign n43319 = ( n4160 & n16900 ) | ( n4160 & n25650 ) | ( n16900 & n25650 ) ;
  assign n43320 = n41692 ^ n39181 ^ 1'b0 ;
  assign n43321 = n23695 ^ n17960 ^ n15936 ;
  assign n43322 = n25309 ^ n15650 ^ n4702 ;
  assign n43323 = n22249 ^ n2947 ^ 1'b0 ;
  assign n43324 = n10540 & n43323 ;
  assign n43325 = ~n8302 & n43324 ;
  assign n43326 = n14054 | n16450 ;
  assign n43327 = n15132 | n43326 ;
  assign n43328 = n18828 | n18976 ;
  assign n43329 = n43328 ^ n22872 ^ 1'b0 ;
  assign n43331 = n5196 & n18184 ;
  assign n43330 = ~n343 & n5899 ;
  assign n43332 = n43331 ^ n43330 ^ 1'b0 ;
  assign n43333 = n34009 ^ n5660 ^ n3399 ;
  assign n43334 = ( ~n14492 & n33395 ) | ( ~n14492 & n43333 ) | ( n33395 & n43333 ) ;
  assign n43337 = n6703 ^ n1539 ^ 1'b0 ;
  assign n43335 = n18689 ^ n7730 ^ n3950 ;
  assign n43336 = ( ~n9675 & n21826 ) | ( ~n9675 & n43335 ) | ( n21826 & n43335 ) ;
  assign n43338 = n43337 ^ n43336 ^ n6853 ;
  assign n43339 = n8718 ^ n1935 ^ 1'b0 ;
  assign n43340 = n18930 | n43339 ;
  assign n43341 = n43340 ^ n30465 ^ n27361 ;
  assign n43342 = n11563 | n19936 ;
  assign n43343 = ( ~n1050 & n32070 ) | ( ~n1050 & n43342 ) | ( n32070 & n43342 ) ;
  assign n43344 = n43343 ^ n12313 ^ n10144 ;
  assign n43345 = n43344 ^ n7063 ^ n593 ;
  assign n43346 = ( n19239 & n31554 ) | ( n19239 & ~n43345 ) | ( n31554 & ~n43345 ) ;
  assign n43347 = n15189 ^ n4000 ^ n961 ;
  assign n43348 = ~n5477 & n41705 ;
  assign n43349 = n29961 & n43348 ;
  assign n43350 = ~n23641 & n43349 ;
  assign n43351 = n15455 | n40252 ;
  assign n43352 = ( n2347 & n2868 ) | ( n2347 & ~n4170 ) | ( n2868 & ~n4170 ) ;
  assign n43353 = n12291 | n43352 ;
  assign n43354 = ~n27836 & n33243 ;
  assign n43355 = n11989 ^ n9149 ^ 1'b0 ;
  assign n43356 = n3998 | n43355 ;
  assign n43357 = n7385 & ~n23884 ;
  assign n43358 = n43357 ^ n23293 ^ 1'b0 ;
  assign n43359 = ( n1266 & n43356 ) | ( n1266 & n43358 ) | ( n43356 & n43358 ) ;
  assign n43360 = ( n8399 & ~n26095 ) | ( n8399 & n36964 ) | ( ~n26095 & n36964 ) ;
  assign n43361 = ( n12335 & n17299 ) | ( n12335 & ~n28149 ) | ( n17299 & ~n28149 ) ;
  assign n43362 = ( n3257 & n12391 ) | ( n3257 & n28320 ) | ( n12391 & n28320 ) ;
  assign n43363 = ( n11256 & n12790 ) | ( n11256 & n43362 ) | ( n12790 & n43362 ) ;
  assign n43364 = n1144 & ~n43363 ;
  assign n43365 = ( ~n4792 & n10921 ) | ( ~n4792 & n18265 ) | ( n10921 & n18265 ) ;
  assign n43366 = n10761 | n43365 ;
  assign n43367 = n8502 & ~n43366 ;
  assign n43368 = n1082 | n26325 ;
  assign n43369 = n43368 ^ n2913 ^ 1'b0 ;
  assign n43370 = n12826 | n28420 ;
  assign n43371 = n11267 & ~n43370 ;
  assign n43372 = n29184 ^ n26341 ^ n11967 ;
  assign n43373 = n24346 ^ n9339 ^ n8239 ;
  assign n43374 = ( n40779 & n42152 ) | ( n40779 & ~n43373 ) | ( n42152 & ~n43373 ) ;
  assign n43377 = n25862 ^ n22713 ^ 1'b0 ;
  assign n43375 = n7749 ^ n5376 ^ 1'b0 ;
  assign n43376 = ( n19210 & n35237 ) | ( n19210 & ~n43375 ) | ( n35237 & ~n43375 ) ;
  assign n43378 = n43377 ^ n43376 ^ 1'b0 ;
  assign n43379 = n34218 ^ n5770 ^ 1'b0 ;
  assign n43380 = n18954 ^ n11781 ^ n8617 ;
  assign n43381 = n14215 & ~n43380 ;
  assign n43382 = n11106 & n37761 ;
  assign n43383 = n28906 & n43382 ;
  assign n43384 = n43383 ^ n9216 ^ n3579 ;
  assign n43385 = n19415 ^ n4215 ^ 1'b0 ;
  assign n43386 = n30596 | n31611 ;
  assign n43388 = n13605 & ~n29372 ;
  assign n43387 = ~n7409 & n7876 ;
  assign n43389 = n43388 ^ n43387 ^ 1'b0 ;
  assign n43390 = ~n7620 & n25297 ;
  assign n43391 = n8262 & n43390 ;
  assign n43393 = ( n8012 & n21174 ) | ( n8012 & n23087 ) | ( n21174 & n23087 ) ;
  assign n43394 = n43393 ^ n22930 ^ x83 ;
  assign n43392 = n8410 | n42786 ;
  assign n43395 = n43394 ^ n43392 ^ n2129 ;
  assign n43396 = n3331 & n7656 ;
  assign n43397 = ( ~n11304 & n28180 ) | ( ~n11304 & n43396 ) | ( n28180 & n43396 ) ;
  assign n43398 = ( ~n4933 & n8580 ) | ( ~n4933 & n16028 ) | ( n8580 & n16028 ) ;
  assign n43399 = n43398 ^ x39 ^ 1'b0 ;
  assign n43400 = ( ~n16720 & n40522 ) | ( ~n16720 & n43399 ) | ( n40522 & n43399 ) ;
  assign n43401 = ~n5357 & n8800 ;
  assign n43402 = ~n41056 & n43401 ;
  assign n43403 = n39065 ^ n3629 ^ 1'b0 ;
  assign n43404 = ~n43402 & n43403 ;
  assign n43407 = n2562 & ~n29981 ;
  assign n43408 = n43407 ^ n1132 ^ 1'b0 ;
  assign n43405 = n34564 ^ n34071 ^ n9200 ;
  assign n43406 = n33055 & n43405 ;
  assign n43409 = n43408 ^ n43406 ^ 1'b0 ;
  assign n43410 = n14163 | n37781 ;
  assign n43411 = n43410 ^ n6843 ^ 1'b0 ;
  assign n43412 = n28335 ^ n14084 ^ n8424 ;
  assign n43413 = n9736 & n43412 ;
  assign n43414 = n43411 & n43413 ;
  assign n43415 = n9526 | n43414 ;
  assign n43416 = n5374 | n43415 ;
  assign n43417 = n17529 & ~n32902 ;
  assign n43421 = n3351 | n14112 ;
  assign n43422 = n43421 ^ n39961 ^ 1'b0 ;
  assign n43418 = n35815 ^ n3813 ^ 1'b0 ;
  assign n43419 = n34469 & ~n43418 ;
  assign n43420 = n13009 & n43419 ;
  assign n43423 = n43422 ^ n43420 ^ n25938 ;
  assign n43424 = n42630 & n43423 ;
  assign n43425 = n26478 ^ n14163 ^ 1'b0 ;
  assign n43426 = ~n5864 & n19064 ;
  assign n43427 = n43426 ^ n39677 ^ n21429 ;
  assign n43428 = ( n30784 & n43425 ) | ( n30784 & ~n43427 ) | ( n43425 & ~n43427 ) ;
  assign n43429 = n29838 ^ n18173 ^ n12622 ;
  assign n43430 = n37158 ^ n17332 ^ 1'b0 ;
  assign n43431 = n40680 ^ n20015 ^ n16048 ;
  assign n43432 = n12181 ^ n1202 ^ 1'b0 ;
  assign n43433 = n39648 ^ n25834 ^ n1887 ;
  assign n43434 = n43433 ^ n21552 ^ n8073 ;
  assign n43435 = n43434 ^ n5338 ^ 1'b0 ;
  assign n43436 = n1369 | n15594 ;
  assign n43437 = n43436 ^ n13504 ^ n4867 ;
  assign n43438 = ( n34608 & n40296 ) | ( n34608 & ~n43437 ) | ( n40296 & ~n43437 ) ;
  assign n43439 = n17226 & n33866 ;
  assign n43440 = n43439 ^ n342 ^ 1'b0 ;
  assign n43442 = n31549 | n34644 ;
  assign n43441 = ( ~n14511 & n17074 ) | ( ~n14511 & n37781 ) | ( n17074 & n37781 ) ;
  assign n43443 = n43442 ^ n43441 ^ n23861 ;
  assign n43444 = n7903 & n11920 ;
  assign n43445 = n43444 ^ n36102 ^ n32186 ;
  assign n43446 = ~n9868 & n43445 ;
  assign n43447 = n43446 ^ n21679 ^ 1'b0 ;
  assign n43448 = ( n43440 & n43443 ) | ( n43440 & ~n43447 ) | ( n43443 & ~n43447 ) ;
  assign n43455 = n19945 ^ n5695 ^ 1'b0 ;
  assign n43456 = ~n15962 & n43455 ;
  assign n43449 = n10991 & ~n28719 ;
  assign n43450 = n43449 ^ n10695 ^ n4942 ;
  assign n43451 = n20958 ^ n13419 ^ 1'b0 ;
  assign n43452 = ( x185 & n733 ) | ( x185 & ~n43451 ) | ( n733 & ~n43451 ) ;
  assign n43453 = ( n36747 & n43450 ) | ( n36747 & ~n43452 ) | ( n43450 & ~n43452 ) ;
  assign n43454 = n43453 ^ n6671 ^ 1'b0 ;
  assign n43457 = n43456 ^ n43454 ^ n40602 ;
  assign n43461 = ~n5670 & n18853 ;
  assign n43458 = n16914 ^ n5022 ^ n325 ;
  assign n43459 = n12087 & n15434 ;
  assign n43460 = ( ~n35971 & n43458 ) | ( ~n35971 & n43459 ) | ( n43458 & n43459 ) ;
  assign n43462 = n43461 ^ n43460 ^ x230 ;
  assign n43463 = n11501 & ~n13517 ;
  assign n43464 = ( n2025 & ~n10454 ) | ( n2025 & n22716 ) | ( ~n10454 & n22716 ) ;
  assign n43465 = n24199 & ~n26798 ;
  assign n43466 = ~n43464 & n43465 ;
  assign n43467 = n17036 & ~n21496 ;
  assign n43468 = n18481 | n43467 ;
  assign n43469 = n31940 ^ n6982 ^ 1'b0 ;
  assign n43470 = n43469 ^ n18239 ^ n11178 ;
  assign n43471 = n23276 & n43470 ;
  assign n43472 = ~n18105 & n32294 ;
  assign n43473 = n43472 ^ n4397 ^ 1'b0 ;
  assign n43474 = n43473 ^ n37529 ^ n7708 ;
  assign n43475 = ( n10523 & n17610 ) | ( n10523 & ~n19711 ) | ( n17610 & ~n19711 ) ;
  assign n43476 = n21725 & ~n43475 ;
  assign n43477 = ( n18497 & n19370 ) | ( n18497 & n43476 ) | ( n19370 & n43476 ) ;
  assign n43478 = n18251 | n22697 ;
  assign n43479 = n26334 & ~n40320 ;
  assign n43480 = n43479 ^ n39827 ^ 1'b0 ;
  assign n43481 = n32923 ^ n25290 ^ n18364 ;
  assign n43482 = ( n10240 & n43480 ) | ( n10240 & ~n43481 ) | ( n43480 & ~n43481 ) ;
  assign n43483 = ( n3571 & n11251 ) | ( n3571 & n22604 ) | ( n11251 & n22604 ) ;
  assign n43484 = n16709 ^ n4094 ^ 1'b0 ;
  assign n43485 = n43483 & ~n43484 ;
  assign n43486 = n43485 ^ n4639 ^ 1'b0 ;
  assign n43487 = n30920 & n43486 ;
  assign n43488 = n20358 | n43084 ;
  assign n43490 = ( ~n5172 & n12539 ) | ( ~n5172 & n42540 ) | ( n12539 & n42540 ) ;
  assign n43489 = ( ~n574 & n6207 ) | ( ~n574 & n39133 ) | ( n6207 & n39133 ) ;
  assign n43491 = n43490 ^ n43489 ^ x82 ;
  assign n43492 = n8875 & ~n32464 ;
  assign n43493 = ~n7922 & n14621 ;
  assign n43494 = n43493 ^ n7671 ^ 1'b0 ;
  assign n43496 = ( n10462 & n25342 ) | ( n10462 & ~n29733 ) | ( n25342 & ~n29733 ) ;
  assign n43497 = n15330 | n43496 ;
  assign n43495 = n3265 & ~n10676 ;
  assign n43498 = n43497 ^ n43495 ^ 1'b0 ;
  assign n43499 = n35719 ^ n14939 ^ 1'b0 ;
  assign n43500 = n30714 & n43499 ;
  assign n43501 = n27125 ^ n15172 ^ n10179 ;
  assign n43502 = ( n7670 & n43067 ) | ( n7670 & n43501 ) | ( n43067 & n43501 ) ;
  assign n43503 = n13280 & ~n13521 ;
  assign n43504 = ( n16354 & n18783 ) | ( n16354 & n43503 ) | ( n18783 & n43503 ) ;
  assign n43505 = n9423 ^ x111 ^ 1'b0 ;
  assign n43506 = n1274 & ~n2506 ;
  assign n43507 = n43506 ^ n17662 ^ 1'b0 ;
  assign n43508 = ~n11448 & n18992 ;
  assign n43509 = ( n13279 & n43507 ) | ( n13279 & n43508 ) | ( n43507 & n43508 ) ;
  assign n43510 = n43509 ^ n21834 ^ n20215 ;
  assign n43511 = n32907 ^ n915 ^ 1'b0 ;
  assign n43512 = n18182 ^ n14306 ^ n12151 ;
  assign n43513 = ( ~n351 & n17289 ) | ( ~n351 & n43512 ) | ( n17289 & n43512 ) ;
  assign n43514 = ~n11172 & n18664 ;
  assign n43515 = n14626 & n43514 ;
  assign n43516 = n43515 ^ n34232 ^ n25044 ;
  assign n43517 = ( n693 & n43513 ) | ( n693 & n43516 ) | ( n43513 & n43516 ) ;
  assign n43518 = n20045 & ~n28491 ;
  assign n43519 = ( ~n6006 & n33478 ) | ( ~n6006 & n43518 ) | ( n33478 & n43518 ) ;
  assign n43520 = ~n12914 & n26629 ;
  assign n43521 = n43520 ^ n3412 ^ 1'b0 ;
  assign n43522 = ( n10256 & n43456 ) | ( n10256 & n43521 ) | ( n43456 & n43521 ) ;
  assign n43523 = n43522 ^ n10715 ^ 1'b0 ;
  assign n43524 = n19984 & n43523 ;
  assign n43525 = n42220 ^ n5558 ^ 1'b0 ;
  assign n43526 = n11759 & ~n43525 ;
  assign n43527 = ~n20314 & n43526 ;
  assign n43531 = n5861 & n10119 ;
  assign n43532 = n43531 ^ n20488 ^ 1'b0 ;
  assign n43528 = n17014 ^ n15873 ^ 1'b0 ;
  assign n43529 = ~n14836 & n43528 ;
  assign n43530 = n8822 & n43529 ;
  assign n43533 = n43532 ^ n43530 ^ 1'b0 ;
  assign n43534 = n8448 | n22279 ;
  assign n43535 = n31076 & n31571 ;
  assign n43536 = n43535 ^ n38833 ^ n6997 ;
  assign n43537 = n42217 ^ n8285 ^ n7432 ;
  assign n43538 = n43537 ^ n19611 ^ n7486 ;
  assign n43539 = ( n269 & n10612 ) | ( n269 & ~n35732 ) | ( n10612 & ~n35732 ) ;
  assign n43540 = ( n14678 & ~n17047 ) | ( n14678 & n23310 ) | ( ~n17047 & n23310 ) ;
  assign n43541 = ~n10033 & n29907 ;
  assign n43542 = ~n5350 & n10487 ;
  assign n43543 = ( n2592 & ~n9047 ) | ( n2592 & n10702 ) | ( ~n9047 & n10702 ) ;
  assign n43544 = n37421 ^ n32740 ^ n2292 ;
  assign n43545 = ( n41436 & n43543 ) | ( n41436 & ~n43544 ) | ( n43543 & ~n43544 ) ;
  assign n43546 = n43545 ^ n36370 ^ n749 ;
  assign n43547 = n26065 & ~n43546 ;
  assign n43548 = n43547 ^ n38464 ^ 1'b0 ;
  assign n43549 = ~n6116 & n31984 ;
  assign n43550 = n43549 ^ n35764 ^ 1'b0 ;
  assign n43551 = n21985 ^ n13163 ^ n1976 ;
  assign n43552 = n43551 ^ n11006 ^ 1'b0 ;
  assign n43553 = n25484 | n43552 ;
  assign n43554 = ~n2699 & n4368 ;
  assign n43555 = n36783 | n43554 ;
  assign n43556 = ( n8885 & n18620 ) | ( n8885 & n30351 ) | ( n18620 & n30351 ) ;
  assign n43557 = n27074 ^ n24995 ^ x53 ;
  assign n43558 = n40549 ^ n36957 ^ n9081 ;
  assign n43559 = ( n742 & n10999 ) | ( n742 & ~n32692 ) | ( n10999 & ~n32692 ) ;
  assign n43560 = n43559 ^ n6740 ^ n539 ;
  assign n43561 = ( n8321 & n43558 ) | ( n8321 & n43560 ) | ( n43558 & n43560 ) ;
  assign n43563 = n20077 ^ n5929 ^ 1'b0 ;
  assign n43564 = n43563 ^ n13844 ^ n1101 ;
  assign n43565 = n43564 ^ n27390 ^ n6678 ;
  assign n43566 = n43565 ^ n31430 ^ n12730 ;
  assign n43567 = ( n29159 & ~n43241 ) | ( n29159 & n43566 ) | ( ~n43241 & n43566 ) ;
  assign n43562 = n3967 | n4178 ;
  assign n43568 = n43567 ^ n43562 ^ 1'b0 ;
  assign n43569 = ( n627 & ~n18316 ) | ( n627 & n39392 ) | ( ~n18316 & n39392 ) ;
  assign n43570 = n43569 ^ n30792 ^ n15141 ;
  assign n43571 = n41114 ^ n30076 ^ 1'b0 ;
  assign n43572 = n1942 | n31124 ;
  assign n43573 = ~n3247 & n28919 ;
  assign n43574 = ( ~n10486 & n20801 ) | ( ~n10486 & n26823 ) | ( n20801 & n26823 ) ;
  assign n43575 = n43574 ^ n38718 ^ n6234 ;
  assign n43577 = ~n2755 & n10658 ;
  assign n43578 = n43577 ^ n11540 ^ 1'b0 ;
  assign n43576 = n7375 & ~n23045 ;
  assign n43579 = n43578 ^ n43576 ^ n14654 ;
  assign n43580 = n36415 ^ n5103 ^ n3918 ;
  assign n43581 = n43580 ^ n42606 ^ 1'b0 ;
  assign n43582 = n22631 & ~n43581 ;
  assign n43583 = n43102 ^ n35728 ^ 1'b0 ;
  assign n43584 = ~n20300 & n43583 ;
  assign n43585 = n9751 | n24981 ;
  assign n43586 = n26088 | n43585 ;
  assign n43587 = ( ~n5607 & n17665 ) | ( ~n5607 & n23518 ) | ( n17665 & n23518 ) ;
  assign n43588 = ( n7089 & ~n42405 ) | ( n7089 & n43587 ) | ( ~n42405 & n43587 ) ;
  assign n43589 = ~n16190 & n43588 ;
  assign n43590 = n27079 ^ n16424 ^ n5311 ;
  assign n43591 = n43590 ^ n34582 ^ n10366 ;
  assign n43592 = n25610 & ~n28547 ;
  assign n43593 = n13003 | n42220 ;
  assign n43594 = n43592 & ~n43593 ;
  assign n43595 = ( n24273 & n36968 ) | ( n24273 & ~n43594 ) | ( n36968 & ~n43594 ) ;
  assign n43596 = ( n13363 & n14279 ) | ( n13363 & ~n19924 ) | ( n14279 & ~n19924 ) ;
  assign n43597 = ( n43591 & n43595 ) | ( n43591 & ~n43596 ) | ( n43595 & ~n43596 ) ;
  assign n43598 = n28910 ^ n18097 ^ n3072 ;
  assign n43600 = n16048 ^ n15437 ^ 1'b0 ;
  assign n43601 = n6052 & ~n43600 ;
  assign n43599 = n32266 ^ n25818 ^ n938 ;
  assign n43602 = n43601 ^ n43599 ^ n18053 ;
  assign n43603 = x25 & n28626 ;
  assign n43604 = ~n6189 & n43603 ;
  assign n43605 = n43604 ^ n37716 ^ n16025 ;
  assign n43606 = n36056 ^ n8224 ^ n2948 ;
  assign n43607 = n43606 ^ n30643 ^ 1'b0 ;
  assign n43608 = ( n2601 & n25752 ) | ( n2601 & ~n43607 ) | ( n25752 & ~n43607 ) ;
  assign n43609 = n9075 ^ n7102 ^ 1'b0 ;
  assign n43610 = ( ~n4182 & n16410 ) | ( ~n4182 & n43609 ) | ( n16410 & n43609 ) ;
  assign n43611 = n11163 ^ n9614 ^ n8109 ;
  assign n43612 = ( n13100 & n43610 ) | ( n13100 & n43611 ) | ( n43610 & n43611 ) ;
  assign n43614 = ( ~x168 & n4207 ) | ( ~x168 & n17421 ) | ( n4207 & n17421 ) ;
  assign n43615 = ( ~n852 & n6422 ) | ( ~n852 & n43614 ) | ( n6422 & n43614 ) ;
  assign n43613 = n21992 ^ n5580 ^ n2590 ;
  assign n43616 = n43615 ^ n43613 ^ n10560 ;
  assign n43617 = n25323 | n43616 ;
  assign n43618 = n43612 & ~n43617 ;
  assign n43619 = n18087 | n31753 ;
  assign n43620 = n17691 & ~n43619 ;
  assign n43621 = n43620 ^ n24574 ^ 1'b0 ;
  assign n43622 = n5504 & ~n15519 ;
  assign n43623 = n43622 ^ n36846 ^ 1'b0 ;
  assign n43624 = n27908 ^ n19957 ^ n3925 ;
  assign n43625 = ( ~n9596 & n26436 ) | ( ~n9596 & n41605 ) | ( n26436 & n41605 ) ;
  assign n43626 = n28311 ^ n12162 ^ 1'b0 ;
  assign n43627 = n39612 ^ n1446 ^ 1'b0 ;
  assign n43628 = ~n14302 & n16284 ;
  assign n43629 = ~n11197 & n13951 ;
  assign n43630 = ~n340 & n43629 ;
  assign n43631 = n6383 & ~n13081 ;
  assign n43632 = ~n5082 & n43631 ;
  assign n43633 = ( n26318 & ~n31281 ) | ( n26318 & n32861 ) | ( ~n31281 & n32861 ) ;
  assign n43634 = n34763 ^ n33080 ^ n24578 ;
  assign n43635 = ( ~n645 & n2794 ) | ( ~n645 & n12032 ) | ( n2794 & n12032 ) ;
  assign n43636 = n43635 ^ n3803 ^ x217 ;
  assign n43637 = n43636 ^ n31698 ^ n27714 ;
  assign n43638 = n32770 ^ n21897 ^ 1'b0 ;
  assign n43639 = n14367 ^ n382 ^ 1'b0 ;
  assign n43640 = n43638 & n43639 ;
  assign n43641 = n36132 ^ n7485 ^ n5613 ;
  assign n43642 = n39033 ^ n22716 ^ n2506 ;
  assign n43643 = n43642 ^ n9272 ^ n7093 ;
  assign n43644 = ( n23539 & n43641 ) | ( n23539 & n43643 ) | ( n43641 & n43643 ) ;
  assign n43645 = n16758 ^ n4685 ^ 1'b0 ;
  assign n43646 = ( ~n5086 & n42278 ) | ( ~n5086 & n43645 ) | ( n42278 & n43645 ) ;
  assign n43647 = ( ~n3160 & n6248 ) | ( ~n3160 & n16999 ) | ( n6248 & n16999 ) ;
  assign n43648 = ( n32065 & ~n36874 ) | ( n32065 & n43647 ) | ( ~n36874 & n43647 ) ;
  assign n43649 = n17834 & ~n43648 ;
  assign n43650 = n1631 ^ n708 ^ 1'b0 ;
  assign n43651 = n31794 | n43650 ;
  assign n43660 = ( n9639 & n10748 ) | ( n9639 & n25376 ) | ( n10748 & n25376 ) ;
  assign n43661 = n2820 ^ x110 ^ 1'b0 ;
  assign n43662 = n43660 | n43661 ;
  assign n43654 = n4035 & ~n17014 ;
  assign n43655 = n43654 ^ n16979 ^ 1'b0 ;
  assign n43656 = n10519 ^ n8625 ^ 1'b0 ;
  assign n43657 = ( n1992 & n43655 ) | ( n1992 & ~n43656 ) | ( n43655 & ~n43656 ) ;
  assign n43658 = ( n18740 & ~n28643 ) | ( n18740 & n43657 ) | ( ~n28643 & n43657 ) ;
  assign n43652 = ( n9396 & n22335 ) | ( n9396 & ~n28263 ) | ( n22335 & ~n28263 ) ;
  assign n43653 = ( n27226 & ~n31034 ) | ( n27226 & n43652 ) | ( ~n31034 & n43652 ) ;
  assign n43659 = n43658 ^ n43653 ^ n38951 ;
  assign n43663 = n43662 ^ n43659 ^ 1'b0 ;
  assign n43664 = n27886 ^ n4828 ^ 1'b0 ;
  assign n43665 = n19773 & ~n43664 ;
  assign n43666 = n39291 ^ n30436 ^ 1'b0 ;
  assign n43667 = ( n22887 & n43665 ) | ( n22887 & ~n43666 ) | ( n43665 & ~n43666 ) ;
  assign n43668 = ( ~n26951 & n36295 ) | ( ~n26951 & n43667 ) | ( n36295 & n43667 ) ;
  assign n43669 = n34623 ^ n28522 ^ n16220 ;
  assign n43670 = n13412 | n43669 ;
  assign n43671 = ~n13432 & n31153 ;
  assign n43672 = n43671 ^ n5192 ^ 1'b0 ;
  assign n43673 = n20430 | n39283 ;
  assign n43674 = n8067 & ~n43673 ;
  assign n43675 = n3595 & n37438 ;
  assign n43676 = n43675 ^ n1100 ^ 1'b0 ;
  assign n43677 = n28474 ^ n12867 ^ n9905 ;
  assign n43680 = n16114 ^ n3567 ^ 1'b0 ;
  assign n43678 = n31790 ^ n15453 ^ 1'b0 ;
  assign n43679 = ~n1681 & n43678 ;
  assign n43681 = n43680 ^ n43679 ^ n12105 ;
  assign n43684 = n11784 ^ n1405 ^ 1'b0 ;
  assign n43685 = n2202 & ~n43684 ;
  assign n43682 = ~n2496 & n14889 ;
  assign n43683 = n43682 ^ n21754 ^ 1'b0 ;
  assign n43686 = n43685 ^ n43683 ^ n16780 ;
  assign n43687 = n38908 ^ n32119 ^ n25883 ;
  assign n43688 = ( n23544 & ~n30760 ) | ( n23544 & n31323 ) | ( ~n30760 & n31323 ) ;
  assign n43689 = n43688 ^ n42814 ^ n20512 ;
  assign n43690 = ( ~n10079 & n16702 ) | ( ~n10079 & n24273 ) | ( n16702 & n24273 ) ;
  assign n43691 = n9854 & ~n20941 ;
  assign n43692 = n43690 & n43691 ;
  assign n43693 = n13255 & ~n26478 ;
  assign n43694 = n43693 ^ n22077 ^ 1'b0 ;
  assign n43695 = n13714 & n43694 ;
  assign n43696 = n37023 & n43695 ;
  assign n43701 = n6768 & ~n24664 ;
  assign n43702 = ~n11611 & n43701 ;
  assign n43697 = n15378 ^ n11363 ^ n2098 ;
  assign n43698 = n43697 ^ n18909 ^ n8047 ;
  assign n43699 = n43698 ^ n40123 ^ n4479 ;
  assign n43700 = ~n3061 & n43699 ;
  assign n43703 = n43702 ^ n43700 ^ n29965 ;
  assign n43704 = ( n9797 & n18060 ) | ( n9797 & n36603 ) | ( n18060 & n36603 ) ;
  assign n43705 = n18626 ^ n17922 ^ n6126 ;
  assign n43706 = n43705 ^ n18705 ^ 1'b0 ;
  assign n43707 = n35216 & ~n43706 ;
  assign n43708 = ( ~n1146 & n43704 ) | ( ~n1146 & n43707 ) | ( n43704 & n43707 ) ;
  assign n43709 = n33119 ^ n18064 ^ 1'b0 ;
  assign n43710 = ( n5717 & ~n8528 ) | ( n5717 & n43709 ) | ( ~n8528 & n43709 ) ;
  assign n43711 = ( n33395 & n40345 ) | ( n33395 & n43710 ) | ( n40345 & n43710 ) ;
  assign n43712 = n5582 & ~n19095 ;
  assign n43713 = ~n16389 & n43712 ;
  assign n43714 = n36442 | n43713 ;
  assign n43715 = n23427 & n41239 ;
  assign n43716 = n43715 ^ n11785 ^ 1'b0 ;
  assign n43717 = n28645 ^ n21227 ^ 1'b0 ;
  assign n43718 = ~n26553 & n43717 ;
  assign n43719 = n39326 ^ n7479 ^ 1'b0 ;
  assign n43720 = n1573 & ~n43719 ;
  assign n43721 = n21584 ^ n17776 ^ 1'b0 ;
  assign n43722 = ( n16925 & ~n19239 ) | ( n16925 & n33192 ) | ( ~n19239 & n33192 ) ;
  assign n43724 = n5058 ^ n3548 ^ 1'b0 ;
  assign n43725 = n14844 & n43724 ;
  assign n43723 = ( n4225 & n22288 ) | ( n4225 & ~n37524 ) | ( n22288 & ~n37524 ) ;
  assign n43726 = n43725 ^ n43723 ^ n2527 ;
  assign n43727 = n34508 ^ n23188 ^ 1'b0 ;
  assign n43728 = n41244 ^ n15289 ^ 1'b0 ;
  assign n43733 = ( ~n883 & n7686 ) | ( ~n883 & n22374 ) | ( n7686 & n22374 ) ;
  assign n43729 = n4350 | n7072 ;
  assign n43730 = n18740 & ~n43729 ;
  assign n43731 = ~n14958 & n40687 ;
  assign n43732 = n43730 & n43731 ;
  assign n43734 = n43733 ^ n43732 ^ n29559 ;
  assign n43735 = n9762 & ~n28271 ;
  assign n43736 = n43734 & n43735 ;
  assign n43737 = ( ~n19413 & n21262 ) | ( ~n19413 & n25794 ) | ( n21262 & n25794 ) ;
  assign n43739 = n16298 & n24889 ;
  assign n43740 = ~n28194 & n43739 ;
  assign n43738 = n14391 ^ n3034 ^ 1'b0 ;
  assign n43741 = n43740 ^ n43738 ^ n5037 ;
  assign n43742 = n27736 ^ n4773 ^ 1'b0 ;
  assign n43743 = n43742 ^ n27368 ^ n26685 ;
  assign n43744 = ( n19034 & ~n25445 ) | ( n19034 & n33183 ) | ( ~n25445 & n33183 ) ;
  assign n43745 = n26742 & n35797 ;
  assign n43746 = n43745 ^ n10497 ^ 1'b0 ;
  assign n43747 = n11080 ^ n10748 ^ 1'b0 ;
  assign n43748 = n17513 & ~n43747 ;
  assign n43749 = ~n30991 & n43748 ;
  assign n43750 = n33973 ^ n19729 ^ n13485 ;
  assign n43751 = ( ~n43412 & n43749 ) | ( ~n43412 & n43750 ) | ( n43749 & n43750 ) ;
  assign n43752 = n37866 ^ n9056 ^ 1'b0 ;
  assign n43753 = n43751 & n43752 ;
  assign n43754 = ( n8636 & n13031 ) | ( n8636 & n20912 ) | ( n13031 & n20912 ) ;
  assign n43755 = n4202 & ~n31550 ;
  assign n43756 = n43755 ^ n7419 ^ 1'b0 ;
  assign n43757 = ( n2542 & n43754 ) | ( n2542 & n43756 ) | ( n43754 & n43756 ) ;
  assign n43758 = ( n20885 & n24003 ) | ( n20885 & ~n43757 ) | ( n24003 & ~n43757 ) ;
  assign n43759 = ( ~n15395 & n32587 ) | ( ~n15395 & n38781 ) | ( n32587 & n38781 ) ;
  assign n43760 = n37984 ^ n22539 ^ n15883 ;
  assign n43761 = n31241 & ~n43760 ;
  assign n43762 = n11005 | n23755 ;
  assign n43763 = n43762 ^ n16395 ^ 1'b0 ;
  assign n43764 = n43763 ^ n22597 ^ n18667 ;
  assign n43765 = n8990 ^ n2955 ^ 1'b0 ;
  assign n43766 = n41571 & n43765 ;
  assign n43767 = n3878 & ~n10004 ;
  assign n43768 = ~n37502 & n43767 ;
  assign n43769 = n33000 ^ n25352 ^ 1'b0 ;
  assign n43770 = ( n14708 & ~n24882 ) | ( n14708 & n43769 ) | ( ~n24882 & n43769 ) ;
  assign n43771 = n37895 ^ n17853 ^ n13483 ;
  assign n43772 = n26814 | n37841 ;
  assign n43775 = n15038 ^ n8798 ^ 1'b0 ;
  assign n43776 = n10573 | n43775 ;
  assign n43773 = n7136 & n33593 ;
  assign n43774 = ( ~n14769 & n28049 ) | ( ~n14769 & n43773 ) | ( n28049 & n43773 ) ;
  assign n43777 = n43776 ^ n43774 ^ n971 ;
  assign n43778 = n37263 ^ n17297 ^ 1'b0 ;
  assign n43779 = n33168 | n43778 ;
  assign n43780 = ( n13002 & n24132 ) | ( n13002 & ~n25319 ) | ( n24132 & ~n25319 ) ;
  assign n43781 = n43780 ^ n43680 ^ 1'b0 ;
  assign n43784 = n9273 ^ n5251 ^ n1359 ;
  assign n43785 = n43784 ^ n33669 ^ n4859 ;
  assign n43782 = n2853 ^ n1535 ^ n702 ;
  assign n43783 = n43782 ^ n18895 ^ n17069 ;
  assign n43786 = n43785 ^ n43783 ^ n27165 ;
  assign n43789 = ( ~n2345 & n6298 ) | ( ~n2345 & n8694 ) | ( n6298 & n8694 ) ;
  assign n43787 = n12685 | n14212 ;
  assign n43788 = n43787 ^ n12818 ^ 1'b0 ;
  assign n43790 = n43789 ^ n43788 ^ n26132 ;
  assign n43791 = n40598 ^ n39432 ^ n23053 ;
  assign n43792 = n6600 & ~n16362 ;
  assign n43793 = ~n24510 & n43792 ;
  assign n43794 = ( ~n3027 & n25368 ) | ( ~n3027 & n39079 ) | ( n25368 & n39079 ) ;
  assign n43795 = n43793 & n43794 ;
  assign n43798 = n13658 ^ n10844 ^ 1'b0 ;
  assign n43796 = n8431 & ~n30970 ;
  assign n43797 = n43796 ^ n18306 ^ 1'b0 ;
  assign n43799 = n43798 ^ n43797 ^ n27427 ;
  assign n43800 = n39498 ^ n6281 ^ 1'b0 ;
  assign n43801 = n29138 & n43800 ;
  assign n43802 = ( n14651 & n20796 ) | ( n14651 & n36000 ) | ( n20796 & n36000 ) ;
  assign n43803 = n36369 ^ n8569 ^ 1'b0 ;
  assign n43804 = n43802 | n43803 ;
  assign n43805 = ( ~n1285 & n28496 ) | ( ~n1285 & n30975 ) | ( n28496 & n30975 ) ;
  assign n43806 = n26754 & ~n43805 ;
  assign n43807 = n16837 & n43806 ;
  assign n43808 = n13486 ^ n9673 ^ 1'b0 ;
  assign n43809 = ~n14208 & n43808 ;
  assign n43810 = n31733 | n43809 ;
  assign n43811 = ( ~n21674 & n38503 ) | ( ~n21674 & n43810 ) | ( n38503 & n43810 ) ;
  assign n43812 = n39998 ^ n12118 ^ 1'b0 ;
  assign n43814 = ( ~n3874 & n21700 ) | ( ~n3874 & n27702 ) | ( n21700 & n27702 ) ;
  assign n43813 = ( n12259 & n24818 ) | ( n12259 & n41444 ) | ( n24818 & n41444 ) ;
  assign n43815 = n43814 ^ n43813 ^ n9494 ;
  assign n43816 = n15100 ^ n7794 ^ n7366 ;
  assign n43817 = ( n16514 & n31255 ) | ( n16514 & n43816 ) | ( n31255 & n43816 ) ;
  assign n43818 = ( ~n14194 & n23085 ) | ( ~n14194 & n43817 ) | ( n23085 & n43817 ) ;
  assign n43819 = ~n12637 & n22770 ;
  assign n43820 = ~n3301 & n43819 ;
  assign n43821 = n30494 | n43820 ;
  assign n43822 = n10423 & ~n14854 ;
  assign n43823 = n43822 ^ n12672 ^ 1'b0 ;
  assign n43824 = n3617 & n11406 ;
  assign n43825 = n3103 | n43824 ;
  assign n43826 = n36304 & ~n43825 ;
  assign n43827 = n16004 ^ n9590 ^ n8965 ;
  assign n43828 = n43827 ^ n3980 ^ n1457 ;
  assign n43829 = n1527 ^ n912 ^ 1'b0 ;
  assign n43830 = n22227 & ~n43829 ;
  assign n43831 = ( n23648 & n36007 ) | ( n23648 & n43830 ) | ( n36007 & n43830 ) ;
  assign n43832 = ( ~n12008 & n26769 ) | ( ~n12008 & n36548 ) | ( n26769 & n36548 ) ;
  assign n43833 = n43832 ^ n17369 ^ n5821 ;
  assign n43834 = ( ~n7475 & n15515 ) | ( ~n7475 & n16756 ) | ( n15515 & n16756 ) ;
  assign n43835 = n14759 ^ n12065 ^ n9170 ;
  assign n43836 = n43835 ^ n22082 ^ 1'b0 ;
  assign n43837 = ~n6394 & n43836 ;
  assign n43838 = n12191 ^ n4104 ^ 1'b0 ;
  assign n43839 = n1192 & n43838 ;
  assign n43840 = n27844 ^ n12689 ^ n4879 ;
  assign n43841 = n14602 & ~n43840 ;
  assign n43842 = n43841 ^ n3975 ^ 1'b0 ;
  assign n43843 = n26778 ^ n9574 ^ 1'b0 ;
  assign n43844 = n41873 & ~n43843 ;
  assign n43845 = n43844 ^ n27566 ^ n15309 ;
  assign n43846 = n36452 ^ n25091 ^ n12483 ;
  assign n43847 = ( ~n34364 & n38365 ) | ( ~n34364 & n38839 ) | ( n38365 & n38839 ) ;
  assign n43848 = n11306 | n25535 ;
  assign n43849 = n43848 ^ n18644 ^ n10845 ;
  assign n43852 = ( n368 & ~n7079 ) | ( n368 & n15228 ) | ( ~n7079 & n15228 ) ;
  assign n43853 = n43852 ^ n11241 ^ 1'b0 ;
  assign n43850 = n5784 & n23309 ;
  assign n43851 = ~n30154 & n43850 ;
  assign n43854 = n43853 ^ n43851 ^ n34058 ;
  assign n43855 = n36078 ^ n23711 ^ 1'b0 ;
  assign n43856 = ~n11991 & n43855 ;
  assign n43857 = n43856 ^ n13121 ^ n8081 ;
  assign n43858 = n35033 ^ n33519 ^ 1'b0 ;
  assign n43859 = n7562 & ~n43858 ;
  assign n43860 = n27765 & n28586 ;
  assign n43861 = n39206 ^ n28181 ^ 1'b0 ;
  assign n43862 = n16971 & n43861 ;
  assign n43863 = n24166 & n28721 ;
  assign n43864 = ~n43862 & n43863 ;
  assign n43865 = n25481 ^ n19869 ^ 1'b0 ;
  assign n43866 = n325 | n43865 ;
  assign n43870 = ( ~x83 & n24492 ) | ( ~x83 & n26573 ) | ( n24492 & n26573 ) ;
  assign n43867 = ( n6026 & ~n14836 ) | ( n6026 & n37930 ) | ( ~n14836 & n37930 ) ;
  assign n43868 = n15983 ^ x96 ^ 1'b0 ;
  assign n43869 = ~n43867 & n43868 ;
  assign n43871 = n43870 ^ n43869 ^ n41353 ;
  assign n43874 = ( ~n8941 & n10589 ) | ( ~n8941 & n20568 ) | ( n10589 & n20568 ) ;
  assign n43872 = n5390 & ~n6693 ;
  assign n43873 = n43872 ^ n5905 ^ 1'b0 ;
  assign n43875 = n43874 ^ n43873 ^ n37229 ;
  assign n43876 = n30924 & n43440 ;
  assign n43877 = n36633 ^ n31616 ^ 1'b0 ;
  assign n43878 = ( n10949 & n14203 ) | ( n10949 & n43877 ) | ( n14203 & n43877 ) ;
  assign n43879 = n13933 ^ n12644 ^ n11024 ;
  assign n43880 = n20052 | n33596 ;
  assign n43881 = n8732 & n22012 ;
  assign n43882 = n7585 | n13397 ;
  assign n43883 = n15690 ^ n14113 ^ n13684 ;
  assign n43884 = n43883 ^ n28772 ^ n26316 ;
  assign n43885 = ( n14909 & n43882 ) | ( n14909 & ~n43884 ) | ( n43882 & ~n43884 ) ;
  assign n43886 = ( ~n1293 & n25328 ) | ( ~n1293 & n25459 ) | ( n25328 & n25459 ) ;
  assign n43887 = ( n25862 & ~n43168 ) | ( n25862 & n43886 ) | ( ~n43168 & n43886 ) ;
  assign n43888 = n39528 ^ n34556 ^ n4063 ;
  assign n43889 = n23567 ^ n19733 ^ n5069 ;
  assign n43890 = n32622 & n43889 ;
  assign n43891 = ( x78 & n1261 ) | ( x78 & ~n8940 ) | ( n1261 & ~n8940 ) ;
  assign n43892 = n43891 ^ n17032 ^ n5617 ;
  assign n43893 = ~n5678 & n9836 ;
  assign n43894 = n43893 ^ n22107 ^ 1'b0 ;
  assign n43895 = n20340 ^ n2785 ^ n1113 ;
  assign n43896 = n43895 ^ n30251 ^ n10652 ;
  assign n43897 = n11576 ^ n11408 ^ 1'b0 ;
  assign n43898 = ( n2530 & n15506 ) | ( n2530 & n43897 ) | ( n15506 & n43897 ) ;
  assign n43899 = ( n11611 & ~n26643 ) | ( n11611 & n43898 ) | ( ~n26643 & n43898 ) ;
  assign n43900 = n43899 ^ n31000 ^ n3556 ;
  assign n43901 = n43900 ^ n25396 ^ n3048 ;
  assign n43902 = n15094 & ~n38282 ;
  assign n43903 = ( n18718 & n30490 ) | ( n18718 & ~n35002 ) | ( n30490 & ~n35002 ) ;
  assign n43904 = n33236 ^ n8188 ^ 1'b0 ;
  assign n43905 = n35994 & ~n43904 ;
  assign n43906 = n43905 ^ n7114 ^ 1'b0 ;
  assign n43907 = ~n14201 & n43906 ;
  assign n43908 = n35208 ^ n33336 ^ n8392 ;
  assign n43909 = ~n25442 & n41969 ;
  assign n43910 = ~n39924 & n43909 ;
  assign n43911 = ~n43908 & n43910 ;
  assign n43912 = n3441 & n7589 ;
  assign n43913 = n25525 ^ n14697 ^ n3601 ;
  assign n43914 = n1692 | n3677 ;
  assign n43915 = n1444 | n14227 ;
  assign n43916 = n24680 & ~n43915 ;
  assign n43917 = ( n9138 & ~n43914 ) | ( n9138 & n43916 ) | ( ~n43914 & n43916 ) ;
  assign n43918 = n25601 ^ n3813 ^ n756 ;
  assign n43919 = n2813 & ~n14478 ;
  assign n43920 = n43919 ^ n5565 ^ 1'b0 ;
  assign n43921 = n43920 ^ n9976 ^ n9065 ;
  assign n43923 = n32663 ^ n24647 ^ 1'b0 ;
  assign n43922 = n3030 & n8847 ;
  assign n43924 = n43923 ^ n43922 ^ 1'b0 ;
  assign n43925 = n5092 | n9285 ;
  assign n43926 = n43925 ^ n16845 ^ 1'b0 ;
  assign n43927 = n2255 | n14653 ;
  assign n43928 = n43927 ^ n27264 ^ n12712 ;
  assign n43929 = ( ~n15647 & n17105 ) | ( ~n15647 & n21737 ) | ( n17105 & n21737 ) ;
  assign n43931 = n18127 ^ n4994 ^ n3221 ;
  assign n43930 = ( n2256 & n28073 ) | ( n2256 & n33219 ) | ( n28073 & n33219 ) ;
  assign n43932 = n43931 ^ n43930 ^ n37382 ;
  assign n43933 = n42625 ^ n11208 ^ 1'b0 ;
  assign n43934 = ~n13742 & n29115 ;
  assign n43935 = n43934 ^ n16697 ^ 1'b0 ;
  assign n43936 = n39816 ^ n28129 ^ n8417 ;
  assign n43937 = n43936 ^ n16721 ^ 1'b0 ;
  assign n43938 = ~n43935 & n43937 ;
  assign n43939 = ~n672 & n6516 ;
  assign n43940 = n37006 & n43939 ;
  assign n43943 = n34340 & n38185 ;
  assign n43944 = n9546 & n43943 ;
  assign n43941 = n12049 & n21723 ;
  assign n43942 = n13169 | n43941 ;
  assign n43945 = n43944 ^ n43942 ^ 1'b0 ;
  assign n43946 = n31346 & ~n42508 ;
  assign n43947 = n43946 ^ n42846 ^ n39874 ;
  assign n43948 = n43947 ^ n17869 ^ n6106 ;
  assign n43950 = n25055 ^ n5935 ^ n3445 ;
  assign n43949 = ~n5328 & n16138 ;
  assign n43951 = n43950 ^ n43949 ^ 1'b0 ;
  assign n43952 = ( n23293 & ~n23676 ) | ( n23293 & n43951 ) | ( ~n23676 & n43951 ) ;
  assign n43953 = n31549 ^ n11365 ^ 1'b0 ;
  assign n43954 = n15686 | n43953 ;
  assign n43955 = ( n9687 & n34864 ) | ( n9687 & ~n43954 ) | ( n34864 & ~n43954 ) ;
  assign n43956 = ( n4000 & ~n18433 ) | ( n4000 & n31559 ) | ( ~n18433 & n31559 ) ;
  assign n43957 = n14341 ^ n1917 ^ n1125 ;
  assign n43958 = n19150 | n43957 ;
  assign n43959 = n37787 | n43958 ;
  assign n43960 = x218 & n40984 ;
  assign n43961 = ( n12212 & ~n16823 ) | ( n12212 & n18378 ) | ( ~n16823 & n18378 ) ;
  assign n43962 = n2158 & n43961 ;
  assign n43963 = n10229 & n43962 ;
  assign n43964 = n12776 | n14332 ;
  assign n43966 = ~n3164 & n18471 ;
  assign n43967 = n43966 ^ n4967 ^ 1'b0 ;
  assign n43965 = ( n3290 & n13896 ) | ( n3290 & n29778 ) | ( n13896 & n29778 ) ;
  assign n43968 = n43967 ^ n43965 ^ n39717 ;
  assign n43969 = ( n8576 & n29162 ) | ( n8576 & ~n37233 ) | ( n29162 & ~n37233 ) ;
  assign n43970 = ( n5246 & ~n26742 ) | ( n5246 & n28131 ) | ( ~n26742 & n28131 ) ;
  assign n43971 = ( ~n9677 & n12518 ) | ( ~n9677 & n15094 ) | ( n12518 & n15094 ) ;
  assign n43972 = n29374 & n43971 ;
  assign n43973 = n38871 ^ n9483 ^ n4815 ;
  assign n43974 = ( n26768 & ~n43972 ) | ( n26768 & n43973 ) | ( ~n43972 & n43973 ) ;
  assign n43975 = n35586 ^ n18983 ^ n13084 ;
  assign n43976 = ( n16573 & ~n23547 ) | ( n16573 & n43975 ) | ( ~n23547 & n43975 ) ;
  assign n43977 = ( n13849 & n14318 ) | ( n13849 & n19258 ) | ( n14318 & n19258 ) ;
  assign n43978 = n7283 ^ n922 ^ n541 ;
  assign n43979 = ( n7318 & ~n7645 ) | ( n7318 & n33712 ) | ( ~n7645 & n33712 ) ;
  assign n43980 = n18156 ^ n12488 ^ n12465 ;
  assign n43981 = ( ~x88 & n19649 ) | ( ~x88 & n29723 ) | ( n19649 & n29723 ) ;
  assign n43982 = n12210 & n37860 ;
  assign n43983 = n43982 ^ n21789 ^ 1'b0 ;
  assign n43984 = n17091 ^ n6364 ^ 1'b0 ;
  assign n43985 = n43984 ^ n8195 ^ 1'b0 ;
  assign n43986 = n31330 & n43985 ;
  assign n43987 = n21142 ^ n1390 ^ 1'b0 ;
  assign n43988 = ~n24665 & n43987 ;
  assign n43989 = ~n24510 & n43988 ;
  assign n43990 = ~n23018 & n43989 ;
  assign n43991 = ( n7551 & n18544 ) | ( n7551 & n24655 ) | ( n18544 & n24655 ) ;
  assign n43992 = n10885 & ~n43991 ;
  assign n43993 = n43992 ^ n37851 ^ 1'b0 ;
  assign n43994 = n14844 ^ n6252 ^ 1'b0 ;
  assign n43995 = ~n40478 & n43994 ;
  assign n43996 = ( n16064 & n26778 ) | ( n16064 & ~n43995 ) | ( n26778 & ~n43995 ) ;
  assign n43997 = n8022 | n43996 ;
  assign n43998 = n2711 & n37192 ;
  assign n43999 = n3227 & n43998 ;
  assign n44000 = ( n8899 & n12243 ) | ( n8899 & ~n43999 ) | ( n12243 & ~n43999 ) ;
  assign n44001 = ( n1527 & n9484 ) | ( n1527 & ~n20333 ) | ( n9484 & ~n20333 ) ;
  assign n44002 = ( ~n18774 & n30848 ) | ( ~n18774 & n44001 ) | ( n30848 & n44001 ) ;
  assign n44003 = x72 & ~n6878 ;
  assign n44004 = n44003 ^ n32528 ^ 1'b0 ;
  assign n44005 = n25756 ^ n14948 ^ 1'b0 ;
  assign n44006 = n22222 ^ n2816 ^ x212 ;
  assign n44007 = n11747 & n17548 ;
  assign n44008 = ~n44006 & n44007 ;
  assign n44009 = ( n14846 & n36539 ) | ( n14846 & ~n40316 ) | ( n36539 & ~n40316 ) ;
  assign n44010 = n44009 ^ n42824 ^ n9209 ;
  assign n44014 = ( ~n1173 & n6214 ) | ( ~n1173 & n6427 ) | ( n6214 & n6427 ) ;
  assign n44011 = n36208 ^ n12229 ^ n4264 ;
  assign n44012 = n20706 ^ n12377 ^ 1'b0 ;
  assign n44013 = n44011 | n44012 ;
  assign n44015 = n44014 ^ n44013 ^ n7402 ;
  assign n44016 = ( n16841 & n44010 ) | ( n16841 & n44015 ) | ( n44010 & n44015 ) ;
  assign n44017 = n30630 ^ n20697 ^ n6991 ;
  assign n44018 = n44017 ^ n33928 ^ 1'b0 ;
  assign n44019 = n3386 & n5149 ;
  assign n44020 = n12115 & n44019 ;
  assign n44021 = ( n7600 & n33845 ) | ( n7600 & ~n44020 ) | ( n33845 & ~n44020 ) ;
  assign n44022 = n13027 | n31223 ;
  assign n44023 = n44022 ^ n3647 ^ 1'b0 ;
  assign n44024 = n11392 & n15431 ;
  assign n44025 = ~n10805 & n17400 ;
  assign n44026 = ( n44023 & n44024 ) | ( n44023 & ~n44025 ) | ( n44024 & ~n44025 ) ;
  assign n44027 = ( n14384 & ~n26240 ) | ( n14384 & n35099 ) | ( ~n26240 & n35099 ) ;
  assign n44028 = ( ~n39497 & n40469 ) | ( ~n39497 & n44027 ) | ( n40469 & n44027 ) ;
  assign n44029 = n16436 ^ n7000 ^ 1'b0 ;
  assign n44030 = n44029 ^ n25447 ^ n1748 ;
  assign n44031 = ( n2960 & n8336 ) | ( n2960 & ~n29937 ) | ( n8336 & ~n29937 ) ;
  assign n44032 = ( n5131 & n29200 ) | ( n5131 & ~n44031 ) | ( n29200 & ~n44031 ) ;
  assign n44033 = ~n1500 & n3538 ;
  assign n44034 = n40758 & n44033 ;
  assign n44035 = n44034 ^ n33995 ^ n28330 ;
  assign n44036 = ~n8736 & n30924 ;
  assign n44037 = n44036 ^ n20698 ^ n11603 ;
  assign n44038 = n39802 ^ n7943 ^ 1'b0 ;
  assign n44039 = ( n4397 & n34990 ) | ( n4397 & ~n44038 ) | ( n34990 & ~n44038 ) ;
  assign n44040 = ~n22064 & n33153 ;
  assign n44041 = n26438 ^ n16432 ^ n3358 ;
  assign n44042 = n44041 ^ n6907 ^ 1'b0 ;
  assign n44043 = n2995 & n9897 ;
  assign n44044 = ~n8722 & n44043 ;
  assign n44045 = n44044 ^ n16431 ^ 1'b0 ;
  assign n44046 = n20529 ^ n2749 ^ 1'b0 ;
  assign n44047 = n27699 ^ n4268 ^ 1'b0 ;
  assign n44048 = n3040 & n44047 ;
  assign n44049 = n44048 ^ n16345 ^ 1'b0 ;
  assign n44050 = n44049 ^ n38469 ^ n29696 ;
  assign n44051 = ( n2994 & ~n6231 ) | ( n2994 & n8203 ) | ( ~n6231 & n8203 ) ;
  assign n44052 = ( ~n16176 & n23746 ) | ( ~n16176 & n44051 ) | ( n23746 & n44051 ) ;
  assign n44053 = ~n8727 & n15776 ;
  assign n44054 = n33957 & n44053 ;
  assign n44055 = ( n28542 & ~n39111 ) | ( n28542 & n44054 ) | ( ~n39111 & n44054 ) ;
  assign n44056 = n24662 ^ n14046 ^ 1'b0 ;
  assign n44057 = n44055 & ~n44056 ;
  assign n44058 = x203 & n38002 ;
  assign n44059 = ~n6054 & n44058 ;
  assign n44060 = n12842 | n17752 ;
  assign n44061 = n44060 ^ n39439 ^ 1'b0 ;
  assign n44062 = n1893 ^ n1188 ^ 1'b0 ;
  assign n44063 = n1745 & n12808 ;
  assign n44064 = n44063 ^ n4671 ^ 1'b0 ;
  assign n44065 = ( n3758 & n31730 ) | ( n3758 & n44064 ) | ( n31730 & n44064 ) ;
  assign n44066 = n38407 & ~n40107 ;
  assign n44067 = ( n1463 & n6139 ) | ( n1463 & n12215 ) | ( n6139 & n12215 ) ;
  assign n44068 = n44067 ^ n37350 ^ n37256 ;
  assign n44069 = ( n438 & ~n3428 ) | ( n438 & n25200 ) | ( ~n3428 & n25200 ) ;
  assign n44070 = n38031 ^ n25425 ^ n22043 ;
  assign n44071 = n44070 ^ n1042 ^ n891 ;
  assign n44072 = n30511 ^ n30263 ^ n14979 ;
  assign n44073 = n4658 & n35316 ;
  assign n44074 = n10423 & n44073 ;
  assign n44075 = ~n44072 & n44074 ;
  assign n44076 = n36150 ^ n18795 ^ 1'b0 ;
  assign n44078 = n3481 | n16814 ;
  assign n44079 = n44078 ^ n10513 ^ 1'b0 ;
  assign n44080 = ( ~n9462 & n36581 ) | ( ~n9462 & n44079 ) | ( n36581 & n44079 ) ;
  assign n44081 = n6241 | n44080 ;
  assign n44077 = n19166 ^ n18330 ^ n14552 ;
  assign n44082 = n44081 ^ n44077 ^ n27650 ;
  assign n44083 = n21044 & ~n44082 ;
  assign n44084 = n44083 ^ n14630 ^ 1'b0 ;
  assign n44085 = n25369 ^ n11327 ^ n3794 ;
  assign n44086 = ( n14934 & ~n17333 ) | ( n14934 & n33362 ) | ( ~n17333 & n33362 ) ;
  assign n44087 = n27486 ^ n24126 ^ n5429 ;
  assign n44088 = ( n3191 & n29633 ) | ( n3191 & n36855 ) | ( n29633 & n36855 ) ;
  assign n44089 = ( n33244 & n44087 ) | ( n33244 & ~n44088 ) | ( n44087 & ~n44088 ) ;
  assign n44091 = n42859 ^ n37877 ^ n34379 ;
  assign n44092 = n1146 | n9947 ;
  assign n44093 = n39466 ^ n27761 ^ n5529 ;
  assign n44094 = n535 | n44093 ;
  assign n44095 = n44092 | n44094 ;
  assign n44096 = ( ~n4131 & n44091 ) | ( ~n4131 & n44095 ) | ( n44091 & n44095 ) ;
  assign n44097 = n44096 ^ n20587 ^ n19708 ;
  assign n44090 = n35475 ^ n34592 ^ 1'b0 ;
  assign n44098 = n44097 ^ n44090 ^ n7483 ;
  assign n44099 = n24069 ^ n16764 ^ n7142 ;
  assign n44100 = n42595 ^ n34554 ^ n11505 ;
  assign n44101 = ( ~n3614 & n34345 ) | ( ~n3614 & n44100 ) | ( n34345 & n44100 ) ;
  assign n44102 = n41131 ^ n32223 ^ n29138 ;
  assign n44103 = n44102 ^ n19609 ^ 1'b0 ;
  assign n44104 = n28271 | n33535 ;
  assign n44105 = n44104 ^ n1602 ^ 1'b0 ;
  assign n44106 = ~n32554 & n41619 ;
  assign n44107 = ~n37645 & n44106 ;
  assign n44108 = ( n5877 & n19290 ) | ( n5877 & n35778 ) | ( n19290 & n35778 ) ;
  assign n44109 = n44108 ^ n18185 ^ 1'b0 ;
  assign n44110 = n35749 ^ n14638 ^ n7178 ;
  assign n44111 = n44110 ^ n37826 ^ 1'b0 ;
  assign n44112 = n30662 ^ n11676 ^ n10761 ;
  assign n44113 = n44112 ^ n2614 ^ 1'b0 ;
  assign n44114 = n32011 | n44113 ;
  assign n44115 = ( n22343 & n23650 ) | ( n22343 & ~n44114 ) | ( n23650 & ~n44114 ) ;
  assign n44116 = ( n1589 & n17935 ) | ( n1589 & n23768 ) | ( n17935 & n23768 ) ;
  assign n44117 = n44116 ^ n42041 ^ n5158 ;
  assign n44118 = ~n15805 & n33824 ;
  assign n44119 = n37246 ^ n31784 ^ 1'b0 ;
  assign n44120 = n31348 & n44119 ;
  assign n44121 = n39920 ^ n12250 ^ n2164 ;
  assign n44122 = ( ~n30370 & n44120 ) | ( ~n30370 & n44121 ) | ( n44120 & n44121 ) ;
  assign n44123 = ( n6092 & n8161 ) | ( n6092 & ~n10303 ) | ( n8161 & ~n10303 ) ;
  assign n44124 = n44123 ^ n39655 ^ n39636 ;
  assign n44125 = n37336 ^ n14580 ^ 1'b0 ;
  assign n44126 = ~n43840 & n44125 ;
  assign n44127 = ( ~n1801 & n18654 ) | ( ~n1801 & n19960 ) | ( n18654 & n19960 ) ;
  assign n44128 = n1034 & n44127 ;
  assign n44129 = n15621 & n44128 ;
  assign n44130 = n42137 ^ n17615 ^ 1'b0 ;
  assign n44131 = ( n6677 & ~n7259 ) | ( n6677 & n44130 ) | ( ~n7259 & n44130 ) ;
  assign n44132 = n24124 | n44131 ;
  assign n44133 = ( n3435 & n23144 ) | ( n3435 & n39584 ) | ( n23144 & n39584 ) ;
  assign n44134 = ( ~n24112 & n27526 ) | ( ~n24112 & n44133 ) | ( n27526 & n44133 ) ;
  assign n44135 = n29109 ^ n17043 ^ 1'b0 ;
  assign n44136 = ( n548 & n18768 ) | ( n548 & ~n33805 ) | ( n18768 & ~n33805 ) ;
  assign n44137 = ~n33695 & n37314 ;
  assign n44138 = ~n44136 & n44137 ;
  assign n44139 = n44135 & ~n44138 ;
  assign n44140 = n24581 ^ n10727 ^ n2974 ;
  assign n44141 = n44140 ^ n6645 ^ n6525 ;
  assign n44142 = n44141 ^ n20736 ^ 1'b0 ;
  assign n44143 = ~n21164 & n39460 ;
  assign n44144 = n32714 ^ n15852 ^ n5948 ;
  assign n44145 = n44143 & ~n44144 ;
  assign n44146 = ~n18473 & n19052 ;
  assign n44147 = n25765 & n44146 ;
  assign n44148 = n7554 & n21648 ;
  assign n44149 = n44148 ^ n28815 ^ 1'b0 ;
  assign n44150 = n39914 ^ n33645 ^ n23982 ;
  assign n44151 = n38954 ^ n21900 ^ n5725 ;
  assign n44152 = n37851 ^ n20741 ^ n19882 ;
  assign n44153 = n39564 ^ n27363 ^ 1'b0 ;
  assign n44154 = n16918 & n44153 ;
  assign n44155 = n44154 ^ n27550 ^ n27033 ;
  assign n44156 = n13355 ^ n6867 ^ n717 ;
  assign n44157 = ( n11210 & n39206 ) | ( n11210 & ~n44156 ) | ( n39206 & ~n44156 ) ;
  assign n44158 = ( n8656 & ~n22500 ) | ( n8656 & n37111 ) | ( ~n22500 & n37111 ) ;
  assign n44159 = ~n44157 & n44158 ;
  assign n44160 = ( n10036 & ~n26919 ) | ( n10036 & n44159 ) | ( ~n26919 & n44159 ) ;
  assign n44161 = ~n16517 & n26351 ;
  assign n44162 = ~n2941 & n44161 ;
  assign n44163 = n20360 ^ n11234 ^ n6327 ;
  assign n44164 = ( ~n33886 & n44162 ) | ( ~n33886 & n44163 ) | ( n44162 & n44163 ) ;
  assign n44165 = n38723 ^ n24303 ^ n16905 ;
  assign n44166 = ( n11837 & n19715 ) | ( n11837 & ~n33622 ) | ( n19715 & ~n33622 ) ;
  assign n44167 = n44166 ^ n17081 ^ 1'b0 ;
  assign n44168 = ( n4059 & n5437 ) | ( n4059 & ~n37180 ) | ( n5437 & ~n37180 ) ;
  assign n44169 = n17580 ^ n5147 ^ 1'b0 ;
  assign n44170 = n33823 & n44169 ;
  assign n44171 = n15205 ^ n7832 ^ 1'b0 ;
  assign n44172 = n11421 | n20672 ;
  assign n44173 = n44172 ^ n2932 ^ 1'b0 ;
  assign n44174 = ( n1688 & n21232 ) | ( n1688 & n27110 ) | ( n21232 & n27110 ) ;
  assign n44175 = n44174 ^ n27491 ^ 1'b0 ;
  assign n44176 = n959 & n44175 ;
  assign n44177 = n44176 ^ n36889 ^ n33573 ;
  assign n44178 = ( n6926 & ~n25542 ) | ( n6926 & n35231 ) | ( ~n25542 & n35231 ) ;
  assign n44179 = ( ~x216 & n31572 ) | ( ~x216 & n35860 ) | ( n31572 & n35860 ) ;
  assign n44180 = n37868 ^ n18976 ^ n8329 ;
  assign n44181 = ( n845 & n12553 ) | ( n845 & n30379 ) | ( n12553 & n30379 ) ;
  assign n44182 = n44181 ^ n10112 ^ n6763 ;
  assign n44183 = n33371 | n44182 ;
  assign n44184 = n24383 ^ n19319 ^ 1'b0 ;
  assign n44185 = n17211 ^ n9929 ^ n5660 ;
  assign n44186 = ( n14757 & n20630 ) | ( n14757 & ~n44185 ) | ( n20630 & ~n44185 ) ;
  assign n44187 = n10832 & n44186 ;
  assign n44188 = ( n3139 & n44184 ) | ( n3139 & n44187 ) | ( n44184 & n44187 ) ;
  assign n44189 = ( n24227 & n29155 ) | ( n24227 & ~n44188 ) | ( n29155 & ~n44188 ) ;
  assign n44190 = ~n31222 & n44189 ;
  assign n44191 = ~n1770 & n44190 ;
  assign n44192 = n32404 ^ n18818 ^ 1'b0 ;
  assign n44193 = n2711 & n44192 ;
  assign n44194 = n13006 & n15729 ;
  assign n44195 = n44194 ^ n12815 ^ 1'b0 ;
  assign n44196 = ( n13299 & ~n22010 ) | ( n13299 & n30611 ) | ( ~n22010 & n30611 ) ;
  assign n44197 = n44196 ^ n17517 ^ n1417 ;
  assign n44198 = ( ~n2081 & n16961 ) | ( ~n2081 & n19163 ) | ( n16961 & n19163 ) ;
  assign n44199 = ~n5151 & n12203 ;
  assign n44200 = ( n14334 & n44198 ) | ( n14334 & ~n44199 ) | ( n44198 & ~n44199 ) ;
  assign n44202 = n37610 ^ n30839 ^ n20506 ;
  assign n44201 = n13261 & ~n16339 ;
  assign n44203 = n44202 ^ n44201 ^ 1'b0 ;
  assign n44204 = n44203 ^ n39017 ^ n30191 ;
  assign n44205 = ( n3669 & n22830 ) | ( n3669 & ~n30563 ) | ( n22830 & ~n30563 ) ;
  assign n44206 = ~n470 & n11312 ;
  assign n44207 = ( n9237 & n14000 ) | ( n9237 & ~n44206 ) | ( n14000 & ~n44206 ) ;
  assign n44208 = ( n5821 & ~n15847 ) | ( n5821 & n17400 ) | ( ~n15847 & n17400 ) ;
  assign n44209 = ( n899 & ~n2019 ) | ( n899 & n3947 ) | ( ~n2019 & n3947 ) ;
  assign n44210 = n44209 ^ n21436 ^ n18479 ;
  assign n44211 = n1602 & n44210 ;
  assign n44212 = ( n4969 & n15560 ) | ( n4969 & ~n37669 ) | ( n15560 & ~n37669 ) ;
  assign n44213 = ( n4306 & n7166 ) | ( n4306 & ~n44212 ) | ( n7166 & ~n44212 ) ;
  assign n44214 = ( ~n271 & n747 ) | ( ~n271 & n36954 ) | ( n747 & n36954 ) ;
  assign n44215 = ~n8662 & n39460 ;
  assign n44216 = ( n16437 & n27350 ) | ( n16437 & n44215 ) | ( n27350 & n44215 ) ;
  assign n44217 = n31556 ^ n15013 ^ n817 ;
  assign n44218 = n10573 | n38789 ;
  assign n44219 = ( n10103 & n31428 ) | ( n10103 & n44218 ) | ( n31428 & n44218 ) ;
  assign n44220 = n21479 ^ n7109 ^ n1571 ;
  assign n44221 = n4863 & n44220 ;
  assign n44222 = ~n5270 & n44221 ;
  assign n44223 = ( n6618 & ~n26301 ) | ( n6618 & n39062 ) | ( ~n26301 & n39062 ) ;
  assign n44224 = ~n44222 & n44223 ;
  assign n44225 = n44224 ^ n29512 ^ 1'b0 ;
  assign n44226 = n44225 ^ n23332 ^ 1'b0 ;
  assign n44227 = ( ~n6501 & n6505 ) | ( ~n6501 & n44226 ) | ( n6505 & n44226 ) ;
  assign n44228 = n36721 ^ n8818 ^ 1'b0 ;
  assign n44229 = n44227 & n44228 ;
  assign n44230 = n9917 ^ n9046 ^ 1'b0 ;
  assign n44231 = n15229 & n44230 ;
  assign n44232 = n15157 ^ n10354 ^ 1'b0 ;
  assign n44233 = n13723 | n44232 ;
  assign n44234 = ( n34489 & ~n38997 ) | ( n34489 & n44233 ) | ( ~n38997 & n44233 ) ;
  assign n44235 = ~n14274 & n22286 ;
  assign n44236 = n44234 & n44235 ;
  assign n44237 = n44236 ^ n35656 ^ 1'b0 ;
  assign n44238 = n2355 | n44237 ;
  assign n44239 = ( n481 & n2024 ) | ( n481 & ~n2533 ) | ( n2024 & ~n2533 ) ;
  assign n44240 = ( ~n3635 & n13210 ) | ( ~n3635 & n44239 ) | ( n13210 & n44239 ) ;
  assign n44241 = ( x215 & ~n12353 ) | ( x215 & n31205 ) | ( ~n12353 & n31205 ) ;
  assign n44242 = n21316 ^ n4800 ^ 1'b0 ;
  assign n44243 = ~n29629 & n44242 ;
  assign n44244 = n19027 | n44243 ;
  assign n44245 = ( ~n4144 & n39816 ) | ( ~n4144 & n44244 ) | ( n39816 & n44244 ) ;
  assign n44246 = n1787 | n14020 ;
  assign n44247 = ( n10995 & n17848 ) | ( n10995 & ~n44246 ) | ( n17848 & ~n44246 ) ;
  assign n44248 = n44247 ^ n1327 ^ 1'b0 ;
  assign n44249 = n31534 ^ n3518 ^ 1'b0 ;
  assign n44250 = ~n33095 & n44249 ;
  assign n44251 = n44250 ^ n17103 ^ 1'b0 ;
  assign n44253 = ~n9107 & n20746 ;
  assign n44254 = n44253 ^ n4072 ^ 1'b0 ;
  assign n44252 = ~n2021 & n35581 ;
  assign n44255 = n44254 ^ n44252 ^ 1'b0 ;
  assign n44256 = n24178 ^ n20585 ^ n6012 ;
  assign n44257 = ( n8891 & ~n23074 ) | ( n8891 & n44256 ) | ( ~n23074 & n44256 ) ;
  assign n44258 = n44257 ^ n40656 ^ 1'b0 ;
  assign n44259 = n5075 ^ n1734 ^ 1'b0 ;
  assign n44260 = n44259 ^ n15030 ^ 1'b0 ;
  assign n44261 = n22161 ^ n10852 ^ 1'b0 ;
  assign n44262 = ( n1927 & ~n28728 ) | ( n1927 & n40957 ) | ( ~n28728 & n40957 ) ;
  assign n44263 = ( n20257 & n42139 ) | ( n20257 & n44262 ) | ( n42139 & n44262 ) ;
  assign n44264 = ( x180 & n8799 ) | ( x180 & ~n15997 ) | ( n8799 & ~n15997 ) ;
  assign n44265 = n20486 ^ n11331 ^ n7118 ;
  assign n44266 = ( n23495 & n44264 ) | ( n23495 & ~n44265 ) | ( n44264 & ~n44265 ) ;
  assign n44267 = n7425 & ~n32564 ;
  assign n44268 = n20282 ^ n10394 ^ 1'b0 ;
  assign n44271 = ~n26218 & n30713 ;
  assign n44272 = ~n30320 & n44271 ;
  assign n44269 = n27099 ^ n11897 ^ n7306 ;
  assign n44270 = n21422 & ~n44269 ;
  assign n44273 = n44272 ^ n44270 ^ 1'b0 ;
  assign n44274 = n27175 ^ n17273 ^ 1'b0 ;
  assign n44275 = n32923 & ~n44274 ;
  assign n44276 = n44273 & n44275 ;
  assign n44277 = n44276 ^ n33089 ^ 1'b0 ;
  assign n44278 = n5860 & ~n11745 ;
  assign n44279 = n1611 & ~n44278 ;
  assign n44280 = n44279 ^ n24935 ^ 1'b0 ;
  assign n44281 = ( ~n2362 & n20199 ) | ( ~n2362 & n24781 ) | ( n20199 & n24781 ) ;
  assign n44282 = ( x92 & ~n11320 ) | ( x92 & n23500 ) | ( ~n11320 & n23500 ) ;
  assign n44283 = n9056 ^ n1748 ^ 1'b0 ;
  assign n44284 = n44283 ^ n39803 ^ x228 ;
  assign n44285 = n16732 & ~n39358 ;
  assign n44286 = ( ~n14986 & n23942 ) | ( ~n14986 & n44285 ) | ( n23942 & n44285 ) ;
  assign n44290 = n29629 ^ n6651 ^ n999 ;
  assign n44287 = n19083 ^ n4108 ^ 1'b0 ;
  assign n44288 = n16655 & ~n44287 ;
  assign n44289 = ( n13448 & n18619 ) | ( n13448 & ~n44288 ) | ( n18619 & ~n44288 ) ;
  assign n44291 = n44290 ^ n44289 ^ n23087 ;
  assign n44292 = n22200 ^ n21808 ^ 1'b0 ;
  assign n44293 = ( n11591 & n15199 ) | ( n11591 & ~n44292 ) | ( n15199 & ~n44292 ) ;
  assign n44294 = n44293 ^ n11219 ^ 1'b0 ;
  assign n44295 = ( n8927 & n35674 ) | ( n8927 & ~n39883 ) | ( n35674 & ~n39883 ) ;
  assign n44296 = ( ~n1899 & n11213 ) | ( ~n1899 & n44295 ) | ( n11213 & n44295 ) ;
  assign n44297 = n16085 ^ n6031 ^ 1'b0 ;
  assign n44298 = ~n44296 & n44297 ;
  assign n44299 = n1014 & n37578 ;
  assign n44300 = n35894 & n44299 ;
  assign n44301 = n40972 ^ n38445 ^ n10527 ;
  assign n44302 = ( ~n9340 & n15678 ) | ( ~n9340 & n30187 ) | ( n15678 & n30187 ) ;
  assign n44303 = n19630 ^ n6596 ^ n3904 ;
  assign n44304 = n24697 ^ n10850 ^ n10597 ;
  assign n44305 = ( n18251 & ~n29270 ) | ( n18251 & n42346 ) | ( ~n29270 & n42346 ) ;
  assign n44306 = n1983 & n31949 ;
  assign n44307 = n44306 ^ n31534 ^ 1'b0 ;
  assign n44308 = n39269 ^ n18797 ^ 1'b0 ;
  assign n44309 = ~n3622 & n44308 ;
  assign n44310 = n12752 ^ n10005 ^ n5938 ;
  assign n44311 = n44310 ^ n12848 ^ 1'b0 ;
  assign n44312 = n44309 & n44311 ;
  assign n44313 = ( n5046 & n20690 ) | ( n5046 & ~n27652 ) | ( n20690 & ~n27652 ) ;
  assign n44314 = n44313 ^ n24075 ^ n6984 ;
  assign n44315 = ( n5598 & ~n9181 ) | ( n5598 & n39124 ) | ( ~n9181 & n39124 ) ;
  assign n44316 = n21752 ^ n17516 ^ n3536 ;
  assign n44317 = n44316 ^ n15123 ^ 1'b0 ;
  assign n44318 = n14014 ^ n11044 ^ n1683 ;
  assign n44319 = n43507 ^ n17188 ^ n11368 ;
  assign n44320 = n44319 ^ n21118 ^ 1'b0 ;
  assign n44321 = ( n13306 & n44318 ) | ( n13306 & ~n44320 ) | ( n44318 & ~n44320 ) ;
  assign n44322 = n29935 ^ n7779 ^ 1'b0 ;
  assign n44323 = n44322 ^ n41274 ^ 1'b0 ;
  assign n44324 = n12648 & n44323 ;
  assign n44325 = n12864 & ~n44324 ;
  assign n44326 = n44325 ^ n2508 ^ 1'b0 ;
  assign n44327 = ( ~n6735 & n20321 ) | ( ~n6735 & n36341 ) | ( n20321 & n36341 ) ;
  assign n44328 = n44327 ^ n28858 ^ n7765 ;
  assign n44329 = n8447 ^ n5757 ^ 1'b0 ;
  assign n44330 = n34620 & n44329 ;
  assign n44331 = n35017 ^ n28813 ^ 1'b0 ;
  assign n44332 = ( n4477 & ~n29135 ) | ( n4477 & n44331 ) | ( ~n29135 & n44331 ) ;
  assign n44333 = n42836 ^ n31995 ^ n23999 ;
  assign n44334 = n19653 ^ n9721 ^ 1'b0 ;
  assign n44335 = n44334 ^ n38213 ^ n15147 ;
  assign n44336 = n24975 ^ n17588 ^ n13019 ;
  assign n44337 = n44336 ^ n28471 ^ n16911 ;
  assign n44338 = ~n6388 & n34071 ;
  assign n44339 = n44338 ^ n7465 ^ n598 ;
  assign n44340 = n8831 | n43824 ;
  assign n44341 = n4314 ^ n2545 ^ 1'b0 ;
  assign n44342 = n4517 | n44341 ;
  assign n44343 = n14327 & ~n44342 ;
  assign n44344 = n44343 ^ n25251 ^ 1'b0 ;
  assign n44345 = n35786 ^ n17614 ^ n14071 ;
  assign n44346 = ~n13226 & n44345 ;
  assign n44347 = n17877 ^ n15876 ^ 1'b0 ;
  assign n44348 = n24816 & n44347 ;
  assign n44355 = n21667 ^ n18598 ^ n15146 ;
  assign n44356 = n2977 | n44355 ;
  assign n44352 = n34807 ^ n21565 ^ n7815 ;
  assign n44353 = n44352 ^ n24346 ^ n20556 ;
  assign n44354 = ( n7465 & n22754 ) | ( n7465 & n44353 ) | ( n22754 & n44353 ) ;
  assign n44349 = n11393 ^ n6675 ^ n558 ;
  assign n44350 = n44349 ^ n35671 ^ n12614 ;
  assign n44351 = ( n10345 & ~n15224 ) | ( n10345 & n44350 ) | ( ~n15224 & n44350 ) ;
  assign n44357 = n44356 ^ n44354 ^ n44351 ;
  assign n44358 = n41103 ^ n23730 ^ 1'b0 ;
  assign n44359 = ( ~n4060 & n4093 ) | ( ~n4060 & n12609 ) | ( n4093 & n12609 ) ;
  assign n44360 = n1886 ^ n574 ^ 1'b0 ;
  assign n44361 = ( n25173 & ~n41717 ) | ( n25173 & n44360 ) | ( ~n41717 & n44360 ) ;
  assign n44362 = ( n19408 & ~n22595 ) | ( n19408 & n44361 ) | ( ~n22595 & n44361 ) ;
  assign n44363 = n40833 ^ n36826 ^ n19846 ;
  assign n44364 = ( n1457 & n3990 ) | ( n1457 & ~n44363 ) | ( n3990 & ~n44363 ) ;
  assign n44366 = n883 & n3131 ;
  assign n44367 = ( ~n1828 & n10890 ) | ( ~n1828 & n44366 ) | ( n10890 & n44366 ) ;
  assign n44365 = n14890 & n35827 ;
  assign n44368 = n44367 ^ n44365 ^ n15227 ;
  assign n44369 = n24390 ^ n22012 ^ n11220 ;
  assign n44370 = n44369 ^ n1665 ^ 1'b0 ;
  assign n44371 = n34155 ^ n13794 ^ n697 ;
  assign n44375 = ~n10172 & n19883 ;
  assign n44376 = n18703 & n44375 ;
  assign n44377 = n6227 | n9952 ;
  assign n44378 = n44376 & ~n44377 ;
  assign n44372 = n14232 ^ n12812 ^ n1269 ;
  assign n44373 = ( n1848 & ~n40638 ) | ( n1848 & n44372 ) | ( ~n40638 & n44372 ) ;
  assign n44374 = ( n6946 & ~n28753 ) | ( n6946 & n44373 ) | ( ~n28753 & n44373 ) ;
  assign n44379 = n44378 ^ n44374 ^ n1420 ;
  assign n44380 = n43302 ^ n32764 ^ n27564 ;
  assign n44381 = n19546 | n29486 ;
  assign n44382 = ( n10307 & n11267 ) | ( n10307 & n44381 ) | ( n11267 & n44381 ) ;
  assign n44383 = ( ~n8478 & n23974 ) | ( ~n8478 & n44382 ) | ( n23974 & n44382 ) ;
  assign n44385 = ( ~n2878 & n5129 ) | ( ~n2878 & n43967 ) | ( n5129 & n43967 ) ;
  assign n44384 = ~n7889 & n36247 ;
  assign n44386 = n44385 ^ n44384 ^ 1'b0 ;
  assign n44387 = n10366 & ~n44386 ;
  assign n44388 = n44387 ^ n34769 ^ 1'b0 ;
  assign n44389 = n4351 | n23072 ;
  assign n44390 = ( n5363 & ~n14394 ) | ( n5363 & n14526 ) | ( ~n14394 & n14526 ) ;
  assign n44391 = ( x202 & ~n1384 ) | ( x202 & n44390 ) | ( ~n1384 & n44390 ) ;
  assign n44392 = n44391 ^ n34765 ^ n30300 ;
  assign n44393 = n40502 ^ n35350 ^ n14048 ;
  assign n44400 = ( n19119 & ~n25624 ) | ( n19119 & n28700 ) | ( ~n25624 & n28700 ) ;
  assign n44395 = n20075 ^ n7013 ^ n4692 ;
  assign n44394 = ( n6676 & ~n7609 ) | ( n6676 & n12918 ) | ( ~n7609 & n12918 ) ;
  assign n44396 = n44395 ^ n44394 ^ n18499 ;
  assign n44397 = n17734 ^ n6363 ^ n1871 ;
  assign n44398 = n44397 ^ n17647 ^ 1'b0 ;
  assign n44399 = n44396 & ~n44398 ;
  assign n44401 = n44400 ^ n44399 ^ n23933 ;
  assign n44404 = ( n6394 & ~n8983 ) | ( n6394 & n43655 ) | ( ~n8983 & n43655 ) ;
  assign n44402 = n40256 ^ n17848 ^ 1'b0 ;
  assign n44403 = ~n23944 & n44402 ;
  assign n44405 = n44404 ^ n44403 ^ n20396 ;
  assign n44406 = n43481 ^ n42599 ^ 1'b0 ;
  assign n44407 = n4689 & ~n44406 ;
  assign n44408 = ( n25123 & n34556 ) | ( n25123 & ~n35636 ) | ( n34556 & ~n35636 ) ;
  assign n44409 = n7430 & ~n14927 ;
  assign n44411 = n15191 ^ n11721 ^ n3595 ;
  assign n44410 = n32366 ^ n22330 ^ n5144 ;
  assign n44412 = n44411 ^ n44410 ^ 1'b0 ;
  assign n44413 = ~n44409 & n44412 ;
  assign n44417 = n834 & ~n15699 ;
  assign n44416 = n24381 ^ n22251 ^ n12798 ;
  assign n44414 = n40357 ^ n27323 ^ n20995 ;
  assign n44415 = n44414 ^ n42075 ^ n14205 ;
  assign n44418 = n44417 ^ n44416 ^ n44415 ;
  assign n44419 = n4229 & n34690 ;
  assign n44420 = n44419 ^ n12598 ^ 1'b0 ;
  assign n44421 = ~n15677 & n16121 ;
  assign n44422 = n44421 ^ n17294 ^ 1'b0 ;
  assign n44423 = n11592 & n22170 ;
  assign n44424 = n9217 | n20104 ;
  assign n44425 = n44424 ^ n23537 ^ 1'b0 ;
  assign n44426 = ( n12618 & n15502 ) | ( n12618 & n44425 ) | ( n15502 & n44425 ) ;
  assign n44427 = ( n9593 & n18729 ) | ( n9593 & ~n44426 ) | ( n18729 & ~n44426 ) ;
  assign n44428 = n27144 ^ n1627 ^ 1'b0 ;
  assign n44430 = n9390 | n31552 ;
  assign n44429 = n38429 ^ n9944 ^ n1879 ;
  assign n44431 = n44430 ^ n44429 ^ n31748 ;
  assign n44432 = n6637 | n28162 ;
  assign n44433 = n37606 ^ n22624 ^ n21832 ;
  assign n44434 = ( ~n1655 & n44432 ) | ( ~n1655 & n44433 ) | ( n44432 & n44433 ) ;
  assign n44435 = n33916 ^ n15526 ^ n12840 ;
  assign n44436 = ( n17352 & n29771 ) | ( n17352 & ~n44435 ) | ( n29771 & ~n44435 ) ;
  assign n44437 = n25549 ^ n25308 ^ 1'b0 ;
  assign n44438 = n22058 & ~n44437 ;
  assign n44439 = n20817 ^ n10850 ^ 1'b0 ;
  assign n44440 = ~n10771 & n44439 ;
  assign n44441 = n36357 ^ n31762 ^ n7682 ;
  assign n44442 = n8234 ^ n1258 ^ 1'b0 ;
  assign n44443 = ( n25946 & ~n30317 ) | ( n25946 & n44442 ) | ( ~n30317 & n44442 ) ;
  assign n44444 = ( n3414 & n10439 ) | ( n3414 & ~n37350 ) | ( n10439 & ~n37350 ) ;
  assign n44445 = n38402 ^ n17486 ^ 1'b0 ;
  assign n44446 = ~n2566 & n44445 ;
  assign n44447 = n44446 ^ n42508 ^ n23816 ;
  assign n44448 = n33729 ^ n2033 ^ 1'b0 ;
  assign n44451 = n19965 ^ n1373 ^ 1'b0 ;
  assign n44449 = ~n18946 & n26745 ;
  assign n44450 = n17697 & n44449 ;
  assign n44452 = n44451 ^ n44450 ^ n18291 ;
  assign n44453 = n16448 ^ n13213 ^ n8628 ;
  assign n44454 = n44453 ^ n13528 ^ 1'b0 ;
  assign n44455 = n42647 & ~n44454 ;
  assign n44456 = ( ~x107 & n6394 ) | ( ~x107 & n27013 ) | ( n6394 & n27013 ) ;
  assign n44457 = ( n7844 & n23685 ) | ( n7844 & n44456 ) | ( n23685 & n44456 ) ;
  assign n44458 = ~n6479 & n44457 ;
  assign n44459 = n1717 & ~n7613 ;
  assign n44460 = n44459 ^ n31922 ^ n9088 ;
  assign n44461 = ~n25955 & n44460 ;
  assign n44462 = n44461 ^ n28790 ^ n28628 ;
  assign n44463 = n19349 ^ n13989 ^ n11838 ;
  assign n44464 = n44463 ^ n30651 ^ n17605 ;
  assign n44465 = ( n12429 & ~n35415 ) | ( n12429 & n44464 ) | ( ~n35415 & n44464 ) ;
  assign n44466 = ~n4819 & n28666 ;
  assign n44467 = n44465 & n44466 ;
  assign n44468 = n7378 | n44467 ;
  assign n44469 = n8777 ^ n6591 ^ x151 ;
  assign n44470 = n44469 ^ n40565 ^ n28507 ;
  assign n44471 = n12564 ^ n5106 ^ n4152 ;
  assign n44472 = ( n4191 & n4712 ) | ( n4191 & ~n30406 ) | ( n4712 & ~n30406 ) ;
  assign n44473 = n27564 & ~n39503 ;
  assign n44474 = n20651 ^ n11236 ^ n6175 ;
  assign n44475 = ( n5121 & n5953 ) | ( n5121 & n24898 ) | ( n5953 & n24898 ) ;
  assign n44476 = n15141 ^ n14106 ^ n7345 ;
  assign n44477 = n31145 ^ n22273 ^ n2470 ;
  assign n44478 = ( n42601 & ~n44476 ) | ( n42601 & n44477 ) | ( ~n44476 & n44477 ) ;
  assign n44479 = ( ~n1577 & n3250 ) | ( ~n1577 & n10372 ) | ( n3250 & n10372 ) ;
  assign n44480 = n39116 | n44479 ;
  assign n44481 = n20058 ^ n17707 ^ n9487 ;
  assign n44482 = n30358 ^ n30337 ^ n28121 ;
  assign n44483 = n18932 & n44482 ;
  assign n44484 = n44483 ^ n33829 ^ 1'b0 ;
  assign n44485 = n37598 ^ n30589 ^ n12930 ;
  assign n44486 = n44485 ^ n39870 ^ 1'b0 ;
  assign n44487 = n25012 ^ n4807 ^ 1'b0 ;
  assign n44488 = ( n28645 & n33747 ) | ( n28645 & n34871 ) | ( n33747 & n34871 ) ;
  assign n44489 = ( n1845 & n4779 ) | ( n1845 & ~n5095 ) | ( n4779 & ~n5095 ) ;
  assign n44490 = n17694 & ~n44489 ;
  assign n44491 = n4969 ^ n3642 ^ 1'b0 ;
  assign n44492 = ~n5109 & n20899 ;
  assign n44493 = n44492 ^ n19067 ^ 1'b0 ;
  assign n44494 = n44493 ^ n23159 ^ n14401 ;
  assign n44495 = ( n17488 & ~n27859 ) | ( n17488 & n33104 ) | ( ~n27859 & n33104 ) ;
  assign n44496 = n22264 | n26132 ;
  assign n44497 = n44496 ^ n30421 ^ 1'b0 ;
  assign n44498 = ( n3802 & n18506 ) | ( n3802 & n36499 ) | ( n18506 & n36499 ) ;
  assign n44499 = n3849 ^ n1172 ^ 1'b0 ;
  assign n44500 = ( n11856 & ~n15568 ) | ( n11856 & n44499 ) | ( ~n15568 & n44499 ) ;
  assign n44501 = n44500 ^ n24752 ^ n2197 ;
  assign n44502 = n44264 ^ n27913 ^ n22278 ;
  assign n44503 = ( n34033 & ~n36663 ) | ( n34033 & n44502 ) | ( ~n36663 & n44502 ) ;
  assign n44504 = n1850 & n10222 ;
  assign n44505 = n5654 & n44504 ;
  assign n44506 = ( n6246 & ~n28058 ) | ( n6246 & n44505 ) | ( ~n28058 & n44505 ) ;
  assign n44507 = n44506 ^ n43497 ^ n11497 ;
  assign n44508 = ~n11675 & n19815 ;
  assign n44509 = n4525 & n44508 ;
  assign n44510 = n44509 ^ n16377 ^ 1'b0 ;
  assign n44511 = n18667 & ~n27625 ;
  assign n44512 = ~n35688 & n44511 ;
  assign n44513 = n37495 ^ n28487 ^ n7147 ;
  assign n44514 = n43645 & ~n44513 ;
  assign n44515 = n655 & n4375 ;
  assign n44516 = ( ~n8456 & n44514 ) | ( ~n8456 & n44515 ) | ( n44514 & n44515 ) ;
  assign n44517 = n44516 ^ n43443 ^ n5417 ;
  assign n44518 = ( n6731 & ~n7451 ) | ( n6731 & n12209 ) | ( ~n7451 & n12209 ) ;
  assign n44519 = ( ~n2123 & n15029 ) | ( ~n2123 & n44518 ) | ( n15029 & n44518 ) ;
  assign n44520 = n44519 ^ n23325 ^ n16922 ;
  assign n44521 = ( n34016 & n35860 ) | ( n34016 & n44520 ) | ( n35860 & n44520 ) ;
  assign n44522 = n4945 ^ n4658 ^ 1'b0 ;
  assign n44523 = n10630 & n44522 ;
  assign n44524 = n44523 ^ n15717 ^ 1'b0 ;
  assign n44525 = n27797 ^ n23540 ^ n758 ;
  assign n44526 = n33735 ^ n27457 ^ n24662 ;
  assign n44527 = n9315 | n14040 ;
  assign n44528 = n44527 ^ n42557 ^ n676 ;
  assign n44529 = n44528 ^ n43660 ^ n26371 ;
  assign n44530 = n38831 ^ n32039 ^ 1'b0 ;
  assign n44531 = n15186 & n44530 ;
  assign n44532 = n1987 & n3176 ;
  assign n44533 = n905 & n44532 ;
  assign n44534 = n31955 ^ n9712 ^ n7594 ;
  assign n44535 = ( ~n16725 & n44533 ) | ( ~n16725 & n44534 ) | ( n44533 & n44534 ) ;
  assign n44536 = n44535 ^ n38744 ^ 1'b0 ;
  assign n44537 = n40507 ^ n28933 ^ n17767 ;
  assign n44538 = n19108 ^ n11198 ^ 1'b0 ;
  assign n44539 = n26647 | n44538 ;
  assign n44540 = n19660 ^ n11055 ^ n1870 ;
  assign n44541 = ( n6455 & n14110 ) | ( n6455 & n30869 ) | ( n14110 & n30869 ) ;
  assign n44542 = n27220 ^ n4805 ^ n1177 ;
  assign n44543 = n44542 ^ n23017 ^ n8645 ;
  assign n44544 = ( ~n1473 & n19396 ) | ( ~n1473 & n34787 ) | ( n19396 & n34787 ) ;
  assign n44545 = ( n21137 & ~n43680 ) | ( n21137 & n44544 ) | ( ~n43680 & n44544 ) ;
  assign n44546 = n36373 ^ n1999 ^ 1'b0 ;
  assign n44547 = n37572 & n44546 ;
  assign n44548 = n44547 ^ n34821 ^ 1'b0 ;
  assign n44549 = n13285 & n44548 ;
  assign n44550 = ~n24327 & n29073 ;
  assign n44551 = n44550 ^ n41740 ^ 1'b0 ;
  assign n44552 = ( n794 & n22602 ) | ( n794 & n34179 ) | ( n22602 & n34179 ) ;
  assign n44553 = n32342 ^ n29357 ^ 1'b0 ;
  assign n44554 = n44552 | n44553 ;
  assign n44555 = ~n18441 & n27964 ;
  assign n44556 = ~n22797 & n44555 ;
  assign n44557 = n5285 ^ n2977 ^ n961 ;
  assign n44558 = n44557 ^ n38194 ^ n11189 ;
  assign n44559 = ( n2012 & n13023 ) | ( n2012 & n44558 ) | ( n13023 & n44558 ) ;
  assign n44560 = ~n15659 & n18403 ;
  assign n44561 = n39612 ^ n6048 ^ n969 ;
  assign n44562 = ( n1037 & ~n44560 ) | ( n1037 & n44561 ) | ( ~n44560 & n44561 ) ;
  assign n44563 = ~n1146 & n21155 ;
  assign n44564 = n44563 ^ n23035 ^ 1'b0 ;
  assign n44565 = ( n600 & n8593 ) | ( n600 & ~n23364 ) | ( n8593 & ~n23364 ) ;
  assign n44566 = n44565 ^ n4009 ^ 1'b0 ;
  assign n44567 = ~n10736 & n44566 ;
  assign n44568 = n44567 ^ n23628 ^ n21664 ;
  assign n44569 = n32521 ^ n11629 ^ n626 ;
  assign n44570 = ( n6872 & n10894 ) | ( n6872 & ~n14594 ) | ( n10894 & ~n14594 ) ;
  assign n44571 = ( n10498 & ~n10862 ) | ( n10498 & n44570 ) | ( ~n10862 & n44570 ) ;
  assign n44572 = n6960 & ~n44571 ;
  assign n44573 = ~n531 & n44572 ;
  assign n44574 = ( n19355 & n44569 ) | ( n19355 & ~n44573 ) | ( n44569 & ~n44573 ) ;
  assign n44575 = n37023 ^ n14355 ^ n6612 ;
  assign n44576 = n44575 ^ n18840 ^ n6972 ;
  assign n44577 = n14350 ^ n12906 ^ 1'b0 ;
  assign n44578 = ~n7125 & n44577 ;
  assign n44579 = n44578 ^ n4264 ^ 1'b0 ;
  assign n44580 = ~n1074 & n44579 ;
  assign n44581 = ( ~n8646 & n8854 ) | ( ~n8646 & n13931 ) | ( n8854 & n13931 ) ;
  assign n44582 = n12848 ^ n2892 ^ 1'b0 ;
  assign n44583 = n44582 ^ n41639 ^ 1'b0 ;
  assign n44584 = ( n2994 & n3367 ) | ( n2994 & ~n21533 ) | ( n3367 & ~n21533 ) ;
  assign n44585 = ( n9048 & ~n18167 ) | ( n9048 & n44584 ) | ( ~n18167 & n44584 ) ;
  assign n44586 = n28711 | n31016 ;
  assign n44587 = ( n8201 & n44585 ) | ( n8201 & ~n44586 ) | ( n44585 & ~n44586 ) ;
  assign n44588 = n21712 & n41462 ;
  assign n44589 = n298 | n22157 ;
  assign n44590 = n26766 & ~n44589 ;
  assign n44591 = n44590 ^ n40007 ^ 1'b0 ;
  assign n44592 = n1418 & n25756 ;
  assign n44593 = n44592 ^ n5906 ^ 1'b0 ;
  assign n44594 = n40258 ^ n36027 ^ 1'b0 ;
  assign n44595 = n44593 & ~n44594 ;
  assign n44596 = n22787 ^ n19379 ^ 1'b0 ;
  assign n44597 = n44596 ^ n22655 ^ n18014 ;
  assign n44598 = ( n4399 & ~n20157 ) | ( n4399 & n44597 ) | ( ~n20157 & n44597 ) ;
  assign n44599 = n44598 ^ n32819 ^ n8265 ;
  assign n44600 = n10802 & n22025 ;
  assign n44601 = ( n21634 & n40948 ) | ( n21634 & n44600 ) | ( n40948 & n44600 ) ;
  assign n44602 = ( n17172 & n27182 ) | ( n17172 & ~n34297 ) | ( n27182 & ~n34297 ) ;
  assign n44603 = n22962 ^ n11790 ^ n9337 ;
  assign n44604 = ( ~n2778 & n31360 ) | ( ~n2778 & n44603 ) | ( n31360 & n44603 ) ;
  assign n44605 = n34076 ^ n9016 ^ 1'b0 ;
  assign n44606 = n11642 ^ n5442 ^ 1'b0 ;
  assign n44607 = n44606 ^ n23248 ^ n22408 ;
  assign n44608 = n10437 ^ n6481 ^ n1098 ;
  assign n44609 = ( n4628 & n19732 ) | ( n4628 & ~n44608 ) | ( n19732 & ~n44608 ) ;
  assign n44610 = ( n2108 & ~n16028 ) | ( n2108 & n36977 ) | ( ~n16028 & n36977 ) ;
  assign n44611 = n42381 ^ n21543 ^ n13578 ;
  assign n44612 = ( ~n14240 & n24039 ) | ( ~n14240 & n40409 ) | ( n24039 & n40409 ) ;
  assign n44613 = n599 | n29861 ;
  assign n44614 = n37938 | n44613 ;
  assign n44615 = n44614 ^ n4471 ^ 1'b0 ;
  assign n44616 = ( ~n2884 & n6048 ) | ( ~n2884 & n18188 ) | ( n6048 & n18188 ) ;
  assign n44617 = ( n26672 & n34274 ) | ( n26672 & n39026 ) | ( n34274 & n39026 ) ;
  assign n44618 = ( n13687 & n44616 ) | ( n13687 & n44617 ) | ( n44616 & n44617 ) ;
  assign n44619 = ~n30019 & n44618 ;
  assign n44620 = n2967 & ~n23754 ;
  assign n44621 = ~n28323 & n44620 ;
  assign n44622 = ~n725 & n44621 ;
  assign n44623 = n12263 ^ n2305 ^ 1'b0 ;
  assign n44624 = ( n10550 & n41692 ) | ( n10550 & ~n44623 ) | ( n41692 & ~n44623 ) ;
  assign n44625 = n44624 ^ n422 ^ 1'b0 ;
  assign n44626 = ~n34205 & n44625 ;
  assign n44627 = n1241 & ~n12610 ;
  assign n44628 = n18718 & n44627 ;
  assign n44629 = ~n36296 & n44628 ;
  assign n44630 = ( n35831 & ~n43027 ) | ( n35831 & n44629 ) | ( ~n43027 & n44629 ) ;
  assign n44631 = n20797 & n22259 ;
  assign n44632 = n14804 & n44631 ;
  assign n44633 = n44632 ^ n20519 ^ n12560 ;
  assign n44634 = n21558 ^ n20126 ^ 1'b0 ;
  assign n44635 = ~n3953 & n25832 ;
  assign n44636 = ( ~n6798 & n10404 ) | ( ~n6798 & n44635 ) | ( n10404 & n44635 ) ;
  assign n44637 = ( n18285 & n44634 ) | ( n18285 & n44636 ) | ( n44634 & n44636 ) ;
  assign n44638 = n5581 & ~n35063 ;
  assign n44639 = n44638 ^ n21382 ^ 1'b0 ;
  assign n44640 = n5133 ^ n2839 ^ n1323 ;
  assign n44641 = n44640 ^ n15034 ^ n4023 ;
  assign n44642 = n44641 ^ n14045 ^ n5608 ;
  assign n44643 = ( n4890 & ~n44639 ) | ( n4890 & n44642 ) | ( ~n44639 & n44642 ) ;
  assign n44644 = n33365 ^ n5006 ^ 1'b0 ;
  assign n44645 = n44644 ^ n29926 ^ 1'b0 ;
  assign n44646 = n14719 ^ n12844 ^ n11080 ;
  assign n44647 = n44646 ^ n29835 ^ 1'b0 ;
  assign n44648 = n44647 ^ n31503 ^ 1'b0 ;
  assign n44649 = n15338 ^ n12922 ^ n3225 ;
  assign n44650 = n44649 ^ n9178 ^ 1'b0 ;
  assign n44651 = n44648 | n44650 ;
  assign n44652 = n15956 ^ n3104 ^ 1'b0 ;
  assign n44653 = x166 & ~n1595 ;
  assign n44654 = n44653 ^ n31722 ^ 1'b0 ;
  assign n44657 = n25350 ^ n14150 ^ n4469 ;
  assign n44658 = n44657 ^ n25769 ^ 1'b0 ;
  assign n44655 = ~n7108 & n26767 ;
  assign n44656 = n44655 ^ n30827 ^ 1'b0 ;
  assign n44659 = n44658 ^ n44656 ^ n41907 ;
  assign n44660 = ( ~n32342 & n44654 ) | ( ~n32342 & n44659 ) | ( n44654 & n44659 ) ;
  assign n44661 = ( n3952 & ~n4371 ) | ( n3952 & n12370 ) | ( ~n4371 & n12370 ) ;
  assign n44662 = n5353 ^ n2889 ^ n943 ;
  assign n44663 = n44662 ^ n6521 ^ n2016 ;
  assign n44664 = n44663 ^ n39211 ^ n16770 ;
  assign n44665 = n9376 ^ n1686 ^ 1'b0 ;
  assign n44666 = ( ~n15997 & n35833 ) | ( ~n15997 & n44665 ) | ( n35833 & n44665 ) ;
  assign n44667 = n44666 ^ n18710 ^ n17103 ;
  assign n44668 = n40343 ^ n25961 ^ n3973 ;
  assign n44669 = n34833 ^ n32591 ^ n9546 ;
  assign n44670 = n7098 & n44669 ;
  assign n44671 = n44670 ^ n15046 ^ 1'b0 ;
  assign n44672 = n44671 ^ n26911 ^ n8321 ;
  assign n44673 = n41809 ^ n21269 ^ 1'b0 ;
  assign n44674 = n988 & n44673 ;
  assign n44675 = n29566 ^ n16940 ^ 1'b0 ;
  assign n44676 = n8155 & n44675 ;
  assign n44677 = ( ~n4419 & n8100 ) | ( ~n4419 & n14712 ) | ( n8100 & n14712 ) ;
  assign n44678 = ( ~x4 & n13460 ) | ( ~x4 & n44677 ) | ( n13460 & n44677 ) ;
  assign n44679 = ( n14232 & ~n16777 ) | ( n14232 & n24769 ) | ( ~n16777 & n24769 ) ;
  assign n44683 = n33843 ^ n19164 ^ n16989 ;
  assign n44680 = n14538 & n21579 ;
  assign n44681 = ~n13457 & n44680 ;
  assign n44682 = ( n22067 & n28918 ) | ( n22067 & n44681 ) | ( n28918 & n44681 ) ;
  assign n44684 = n44683 ^ n44682 ^ n13020 ;
  assign n44686 = n7857 ^ n5165 ^ 1'b0 ;
  assign n44685 = n29285 ^ n15531 ^ n7390 ;
  assign n44687 = n44686 ^ n44685 ^ n15322 ;
  assign n44688 = ( ~x247 & n5194 ) | ( ~x247 & n17100 ) | ( n5194 & n17100 ) ;
  assign n44689 = ( ~x67 & n3430 ) | ( ~x67 & n44688 ) | ( n3430 & n44688 ) ;
  assign n44690 = n44689 ^ n28193 ^ n10823 ;
  assign n44691 = n11037 ^ n2465 ^ 1'b0 ;
  assign n44692 = n44691 ^ n25520 ^ n3251 ;
  assign n44693 = n4424 & n22617 ;
  assign n44694 = n44693 ^ x107 ^ 1'b0 ;
  assign n44695 = ~n6067 & n24270 ;
  assign n44696 = n27468 | n44695 ;
  assign n44697 = n44696 ^ n27145 ^ 1'b0 ;
  assign n44698 = ~n23099 & n44697 ;
  assign n44699 = n41025 ^ n19354 ^ n7798 ;
  assign n44700 = ~n14511 & n16515 ;
  assign n44701 = ( n1901 & ~n4219 ) | ( n1901 & n17743 ) | ( ~n4219 & n17743 ) ;
  assign n44702 = n14359 ^ n11071 ^ n1931 ;
  assign n44703 = ( n44700 & ~n44701 ) | ( n44700 & n44702 ) | ( ~n44701 & n44702 ) ;
  assign n44704 = n21327 ^ n19425 ^ 1'b0 ;
  assign n44705 = ( n3726 & n13423 ) | ( n3726 & ~n26051 ) | ( n13423 & ~n26051 ) ;
  assign n44706 = ~n1748 & n44705 ;
  assign n44707 = n44706 ^ n17857 ^ 1'b0 ;
  assign n44708 = ( n35333 & ~n44704 ) | ( n35333 & n44707 ) | ( ~n44704 & n44707 ) ;
  assign n44709 = n14376 ^ n12796 ^ n3708 ;
  assign n44710 = n19552 ^ n15224 ^ n11840 ;
  assign n44711 = ( n2208 & ~n9681 ) | ( n2208 & n44710 ) | ( ~n9681 & n44710 ) ;
  assign n44712 = ~n10504 & n44711 ;
  assign n44713 = ( n24897 & n44709 ) | ( n24897 & ~n44712 ) | ( n44709 & ~n44712 ) ;
  assign n44714 = n13562 & ~n37218 ;
  assign n44715 = n3294 | n27600 ;
  assign n44716 = n15251 & ~n44715 ;
  assign n44717 = n41154 | n44716 ;
  assign n44718 = n29182 | n44717 ;
  assign n44719 = n38567 ^ n18785 ^ n11634 ;
  assign n44720 = n28443 & ~n29681 ;
  assign n44721 = n44720 ^ n32926 ^ n1280 ;
  assign n44722 = ( n8895 & n20396 ) | ( n8895 & n38026 ) | ( n20396 & n38026 ) ;
  assign n44723 = n39418 ^ n17404 ^ n15415 ;
  assign n44724 = ~n15507 & n17976 ;
  assign n44725 = n7153 ^ n2164 ^ 1'b0 ;
  assign n44726 = n10085 & ~n21510 ;
  assign n44727 = n7435 & n44726 ;
  assign n44728 = n3445 & n23161 ;
  assign n44729 = ~n5204 & n44728 ;
  assign n44730 = n44729 ^ n30470 ^ 1'b0 ;
  assign n44731 = n25016 ^ n4603 ^ 1'b0 ;
  assign n44732 = n44730 & ~n44731 ;
  assign n44733 = n4017 & n19198 ;
  assign n44734 = n41639 & n44733 ;
  assign n44735 = n18432 ^ n18073 ^ n6342 ;
  assign n44736 = ( n2198 & n16538 ) | ( n2198 & n44735 ) | ( n16538 & n44735 ) ;
  assign n44737 = ( n4886 & n23318 ) | ( n4886 & n35441 ) | ( n23318 & n35441 ) ;
  assign n44738 = ( n12858 & n16621 ) | ( n12858 & ~n44737 ) | ( n16621 & ~n44737 ) ;
  assign n44739 = n25077 ^ n24161 ^ 1'b0 ;
  assign n44740 = n44739 ^ n25778 ^ n7053 ;
  assign n44741 = ( n9952 & n12762 ) | ( n9952 & n21061 ) | ( n12762 & n21061 ) ;
  assign n44742 = n35518 ^ n13866 ^ n9366 ;
  assign n44743 = n14424 & ~n44742 ;
  assign n44744 = ~n12320 & n21667 ;
  assign n44745 = ( n44741 & n44743 ) | ( n44741 & n44744 ) | ( n44743 & n44744 ) ;
  assign n44746 = n23549 ^ n15491 ^ n13077 ;
  assign n44747 = n14438 | n30096 ;
  assign n44748 = n44747 ^ n42324 ^ 1'b0 ;
  assign n44749 = ( ~n1740 & n15592 ) | ( ~n1740 & n44748 ) | ( n15592 & n44748 ) ;
  assign n44750 = ( ~n6237 & n6742 ) | ( ~n6237 & n12876 ) | ( n6742 & n12876 ) ;
  assign n44751 = n2958 | n16596 ;
  assign n44752 = n8255 | n44751 ;
  assign n44753 = n43569 & ~n44752 ;
  assign n44754 = ( n27749 & ~n44750 ) | ( n27749 & n44753 ) | ( ~n44750 & n44753 ) ;
  assign n44755 = n8284 | n20691 ;
  assign n44756 = n44755 ^ n28854 ^ 1'b0 ;
  assign n44757 = n23873 & n31358 ;
  assign n44758 = ~n44159 & n44757 ;
  assign n44759 = n24356 ^ n13209 ^ n11340 ;
  assign n44760 = n25219 ^ n21543 ^ n6883 ;
  assign n44761 = n44760 ^ n29285 ^ 1'b0 ;
  assign n44762 = ( n43058 & ~n44759 ) | ( n43058 & n44761 ) | ( ~n44759 & n44761 ) ;
  assign n44763 = n26001 ^ n19437 ^ n8169 ;
  assign n44764 = ( n7346 & ~n22819 ) | ( n7346 & n44763 ) | ( ~n22819 & n44763 ) ;
  assign n44765 = ( n594 & ~n29893 ) | ( n594 & n34569 ) | ( ~n29893 & n34569 ) ;
  assign n44766 = n20345 ^ n15911 ^ 1'b0 ;
  assign n44767 = ( ~n1502 & n17189 ) | ( ~n1502 & n26911 ) | ( n17189 & n26911 ) ;
  assign n44770 = ( n772 & n18680 ) | ( n772 & n22642 ) | ( n18680 & n22642 ) ;
  assign n44768 = n3681 & ~n5197 ;
  assign n44769 = n44768 ^ n44385 ^ n19826 ;
  assign n44771 = n44770 ^ n44769 ^ 1'b0 ;
  assign n44772 = n11287 & ~n44771 ;
  assign n44773 = n10101 ^ n3989 ^ n1555 ;
  assign n44774 = n15992 & n19287 ;
  assign n44775 = ~n44773 & n44774 ;
  assign n44776 = n8687 | n37119 ;
  assign n44777 = n44776 ^ n13489 ^ 1'b0 ;
  assign n44778 = ( n14584 & n18772 ) | ( n14584 & n23332 ) | ( n18772 & n23332 ) ;
  assign n44779 = ( ~n28917 & n30121 ) | ( ~n28917 & n44778 ) | ( n30121 & n44778 ) ;
  assign n44780 = n44779 ^ n18685 ^ n7618 ;
  assign n44781 = n4555 | n35411 ;
  assign n44782 = n44781 ^ n40940 ^ 1'b0 ;
  assign n44784 = n4801 ^ n1582 ^ 1'b0 ;
  assign n44783 = n44432 ^ n34818 ^ n834 ;
  assign n44785 = n44784 ^ n44783 ^ n10933 ;
  assign n44786 = ( ~n5693 & n17499 ) | ( ~n5693 & n20283 ) | ( n17499 & n20283 ) ;
  assign n44787 = ( n2638 & n27650 ) | ( n2638 & ~n44786 ) | ( n27650 & ~n44786 ) ;
  assign n44788 = n30893 ^ n17196 ^ n6085 ;
  assign n44789 = n7036 ^ n1976 ^ 1'b0 ;
  assign n44790 = n24537 & n44789 ;
  assign n44791 = n30906 ^ n22503 ^ 1'b0 ;
  assign n44792 = n13891 ^ n7039 ^ 1'b0 ;
  assign n44793 = n26789 | n44792 ;
  assign n44794 = n2941 & n44793 ;
  assign n44795 = ( n3170 & n36826 ) | ( n3170 & ~n44794 ) | ( n36826 & ~n44794 ) ;
  assign n44796 = n44795 ^ n41705 ^ n32692 ;
  assign n44797 = n44796 ^ n337 ^ 1'b0 ;
  assign n44798 = n42124 ^ n18722 ^ 1'b0 ;
  assign n44799 = n40992 ^ n15556 ^ 1'b0 ;
  assign n44803 = n16654 ^ n10380 ^ n8902 ;
  assign n44800 = n14673 | n23233 ;
  assign n44801 = n24600 | n44800 ;
  assign n44802 = n44801 ^ n34600 ^ n15291 ;
  assign n44804 = n44803 ^ n44802 ^ n16585 ;
  assign n44805 = ( n6404 & n6474 ) | ( n6404 & n11497 ) | ( n6474 & n11497 ) ;
  assign n44806 = ( n23416 & n42261 ) | ( n23416 & n44805 ) | ( n42261 & n44805 ) ;
  assign n44807 = n44806 ^ n19491 ^ n17534 ;
  assign n44808 = ( ~n22807 & n33656 ) | ( ~n22807 & n43067 ) | ( n33656 & n43067 ) ;
  assign n44809 = n27330 ^ n20167 ^ n6235 ;
  assign n44810 = n6494 | n36086 ;
  assign n44811 = n10346 ^ n3630 ^ n699 ;
  assign n44812 = n44811 ^ n27090 ^ n26340 ;
  assign n44813 = n36631 ^ n32333 ^ 1'b0 ;
  assign n44814 = ~n44812 & n44813 ;
  assign n44817 = ~n313 & n2125 ;
  assign n44818 = n44817 ^ n35733 ^ 1'b0 ;
  assign n44815 = n7414 | n17332 ;
  assign n44816 = n20774 | n44815 ;
  assign n44819 = n44818 ^ n44816 ^ 1'b0 ;
  assign n44820 = ( n8117 & n19870 ) | ( n8117 & ~n44819 ) | ( n19870 & ~n44819 ) ;
  assign n44821 = n28367 ^ n26846 ^ n18694 ;
  assign n44822 = ( n11545 & ~n30163 ) | ( n11545 & n39695 ) | ( ~n30163 & n39695 ) ;
  assign n44823 = n11505 & ~n35725 ;
  assign n44824 = n44823 ^ n21900 ^ n20945 ;
  assign n44825 = ( n13798 & n16911 ) | ( n13798 & ~n41452 ) | ( n16911 & ~n41452 ) ;
  assign n44826 = n44048 ^ n19502 ^ n12105 ;
  assign n44827 = ( n31236 & n44825 ) | ( n31236 & n44826 ) | ( n44825 & n44826 ) ;
  assign n44828 = n44827 ^ n44406 ^ 1'b0 ;
  assign n44831 = n36608 ^ n31016 ^ n7151 ;
  assign n44832 = n44831 ^ n40505 ^ n25423 ;
  assign n44829 = ( n1641 & ~n2685 ) | ( n1641 & n5010 ) | ( ~n2685 & n5010 ) ;
  assign n44830 = n18154 | n44829 ;
  assign n44833 = n44832 ^ n44830 ^ 1'b0 ;
  assign n44834 = n26281 ^ n22013 ^ n6427 ;
  assign n44835 = n32367 & ~n44834 ;
  assign n44836 = n36781 ^ n7275 ^ 1'b0 ;
  assign n44837 = n6503 & n44836 ;
  assign n44838 = ( ~x227 & n10609 ) | ( ~x227 & n29378 ) | ( n10609 & n29378 ) ;
  assign n44839 = n44838 ^ n18996 ^ n17770 ;
  assign n44840 = n40133 ^ n29964 ^ 1'b0 ;
  assign n44841 = n16310 ^ n14046 ^ n13380 ;
  assign n44842 = n42616 ^ n38479 ^ n22498 ;
  assign n44843 = ( n11084 & n15145 ) | ( n11084 & ~n18549 ) | ( n15145 & ~n18549 ) ;
  assign n44844 = n44843 ^ n5332 ^ 1'b0 ;
  assign n44845 = ( n7284 & ~n44842 ) | ( n7284 & n44844 ) | ( ~n44842 & n44844 ) ;
  assign n44846 = ( n16558 & ~n22532 ) | ( n16558 & n26196 ) | ( ~n22532 & n26196 ) ;
  assign n44847 = n44846 ^ n22339 ^ n13071 ;
  assign n44848 = n44847 ^ n19679 ^ n9843 ;
  assign n44852 = n13660 ^ n8095 ^ 1'b0 ;
  assign n44851 = ( ~n10784 & n34127 ) | ( ~n10784 & n40018 ) | ( n34127 & n40018 ) ;
  assign n44853 = n44852 ^ n44851 ^ 1'b0 ;
  assign n44854 = n44853 ^ n11308 ^ 1'b0 ;
  assign n44855 = n14270 & n44854 ;
  assign n44849 = n8676 & n14651 ;
  assign n44850 = n44849 ^ n1612 ^ 1'b0 ;
  assign n44856 = n44855 ^ n44850 ^ n8887 ;
  assign n44857 = n41040 ^ n39459 ^ n18907 ;
  assign n44858 = n5123 & n6537 ;
  assign n44859 = n44857 & n44858 ;
  assign n44860 = n10245 & n26727 ;
  assign n44861 = n44860 ^ n10841 ^ 1'b0 ;
  assign n44863 = n15330 ^ n7705 ^ 1'b0 ;
  assign n44864 = n36417 & n44863 ;
  assign n44865 = ( x52 & n16421 ) | ( x52 & n44864 ) | ( n16421 & n44864 ) ;
  assign n44862 = ~n599 & n20738 ;
  assign n44866 = n44865 ^ n44862 ^ 1'b0 ;
  assign n44867 = ( n7570 & ~n8515 ) | ( n7570 & n39239 ) | ( ~n8515 & n39239 ) ;
  assign n44868 = n31785 ^ n15857 ^ 1'b0 ;
  assign n44869 = n44584 ^ n20508 ^ n834 ;
  assign n44870 = n44869 ^ n39213 ^ n7178 ;
  assign n44871 = n22156 ^ n20853 ^ 1'b0 ;
  assign n44872 = n8893 & ~n44871 ;
  assign n44873 = ( n13206 & ~n38307 ) | ( n13206 & n44872 ) | ( ~n38307 & n44872 ) ;
  assign n44874 = ( ~n4567 & n25222 ) | ( ~n4567 & n33248 ) | ( n25222 & n33248 ) ;
  assign n44875 = n43869 ^ n32927 ^ 1'b0 ;
  assign n44876 = n27368 ^ n5627 ^ 1'b0 ;
  assign n44877 = n38850 & ~n44876 ;
  assign n44880 = ( n5275 & n8191 ) | ( n5275 & ~n31760 ) | ( n8191 & ~n31760 ) ;
  assign n44881 = ( n3878 & n14712 ) | ( n3878 & n44880 ) | ( n14712 & n44880 ) ;
  assign n44878 = n2998 & n10038 ;
  assign n44879 = n7822 | n44878 ;
  assign n44882 = n44881 ^ n44879 ^ n6724 ;
  assign n44883 = n15296 | n16543 ;
  assign n44884 = n44882 | n44883 ;
  assign n44885 = n30651 ^ n29038 ^ n24312 ;
  assign n44886 = ( n6892 & ~n14727 ) | ( n6892 & n18735 ) | ( ~n14727 & n18735 ) ;
  assign n44887 = n44886 ^ n11726 ^ n6801 ;
  assign n44888 = n7482 | n25378 ;
  assign n44889 = n44888 ^ n21368 ^ 1'b0 ;
  assign n44890 = ( n19715 & n31587 ) | ( n19715 & ~n44889 ) | ( n31587 & ~n44889 ) ;
  assign n44891 = ( ~n18101 & n28042 ) | ( ~n18101 & n43641 ) | ( n28042 & n43641 ) ;
  assign n44892 = n11232 ^ n6029 ^ 1'b0 ;
  assign n44893 = n15658 & ~n44892 ;
  assign n44894 = n44893 ^ n27242 ^ n26831 ;
  assign n44895 = x194 & n31598 ;
  assign n44896 = n31593 ^ n24492 ^ n14078 ;
  assign n44897 = n44896 ^ n38895 ^ n29364 ;
  assign n44899 = n42926 ^ n20113 ^ n7013 ;
  assign n44898 = ( ~n5109 & n8099 ) | ( ~n5109 & n14512 ) | ( n8099 & n14512 ) ;
  assign n44900 = n44899 ^ n44898 ^ n17526 ;
  assign n44901 = n40266 ^ n26798 ^ n4787 ;
  assign n44902 = n44901 ^ n44417 ^ n23708 ;
  assign n44903 = n41279 & n44902 ;
  assign n44904 = ~n2224 & n10342 ;
  assign n44905 = n44904 ^ n20212 ^ 1'b0 ;
  assign n44906 = ( n7299 & ~n12949 ) | ( n7299 & n20673 ) | ( ~n12949 & n20673 ) ;
  assign n44907 = ( n26954 & n34274 ) | ( n26954 & n44906 ) | ( n34274 & n44906 ) ;
  assign n44908 = ( n5632 & ~n9162 ) | ( n5632 & n9295 ) | ( ~n9162 & n9295 ) ;
  assign n44909 = n39196 ^ n28644 ^ 1'b0 ;
  assign n44910 = ~n38000 & n44909 ;
  assign n44911 = ( n28547 & ~n44908 ) | ( n28547 & n44910 ) | ( ~n44908 & n44910 ) ;
  assign n44912 = ( n44905 & ~n44907 ) | ( n44905 & n44911 ) | ( ~n44907 & n44911 ) ;
  assign n44913 = ~n6523 & n8365 ;
  assign n44914 = n44913 ^ n16256 ^ 1'b0 ;
  assign n44915 = n621 | n44914 ;
  assign n44916 = n19993 & ~n23698 ;
  assign n44917 = n44916 ^ n8522 ^ n1365 ;
  assign n44918 = ~n8152 & n13555 ;
  assign n44919 = n4693 & n44918 ;
  assign n44920 = ~n3697 & n31928 ;
  assign n44921 = n26513 ^ n14883 ^ 1'b0 ;
  assign n44922 = n44920 & ~n44921 ;
  assign n44923 = ~n9017 & n27766 ;
  assign n44924 = ~n44922 & n44923 ;
  assign n44925 = n25643 ^ x230 ^ 1'b0 ;
  assign n44926 = n35188 | n44925 ;
  assign n44927 = n24365 & n28721 ;
  assign n44928 = ~n5511 & n9747 ;
  assign n44929 = n44928 ^ n25482 ^ 1'b0 ;
  assign n44930 = ( ~n34496 & n40036 ) | ( ~n34496 & n44929 ) | ( n40036 & n44929 ) ;
  assign n44931 = n26778 ^ n17677 ^ n14000 ;
  assign n44932 = ( n16507 & ~n44930 ) | ( n16507 & n44931 ) | ( ~n44930 & n44931 ) ;
  assign n44933 = n20924 & n31482 ;
  assign n44934 = n44933 ^ n23498 ^ 1'b0 ;
  assign n44935 = n44934 ^ n23565 ^ n6903 ;
  assign n44936 = ( n24693 & n27407 ) | ( n24693 & n44935 ) | ( n27407 & n44935 ) ;
  assign n44937 = n23460 ^ n13744 ^ 1'b0 ;
  assign n44938 = ~n482 & n7004 ;
  assign n44939 = n14722 & n44938 ;
  assign n44940 = n24043 & ~n44939 ;
  assign n44941 = ( ~n1130 & n36491 ) | ( ~n1130 & n44940 ) | ( n36491 & n44940 ) ;
  assign n44942 = n9492 & n11383 ;
  assign n44943 = ( ~n690 & n42640 ) | ( ~n690 & n44942 ) | ( n42640 & n44942 ) ;
  assign n44944 = n35725 ^ n27037 ^ n14817 ;
  assign n44945 = n2311 | n44944 ;
  assign n44946 = n44945 ^ n13990 ^ 1'b0 ;
  assign n44947 = n35352 & ~n41498 ;
  assign n44948 = ( n6503 & ~n8081 ) | ( n6503 & n18708 ) | ( ~n8081 & n18708 ) ;
  assign n44949 = n36255 ^ n17965 ^ n16621 ;
  assign n44950 = n44949 ^ n31226 ^ n1703 ;
  assign n44955 = n6975 & ~n10369 ;
  assign n44956 = n8750 & n44955 ;
  assign n44951 = n8184 ^ n4649 ^ 1'b0 ;
  assign n44952 = ~n19240 & n44951 ;
  assign n44953 = n16343 ^ n14635 ^ 1'b0 ;
  assign n44954 = ( ~n32238 & n44952 ) | ( ~n32238 & n44953 ) | ( n44952 & n44953 ) ;
  assign n44957 = n44956 ^ n44954 ^ n11470 ;
  assign n44958 = n40644 ^ n19863 ^ n4003 ;
  assign n44959 = n32751 ^ n12067 ^ n5630 ;
  assign n44960 = n1605 & n3180 ;
  assign n44961 = n44960 ^ n14700 ^ 1'b0 ;
  assign n44962 = n9486 ^ n4630 ^ 1'b0 ;
  assign n44963 = ~n9484 & n44962 ;
  assign n44965 = n8711 | n37745 ;
  assign n44966 = ( n20221 & n40452 ) | ( n20221 & ~n44965 ) | ( n40452 & ~n44965 ) ;
  assign n44964 = n706 & n4369 ;
  assign n44967 = n44966 ^ n44964 ^ x96 ;
  assign n44968 = n39914 ^ n16897 ^ n10271 ;
  assign n44969 = n44968 ^ n3092 ^ 1'b0 ;
  assign n44970 = n1574 & n44969 ;
  assign n44971 = n35294 ^ n13149 ^ x176 ;
  assign n44972 = ( n3733 & n19579 ) | ( n3733 & n44971 ) | ( n19579 & n44971 ) ;
  assign n44973 = n44972 ^ n30647 ^ 1'b0 ;
  assign n44974 = ( ~n23780 & n24072 ) | ( ~n23780 & n33728 ) | ( n24072 & n33728 ) ;
  assign n44975 = ( n13789 & n22344 ) | ( n13789 & ~n33937 ) | ( n22344 & ~n33937 ) ;
  assign n44976 = ( ~n16027 & n26531 ) | ( ~n16027 & n31929 ) | ( n26531 & n31929 ) ;
  assign n44977 = ( ~n23542 & n44975 ) | ( ~n23542 & n44976 ) | ( n44975 & n44976 ) ;
  assign n44978 = n24910 ^ n8504 ^ 1'b0 ;
  assign n44979 = n28983 ^ n23267 ^ n21750 ;
  assign n44980 = ( ~x10 & n25391 ) | ( ~x10 & n43066 ) | ( n25391 & n43066 ) ;
  assign n44981 = ( n1207 & n6029 ) | ( n1207 & n44980 ) | ( n6029 & n44980 ) ;
  assign n44982 = n44981 ^ n32849 ^ 1'b0 ;
  assign n44983 = n44979 & n44982 ;
  assign n44984 = ( ~n21822 & n22865 ) | ( ~n21822 & n27921 ) | ( n22865 & n27921 ) ;
  assign n44985 = n44984 ^ n29075 ^ n20861 ;
  assign n44986 = ( n11989 & n16702 ) | ( n11989 & n21326 ) | ( n16702 & n21326 ) ;
  assign n44987 = n38757 & n44986 ;
  assign n44988 = ( n15573 & ~n25772 ) | ( n15573 & n26882 ) | ( ~n25772 & n26882 ) ;
  assign n44989 = n44988 ^ n43168 ^ n25962 ;
  assign n44990 = n44989 ^ n42255 ^ n34592 ;
  assign n44991 = ( n11614 & n44987 ) | ( n11614 & ~n44990 ) | ( n44987 & ~n44990 ) ;
  assign n44992 = n44991 ^ n13341 ^ n337 ;
  assign n44993 = n1070 & n2618 ;
  assign n44994 = n44993 ^ n31455 ^ 1'b0 ;
  assign n44995 = n44994 ^ n8109 ^ 1'b0 ;
  assign n44996 = n31089 ^ n17111 ^ n13988 ;
  assign n44997 = n41673 ^ n11089 ^ 1'b0 ;
  assign n44998 = ~n19834 & n26835 ;
  assign n45003 = n15574 ^ n781 ^ 1'b0 ;
  assign n45004 = n1162 & n45003 ;
  assign n44999 = ( ~n766 & n2828 ) | ( ~n766 & n5830 ) | ( n2828 & n5830 ) ;
  assign n45000 = ( n9983 & ~n39914 ) | ( n9983 & n44999 ) | ( ~n39914 & n44999 ) ;
  assign n45001 = ( n23383 & n41232 ) | ( n23383 & n45000 ) | ( n41232 & n45000 ) ;
  assign n45002 = ( n16004 & ~n32120 ) | ( n16004 & n45001 ) | ( ~n32120 & n45001 ) ;
  assign n45005 = n45004 ^ n45002 ^ 1'b0 ;
  assign n45006 = n27523 | n45005 ;
  assign n45007 = n25422 ^ n13213 ^ n7440 ;
  assign n45008 = ( ~n4045 & n15978 ) | ( ~n4045 & n34613 ) | ( n15978 & n34613 ) ;
  assign n45009 = n45008 ^ n18967 ^ 1'b0 ;
  assign n45010 = n4605 & ~n9608 ;
  assign n45011 = ~n23371 & n25115 ;
  assign n45012 = ~n45010 & n45011 ;
  assign n45013 = ( n18037 & n35170 ) | ( n18037 & ~n45012 ) | ( n35170 & ~n45012 ) ;
  assign n45014 = ~n21525 & n22456 ;
  assign n45017 = n23681 ^ n7145 ^ n5166 ;
  assign n45018 = ( ~n2475 & n7661 ) | ( ~n2475 & n45017 ) | ( n7661 & n45017 ) ;
  assign n45019 = ( n10999 & n23662 ) | ( n10999 & ~n45018 ) | ( n23662 & ~n45018 ) ;
  assign n45015 = ( n11292 & n15779 ) | ( n11292 & n44198 ) | ( n15779 & n44198 ) ;
  assign n45016 = n26188 & ~n45015 ;
  assign n45020 = n45019 ^ n45016 ^ 1'b0 ;
  assign n45021 = ~n38927 & n45020 ;
  assign n45022 = n35025 ^ n32771 ^ n21154 ;
  assign n45023 = ( x19 & ~n20038 ) | ( x19 & n31577 ) | ( ~n20038 & n31577 ) ;
  assign n45024 = n10492 & n14660 ;
  assign n45025 = ~n16889 & n45024 ;
  assign n45026 = n24548 ^ n3175 ^ 1'b0 ;
  assign n45027 = n35310 ^ n19900 ^ n19415 ;
  assign n45028 = n45027 ^ n24847 ^ 1'b0 ;
  assign n45029 = n41495 ^ n18050 ^ n12599 ;
  assign n45030 = ~x140 & n14660 ;
  assign n45031 = ( ~n24252 & n28669 ) | ( ~n24252 & n45030 ) | ( n28669 & n45030 ) ;
  assign n45032 = n45031 ^ n12307 ^ n10289 ;
  assign n45033 = n14652 ^ n8783 ^ 1'b0 ;
  assign n45034 = ( n21079 & n29021 ) | ( n21079 & ~n45033 ) | ( n29021 & ~n45033 ) ;
  assign n45035 = ( ~n9039 & n18059 ) | ( ~n9039 & n42481 ) | ( n18059 & n42481 ) ;
  assign n45036 = n45035 ^ n23282 ^ n8119 ;
  assign n45037 = n12034 & n45036 ;
  assign n45038 = ( n700 & ~n41117 ) | ( n700 & n43172 ) | ( ~n41117 & n43172 ) ;
  assign n45039 = n1084 & n1869 ;
  assign n45040 = ( n14773 & n20492 ) | ( n14773 & n28174 ) | ( n20492 & n28174 ) ;
  assign n45041 = n45039 & n45040 ;
  assign n45042 = n45041 ^ n13078 ^ n2329 ;
  assign n45043 = ( n12965 & ~n16615 ) | ( n12965 & n32303 ) | ( ~n16615 & n32303 ) ;
  assign n45044 = n10566 ^ n5806 ^ 1'b0 ;
  assign n45045 = ( ~n4407 & n5500 ) | ( ~n4407 & n13890 ) | ( n5500 & n13890 ) ;
  assign n45046 = n45045 ^ n11108 ^ 1'b0 ;
  assign n45047 = n8734 & n44964 ;
  assign n45048 = n21993 & n45047 ;
  assign n45049 = ( n37376 & n43516 ) | ( n37376 & ~n45048 ) | ( n43516 & ~n45048 ) ;
  assign n45050 = ( ~n9180 & n14000 ) | ( ~n9180 & n31438 ) | ( n14000 & n31438 ) ;
  assign n45051 = n16564 ^ n10639 ^ n2288 ;
  assign n45052 = ( ~n35768 & n45050 ) | ( ~n35768 & n45051 ) | ( n45050 & n45051 ) ;
  assign n45053 = n35316 ^ n11042 ^ n2683 ;
  assign n45054 = n45053 ^ n35962 ^ n24709 ;
  assign n45055 = n45054 ^ n19583 ^ 1'b0 ;
  assign n45056 = n18253 & ~n29326 ;
  assign n45057 = n2400 & n45056 ;
  assign n45058 = n35837 ^ n29773 ^ n27414 ;
  assign n45059 = n43713 ^ n23724 ^ n12850 ;
  assign n45060 = n28911 ^ n11726 ^ n5386 ;
  assign n45061 = ~n22494 & n25422 ;
  assign n45062 = n45061 ^ n10125 ^ 1'b0 ;
  assign n45063 = ( n2899 & ~n10963 ) | ( n2899 & n14653 ) | ( ~n10963 & n14653 ) ;
  assign n45065 = n21930 ^ n14405 ^ n9600 ;
  assign n45064 = n27455 ^ n9638 ^ n798 ;
  assign n45066 = n45065 ^ n45064 ^ n31448 ;
  assign n45069 = n16993 ^ n13138 ^ n3800 ;
  assign n45067 = n34984 ^ n12296 ^ 1'b0 ;
  assign n45068 = n45067 ^ n15610 ^ n269 ;
  assign n45070 = n45069 ^ n45068 ^ n35063 ;
  assign n45071 = n3390 | n15438 ;
  assign n45072 = n8902 | n45071 ;
  assign n45073 = n546 & ~n19259 ;
  assign n45074 = n45072 & n45073 ;
  assign n45075 = n45074 ^ n33117 ^ 1'b0 ;
  assign n45076 = n9540 ^ n4684 ^ n1379 ;
  assign n45077 = n8105 & n45076 ;
  assign n45078 = ~n18972 & n23045 ;
  assign n45079 = n5675 ^ n5176 ^ n3939 ;
  assign n45080 = ( n11756 & n23023 ) | ( n11756 & ~n45079 ) | ( n23023 & ~n45079 ) ;
  assign n45081 = n38567 ^ n37337 ^ n30911 ;
  assign n45082 = ( n35552 & ~n41089 ) | ( n35552 & n45081 ) | ( ~n41089 & n45081 ) ;
  assign n45083 = n9785 & ~n31557 ;
  assign n45084 = n45083 ^ n15361 ^ n11144 ;
  assign n45085 = ( n10612 & n35357 ) | ( n10612 & n45084 ) | ( n35357 & n45084 ) ;
  assign n45086 = n40971 ^ n38287 ^ 1'b0 ;
  assign n45087 = n5975 ^ n5370 ^ 1'b0 ;
  assign n45088 = n18869 & n45087 ;
  assign n45089 = n3766 & ~n22481 ;
  assign n45090 = ~n3341 & n45089 ;
  assign n45091 = n7961 | n45090 ;
  assign n45092 = n45091 ^ n15761 ^ 1'b0 ;
  assign n45093 = n15891 ^ n11811 ^ 1'b0 ;
  assign n45094 = n45093 ^ n24471 ^ 1'b0 ;
  assign n45095 = n45092 | n45094 ;
  assign n45096 = n14389 ^ n7448 ^ n5812 ;
  assign n45097 = n45096 ^ n39612 ^ 1'b0 ;
  assign n45098 = ~n16074 & n22506 ;
  assign n45099 = n45098 ^ n14544 ^ 1'b0 ;
  assign n45100 = n23086 | n45099 ;
  assign n45101 = n26716 | n45100 ;
  assign n45102 = n45101 ^ n41848 ^ 1'b0 ;
  assign n45103 = ~n12952 & n15676 ;
  assign n45104 = ~n12985 & n45103 ;
  assign n45105 = ( n23749 & ~n32420 ) | ( n23749 & n45104 ) | ( ~n32420 & n45104 ) ;
  assign n45109 = ~n6451 & n16754 ;
  assign n45110 = n45109 ^ n12115 ^ 1'b0 ;
  assign n45111 = n45110 ^ n9439 ^ n6336 ;
  assign n45112 = n26288 ^ n10027 ^ 1'b0 ;
  assign n45113 = ~n26956 & n45112 ;
  assign n45114 = ( n2668 & n45111 ) | ( n2668 & n45113 ) | ( n45111 & n45113 ) ;
  assign n45106 = x5 & ~n6871 ;
  assign n45107 = ( n840 & ~n29569 ) | ( n840 & n45106 ) | ( ~n29569 & n45106 ) ;
  assign n45108 = n20040 | n45107 ;
  assign n45115 = n45114 ^ n45108 ^ n36603 ;
  assign n45116 = ( ~n24012 & n45105 ) | ( ~n24012 & n45115 ) | ( n45105 & n45115 ) ;
  assign n45117 = ( n13632 & ~n21738 ) | ( n13632 & n29702 ) | ( ~n21738 & n29702 ) ;
  assign n45118 = n31561 ^ n22464 ^ n21898 ;
  assign n45119 = n14105 ^ n2341 ^ n766 ;
  assign n45120 = n45119 ^ n2704 ^ n715 ;
  assign n45121 = n44417 ^ n38779 ^ n2452 ;
  assign n45122 = n1057 | n16047 ;
  assign n45123 = n45122 ^ n10538 ^ 1'b0 ;
  assign n45124 = n36601 ^ n27406 ^ n22408 ;
  assign n45125 = n36184 ^ n33956 ^ n15033 ;
  assign n45126 = n45125 ^ n30330 ^ n18666 ;
  assign n45127 = ( n16128 & n27135 ) | ( n16128 & n45126 ) | ( n27135 & n45126 ) ;
  assign n45128 = n28419 ^ n17612 ^ 1'b0 ;
  assign n45129 = n45128 ^ n18679 ^ n15962 ;
  assign n45130 = ( n2833 & ~n17399 ) | ( n2833 & n45129 ) | ( ~n17399 & n45129 ) ;
  assign n45131 = n42124 ^ n26775 ^ n11012 ;
  assign n45132 = ( ~n13779 & n28180 ) | ( ~n13779 & n38155 ) | ( n28180 & n38155 ) ;
  assign n45133 = n40648 ^ n39738 ^ n4904 ;
  assign n45134 = n34563 ^ n30216 ^ n1883 ;
  assign n45135 = n6499 | n40473 ;
  assign n45136 = n45134 | n45135 ;
  assign n45137 = n8856 & n17913 ;
  assign n45138 = n45137 ^ n5236 ^ 1'b0 ;
  assign n45140 = ( n27553 & n38221 ) | ( n27553 & n40282 ) | ( n38221 & n40282 ) ;
  assign n45141 = ( n29079 & ~n31936 ) | ( n29079 & n45140 ) | ( ~n31936 & n45140 ) ;
  assign n45139 = n1555 & ~n2929 ;
  assign n45142 = n45141 ^ n45139 ^ 1'b0 ;
  assign n45145 = n31111 ^ n6199 ^ 1'b0 ;
  assign n45143 = ~n20423 & n28731 ;
  assign n45144 = n45143 ^ x40 ^ 1'b0 ;
  assign n45146 = n45145 ^ n45144 ^ x42 ;
  assign n45147 = n24741 ^ n14673 ^ n2435 ;
  assign n45148 = ( ~n34118 & n37692 ) | ( ~n34118 & n45147 ) | ( n37692 & n45147 ) ;
  assign n45149 = n45148 ^ n26892 ^ n14870 ;
  assign n45150 = n32593 ^ n11414 ^ 1'b0 ;
  assign n45151 = n45150 ^ n14528 ^ n6987 ;
  assign n45152 = n42497 ^ n14606 ^ n10590 ;
  assign n45153 = ( n6411 & ~n17567 ) | ( n6411 & n42379 ) | ( ~n17567 & n42379 ) ;
  assign n45154 = n45153 ^ n21823 ^ n2644 ;
  assign n45155 = ~n11012 & n14026 ;
  assign n45156 = n45155 ^ n17935 ^ 1'b0 ;
  assign n45157 = ~n8643 & n31562 ;
  assign n45158 = n15851 | n22060 ;
  assign n45159 = n45158 ^ n7062 ^ 1'b0 ;
  assign n45160 = ( ~n11071 & n23666 ) | ( ~n11071 & n45159 ) | ( n23666 & n45159 ) ;
  assign n45161 = n45160 ^ n9569 ^ 1'b0 ;
  assign n45162 = n34580 & n45161 ;
  assign n45163 = n36949 ^ n19609 ^ 1'b0 ;
  assign n45164 = n36082 & ~n45163 ;
  assign n45165 = n9929 | n27951 ;
  assign n45166 = ( n21354 & n40808 ) | ( n21354 & n45165 ) | ( n40808 & n45165 ) ;
  assign n45167 = ( ~n9067 & n19239 ) | ( ~n9067 & n34346 ) | ( n19239 & n34346 ) ;
  assign n45168 = n527 | n7852 ;
  assign n45169 = n11703 ^ n7367 ^ 1'b0 ;
  assign n45170 = n644 & ~n45169 ;
  assign n45171 = n45170 ^ n35563 ^ n20130 ;
  assign n45172 = ( n42624 & n45168 ) | ( n42624 & ~n45171 ) | ( n45168 & ~n45171 ) ;
  assign n45173 = n29907 ^ n7815 ^ 1'b0 ;
  assign n45174 = n12142 ^ n5888 ^ 1'b0 ;
  assign n45175 = ( n42060 & n45173 ) | ( n42060 & ~n45174 ) | ( n45173 & ~n45174 ) ;
  assign n45177 = ( x76 & n1848 ) | ( x76 & n18346 ) | ( n1848 & n18346 ) ;
  assign n45178 = x86 & n45177 ;
  assign n45179 = n26345 & n45178 ;
  assign n45176 = ~n7765 & n36149 ;
  assign n45180 = n45179 ^ n45176 ^ 1'b0 ;
  assign n45182 = n30450 ^ n23486 ^ n20911 ;
  assign n45181 = ~n18204 & n38413 ;
  assign n45183 = n45182 ^ n45181 ^ 1'b0 ;
  assign n45184 = n3954 & ~n27501 ;
  assign n45188 = n31760 ^ n12121 ^ n5575 ;
  assign n45185 = ( n10172 & ~n10985 ) | ( n10172 & n20307 ) | ( ~n10985 & n20307 ) ;
  assign n45186 = ( n10212 & n16333 ) | ( n10212 & n45185 ) | ( n16333 & n45185 ) ;
  assign n45187 = n45186 ^ n23942 ^ n19561 ;
  assign n45189 = n45188 ^ n45187 ^ n40951 ;
  assign n45190 = n45189 ^ n34851 ^ n3091 ;
  assign n45191 = ( n34601 & ~n39324 ) | ( n34601 & n43100 ) | ( ~n39324 & n43100 ) ;
  assign n45192 = ( ~n21373 & n29143 ) | ( ~n21373 & n35907 ) | ( n29143 & n35907 ) ;
  assign n45193 = n30244 ^ n2150 ^ 1'b0 ;
  assign n45194 = n37874 & n45193 ;
  assign n45195 = n30611 ^ n13493 ^ n2592 ;
  assign n45196 = n27485 ^ n8907 ^ 1'b0 ;
  assign n45197 = n10049 ^ n3599 ^ 1'b0 ;
  assign n45198 = ( n7259 & ~n28397 ) | ( n7259 & n39652 ) | ( ~n28397 & n39652 ) ;
  assign n45199 = ~n9139 & n45198 ;
  assign n45200 = ( n27705 & n35458 ) | ( n27705 & n45199 ) | ( n35458 & n45199 ) ;
  assign n45201 = n27734 | n35804 ;
  assign n45202 = n24204 ^ n14563 ^ 1'b0 ;
  assign n45203 = ~n44620 & n45202 ;
  assign n45204 = n45203 ^ n16377 ^ n1863 ;
  assign n45205 = n20576 ^ n18884 ^ n7738 ;
  assign n45206 = n15944 & ~n23979 ;
  assign n45207 = n45206 ^ n16819 ^ 1'b0 ;
  assign n45208 = n23286 ^ n11152 ^ 1'b0 ;
  assign n45209 = n35749 ^ n31773 ^ 1'b0 ;
  assign n45210 = n45208 & n45209 ;
  assign n45211 = n17621 ^ n14359 ^ 1'b0 ;
  assign n45212 = n45211 ^ n1448 ^ 1'b0 ;
  assign n45213 = n16562 & n45212 ;
  assign n45214 = ~n45210 & n45213 ;
  assign n45215 = n40406 ^ n34624 ^ n25334 ;
  assign n45216 = ( n3581 & n15469 ) | ( n3581 & n45215 ) | ( n15469 & n45215 ) ;
  assign n45217 = ~n857 & n1537 ;
  assign n45218 = ~n23239 & n45217 ;
  assign n45219 = n6652 & n15944 ;
  assign n45220 = n45219 ^ n28995 ^ 1'b0 ;
  assign n45221 = ( n45216 & n45218 ) | ( n45216 & n45220 ) | ( n45218 & n45220 ) ;
  assign n45224 = n36341 ^ n32084 ^ 1'b0 ;
  assign n45222 = n22527 ^ n10170 ^ 1'b0 ;
  assign n45223 = ( n39366 & ~n40909 ) | ( n39366 & n45222 ) | ( ~n40909 & n45222 ) ;
  assign n45225 = n45224 ^ n45223 ^ n21976 ;
  assign n45230 = n10869 ^ n3435 ^ 1'b0 ;
  assign n45231 = n22536 & n45230 ;
  assign n45226 = ~n14667 & n26530 ;
  assign n45227 = n33451 ^ n1632 ^ x232 ;
  assign n45228 = n45226 | n45227 ;
  assign n45229 = n18986 & ~n45228 ;
  assign n45232 = n45231 ^ n45229 ^ n30057 ;
  assign n45233 = ( n15114 & n17589 ) | ( n15114 & ~n42251 ) | ( n17589 & ~n42251 ) ;
  assign n45234 = n8882 | n12298 ;
  assign n45235 = n45234 ^ n3318 ^ 1'b0 ;
  assign n45236 = n31164 | n45235 ;
  assign n45237 = n45236 ^ n6590 ^ 1'b0 ;
  assign n45238 = n3062 & ~n30825 ;
  assign n45239 = ( x99 & n9103 ) | ( x99 & n9846 ) | ( n9103 & n9846 ) ;
  assign n45240 = n45239 ^ n33387 ^ n24825 ;
  assign n45241 = n21102 ^ n9152 ^ n4407 ;
  assign n45242 = ( n8229 & n32351 ) | ( n8229 & n45241 ) | ( n32351 & n45241 ) ;
  assign n45243 = ( ~n1151 & n14391 ) | ( ~n1151 & n28672 ) | ( n14391 & n28672 ) ;
  assign n45244 = n45243 ^ n4838 ^ n4362 ;
  assign n45245 = n12334 & ~n45244 ;
  assign n45246 = n45242 & ~n45245 ;
  assign n45247 = n18092 ^ n13062 ^ n10503 ;
  assign n45248 = n28945 | n45247 ;
  assign n45249 = ( n11241 & n12701 ) | ( n11241 & n40059 ) | ( n12701 & n40059 ) ;
  assign n45250 = n31422 ^ n11475 ^ n8814 ;
  assign n45251 = n8730 & n32369 ;
  assign n45252 = n45250 & n45251 ;
  assign n45253 = n17869 & ~n18356 ;
  assign n45254 = ( n29184 & n35636 ) | ( n29184 & ~n45253 ) | ( n35636 & ~n45253 ) ;
  assign n45255 = x34 & ~n45254 ;
  assign n45256 = n2540 & n16072 ;
  assign n45257 = n45256 ^ n13169 ^ 1'b0 ;
  assign n45258 = n8205 ^ n4216 ^ 1'b0 ;
  assign n45268 = n4704 ^ n971 ^ 1'b0 ;
  assign n45269 = ~n4223 & n45268 ;
  assign n45270 = n14319 ^ n3206 ^ 1'b0 ;
  assign n45271 = n45269 & n45270 ;
  assign n45265 = n33842 ^ n25205 ^ n22833 ;
  assign n45266 = n45265 ^ n20380 ^ 1'b0 ;
  assign n45259 = ( n2740 & ~n7403 ) | ( n2740 & n16526 ) | ( ~n7403 & n16526 ) ;
  assign n45260 = ( ~n4051 & n6025 ) | ( ~n4051 & n45259 ) | ( n6025 & n45259 ) ;
  assign n45261 = n32790 ^ n31254 ^ n11446 ;
  assign n45262 = n45261 ^ n16246 ^ 1'b0 ;
  assign n45263 = n45260 & ~n45262 ;
  assign n45264 = n14231 & n45263 ;
  assign n45267 = n45266 ^ n45264 ^ 1'b0 ;
  assign n45272 = n45271 ^ n45267 ^ 1'b0 ;
  assign n45273 = ( n38538 & n42159 ) | ( n38538 & n45272 ) | ( n42159 & n45272 ) ;
  assign n45274 = n5064 ^ n536 ^ x126 ;
  assign n45275 = n16172 ^ n14582 ^ n9398 ;
  assign n45276 = n45274 & ~n45275 ;
  assign n45277 = ( n2607 & n8970 ) | ( n2607 & n38533 ) | ( n8970 & n38533 ) ;
  assign n45278 = n45277 ^ n15221 ^ n8020 ;
  assign n45279 = n45278 ^ n40256 ^ n10672 ;
  assign n45280 = n6919 ^ n3661 ^ 1'b0 ;
  assign n45281 = n36198 ^ n24461 ^ 1'b0 ;
  assign n45282 = n5962 & ~n45281 ;
  assign n45283 = n5686 & ~n34694 ;
  assign n45284 = n45283 ^ n19640 ^ 1'b0 ;
  assign n45285 = n45284 ^ n28269 ^ n11351 ;
  assign n45286 = n29229 & ~n45285 ;
  assign n45287 = n27999 ^ n20263 ^ 1'b0 ;
  assign n45288 = ~n17767 & n45287 ;
  assign n45289 = ~n12074 & n22690 ;
  assign n45290 = n45289 ^ n21321 ^ n3460 ;
  assign n45291 = n11448 ^ n3677 ^ 1'b0 ;
  assign n45292 = ~n8745 & n45291 ;
  assign n45293 = n40165 ^ n17092 ^ n6307 ;
  assign n45294 = ( n31442 & n45292 ) | ( n31442 & ~n45293 ) | ( n45292 & ~n45293 ) ;
  assign n45295 = n8100 | n20946 ;
  assign n45296 = ( ~n13828 & n29398 ) | ( ~n13828 & n45295 ) | ( n29398 & n45295 ) ;
  assign n45297 = n11792 ^ n7735 ^ 1'b0 ;
  assign n45298 = n36353 & n45297 ;
  assign n45299 = n45298 ^ n2923 ^ 1'b0 ;
  assign n45300 = n45299 ^ n6110 ^ 1'b0 ;
  assign n45301 = ( n7302 & n17667 ) | ( n7302 & ~n19848 ) | ( n17667 & ~n19848 ) ;
  assign n45302 = n45301 ^ n13209 ^ 1'b0 ;
  assign n45303 = ( n23376 & n26066 ) | ( n23376 & ~n32834 ) | ( n26066 & ~n32834 ) ;
  assign n45304 = n24566 ^ n12524 ^ 1'b0 ;
  assign n45305 = n18166 & n22016 ;
  assign n45306 = ~n32099 & n45305 ;
  assign n45307 = n3106 | n12701 ;
  assign n45308 = ( n4067 & n7686 ) | ( n4067 & ~n45307 ) | ( n7686 & ~n45307 ) ;
  assign n45309 = ( n9608 & n45293 ) | ( n9608 & ~n45308 ) | ( n45293 & ~n45308 ) ;
  assign n45310 = n22762 ^ n17931 ^ 1'b0 ;
  assign n45311 = n9674 & ~n45310 ;
  assign n45312 = ( n14150 & ~n17691 ) | ( n14150 & n45311 ) | ( ~n17691 & n45311 ) ;
  assign n45315 = n28889 ^ n15836 ^ n8924 ;
  assign n45314 = ( n2984 & ~n18670 ) | ( n2984 & n33516 ) | ( ~n18670 & n33516 ) ;
  assign n45313 = ( n11440 & ~n14290 ) | ( n11440 & n31587 ) | ( ~n14290 & n31587 ) ;
  assign n45316 = n45315 ^ n45314 ^ n45313 ;
  assign n45320 = n20126 ^ n12132 ^ n4901 ;
  assign n45317 = ( n2750 & n9565 ) | ( n2750 & n10045 ) | ( n9565 & n10045 ) ;
  assign n45318 = n40552 | n45317 ;
  assign n45319 = n9670 & ~n45318 ;
  assign n45321 = n45320 ^ n45319 ^ 1'b0 ;
  assign n45322 = n45321 ^ n40647 ^ n9138 ;
  assign n45323 = ( ~n17595 & n36121 ) | ( ~n17595 & n42237 ) | ( n36121 & n42237 ) ;
  assign n45324 = n45323 ^ n37643 ^ n3053 ;
  assign n45325 = n39526 ^ n32468 ^ 1'b0 ;
  assign n45326 = ( ~n24046 & n43656 ) | ( ~n24046 & n45325 ) | ( n43656 & n45325 ) ;
  assign n45328 = ( ~n23030 & n23057 ) | ( ~n23030 & n28690 ) | ( n23057 & n28690 ) ;
  assign n45327 = ~n32642 & n37955 ;
  assign n45329 = n45328 ^ n45327 ^ 1'b0 ;
  assign n45330 = n9584 ^ n2457 ^ 1'b0 ;
  assign n45331 = ~n37896 & n45330 ;
  assign n45332 = ( n9686 & n11711 ) | ( n9686 & n12105 ) | ( n11711 & n12105 ) ;
  assign n45333 = n45332 ^ n40259 ^ n6423 ;
  assign n45334 = ( ~n1632 & n2406 ) | ( ~n1632 & n32301 ) | ( n2406 & n32301 ) ;
  assign n45335 = n45334 ^ n21200 ^ n20915 ;
  assign n45336 = n39223 ^ n22989 ^ n20202 ;
  assign n45342 = n28586 ^ n22273 ^ 1'b0 ;
  assign n45343 = ~n6624 & n45342 ;
  assign n45340 = n8232 ^ n7980 ^ n4952 ;
  assign n45337 = n3171 ^ n796 ^ 1'b0 ;
  assign n45338 = n8083 | n45337 ;
  assign n45339 = ( ~n1100 & n6031 ) | ( ~n1100 & n45338 ) | ( n6031 & n45338 ) ;
  assign n45341 = n45340 ^ n45339 ^ n13327 ;
  assign n45344 = n45343 ^ n45341 ^ n18990 ;
  assign n45345 = n42124 ^ n11117 ^ n7430 ;
  assign n45346 = n12258 ^ n9884 ^ n5974 ;
  assign n45347 = n13275 | n23379 ;
  assign n45348 = n45347 ^ n41441 ^ 1'b0 ;
  assign n45349 = n2753 & n8197 ;
  assign n45350 = n45349 ^ n21176 ^ 1'b0 ;
  assign n45351 = n24811 | n45350 ;
  assign n45352 = n28221 ^ n23950 ^ n10318 ;
  assign n45353 = ( n15548 & n39139 ) | ( n15548 & ~n45352 ) | ( n39139 & ~n45352 ) ;
  assign n45354 = ( n6283 & n16377 ) | ( n6283 & n39084 ) | ( n16377 & n39084 ) ;
  assign n45355 = n45354 ^ n34253 ^ n26478 ;
  assign n45356 = n21165 ^ n7798 ^ 1'b0 ;
  assign n45357 = n26216 & n45356 ;
  assign n45358 = ( n17230 & n23724 ) | ( n17230 & ~n45357 ) | ( n23724 & ~n45357 ) ;
  assign n45359 = n17951 ^ n11286 ^ 1'b0 ;
  assign n45360 = ( n7635 & n8197 ) | ( n7635 & ~n11021 ) | ( n8197 & ~n11021 ) ;
  assign n45361 = ( n4584 & n16640 ) | ( n4584 & n45360 ) | ( n16640 & n45360 ) ;
  assign n45362 = n45361 ^ n17671 ^ 1'b0 ;
  assign n45363 = n45359 & ~n45362 ;
  assign n45364 = ~n7333 & n45363 ;
  assign n45365 = ( n4872 & ~n12194 ) | ( n4872 & n18577 ) | ( ~n12194 & n18577 ) ;
  assign n45366 = ~n19872 & n45365 ;
  assign n45368 = ( ~n540 & n2629 ) | ( ~n540 & n9593 ) | ( n2629 & n9593 ) ;
  assign n45369 = n1476 & ~n45368 ;
  assign n45367 = ~n12842 & n20119 ;
  assign n45370 = n45369 ^ n45367 ^ n31015 ;
  assign n45371 = n6272 ^ n4657 ^ n563 ;
  assign n45372 = ( n16355 & n24892 ) | ( n16355 & ~n45371 ) | ( n24892 & ~n45371 ) ;
  assign n45373 = n38971 ^ n14950 ^ n606 ;
  assign n45374 = ( n19929 & n45372 ) | ( n19929 & ~n45373 ) | ( n45372 & ~n45373 ) ;
  assign n45375 = n45374 ^ n28434 ^ 1'b0 ;
  assign n45376 = n16360 & ~n45375 ;
  assign n45377 = n11966 | n24025 ;
  assign n45378 = n13647 ^ n6632 ^ n797 ;
  assign n45379 = n45378 ^ n36380 ^ n12346 ;
  assign n45380 = n18574 ^ n14507 ^ 1'b0 ;
  assign n45381 = n15626 | n37558 ;
  assign n45382 = n40850 ^ n5457 ^ n4467 ;
  assign n45383 = n45382 ^ n31801 ^ n3820 ;
  assign n45385 = ( n11417 & n16524 ) | ( n11417 & ~n22622 ) | ( n16524 & ~n22622 ) ;
  assign n45384 = n35947 ^ n5202 ^ 1'b0 ;
  assign n45386 = n45385 ^ n45384 ^ n6279 ;
  assign n45387 = ( n20677 & n20986 ) | ( n20677 & n45386 ) | ( n20986 & n45386 ) ;
  assign n45388 = n29021 & n35271 ;
  assign n45389 = n45388 ^ n30330 ^ 1'b0 ;
  assign n45390 = n15616 & ~n45389 ;
  assign n45391 = ~n36806 & n45390 ;
  assign n45392 = ~n1434 & n21167 ;
  assign n45393 = n27546 & n33244 ;
  assign n45394 = n45393 ^ n35524 ^ 1'b0 ;
  assign n45395 = n45392 | n45394 ;
  assign n45396 = n45395 ^ n9930 ^ 1'b0 ;
  assign n45398 = ~n1705 & n9980 ;
  assign n45397 = n27672 ^ n12370 ^ 1'b0 ;
  assign n45399 = n45398 ^ n45397 ^ n3717 ;
  assign n45400 = n45399 ^ n30583 ^ 1'b0 ;
  assign n45401 = ~n40672 & n45400 ;
  assign n45402 = n2101 & n3591 ;
  assign n45408 = n6336 ^ n3006 ^ 1'b0 ;
  assign n45409 = ~n7467 & n45408 ;
  assign n45406 = n14850 ^ n7944 ^ n4610 ;
  assign n45403 = n11075 | n12579 ;
  assign n45404 = n8944 & n45403 ;
  assign n45405 = n45404 ^ n11198 ^ 1'b0 ;
  assign n45407 = n45406 ^ n45405 ^ n26640 ;
  assign n45410 = n45409 ^ n45407 ^ n7202 ;
  assign n45413 = ( ~n3844 & n4649 ) | ( ~n3844 & n24516 ) | ( n4649 & n24516 ) ;
  assign n45414 = n45413 ^ n34063 ^ n8928 ;
  assign n45411 = n19179 ^ n12954 ^ n9002 ;
  assign n45412 = n45411 ^ n32651 ^ n31639 ;
  assign n45415 = n45414 ^ n45412 ^ 1'b0 ;
  assign n45416 = n31301 ^ n18004 ^ n11039 ;
  assign n45417 = n45416 ^ n39105 ^ 1'b0 ;
  assign n45418 = n12950 & ~n45417 ;
  assign n45419 = n1860 & n5572 ;
  assign n45420 = ~n44870 & n45419 ;
  assign n45421 = ~n7451 & n45420 ;
  assign n45422 = n30588 ^ n20804 ^ 1'b0 ;
  assign n45423 = ~n8015 & n45422 ;
  assign n45424 = ( n7432 & n9560 ) | ( n7432 & ~n13817 ) | ( n9560 & ~n13817 ) ;
  assign n45425 = n45424 ^ n6089 ^ n4826 ;
  assign n45426 = ~n7148 & n24526 ;
  assign n45427 = ( n1947 & n42847 ) | ( n1947 & ~n45426 ) | ( n42847 & ~n45426 ) ;
  assign n45428 = ~n11530 & n44188 ;
  assign n45429 = ( n1645 & n44907 ) | ( n1645 & ~n45428 ) | ( n44907 & ~n45428 ) ;
  assign n45430 = n17186 ^ n9432 ^ n8090 ;
  assign n45431 = n4574 & ~n45430 ;
  assign n45432 = n1790 | n30445 ;
  assign n45433 = ( n15017 & n38862 ) | ( n15017 & n45432 ) | ( n38862 & n45432 ) ;
  assign n45434 = ( n2051 & n10294 ) | ( n2051 & ~n13418 ) | ( n10294 & ~n13418 ) ;
  assign n45435 = n45434 ^ n7264 ^ n6157 ;
  assign n45436 = n24635 ^ n14528 ^ 1'b0 ;
  assign n45437 = n25512 & n45436 ;
  assign n45438 = n32877 ^ n8413 ^ 1'b0 ;
  assign n45439 = ~n31782 & n45438 ;
  assign n45440 = ~n21963 & n37561 ;
  assign n45441 = ~n38150 & n45440 ;
  assign n45442 = n17204 & n37180 ;
  assign n45443 = n45441 & n45442 ;
  assign n45444 = ( ~n12167 & n17005 ) | ( ~n12167 & n19964 ) | ( n17005 & n19964 ) ;
  assign n45445 = n45444 ^ n41986 ^ 1'b0 ;
  assign n45446 = n24922 & ~n45445 ;
  assign n45449 = ( n18316 & n18555 ) | ( n18316 & ~n19399 ) | ( n18555 & ~n19399 ) ;
  assign n45447 = n5256 & ~n31174 ;
  assign n45448 = n41099 & n45447 ;
  assign n45450 = n45449 ^ n45448 ^ n37978 ;
  assign n45451 = n9861 ^ n6737 ^ n5628 ;
  assign n45452 = ~n24320 & n45451 ;
  assign n45453 = n45452 ^ n23253 ^ n4901 ;
  assign n45454 = n36799 | n45453 ;
  assign n45455 = n45454 ^ n12776 ^ 1'b0 ;
  assign n45456 = n45455 ^ n4154 ^ 1'b0 ;
  assign n45457 = n12282 & ~n12807 ;
  assign n45458 = ( ~n1001 & n2260 ) | ( ~n1001 & n16654 ) | ( n2260 & n16654 ) ;
  assign n45459 = n27242 ^ n18699 ^ 1'b0 ;
  assign n45460 = n45459 ^ n15493 ^ n8977 ;
  assign n45461 = ( n15033 & ~n29031 ) | ( n15033 & n41195 ) | ( ~n29031 & n41195 ) ;
  assign n45462 = ( ~n9341 & n21359 ) | ( ~n9341 & n33898 ) | ( n21359 & n33898 ) ;
  assign n45463 = n45431 ^ n17478 ^ 1'b0 ;
  assign n45464 = n25439 ^ n12593 ^ n4517 ;
  assign n45465 = ( ~n3104 & n11301 ) | ( ~n3104 & n27490 ) | ( n11301 & n27490 ) ;
  assign n45466 = n37805 ^ n14205 ^ 1'b0 ;
  assign n45467 = n45466 ^ n23501 ^ n16439 ;
  assign n45468 = ( n3596 & ~n9609 ) | ( n3596 & n9674 ) | ( ~n9609 & n9674 ) ;
  assign n45469 = n45468 ^ n35620 ^ 1'b0 ;
  assign n45470 = n45072 ^ n43897 ^ n4642 ;
  assign n45471 = n45470 ^ n24604 ^ n8897 ;
  assign n45472 = n45471 ^ n14146 ^ 1'b0 ;
  assign n45473 = n16834 ^ n12461 ^ 1'b0 ;
  assign n45474 = n28255 | n45473 ;
  assign n45475 = n3137 & ~n45474 ;
  assign n45476 = n45475 ^ n24228 ^ 1'b0 ;
  assign n45477 = n23315 ^ n12887 ^ n5696 ;
  assign n45478 = n38967 & n44457 ;
  assign n45479 = n45477 & n45478 ;
  assign n45480 = n45479 ^ n42274 ^ n32461 ;
  assign n45481 = ( n19842 & n37725 ) | ( n19842 & n40202 ) | ( n37725 & n40202 ) ;
  assign n45482 = n3917 & n33830 ;
  assign n45483 = ( n17458 & n24709 ) | ( n17458 & n45482 ) | ( n24709 & n45482 ) ;
  assign n45485 = n20008 | n36892 ;
  assign n45484 = ( n6687 & n19894 ) | ( n6687 & n42906 ) | ( n19894 & n42906 ) ;
  assign n45486 = n45485 ^ n45484 ^ n33273 ;
  assign n45487 = ( ~n956 & n11507 ) | ( ~n956 & n20525 ) | ( n11507 & n20525 ) ;
  assign n45488 = ( n24758 & n26431 ) | ( n24758 & ~n45487 ) | ( n26431 & ~n45487 ) ;
  assign n45489 = ( n7305 & n23190 ) | ( n7305 & n45488 ) | ( n23190 & n45488 ) ;
  assign n45490 = n14361 ^ x226 ^ 1'b0 ;
  assign n45491 = ( ~n2737 & n20030 ) | ( ~n2737 & n39008 ) | ( n20030 & n39008 ) ;
  assign n45492 = n10591 & n45491 ;
  assign n45493 = n26817 & n45492 ;
  assign n45494 = ( n8686 & n22646 ) | ( n8686 & ~n24573 ) | ( n22646 & ~n24573 ) ;
  assign n45495 = n45494 ^ n14029 ^ n8160 ;
  assign n45496 = ( ~n310 & n8955 ) | ( ~n310 & n38899 ) | ( n8955 & n38899 ) ;
  assign n45497 = ~n1339 & n7979 ;
  assign n45498 = n21570 | n28696 ;
  assign n45499 = n27474 ^ n6141 ^ 1'b0 ;
  assign n45500 = n26758 | n45499 ;
  assign n45501 = n14105 ^ n4575 ^ 1'b0 ;
  assign n45502 = n24655 & n45501 ;
  assign n45503 = n43219 ^ n8716 ^ n2795 ;
  assign n45504 = n45503 ^ n21107 ^ n7786 ;
  assign n45505 = n28798 ^ n20515 ^ 1'b0 ;
  assign n45506 = ( n45277 & ~n45504 ) | ( n45277 & n45505 ) | ( ~n45504 & n45505 ) ;
  assign n45507 = n4554 ^ n4137 ^ 1'b0 ;
  assign n45508 = n43946 ^ n9810 ^ 1'b0 ;
  assign n45509 = n3131 | n45508 ;
  assign n45510 = ( n13567 & n45507 ) | ( n13567 & n45509 ) | ( n45507 & n45509 ) ;
  assign n45511 = n11779 & n14793 ;
  assign n45512 = n10532 & n45511 ;
  assign n45513 = n45512 ^ n19051 ^ n6635 ;
  assign n45514 = n31036 ^ n10726 ^ n6735 ;
  assign n45515 = n14202 ^ n13176 ^ n340 ;
  assign n45517 = ( n2380 & n21113 ) | ( n2380 & n40501 ) | ( n21113 & n40501 ) ;
  assign n45516 = ~n4350 & n8623 ;
  assign n45518 = n45517 ^ n45516 ^ 1'b0 ;
  assign n45519 = n30423 ^ n22399 ^ n1594 ;
  assign n45520 = n26494 ^ n5420 ^ 1'b0 ;
  assign n45521 = ~n19573 & n24741 ;
  assign n45522 = ~n30594 & n45521 ;
  assign n45523 = ( n6497 & n38888 ) | ( n6497 & n45522 ) | ( n38888 & n45522 ) ;
  assign n45524 = n35112 ^ n20234 ^ n1647 ;
  assign n45528 = ( ~n14318 & n19038 ) | ( ~n14318 & n21189 ) | ( n19038 & n21189 ) ;
  assign n45526 = n18215 & n38236 ;
  assign n45527 = n45526 ^ n24442 ^ n3000 ;
  assign n45525 = ( n5652 & n9725 ) | ( n5652 & n15424 ) | ( n9725 & n15424 ) ;
  assign n45529 = n45528 ^ n45527 ^ n45525 ;
  assign n45530 = n3545 & ~n40625 ;
  assign n45531 = n34545 & n45530 ;
  assign n45532 = n17024 ^ n6786 ^ 1'b0 ;
  assign n45533 = n3507 & n22174 ;
  assign n45534 = ( n26195 & ~n35425 ) | ( n26195 & n42996 ) | ( ~n35425 & n42996 ) ;
  assign n45536 = n15526 ^ n2450 ^ 1'b0 ;
  assign n45537 = n22690 & ~n45536 ;
  assign n45538 = ( n8769 & n11955 ) | ( n8769 & n45537 ) | ( n11955 & n45537 ) ;
  assign n45535 = n30320 ^ n22797 ^ n9848 ;
  assign n45539 = n45538 ^ n45535 ^ n32788 ;
  assign n45540 = n17038 ^ n15809 ^ n14881 ;
  assign n45541 = n28402 ^ n17413 ^ n12217 ;
  assign n45542 = n45541 ^ n22969 ^ n5611 ;
  assign n45543 = n24075 ^ n14394 ^ 1'b0 ;
  assign n45544 = ( ~n1690 & n45542 ) | ( ~n1690 & n45543 ) | ( n45542 & n45543 ) ;
  assign n45545 = n30953 ^ n11267 ^ n8639 ;
  assign n45546 = n6475 ^ n6197 ^ 1'b0 ;
  assign n45547 = n35194 ^ n19078 ^ n1384 ;
  assign n45548 = ( n6991 & ~n15280 ) | ( n6991 & n17653 ) | ( ~n15280 & n17653 ) ;
  assign n45549 = n45548 ^ n10528 ^ 1'b0 ;
  assign n45550 = n45547 & ~n45549 ;
  assign n45551 = n14963 ^ n1503 ^ 1'b0 ;
  assign n45552 = n22595 ^ n11236 ^ n1589 ;
  assign n45553 = n11552 | n45552 ;
  assign n45554 = n45553 ^ n13828 ^ 1'b0 ;
  assign n45555 = n25636 ^ n14678 ^ n9205 ;
  assign n45559 = ~n18496 & n38968 ;
  assign n45556 = n39671 ^ n6046 ^ 1'b0 ;
  assign n45557 = n31504 & ~n45556 ;
  assign n45558 = ( n7288 & n12630 ) | ( n7288 & n45557 ) | ( n12630 & n45557 ) ;
  assign n45560 = n45559 ^ n45558 ^ n27635 ;
  assign n45561 = ( ~n3068 & n9634 ) | ( ~n3068 & n12187 ) | ( n9634 & n12187 ) ;
  assign n45562 = n45561 ^ n18252 ^ n4608 ;
  assign n45563 = n45562 ^ n34257 ^ n32242 ;
  assign n45564 = n25320 ^ n23315 ^ 1'b0 ;
  assign n45565 = n26313 ^ n2932 ^ n517 ;
  assign n45566 = n36044 ^ n16352 ^ 1'b0 ;
  assign n45567 = n37740 & ~n45566 ;
  assign n45568 = ( n3787 & n10594 ) | ( n3787 & n32615 ) | ( n10594 & n32615 ) ;
  assign n45569 = n9289 ^ n8275 ^ 1'b0 ;
  assign n45570 = n45568 & ~n45569 ;
  assign n45571 = ( ~n8105 & n12988 ) | ( ~n8105 & n18798 ) | ( n12988 & n18798 ) ;
  assign n45572 = n45571 ^ n13720 ^ n3820 ;
  assign n45573 = ( ~n4545 & n19473 ) | ( ~n4545 & n31829 ) | ( n19473 & n31829 ) ;
  assign n45574 = ( n16749 & n45572 ) | ( n16749 & n45573 ) | ( n45572 & n45573 ) ;
  assign n45575 = n1997 | n19808 ;
  assign n45576 = n36238 ^ n15004 ^ 1'b0 ;
  assign n45577 = n45576 ^ n35430 ^ 1'b0 ;
  assign n45578 = ( n6465 & n13718 ) | ( n6465 & ~n45577 ) | ( n13718 & ~n45577 ) ;
  assign n45579 = n44770 | n45578 ;
  assign n45580 = ( n2847 & ~n3828 ) | ( n2847 & n22788 ) | ( ~n3828 & n22788 ) ;
  assign n45581 = n16964 ^ n5046 ^ 1'b0 ;
  assign n45582 = n45580 & ~n45581 ;
  assign n45583 = n2985 ^ n662 ^ 1'b0 ;
  assign n45584 = ( ~n5032 & n11928 ) | ( ~n5032 & n45583 ) | ( n11928 & n45583 ) ;
  assign n45585 = n36620 ^ n23260 ^ n5080 ;
  assign n45586 = ~n12140 & n31590 ;
  assign n45587 = n45586 ^ n22308 ^ 1'b0 ;
  assign n45588 = ( n1115 & ~n23147 ) | ( n1115 & n41020 ) | ( ~n23147 & n41020 ) ;
  assign n45589 = n45588 ^ n37569 ^ n24076 ;
  assign n45590 = ( n9304 & n9757 ) | ( n9304 & n29662 ) | ( n9757 & n29662 ) ;
  assign n45591 = ( ~n5052 & n19773 ) | ( ~n5052 & n45590 ) | ( n19773 & n45590 ) ;
  assign n45592 = n45591 ^ n42099 ^ n4568 ;
  assign n45593 = n7944 | n11933 ;
  assign n45594 = ( n9802 & n19596 ) | ( n9802 & ~n45593 ) | ( n19596 & ~n45593 ) ;
  assign n45595 = ( ~n3612 & n3938 ) | ( ~n3612 & n23333 ) | ( n3938 & n23333 ) ;
  assign n45596 = n26823 & n32429 ;
  assign n45597 = ( n21815 & n31728 ) | ( n21815 & n45596 ) | ( n31728 & n45596 ) ;
  assign n45598 = ( n32173 & n40479 ) | ( n32173 & n45597 ) | ( n40479 & n45597 ) ;
  assign n45599 = ( n10019 & n45595 ) | ( n10019 & ~n45598 ) | ( n45595 & ~n45598 ) ;
  assign n45606 = ( n11007 & n11232 ) | ( n11007 & n19617 ) | ( n11232 & n19617 ) ;
  assign n45607 = ( n9848 & n13455 ) | ( n9848 & ~n45606 ) | ( n13455 & ~n45606 ) ;
  assign n45604 = n31484 ^ n726 ^ n666 ;
  assign n45600 = n15439 ^ n9983 ^ n1211 ;
  assign n45601 = n45600 ^ n7360 ^ n3793 ;
  assign n45602 = n45601 ^ n16489 ^ 1'b0 ;
  assign n45603 = n45602 ^ n13900 ^ n5655 ;
  assign n45605 = n45604 ^ n45603 ^ n31221 ;
  assign n45608 = n45607 ^ n45605 ^ n27280 ;
  assign n45609 = ~n10516 & n13059 ;
  assign n45610 = n7795 & n45609 ;
  assign n45611 = n45610 ^ n26281 ^ n1728 ;
  assign n45612 = ( n5847 & ~n8143 ) | ( n5847 & n22822 ) | ( ~n8143 & n22822 ) ;
  assign n45613 = ~n35206 & n45612 ;
  assign n45614 = n45613 ^ n4035 ^ 1'b0 ;
  assign n45615 = n41911 ^ n27446 ^ n872 ;
  assign n45616 = n352 | n29872 ;
  assign n45617 = n45615 | n45616 ;
  assign n45618 = n9800 & n17613 ;
  assign n45619 = n45618 ^ n19063 ^ 1'b0 ;
  assign n45620 = ( n6235 & n33436 ) | ( n6235 & n45619 ) | ( n33436 & n45619 ) ;
  assign n45621 = n45620 ^ n18400 ^ 1'b0 ;
  assign n45622 = n45621 ^ n25697 ^ n2793 ;
  assign n45624 = n12312 | n17132 ;
  assign n45623 = ( n1237 & n22081 ) | ( n1237 & n22925 ) | ( n22081 & n22925 ) ;
  assign n45625 = n45624 ^ n45623 ^ n23739 ;
  assign n45626 = n20090 ^ n15274 ^ n13387 ;
  assign n45627 = ( ~n30950 & n31785 ) | ( ~n30950 & n45615 ) | ( n31785 & n45615 ) ;
  assign n45628 = n45627 ^ n38757 ^ n27129 ;
  assign n45629 = n40357 ^ n30811 ^ n24662 ;
  assign n45630 = ( n8899 & ~n23724 ) | ( n8899 & n41483 ) | ( ~n23724 & n41483 ) ;
  assign n45631 = n8392 & ~n31191 ;
  assign n45632 = n14150 & n45631 ;
  assign n45633 = n3207 & ~n45632 ;
  assign n45634 = n11062 ^ n2594 ^ n830 ;
  assign n45635 = n27072 | n45634 ;
  assign n45636 = n24236 & ~n45635 ;
  assign n45637 = ( ~n1915 & n2619 ) | ( ~n1915 & n45636 ) | ( n2619 & n45636 ) ;
  assign n45638 = n45637 ^ n28097 ^ 1'b0 ;
  assign n45643 = n27117 | n37851 ;
  assign n45644 = n13914 ^ n13587 ^ 1'b0 ;
  assign n45645 = n45643 & n45644 ;
  assign n45639 = n2089 & ~n8279 ;
  assign n45640 = ~n30430 & n45639 ;
  assign n45641 = n45640 ^ n37810 ^ n30830 ;
  assign n45642 = n35096 & n45641 ;
  assign n45646 = n45645 ^ n45642 ^ 1'b0 ;
  assign n45647 = ~n621 & n1460 ;
  assign n45648 = n45647 ^ n20576 ^ 1'b0 ;
  assign n45649 = ( ~n9477 & n19426 ) | ( ~n9477 & n41809 ) | ( n19426 & n41809 ) ;
  assign n45650 = n45649 ^ n27405 ^ n1562 ;
  assign n45651 = n2057 & n9385 ;
  assign n45652 = n30061 ^ n16220 ^ n8934 ;
  assign n45653 = n45652 ^ n26512 ^ n2564 ;
  assign n45654 = n5311 & ~n11737 ;
  assign n45655 = n12158 & n45654 ;
  assign n45656 = n45655 ^ n25637 ^ n23121 ;
  assign n45657 = n20102 ^ n11524 ^ n7567 ;
  assign n45658 = n43991 ^ n27626 ^ n2625 ;
  assign n45659 = n45658 ^ n21995 ^ n12206 ;
  assign n45660 = ~n10277 & n13807 ;
  assign n45661 = n45660 ^ n23363 ^ 1'b0 ;
  assign n45662 = n33201 ^ n29013 ^ 1'b0 ;
  assign n45663 = n45661 & ~n45662 ;
  assign n45664 = n12037 & ~n32755 ;
  assign n45665 = n45664 ^ x133 ^ 1'b0 ;
  assign n45666 = n26856 & ~n45665 ;
  assign n45669 = ( n2348 & n2454 ) | ( n2348 & ~n10644 ) | ( n2454 & ~n10644 ) ;
  assign n45667 = n6223 & ~n18813 ;
  assign n45668 = n45667 ^ n28332 ^ 1'b0 ;
  assign n45670 = n45669 ^ n45668 ^ n34199 ;
  assign n45671 = n45670 ^ n3686 ^ 1'b0 ;
  assign n45672 = ~n9120 & n41601 ;
  assign n45673 = n29076 & n45672 ;
  assign n45674 = n45673 ^ n14760 ^ 1'b0 ;
  assign n45675 = n14424 & n15343 ;
  assign n45676 = n11073 ^ n7635 ^ n6652 ;
  assign n45677 = ( n6653 & n17189 ) | ( n6653 & ~n45676 ) | ( n17189 & ~n45676 ) ;
  assign n45678 = n17795 ^ n9185 ^ 1'b0 ;
  assign n45679 = ( n40642 & n41632 ) | ( n40642 & ~n43535 ) | ( n41632 & ~n43535 ) ;
  assign n45680 = n10683 & n11802 ;
  assign n45681 = n45680 ^ n18201 ^ 1'b0 ;
  assign n45682 = n27857 ^ n25228 ^ x226 ;
  assign n45683 = n30158 ^ n22094 ^ n7135 ;
  assign n45684 = n45683 ^ n9122 ^ 1'b0 ;
  assign n45685 = ( n2161 & n45682 ) | ( n2161 & ~n45684 ) | ( n45682 & ~n45684 ) ;
  assign n45686 = ( n43242 & ~n45681 ) | ( n43242 & n45685 ) | ( ~n45681 & n45685 ) ;
  assign n45687 = n39146 ^ n19826 ^ n1902 ;
  assign n45688 = n45687 ^ n24621 ^ n812 ;
  assign n45689 = ( n34821 & n36818 ) | ( n34821 & ~n45688 ) | ( n36818 & ~n45688 ) ;
  assign n45691 = n43445 ^ n42919 ^ n32772 ;
  assign n45690 = n17049 & ~n42191 ;
  assign n45692 = n45691 ^ n45690 ^ 1'b0 ;
  assign n45693 = ~n12124 & n28052 ;
  assign n45694 = n45693 ^ n13626 ^ 1'b0 ;
  assign n45695 = n17445 | n45694 ;
  assign n45696 = ( n5737 & n26994 ) | ( n5737 & ~n39838 ) | ( n26994 & ~n39838 ) ;
  assign n45697 = ( n11915 & n30558 ) | ( n11915 & n45696 ) | ( n30558 & n45696 ) ;
  assign n45698 = n9251 ^ n5773 ^ 1'b0 ;
  assign n45699 = n45698 ^ n6806 ^ n6433 ;
  assign n45700 = n45699 ^ n1845 ^ 1'b0 ;
  assign n45701 = n1153 | n45700 ;
  assign n45702 = n2745 & ~n5222 ;
  assign n45705 = n12371 ^ n6944 ^ n4154 ;
  assign n45706 = n20630 & n45705 ;
  assign n45703 = n13971 ^ n12722 ^ n9995 ;
  assign n45704 = ( n9492 & n19713 ) | ( n9492 & ~n45703 ) | ( n19713 & ~n45703 ) ;
  assign n45707 = n45706 ^ n45704 ^ 1'b0 ;
  assign n45711 = n11011 ^ n9868 ^ 1'b0 ;
  assign n45712 = ~n25621 & n45711 ;
  assign n45709 = n43975 ^ n30899 ^ n18149 ;
  assign n45708 = n1332 & n17020 ;
  assign n45710 = n45709 ^ n45708 ^ 1'b0 ;
  assign n45713 = n45712 ^ n45710 ^ n6368 ;
  assign n45721 = n44233 ^ n7216 ^ 1'b0 ;
  assign n45719 = ~n28572 & n29327 ;
  assign n45720 = n45719 ^ n9168 ^ 1'b0 ;
  assign n45714 = n18439 ^ n3064 ^ 1'b0 ;
  assign n45715 = ( n6567 & n20590 ) | ( n6567 & ~n45714 ) | ( n20590 & ~n45714 ) ;
  assign n45716 = n1516 & n45715 ;
  assign n45717 = n9619 & ~n17769 ;
  assign n45718 = n45716 & n45717 ;
  assign n45722 = n45721 ^ n45720 ^ n45718 ;
  assign n45723 = n45722 ^ n44707 ^ 1'b0 ;
  assign n45724 = ~n2372 & n44116 ;
  assign n45725 = n12041 ^ n3557 ^ 1'b0 ;
  assign n45726 = ( n7237 & ~n10051 ) | ( n7237 & n13666 ) | ( ~n10051 & n13666 ) ;
  assign n45727 = n45726 ^ n11308 ^ n9177 ;
  assign n45728 = n45727 ^ n24108 ^ 1'b0 ;
  assign n45729 = n45728 ^ n16213 ^ n4923 ;
  assign n45730 = n9007 ^ n6048 ^ n750 ;
  assign n45731 = n12191 & n28465 ;
  assign n45732 = n4897 | n6221 ;
  assign n45733 = n25442 | n45732 ;
  assign n45734 = ( ~n563 & n18837 ) | ( ~n563 & n45733 ) | ( n18837 & n45733 ) ;
  assign n45735 = ~n2164 & n40800 ;
  assign n45736 = ~n12502 & n45735 ;
  assign n45737 = n18262 & n44127 ;
  assign n45738 = n16788 & n45737 ;
  assign n45739 = ( n2152 & n9113 ) | ( n2152 & ~n10259 ) | ( n9113 & ~n10259 ) ;
  assign n45740 = n15088 & n45739 ;
  assign n45741 = n45740 ^ n6395 ^ 1'b0 ;
  assign n45744 = ( n1682 & n21235 ) | ( n1682 & ~n27457 ) | ( n21235 & ~n27457 ) ;
  assign n45742 = n10012 & n15754 ;
  assign n45743 = n32212 & n45742 ;
  assign n45745 = n45744 ^ n45743 ^ n1242 ;
  assign n45746 = n25882 & n41406 ;
  assign n45747 = n44247 ^ n24163 ^ n8699 ;
  assign n45748 = n45747 ^ n26254 ^ n17127 ;
  assign n45749 = ( ~n31635 & n45746 ) | ( ~n31635 & n45748 ) | ( n45746 & n45748 ) ;
  assign n45750 = ( n45741 & n45745 ) | ( n45741 & ~n45749 ) | ( n45745 & ~n45749 ) ;
  assign n45751 = ( ~n6499 & n19606 ) | ( ~n6499 & n42654 ) | ( n19606 & n42654 ) ;
  assign n45752 = ( n4581 & ~n38281 ) | ( n4581 & n45751 ) | ( ~n38281 & n45751 ) ;
  assign n45753 = n44644 & n45752 ;
  assign n45755 = ( n17058 & ~n22719 ) | ( n17058 & n25055 ) | ( ~n22719 & n25055 ) ;
  assign n45754 = n14715 ^ n10409 ^ n8743 ;
  assign n45756 = n45755 ^ n45754 ^ n37863 ;
  assign n45757 = n5754 | n19820 ;
  assign n45758 = n28257 ^ n25179 ^ n6543 ;
  assign n45759 = ~n35069 & n43607 ;
  assign n45760 = n45759 ^ n6955 ^ 1'b0 ;
  assign n45761 = n7385 & n27436 ;
  assign n45762 = ~n38899 & n45761 ;
  assign n45763 = n21076 ^ n4174 ^ n2358 ;
  assign n45764 = ( n7778 & n11943 ) | ( n7778 & n45763 ) | ( n11943 & n45763 ) ;
  assign n45765 = n31274 ^ n5496 ^ 1'b0 ;
  assign n45766 = n16372 ^ n15406 ^ n14708 ;
  assign n45767 = n11058 ^ n9146 ^ 1'b0 ;
  assign n45768 = ( n5579 & n5687 ) | ( n5579 & ~n8165 ) | ( n5687 & ~n8165 ) ;
  assign n45769 = n45768 ^ n3469 ^ 1'b0 ;
  assign n45770 = ( ~n9117 & n43309 ) | ( ~n9117 & n45769 ) | ( n43309 & n45769 ) ;
  assign n45771 = ~n5668 & n45770 ;
  assign n45772 = n27271 ^ n21995 ^ n16322 ;
  assign n45773 = ( n1156 & n4421 ) | ( n1156 & n8142 ) | ( n4421 & n8142 ) ;
  assign n45774 = n24744 ^ n23103 ^ n371 ;
  assign n45775 = n45774 ^ n17465 ^ n1061 ;
  assign n45776 = n45773 & n45775 ;
  assign n45777 = n3820 & n4818 ;
  assign n45778 = n45777 ^ n45673 ^ n45394 ;
  assign n45779 = ( ~n17627 & n21101 ) | ( ~n17627 & n35947 ) | ( n21101 & n35947 ) ;
  assign n45780 = n25261 ^ n3959 ^ n368 ;
  assign n45783 = ( n5875 & n9120 ) | ( n5875 & n18854 ) | ( n9120 & n18854 ) ;
  assign n45781 = n9800 ^ n3362 ^ 1'b0 ;
  assign n45782 = ~n25206 & n45781 ;
  assign n45784 = n45783 ^ n45782 ^ n3654 ;
  assign n45785 = ( n14340 & ~n14406 ) | ( n14340 & n41344 ) | ( ~n14406 & n41344 ) ;
  assign n45786 = n14131 & ~n30893 ;
  assign n45787 = ~n1048 & n45786 ;
  assign n45788 = ( n4651 & n29246 ) | ( n4651 & n38651 ) | ( n29246 & n38651 ) ;
  assign n45789 = ~n37988 & n45788 ;
  assign n45790 = n45789 ^ n28321 ^ 1'b0 ;
  assign n45791 = ( n30305 & ~n45787 ) | ( n30305 & n45790 ) | ( ~n45787 & n45790 ) ;
  assign n45792 = n1449 & ~n6917 ;
  assign n45793 = ~x173 & n45792 ;
  assign n45794 = n2302 & ~n45793 ;
  assign n45795 = n45794 ^ n23290 ^ 1'b0 ;
  assign n45796 = n34926 ^ n12606 ^ 1'b0 ;
  assign n45797 = n13807 & n45796 ;
  assign n45798 = n431 | n2964 ;
  assign n45799 = ( n9496 & ~n11797 ) | ( n9496 & n17730 ) | ( ~n11797 & n17730 ) ;
  assign n45800 = n14948 ^ n8983 ^ 1'b0 ;
  assign n45801 = n26216 & n45800 ;
  assign n45802 = n14420 ^ n8869 ^ n6110 ;
  assign n45803 = ( n9704 & n29867 ) | ( n9704 & ~n45802 ) | ( n29867 & ~n45802 ) ;
  assign n45804 = ( ~n10346 & n11171 ) | ( ~n10346 & n19993 ) | ( n11171 & n19993 ) ;
  assign n45805 = ( n10840 & n15945 ) | ( n10840 & n45804 ) | ( n15945 & n45804 ) ;
  assign n45806 = n27048 ^ n14419 ^ n11845 ;
  assign n45808 = n8826 ^ n3420 ^ n527 ;
  assign n45807 = n13260 | n43951 ;
  assign n45809 = n45808 ^ n45807 ^ 1'b0 ;
  assign n45810 = n5478 | n22453 ;
  assign n45811 = n45810 ^ n7682 ^ 1'b0 ;
  assign n45812 = ~n852 & n30788 ;
  assign n45813 = n19580 ^ n12894 ^ n11962 ;
  assign n45814 = n37392 ^ n30666 ^ n13119 ;
  assign n45815 = ( n13221 & ~n39603 ) | ( n13221 & n45814 ) | ( ~n39603 & n45814 ) ;
  assign n45816 = n45815 ^ n19960 ^ n9655 ;
  assign n45817 = ( n3639 & ~n3878 ) | ( n3639 & n19128 ) | ( ~n3878 & n19128 ) ;
  assign n45818 = n32389 | n45817 ;
  assign n45819 = ( n22097 & ~n22843 ) | ( n22097 & n42731 ) | ( ~n22843 & n42731 ) ;
  assign n45820 = n15720 ^ n3271 ^ n680 ;
  assign n45821 = ( n3786 & n31727 ) | ( n3786 & n41216 ) | ( n31727 & n41216 ) ;
  assign n45822 = ( ~n6362 & n6990 ) | ( ~n6362 & n8071 ) | ( n6990 & n8071 ) ;
  assign n45823 = n45822 ^ n4363 ^ 1'b0 ;
  assign n45824 = n45821 & n45823 ;
  assign n45825 = n45824 ^ n32425 ^ n2636 ;
  assign n45826 = ( ~n35109 & n45820 ) | ( ~n35109 & n45825 ) | ( n45820 & n45825 ) ;
  assign n45827 = ~n10238 & n45826 ;
  assign n45828 = n9274 & n12912 ;
  assign n45829 = n24165 & n45828 ;
  assign n45830 = n33685 ^ n7229 ^ 1'b0 ;
  assign n45831 = n30358 ^ n5579 ^ 1'b0 ;
  assign n45832 = n45831 ^ n6757 ^ n4523 ;
  assign n45833 = n45832 ^ n34097 ^ n25965 ;
  assign n45834 = ( ~n2373 & n11446 ) | ( ~n2373 & n36371 ) | ( n11446 & n36371 ) ;
  assign n45836 = n17090 ^ n3997 ^ 1'b0 ;
  assign n45837 = n45836 ^ n16540 ^ n6285 ;
  assign n45838 = ( n2209 & n16284 ) | ( n2209 & ~n45837 ) | ( n16284 & ~n45837 ) ;
  assign n45835 = ( n2438 & n21450 ) | ( n2438 & n36570 ) | ( n21450 & n36570 ) ;
  assign n45839 = n45838 ^ n45835 ^ n35178 ;
  assign n45840 = ( n1267 & n5358 ) | ( n1267 & n33736 ) | ( n5358 & n33736 ) ;
  assign n45841 = n45840 ^ n23037 ^ n5158 ;
  assign n45842 = n4960 | n37863 ;
  assign n45844 = n1337 & ~n25685 ;
  assign n45843 = n42390 ^ n13807 ^ n7632 ;
  assign n45845 = n45844 ^ n45843 ^ n15249 ;
  assign n45846 = ( n33585 & n38111 ) | ( n33585 & ~n45845 ) | ( n38111 & ~n45845 ) ;
  assign n45847 = n30322 ^ n13309 ^ n7662 ;
  assign n45848 = n19309 ^ n10373 ^ n10329 ;
  assign n45849 = ( ~n13257 & n45847 ) | ( ~n13257 & n45848 ) | ( n45847 & n45848 ) ;
  assign n45850 = n4158 | n45849 ;
  assign n45851 = n45850 ^ n10966 ^ 1'b0 ;
  assign n45852 = x88 & n4467 ;
  assign n45853 = ~n17580 & n45852 ;
  assign n45854 = n14277 ^ n2607 ^ 1'b0 ;
  assign n45855 = n11302 | n45854 ;
  assign n45856 = n45855 ^ n469 ^ n343 ;
  assign n45857 = n21959 & ~n22171 ;
  assign n45858 = ~n45856 & n45857 ;
  assign n45859 = n8722 & n32502 ;
  assign n45860 = n45859 ^ n40760 ^ n5587 ;
  assign n45861 = n39778 ^ n3909 ^ n1469 ;
  assign n45862 = ~n4309 & n23896 ;
  assign n45863 = ~n45861 & n45862 ;
  assign n45864 = ( n12132 & ~n19767 ) | ( n12132 & n45863 ) | ( ~n19767 & n45863 ) ;
  assign n45872 = n3847 ^ n575 ^ 1'b0 ;
  assign n45865 = n668 | n36236 ;
  assign n45866 = n20612 & ~n45865 ;
  assign n45867 = n3726 & ~n45866 ;
  assign n45868 = n45867 ^ n16813 ^ 1'b0 ;
  assign n45869 = ( ~n6550 & n40215 ) | ( ~n6550 & n45868 ) | ( n40215 & n45868 ) ;
  assign n45870 = n45869 ^ n28290 ^ 1'b0 ;
  assign n45871 = n4645 | n45870 ;
  assign n45873 = n45872 ^ n45871 ^ n6408 ;
  assign n45874 = ~n16956 & n22405 ;
  assign n45875 = n9162 & n45874 ;
  assign n45876 = ~n23221 & n36041 ;
  assign n45877 = n45876 ^ n45507 ^ 1'b0 ;
  assign n45878 = ( n32398 & n45875 ) | ( n32398 & n45877 ) | ( n45875 & n45877 ) ;
  assign n45879 = n13008 ^ n11233 ^ 1'b0 ;
  assign n45880 = ~n15199 & n18114 ;
  assign n45881 = ~x125 & n45880 ;
  assign n45882 = n45879 & ~n45881 ;
  assign n45883 = ( ~n4749 & n22743 ) | ( ~n4749 & n45882 ) | ( n22743 & n45882 ) ;
  assign n45884 = n25716 | n45883 ;
  assign n45885 = ( n1840 & ~n7857 ) | ( n1840 & n11117 ) | ( ~n7857 & n11117 ) ;
  assign n45886 = n22983 & ~n45885 ;
  assign n45887 = ~n27434 & n45886 ;
  assign n45888 = n24044 ^ n17171 ^ 1'b0 ;
  assign n45889 = n45888 ^ n33370 ^ 1'b0 ;
  assign n45890 = n39621 & ~n45889 ;
  assign n45891 = ~n3646 & n31136 ;
  assign n45892 = n45891 ^ n29857 ^ n29261 ;
  assign n45893 = ( ~n5352 & n13186 ) | ( ~n5352 & n45892 ) | ( n13186 & n45892 ) ;
  assign n45894 = n18742 & n24957 ;
  assign n45895 = ~n33279 & n45894 ;
  assign n45896 = ( n11207 & n17498 ) | ( n11207 & n45895 ) | ( n17498 & n45895 ) ;
  assign n45897 = ( n9301 & n32846 ) | ( n9301 & ~n45896 ) | ( n32846 & ~n45896 ) ;
  assign n45898 = n30973 ^ n26771 ^ 1'b0 ;
  assign n45899 = n5987 | n38281 ;
  assign n45900 = n3169 | n45899 ;
  assign n45901 = n45900 ^ n28094 ^ 1'b0 ;
  assign n45902 = n15986 ^ n15968 ^ 1'b0 ;
  assign n45903 = n2570 & n4037 ;
  assign n45904 = n45903 ^ n3934 ^ 1'b0 ;
  assign n45905 = n45904 ^ n6498 ^ 1'b0 ;
  assign n45906 = ~n1656 & n9792 ;
  assign n45907 = ~n45558 & n45906 ;
  assign n45912 = ( n7106 & n12948 ) | ( n7106 & n13876 ) | ( n12948 & n13876 ) ;
  assign n45913 = ( n41244 & n43268 ) | ( n41244 & ~n45912 ) | ( n43268 & ~n45912 ) ;
  assign n45908 = n13071 & n35555 ;
  assign n45909 = n17641 ^ n13807 ^ n9067 ;
  assign n45910 = ( n7206 & n17007 ) | ( n7206 & ~n45909 ) | ( n17007 & ~n45909 ) ;
  assign n45911 = ( n580 & ~n45908 ) | ( n580 & n45910 ) | ( ~n45908 & n45910 ) ;
  assign n45914 = n45913 ^ n45911 ^ n33292 ;
  assign n45915 = ( n12103 & ~n17141 ) | ( n12103 & n22953 ) | ( ~n17141 & n22953 ) ;
  assign n45916 = ~n24763 & n29717 ;
  assign n45917 = n26937 & ~n45916 ;
  assign n45918 = ( n29024 & n45915 ) | ( n29024 & ~n45917 ) | ( n45915 & ~n45917 ) ;
  assign n45920 = n13949 | n36132 ;
  assign n45921 = n13941 | n45920 ;
  assign n45919 = ~n9180 & n22562 ;
  assign n45922 = n45921 ^ n45919 ^ n3157 ;
  assign n45923 = n23234 ^ n6947 ^ n3184 ;
  assign n45924 = n45923 ^ n3041 ^ n2198 ;
  assign n45925 = n4607 | n16692 ;
  assign n45926 = n45925 ^ n22474 ^ 1'b0 ;
  assign n45927 = n4908 | n5396 ;
  assign n45928 = n45927 ^ n22422 ^ 1'b0 ;
  assign n45929 = n45928 ^ n2890 ^ 1'b0 ;
  assign n45930 = n42791 & ~n45929 ;
  assign n45931 = n21160 ^ n11752 ^ 1'b0 ;
  assign n45932 = n22950 & ~n45931 ;
  assign n45933 = n45932 ^ n2942 ^ 1'b0 ;
  assign n45935 = n25844 | n43975 ;
  assign n45936 = n16433 & ~n45935 ;
  assign n45934 = n22106 & n35918 ;
  assign n45937 = n45936 ^ n45934 ^ 1'b0 ;
  assign n45938 = n32278 ^ n11621 ^ 1'b0 ;
  assign n45940 = ( n13181 & n15375 ) | ( n13181 & ~n22665 ) | ( n15375 & ~n22665 ) ;
  assign n45941 = ( n19382 & n21113 ) | ( n19382 & n45940 ) | ( n21113 & n45940 ) ;
  assign n45939 = ( n1616 & n19995 ) | ( n1616 & ~n36883 ) | ( n19995 & ~n36883 ) ;
  assign n45942 = n45941 ^ n45939 ^ n20904 ;
  assign n45943 = n12379 ^ n9997 ^ n835 ;
  assign n45944 = n14379 & n19019 ;
  assign n45946 = n41216 ^ n24310 ^ 1'b0 ;
  assign n45945 = n26356 & n40760 ;
  assign n45947 = n45946 ^ n45945 ^ 1'b0 ;
  assign n45948 = n44795 ^ n9041 ^ 1'b0 ;
  assign n45949 = n33256 ^ n270 ^ 1'b0 ;
  assign n45950 = n4603 | n45949 ;
  assign n45951 = ( n17562 & n22549 ) | ( n17562 & n25819 ) | ( n22549 & n25819 ) ;
  assign n45952 = ( n14069 & n38802 ) | ( n14069 & ~n42955 ) | ( n38802 & ~n42955 ) ;
  assign n45953 = n7246 | n30868 ;
  assign n45954 = n16976 & ~n45953 ;
  assign n45955 = ( n16240 & n37396 ) | ( n16240 & ~n45954 ) | ( n37396 & ~n45954 ) ;
  assign n45956 = n45955 ^ n26668 ^ n3717 ;
  assign n45957 = n9096 | n31229 ;
  assign n45958 = n45956 & ~n45957 ;
  assign n45961 = n7891 | n9719 ;
  assign n45962 = n45961 ^ n9261 ^ 1'b0 ;
  assign n45963 = n992 & n45962 ;
  assign n45964 = n45963 ^ n15172 ^ n8200 ;
  assign n45959 = ( ~n18771 & n31839 ) | ( ~n18771 & n42070 ) | ( n31839 & n42070 ) ;
  assign n45960 = n10991 & ~n45959 ;
  assign n45965 = n45964 ^ n45960 ^ 1'b0 ;
  assign n45967 = n6366 & n26381 ;
  assign n45968 = n45967 ^ n3617 ^ 1'b0 ;
  assign n45966 = n42142 ^ n35231 ^ n5157 ;
  assign n45969 = n45968 ^ n45966 ^ 1'b0 ;
  assign n45970 = n42886 ^ n21255 ^ 1'b0 ;
  assign n45971 = ( n8723 & n15218 ) | ( n8723 & ~n20542 ) | ( n15218 & ~n20542 ) ;
  assign n45972 = ( ~n25284 & n28351 ) | ( ~n25284 & n32664 ) | ( n28351 & n32664 ) ;
  assign n45975 = n3932 & n18372 ;
  assign n45973 = n536 | n10370 ;
  assign n45974 = n34275 | n45973 ;
  assign n45976 = n45975 ^ n45974 ^ n35227 ;
  assign n45977 = n7070 & n14541 ;
  assign n45978 = ( n10060 & n28492 ) | ( n10060 & ~n40808 ) | ( n28492 & ~n40808 ) ;
  assign n45979 = ( ~n12150 & n25188 ) | ( ~n12150 & n45978 ) | ( n25188 & n45978 ) ;
  assign n45980 = n15174 ^ n8200 ^ n1992 ;
  assign n45981 = n21538 ^ n17673 ^ n12031 ;
  assign n45982 = ( n33156 & n45980 ) | ( n33156 & n45981 ) | ( n45980 & n45981 ) ;
  assign n45989 = n19494 ^ n7880 ^ 1'b0 ;
  assign n45984 = n2737 ^ n2174 ^ 1'b0 ;
  assign n45985 = n3838 & n45984 ;
  assign n45986 = n28239 ^ n14157 ^ n9602 ;
  assign n45987 = n45985 & ~n45986 ;
  assign n45983 = n16767 | n44735 ;
  assign n45988 = n45987 ^ n45983 ^ 1'b0 ;
  assign n45990 = n45989 ^ n45988 ^ n7551 ;
  assign n45991 = n45990 ^ n17736 ^ n860 ;
  assign n45992 = n25400 ^ n1768 ^ 1'b0 ;
  assign n45993 = n35689 & n45992 ;
  assign n45994 = n21292 ^ n4383 ^ n1528 ;
  assign n45995 = ~n10723 & n13936 ;
  assign n45996 = n5104 | n45995 ;
  assign n45997 = n41485 ^ n4277 ^ 1'b0 ;
  assign n45998 = n24644 | n45997 ;
  assign n45999 = ( ~n19503 & n29497 ) | ( ~n19503 & n30330 ) | ( n29497 & n30330 ) ;
  assign n46000 = n9350 & ~n10285 ;
  assign n46001 = ( ~n22831 & n36675 ) | ( ~n22831 & n46000 ) | ( n36675 & n46000 ) ;
  assign n46002 = n45999 | n46001 ;
  assign n46003 = n43784 ^ n20074 ^ 1'b0 ;
  assign n46004 = n23088 ^ n4743 ^ n2058 ;
  assign n46005 = n35283 & n46004 ;
  assign n46006 = n46005 ^ n30404 ^ 1'b0 ;
  assign n46007 = n32405 ^ n20062 ^ n12192 ;
  assign n46008 = n21039 ^ n20421 ^ 1'b0 ;
  assign n46009 = n40308 & n43317 ;
  assign n46010 = n41239 ^ n17130 ^ n12319 ;
  assign n46011 = n15856 | n46010 ;
  assign n46012 = n27997 ^ n12825 ^ n7128 ;
  assign n46013 = n46011 | n46012 ;
  assign n46014 = n18467 & ~n45165 ;
  assign n46015 = ~n416 & n46014 ;
  assign n46016 = ( n20870 & n31467 ) | ( n20870 & ~n38890 ) | ( n31467 & ~n38890 ) ;
  assign n46017 = n42020 ^ n9183 ^ 1'b0 ;
  assign n46018 = n7445 & n46017 ;
  assign n46019 = ( n18253 & n26322 ) | ( n18253 & ~n46018 ) | ( n26322 & ~n46018 ) ;
  assign n46020 = n4679 & ~n11052 ;
  assign n46021 = ~n12189 & n46020 ;
  assign n46022 = n46021 ^ n18014 ^ 1'b0 ;
  assign n46023 = n27257 ^ n10557 ^ 1'b0 ;
  assign n46026 = ( ~n745 & n6324 ) | ( ~n745 & n13117 ) | ( n6324 & n13117 ) ;
  assign n46027 = n46026 ^ n20373 ^ n14644 ;
  assign n46028 = n46027 ^ n45292 ^ n26610 ;
  assign n46024 = n23698 | n37248 ;
  assign n46025 = ( n7270 & ~n9315 ) | ( n7270 & n46024 ) | ( ~n9315 & n46024 ) ;
  assign n46029 = n46028 ^ n46025 ^ n16373 ;
  assign n46030 = n22593 | n46029 ;
  assign n46034 = n2542 & n4635 ;
  assign n46031 = n8588 & n10130 ;
  assign n46032 = n46031 ^ n15100 ^ n11983 ;
  assign n46033 = n46032 ^ n1534 ^ 1'b0 ;
  assign n46035 = n46034 ^ n46033 ^ n6763 ;
  assign n46036 = n8520 ^ n6682 ^ 1'b0 ;
  assign n46037 = n17182 & ~n46036 ;
  assign n46038 = ( n13265 & n18469 ) | ( n13265 & ~n36808 ) | ( n18469 & ~n36808 ) ;
  assign n46039 = n37043 ^ n6775 ^ 1'b0 ;
  assign n46040 = n46038 | n46039 ;
  assign n46041 = n26558 & n45072 ;
  assign n46042 = ~n15062 & n22540 ;
  assign n46043 = ~n9914 & n46042 ;
  assign n46044 = n37183 ^ n31893 ^ n29595 ;
  assign n46046 = n32354 ^ n29304 ^ n2847 ;
  assign n46045 = n42252 ^ n38632 ^ 1'b0 ;
  assign n46047 = n46046 ^ n46045 ^ n9159 ;
  assign n46048 = n13747 ^ n13562 ^ n9278 ;
  assign n46051 = n20002 ^ n9019 ^ 1'b0 ;
  assign n46049 = n24228 | n29393 ;
  assign n46050 = n46049 ^ n42488 ^ n18234 ;
  assign n46052 = n46051 ^ n46050 ^ n3138 ;
  assign n46053 = n17062 & n33848 ;
  assign n46054 = ( n28446 & n29847 ) | ( n28446 & n46053 ) | ( n29847 & n46053 ) ;
  assign n46055 = n46054 ^ n32282 ^ n24823 ;
  assign n46056 = n15638 ^ n14073 ^ 1'b0 ;
  assign n46057 = n12296 & ~n46056 ;
  assign n46058 = ( n1058 & n21870 ) | ( n1058 & ~n46057 ) | ( n21870 & ~n46057 ) ;
  assign n46059 = ( n7144 & ~n13916 ) | ( n7144 & n24390 ) | ( ~n13916 & n24390 ) ;
  assign n46060 = n17009 & n46059 ;
  assign n46061 = n46060 ^ n17357 ^ 1'b0 ;
  assign n46062 = n12485 ^ n944 ^ 1'b0 ;
  assign n46063 = n20077 ^ n9885 ^ 1'b0 ;
  assign n46064 = n46062 & ~n46063 ;
  assign n46065 = n29271 ^ n6238 ^ 1'b0 ;
  assign n46067 = n12819 | n18531 ;
  assign n46068 = n19967 & ~n46067 ;
  assign n46066 = n42062 ^ n18775 ^ n16736 ;
  assign n46069 = n46068 ^ n46066 ^ n25882 ;
  assign n46070 = n42237 ^ n19666 ^ n2362 ;
  assign n46071 = ( n2077 & n9070 ) | ( n2077 & ~n35886 ) | ( n9070 & ~n35886 ) ;
  assign n46072 = ( n15825 & ~n42162 ) | ( n15825 & n46071 ) | ( ~n42162 & n46071 ) ;
  assign n46073 = n25555 ^ n4391 ^ 1'b0 ;
  assign n46074 = n28997 ^ n19409 ^ n6608 ;
  assign n46075 = n6409 ^ n1748 ^ 1'b0 ;
  assign n46076 = n14933 & n46075 ;
  assign n46078 = ( n21056 & n32999 ) | ( n21056 & n36868 ) | ( n32999 & n36868 ) ;
  assign n46079 = n18246 & n46078 ;
  assign n46077 = n21978 & ~n27780 ;
  assign n46080 = n46079 ^ n46077 ^ 1'b0 ;
  assign n46081 = n16991 ^ n14271 ^ 1'b0 ;
  assign n46082 = n32819 ^ n10566 ^ 1'b0 ;
  assign n46083 = n46081 & n46082 ;
  assign n46084 = n22288 ^ n9679 ^ 1'b0 ;
  assign n46086 = n38894 ^ n32882 ^ n9117 ;
  assign n46085 = ( n736 & n26663 ) | ( n736 & n40521 ) | ( n26663 & n40521 ) ;
  assign n46087 = n46086 ^ n46085 ^ 1'b0 ;
  assign n46088 = n4336 ^ x133 ^ 1'b0 ;
  assign n46089 = ~n18636 & n46088 ;
  assign n46090 = n46089 ^ n45987 ^ n25729 ;
  assign n46091 = n21842 ^ n3965 ^ 1'b0 ;
  assign n46092 = n45284 ^ n37341 ^ 1'b0 ;
  assign n46093 = n36757 ^ n13199 ^ 1'b0 ;
  assign n46094 = ~n46092 & n46093 ;
  assign n46095 = ( n12830 & ~n46091 ) | ( n12830 & n46094 ) | ( ~n46091 & n46094 ) ;
  assign n46096 = n36690 ^ n32643 ^ n30752 ;
  assign n46097 = n32322 & ~n41244 ;
  assign n46098 = n1725 & n46097 ;
  assign n46099 = n8881 ^ n6670 ^ n4142 ;
  assign n46100 = n15705 & ~n46099 ;
  assign n46101 = n41370 & n46100 ;
  assign n46102 = ( n5411 & ~n10414 ) | ( n5411 & n19241 ) | ( ~n10414 & n19241 ) ;
  assign n46103 = n37672 ^ n19584 ^ n5719 ;
  assign n46104 = n11110 & n17426 ;
  assign n46105 = n22710 & n46104 ;
  assign n46106 = n42709 ^ n10972 ^ n275 ;
  assign n46107 = ~n46105 & n46106 ;
  assign n46108 = n9323 & ~n41509 ;
  assign n46109 = n23343 ^ n22907 ^ n16104 ;
  assign n46110 = n46109 ^ n39880 ^ n7068 ;
  assign n46111 = ( ~n23473 & n46108 ) | ( ~n23473 & n46110 ) | ( n46108 & n46110 ) ;
  assign n46112 = ~n434 & n3188 ;
  assign n46113 = n329 & n46112 ;
  assign n46114 = n17203 & n24922 ;
  assign n46115 = ~n2659 & n46114 ;
  assign n46116 = ( n11055 & n46113 ) | ( n11055 & ~n46115 ) | ( n46113 & ~n46115 ) ;
  assign n46118 = n8867 | n9254 ;
  assign n46119 = n46118 ^ n33935 ^ 1'b0 ;
  assign n46120 = n19112 & ~n46119 ;
  assign n46117 = n37179 ^ n23737 ^ 1'b0 ;
  assign n46121 = n46120 ^ n46117 ^ 1'b0 ;
  assign n46122 = n24976 | n46121 ;
  assign n46126 = ( n13139 & n28234 ) | ( n13139 & n34493 ) | ( n28234 & n34493 ) ;
  assign n46123 = n38449 ^ n25128 ^ n21491 ;
  assign n46124 = n36621 & n46123 ;
  assign n46125 = n31283 & n46124 ;
  assign n46127 = n46126 ^ n46125 ^ 1'b0 ;
  assign n46128 = n15659 ^ n1035 ^ 1'b0 ;
  assign n46129 = n46128 ^ n44319 ^ n22898 ;
  assign n46130 = n36237 ^ n35480 ^ n7761 ;
  assign n46131 = ( n9036 & n14668 ) | ( n9036 & n33543 ) | ( n14668 & n33543 ) ;
  assign n46132 = n17069 & n20728 ;
  assign n46133 = n46132 ^ n5457 ^ 1'b0 ;
  assign n46134 = n24711 ^ n19971 ^ 1'b0 ;
  assign n46135 = ~n46133 & n46134 ;
  assign n46136 = n46135 ^ n7730 ^ n4798 ;
  assign n46137 = n24321 ^ n23364 ^ n18762 ;
  assign n46138 = ( n4099 & n46136 ) | ( n4099 & n46137 ) | ( n46136 & n46137 ) ;
  assign n46139 = ~n16071 & n16587 ;
  assign n46140 = n46139 ^ n44290 ^ 1'b0 ;
  assign n46141 = ( n1467 & n39930 ) | ( n1467 & n46140 ) | ( n39930 & n46140 ) ;
  assign n46142 = n46141 ^ n30821 ^ 1'b0 ;
  assign n46143 = ~n26007 & n40580 ;
  assign n46145 = n19756 ^ n1162 ^ 1'b0 ;
  assign n46144 = n15819 & n24000 ;
  assign n46146 = n46145 ^ n46144 ^ n24166 ;
  assign n46147 = n21687 ^ n13273 ^ 1'b0 ;
  assign n46148 = n6984 & ~n46147 ;
  assign n46149 = n46148 ^ n38365 ^ n3663 ;
  assign n46150 = n32173 ^ n861 ^ 1'b0 ;
  assign n46151 = n25849 ^ n7905 ^ 1'b0 ;
  assign n46152 = n46151 ^ n41397 ^ n23157 ;
  assign n46153 = ( n28721 & n31566 ) | ( n28721 & n33216 ) | ( n31566 & n33216 ) ;
  assign n46154 = ( n17002 & ~n18170 ) | ( n17002 & n46153 ) | ( ~n18170 & n46153 ) ;
  assign n46155 = n38818 ^ n36167 ^ 1'b0 ;
  assign n46156 = n22376 & ~n46155 ;
  assign n46157 = n14471 ^ n5824 ^ n603 ;
  assign n46158 = n4923 & ~n46157 ;
  assign n46159 = n42099 & n46158 ;
  assign n46161 = n26653 ^ n9542 ^ n8977 ;
  assign n46160 = n3774 & ~n15271 ;
  assign n46162 = n46161 ^ n46160 ^ 1'b0 ;
  assign n46163 = ( n9079 & n26969 ) | ( n9079 & ~n45278 ) | ( n26969 & ~n45278 ) ;
  assign n46164 = ( ~n4712 & n4853 ) | ( ~n4712 & n32746 ) | ( n4853 & n32746 ) ;
  assign n46165 = n46164 ^ n42642 ^ n27662 ;
  assign n46166 = n41198 ^ n32659 ^ n4480 ;
  assign n46167 = n28101 & n28397 ;
  assign n46168 = ( n3200 & ~n3767 ) | ( n3200 & n46167 ) | ( ~n3767 & n46167 ) ;
  assign n46169 = n38713 ^ n20412 ^ n19603 ;
  assign n46170 = n46169 ^ n1125 ^ x135 ;
  assign n46172 = n17889 ^ n13217 ^ n4707 ;
  assign n46171 = n21100 & ~n27248 ;
  assign n46173 = n46172 ^ n46171 ^ 1'b0 ;
  assign n46174 = n9533 | n24675 ;
  assign n46175 = n46174 ^ n11082 ^ 1'b0 ;
  assign n46176 = n21265 & ~n46175 ;
  assign n46177 = n10411 & ~n17885 ;
  assign n46178 = n26308 & n46177 ;
  assign n46179 = n8932 & ~n35450 ;
  assign n46180 = n46178 & n46179 ;
  assign n46181 = ( ~n22685 & n26637 ) | ( ~n22685 & n34780 ) | ( n26637 & n34780 ) ;
  assign n46182 = n45669 ^ n26864 ^ n22524 ;
  assign n46183 = ( ~n1453 & n7672 ) | ( ~n1453 & n46182 ) | ( n7672 & n46182 ) ;
  assign n46184 = n32402 & ~n46183 ;
  assign n46185 = ( n34853 & n43114 ) | ( n34853 & n46184 ) | ( n43114 & n46184 ) ;
  assign n46186 = ~n3019 & n6577 ;
  assign n46187 = ~n1817 & n46186 ;
  assign n46188 = ( n13232 & n42041 ) | ( n13232 & n46187 ) | ( n42041 & n46187 ) ;
  assign n46189 = ~n10256 & n40647 ;
  assign n46190 = n46189 ^ n5214 ^ 1'b0 ;
  assign n46191 = n46190 ^ n44278 ^ n11637 ;
  assign n46192 = n36277 ^ n34367 ^ n32653 ;
  assign n46193 = n5684 ^ n3060 ^ 1'b0 ;
  assign n46194 = n46193 ^ n29983 ^ n25004 ;
  assign n46195 = ( ~n44649 & n46192 ) | ( ~n44649 & n46194 ) | ( n46192 & n46194 ) ;
  assign n46196 = n9666 & n25791 ;
  assign n46197 = n46196 ^ n1015 ^ 1'b0 ;
  assign n46198 = ~n6978 & n46197 ;
  assign n46199 = ( n1218 & ~n16255 ) | ( n1218 & n32304 ) | ( ~n16255 & n32304 ) ;
  assign n46200 = n46199 ^ n12955 ^ 1'b0 ;
  assign n46201 = n46198 & n46200 ;
  assign n46202 = n25775 ^ n24891 ^ n24204 ;
  assign n46203 = n42078 ^ n25971 ^ 1'b0 ;
  assign n46204 = n46202 & n46203 ;
  assign n46205 = n4375 & ~n40656 ;
  assign n46206 = n30601 & n46205 ;
  assign n46209 = n39868 ^ n16336 ^ n5107 ;
  assign n46207 = n28194 ^ n18377 ^ n8297 ;
  assign n46208 = n3142 & n46207 ;
  assign n46210 = n46209 ^ n46208 ^ 1'b0 ;
  assign n46211 = ~n5796 & n38026 ;
  assign n46212 = ( n18462 & ~n39602 ) | ( n18462 & n43666 ) | ( ~n39602 & n43666 ) ;
  assign n46213 = ( n30191 & n32536 ) | ( n30191 & ~n45558 ) | ( n32536 & ~n45558 ) ;
  assign n46214 = ( ~n9877 & n17917 ) | ( ~n9877 & n27218 ) | ( n17917 & n27218 ) ;
  assign n46215 = n6131 | n28561 ;
  assign n46216 = ( n5609 & ~n18352 ) | ( n5609 & n23707 ) | ( ~n18352 & n23707 ) ;
  assign n46217 = ( n2113 & n16893 ) | ( n2113 & ~n46216 ) | ( n16893 & ~n46216 ) ;
  assign n46218 = n46217 ^ n829 ^ 1'b0 ;
  assign n46219 = n46215 & n46218 ;
  assign n46220 = n46219 ^ n16745 ^ n14863 ;
  assign n46221 = ( n5578 & n8462 ) | ( n5578 & n41274 ) | ( n8462 & n41274 ) ;
  assign n46222 = n24265 & n46221 ;
  assign n46223 = n22048 & ~n22559 ;
  assign n46224 = n46223 ^ n6685 ^ 1'b0 ;
  assign n46225 = n46224 ^ n7685 ^ 1'b0 ;
  assign n46226 = ~n30444 & n46225 ;
  assign n46227 = n20431 & ~n29530 ;
  assign n46228 = n40220 & ~n46227 ;
  assign n46229 = n25034 & n46228 ;
  assign n46231 = n38158 ^ n32476 ^ n2145 ;
  assign n46230 = ~n7235 & n31030 ;
  assign n46232 = n46231 ^ n46230 ^ 1'b0 ;
  assign n46233 = ( n1991 & n5950 ) | ( n1991 & ~n37609 ) | ( n5950 & ~n37609 ) ;
  assign n46234 = n38990 ^ n29835 ^ n22481 ;
  assign n46239 = n34665 ^ n7514 ^ n5938 ;
  assign n46238 = ( ~n1952 & n15839 ) | ( ~n1952 & n38781 ) | ( n15839 & n38781 ) ;
  assign n46237 = ( n3798 & n7700 ) | ( n3798 & n10549 ) | ( n7700 & n10549 ) ;
  assign n46240 = n46239 ^ n46238 ^ n46237 ;
  assign n46235 = n6356 ^ n3897 ^ 1'b0 ;
  assign n46236 = ~n37525 & n46235 ;
  assign n46241 = n46240 ^ n46236 ^ 1'b0 ;
  assign n46242 = ( n46233 & n46234 ) | ( n46233 & ~n46241 ) | ( n46234 & ~n46241 ) ;
  assign n46244 = n4850 | n13163 ;
  assign n46245 = n13342 & ~n46244 ;
  assign n46243 = ( n7056 & ~n25655 ) | ( n7056 & n30526 ) | ( ~n25655 & n30526 ) ;
  assign n46246 = n46245 ^ n46243 ^ 1'b0 ;
  assign n46247 = n42096 ^ n32769 ^ n5588 ;
  assign n46248 = n2258 & n46247 ;
  assign n46249 = n46248 ^ n30891 ^ 1'b0 ;
  assign n46250 = n13684 & n46249 ;
  assign n46251 = ( n25535 & n37414 ) | ( n25535 & ~n39103 ) | ( n37414 & ~n39103 ) ;
  assign n46252 = ( n1996 & ~n14352 ) | ( n1996 & n18944 ) | ( ~n14352 & n18944 ) ;
  assign n46253 = n26176 | n46252 ;
  assign n46254 = n7313 | n46253 ;
  assign n46255 = n11155 | n46254 ;
  assign n46256 = ( n2357 & n2759 ) | ( n2357 & ~n43133 ) | ( n2759 & ~n43133 ) ;
  assign n46257 = ( n22816 & n43007 ) | ( n22816 & ~n46256 ) | ( n43007 & ~n46256 ) ;
  assign n46258 = n43889 ^ n34110 ^ n23537 ;
  assign n46259 = n12306 & n21810 ;
  assign n46260 = ~n11693 & n46259 ;
  assign n46261 = ( n8669 & n41431 ) | ( n8669 & n46260 ) | ( n41431 & n46260 ) ;
  assign n46262 = x243 & ~n46261 ;
  assign n46263 = n46262 ^ n43302 ^ 1'b0 ;
  assign n46264 = n9611 ^ n5312 ^ n4859 ;
  assign n46265 = n28424 ^ n3876 ^ 1'b0 ;
  assign n46266 = n46264 | n46265 ;
  assign n46267 = n14062 | n46266 ;
  assign n46268 = n11798 | n19294 ;
  assign n46269 = n24175 ^ n15315 ^ n14538 ;
  assign n46270 = n46269 ^ n22310 ^ n6985 ;
  assign n46271 = ~n5039 & n46270 ;
  assign n46272 = n37245 ^ n35194 ^ n18149 ;
  assign n46273 = ~n13452 & n18200 ;
  assign n46274 = n12316 & n17867 ;
  assign n46275 = ( n3502 & n22230 ) | ( n3502 & ~n46274 ) | ( n22230 & ~n46274 ) ;
  assign n46276 = n4516 & n35917 ;
  assign n46277 = n3487 & n46276 ;
  assign n46278 = n42547 ^ n18175 ^ 1'b0 ;
  assign n46279 = n4417 ^ n592 ^ 1'b0 ;
  assign n46280 = n46278 | n46279 ;
  assign n46281 = n43827 ^ n33787 ^ n1376 ;
  assign n46282 = ( n40737 & ~n40783 ) | ( n40737 & n46281 ) | ( ~n40783 & n46281 ) ;
  assign n46283 = n27807 ^ n4340 ^ 1'b0 ;
  assign n46284 = ( n1651 & ~n7172 ) | ( n1651 & n13325 ) | ( ~n7172 & n13325 ) ;
  assign n46285 = ( ~n9920 & n37788 ) | ( ~n9920 & n46284 ) | ( n37788 & n46284 ) ;
  assign n46286 = ( n19729 & n34887 ) | ( n19729 & ~n41425 ) | ( n34887 & ~n41425 ) ;
  assign n46287 = ( n6745 & n6898 ) | ( n6745 & ~n13799 ) | ( n6898 & ~n13799 ) ;
  assign n46288 = n46287 ^ n39947 ^ 1'b0 ;
  assign n46289 = n28301 ^ n1664 ^ 1'b0 ;
  assign n46290 = n39979 & n46289 ;
  assign n46291 = ( ~n4346 & n4853 ) | ( ~n4346 & n34433 ) | ( n4853 & n34433 ) ;
  assign n46292 = n45513 ^ n33476 ^ 1'b0 ;
  assign n46293 = n46291 & ~n46292 ;
  assign n46294 = n42509 ^ n34699 ^ n21584 ;
  assign n46295 = n43635 ^ n36984 ^ n4003 ;
  assign n46296 = n46295 ^ n21075 ^ n7774 ;
  assign n46297 = n39883 ^ n36353 ^ n600 ;
  assign n46298 = n44831 ^ n29911 ^ 1'b0 ;
  assign n46299 = n46298 ^ n15049 ^ n2309 ;
  assign n46300 = ( ~n2123 & n31628 ) | ( ~n2123 & n39213 ) | ( n31628 & n39213 ) ;
  assign n46301 = n1709 | n37338 ;
  assign n46302 = n46300 & ~n46301 ;
  assign n46303 = n45912 ^ x67 ^ 1'b0 ;
  assign n46304 = n35797 ^ n11910 ^ 1'b0 ;
  assign n46305 = ( ~n33245 & n46303 ) | ( ~n33245 & n46304 ) | ( n46303 & n46304 ) ;
  assign n46306 = ~n1088 & n1090 ;
  assign n46307 = ~n16186 & n46306 ;
  assign n46308 = ~n4069 & n46307 ;
  assign n46309 = ( ~n14653 & n34316 ) | ( ~n14653 & n39495 ) | ( n34316 & n39495 ) ;
  assign n46310 = n38415 ^ n33903 ^ n578 ;
  assign n46311 = ( n20594 & ~n45231 ) | ( n20594 & n46310 ) | ( ~n45231 & n46310 ) ;
  assign n46312 = ~n11511 & n14439 ;
  assign n46313 = n10465 & n46312 ;
  assign n46314 = n46313 ^ n13639 ^ n6218 ;
  assign n46315 = n18971 ^ n11845 ^ n5705 ;
  assign n46316 = ( n18206 & n22595 ) | ( n18206 & n46315 ) | ( n22595 & n46315 ) ;
  assign n46317 = n4351 & ~n32922 ;
  assign n46318 = ( n7700 & n9913 ) | ( n7700 & n31646 ) | ( n9913 & n31646 ) ;
  assign n46319 = n46318 ^ n23045 ^ 1'b0 ;
  assign n46320 = n11553 & ~n46319 ;
  assign n46321 = n34293 ^ n15217 ^ 1'b0 ;
  assign n46322 = n5446 | n46321 ;
  assign n46323 = n7137 & ~n46322 ;
  assign n46324 = n46323 ^ n16197 ^ 1'b0 ;
  assign n46326 = ~n517 & n13789 ;
  assign n46325 = ( n23363 & n36248 ) | ( n23363 & n37495 ) | ( n36248 & n37495 ) ;
  assign n46327 = n46326 ^ n46325 ^ n7329 ;
  assign n46328 = ( n9605 & n11167 ) | ( n9605 & ~n20657 ) | ( n11167 & ~n20657 ) ;
  assign n46329 = ~n8116 & n35671 ;
  assign n46330 = n46329 ^ n41800 ^ n8071 ;
  assign n46331 = ( ~n2501 & n46328 ) | ( ~n2501 & n46330 ) | ( n46328 & n46330 ) ;
  assign n46332 = n28487 ^ n3372 ^ 1'b0 ;
  assign n46333 = n16223 ^ n14336 ^ 1'b0 ;
  assign n46334 = n24018 | n46333 ;
  assign n46335 = ~n21540 & n46334 ;
  assign n46336 = n18069 & ~n19962 ;
  assign n46337 = n46336 ^ n30345 ^ 1'b0 ;
  assign n46338 = ( n11428 & n41509 ) | ( n11428 & ~n46337 ) | ( n41509 & ~n46337 ) ;
  assign n46339 = ( n5529 & n24642 ) | ( n5529 & ~n44342 ) | ( n24642 & ~n44342 ) ;
  assign n46340 = n46339 ^ n32405 ^ n4600 ;
  assign n46341 = n46340 ^ n36239 ^ 1'b0 ;
  assign n46342 = ~n16919 & n17121 ;
  assign n46345 = ( ~n7152 & n17241 ) | ( ~n7152 & n18751 ) | ( n17241 & n18751 ) ;
  assign n46344 = n9703 | n25599 ;
  assign n46346 = n46345 ^ n46344 ^ 1'b0 ;
  assign n46343 = n7491 | n32764 ;
  assign n46347 = n46346 ^ n46343 ^ 1'b0 ;
  assign n46348 = n12271 & ~n38068 ;
  assign n46349 = ~n15608 & n46348 ;
  assign n46350 = n27202 ^ n3606 ^ 1'b0 ;
  assign n46351 = n23539 | n46350 ;
  assign n46352 = ( n13176 & ~n15215 ) | ( n13176 & n32031 ) | ( ~n15215 & n32031 ) ;
  assign n46353 = ( n3844 & ~n9742 ) | ( n3844 & n46352 ) | ( ~n9742 & n46352 ) ;
  assign n46354 = ~n5021 & n27965 ;
  assign n46355 = n46354 ^ n20427 ^ n7901 ;
  assign n46356 = ( n7147 & n10430 ) | ( n7147 & ~n31746 ) | ( n10430 & ~n31746 ) ;
  assign n46357 = n634 & ~n9605 ;
  assign n46358 = ~n32971 & n46357 ;
  assign n46359 = n46358 ^ n29546 ^ n20463 ;
  assign n46360 = ( n3932 & ~n17040 ) | ( n3932 & n29760 ) | ( ~n17040 & n29760 ) ;
  assign n46361 = n32200 ^ n29506 ^ n15033 ;
  assign n46362 = n30285 ^ n24827 ^ 1'b0 ;
  assign n46363 = n1980 | n46362 ;
  assign n46364 = n16739 & ~n46363 ;
  assign n46365 = n34323 ^ n16437 ^ 1'b0 ;
  assign n46366 = n9471 | n46365 ;
  assign n46367 = n15425 | n46366 ;
  assign n46368 = ( ~n5340 & n17621 ) | ( ~n5340 & n46367 ) | ( n17621 & n46367 ) ;
  assign n46369 = n34127 ^ n10405 ^ n9712 ;
  assign n46370 = ( n379 & n4834 ) | ( n379 & n38617 ) | ( n4834 & n38617 ) ;
  assign n46371 = n29625 ^ n1956 ^ 1'b0 ;
  assign n46372 = n46370 | n46371 ;
  assign n46373 = n46372 ^ n39722 ^ n6951 ;
  assign n46374 = n21055 ^ n5632 ^ 1'b0 ;
  assign n46375 = ~n44110 & n46374 ;
  assign n46376 = n25410 & n41206 ;
  assign n46377 = ~n46375 & n46376 ;
  assign n46378 = n14490 & ~n40050 ;
  assign n46379 = n8780 & n46378 ;
  assign n46380 = n31514 ^ n2975 ^ 1'b0 ;
  assign n46381 = n14346 & n46380 ;
  assign n46382 = ~n46379 & n46381 ;
  assign n46383 = n46382 ^ n17664 ^ 1'b0 ;
  assign n46384 = ( ~n2705 & n12699 ) | ( ~n2705 & n14787 ) | ( n12699 & n14787 ) ;
  assign n46385 = n46384 ^ n22096 ^ n488 ;
  assign n46386 = n3792 & n24829 ;
  assign n46387 = n46385 & n46386 ;
  assign n46388 = n33638 ^ n6331 ^ n359 ;
  assign n46389 = n34620 ^ n12227 ^ n11892 ;
  assign n46390 = n46389 ^ n27106 ^ n8037 ;
  assign n46391 = n31881 ^ n22913 ^ n19261 ;
  assign n46396 = ( n4997 & n14929 ) | ( n4997 & n17027 ) | ( n14929 & n17027 ) ;
  assign n46397 = ( n869 & ~n40081 ) | ( n869 & n46396 ) | ( ~n40081 & n46396 ) ;
  assign n46392 = ( n9042 & n15172 ) | ( n9042 & n20392 ) | ( n15172 & n20392 ) ;
  assign n46393 = n46392 ^ n39605 ^ n35481 ;
  assign n46394 = n46393 ^ n26574 ^ n21320 ;
  assign n46395 = ( n17917 & n38662 ) | ( n17917 & n46394 ) | ( n38662 & n46394 ) ;
  assign n46398 = n46397 ^ n46395 ^ n21543 ;
  assign n46399 = n33633 & ~n45771 ;
  assign n46400 = n39350 ^ n5632 ^ 1'b0 ;
  assign n46401 = n26193 & ~n46400 ;
  assign n46402 = n46401 ^ n23465 ^ 1'b0 ;
  assign n46403 = ( n4934 & n11430 ) | ( n4934 & n46402 ) | ( n11430 & n46402 ) ;
  assign n46404 = n6739 & ~n25026 ;
  assign n46405 = n46404 ^ n22233 ^ 1'b0 ;
  assign n46406 = n46405 ^ n44632 ^ n11518 ;
  assign n46407 = ~n8618 & n44375 ;
  assign n46408 = ( n26778 & n28530 ) | ( n26778 & n34294 ) | ( n28530 & n34294 ) ;
  assign n46409 = ( n40741 & n46407 ) | ( n40741 & n46408 ) | ( n46407 & n46408 ) ;
  assign n46410 = n30416 ^ n6554 ^ 1'b0 ;
  assign n46411 = n46409 & n46410 ;
  assign n46412 = n7476 & ~n29193 ;
  assign n46413 = ~n969 & n46412 ;
  assign n46414 = ( ~n10835 & n26085 ) | ( ~n10835 & n33056 ) | ( n26085 & n33056 ) ;
  assign n46415 = n31561 ^ n28247 ^ n570 ;
  assign n46416 = ~n5718 & n46415 ;
  assign n46417 = ~n14568 & n46416 ;
  assign n46418 = ( ~n9793 & n25193 ) | ( ~n9793 & n46417 ) | ( n25193 & n46417 ) ;
  assign n46419 = n24813 ^ n7467 ^ n691 ;
  assign n46420 = n26216 ^ n6682 ^ 1'b0 ;
  assign n46421 = n4372 | n46420 ;
  assign n46422 = n46421 ^ n37644 ^ n7056 ;
  assign n46423 = n31603 ^ n14280 ^ n5849 ;
  assign n46424 = n46423 ^ n37641 ^ n3636 ;
  assign n46425 = ( ~n722 & n10217 ) | ( ~n722 & n46424 ) | ( n10217 & n46424 ) ;
  assign n46426 = n33557 ^ n10346 ^ 1'b0 ;
  assign n46427 = n34214 & n46426 ;
  assign n46428 = n13374 ^ n8892 ^ n2883 ;
  assign n46429 = n46428 ^ n16362 ^ n10318 ;
  assign n46430 = n9550 | n41012 ;
  assign n46431 = n46430 ^ n2053 ^ 1'b0 ;
  assign n46432 = ( n13558 & n32398 ) | ( n13558 & n46431 ) | ( n32398 & n46431 ) ;
  assign n46433 = n7706 & n20641 ;
  assign n46434 = n46433 ^ n40255 ^ n1254 ;
  assign n46435 = n664 | n2014 ;
  assign n46436 = n28984 & n38827 ;
  assign n46437 = n46436 ^ n17800 ^ n14159 ;
  assign n46438 = ( n7736 & ~n8634 ) | ( n7736 & n25809 ) | ( ~n8634 & n25809 ) ;
  assign n46439 = ( n11151 & n15045 ) | ( n11151 & n42138 ) | ( n15045 & n42138 ) ;
  assign n46440 = n37200 ^ n10753 ^ 1'b0 ;
  assign n46441 = ( n1560 & ~n46439 ) | ( n1560 & n46440 ) | ( ~n46439 & n46440 ) ;
  assign n46442 = ( ~n42241 & n46438 ) | ( ~n42241 & n46441 ) | ( n46438 & n46441 ) ;
  assign n46443 = n43074 ^ n42294 ^ n21461 ;
  assign n46444 = ( n1763 & ~n30997 ) | ( n1763 & n46443 ) | ( ~n30997 & n46443 ) ;
  assign n46445 = ~n1515 & n4489 ;
  assign n46446 = n46445 ^ n20291 ^ 1'b0 ;
  assign n46448 = n23865 ^ n19917 ^ n5554 ;
  assign n46447 = n8325 & n38596 ;
  assign n46449 = n46448 ^ n46447 ^ 1'b0 ;
  assign n46450 = n9838 & ~n35228 ;
  assign n46451 = ~n17469 & n46450 ;
  assign n46452 = n5684 & ~n12551 ;
  assign n46453 = n44223 ^ n10111 ^ n9170 ;
  assign n46454 = n36134 ^ n10133 ^ 1'b0 ;
  assign n46455 = ( n9109 & n46453 ) | ( n9109 & ~n46454 ) | ( n46453 & ~n46454 ) ;
  assign n46456 = n4551 ^ n758 ^ x50 ;
  assign n46457 = n46456 ^ n14095 ^ n7740 ;
  assign n46458 = n5162 & n8089 ;
  assign n46459 = ( n30274 & n46457 ) | ( n30274 & n46458 ) | ( n46457 & n46458 ) ;
  assign n46460 = ( ~n6887 & n8645 ) | ( ~n6887 & n17513 ) | ( n8645 & n17513 ) ;
  assign n46461 = n46460 ^ n3583 ^ n1702 ;
  assign n46462 = ( ~n1945 & n8104 ) | ( ~n1945 & n46461 ) | ( n8104 & n46461 ) ;
  assign n46463 = n40022 ^ n36296 ^ n17759 ;
  assign n46464 = n21119 & ~n25730 ;
  assign n46465 = n46464 ^ n22947 ^ n14599 ;
  assign n46466 = ~n3932 & n33384 ;
  assign n46467 = n46466 ^ n5475 ^ 1'b0 ;
  assign n46469 = n16091 ^ n15124 ^ n11072 ;
  assign n46468 = n24941 & ~n25127 ;
  assign n46470 = n46469 ^ n46468 ^ 1'b0 ;
  assign n46471 = ( n5802 & n7463 ) | ( n5802 & ~n39197 ) | ( n7463 & ~n39197 ) ;
  assign n46472 = n41935 ^ n7792 ^ 1'b0 ;
  assign n46473 = n46471 & n46472 ;
  assign n46474 = n10812 | n25055 ;
  assign n46475 = n46474 ^ n4192 ^ 1'b0 ;
  assign n46476 = ( n15669 & ~n16681 ) | ( n15669 & n46475 ) | ( ~n16681 & n46475 ) ;
  assign n46477 = ( n12163 & ~n14398 ) | ( n12163 & n14742 ) | ( ~n14398 & n14742 ) ;
  assign n46478 = n46477 ^ n14620 ^ n3284 ;
  assign n46479 = n46478 ^ n7513 ^ x192 ;
  assign n46480 = n6652 ^ n6068 ^ n5418 ;
  assign n46481 = n3045 & ~n46480 ;
  assign n46482 = n24521 & n46481 ;
  assign n46483 = n7911 ^ n5815 ^ n5394 ;
  assign n46484 = ( n36470 & n46482 ) | ( n36470 & ~n46483 ) | ( n46482 & ~n46483 ) ;
  assign n46485 = ( n2463 & n4746 ) | ( n2463 & n27551 ) | ( n4746 & n27551 ) ;
  assign n46486 = n10851 & ~n15553 ;
  assign n46487 = n2091 & n46486 ;
  assign n46488 = ( n12681 & ~n46485 ) | ( n12681 & n46487 ) | ( ~n46485 & n46487 ) ;
  assign n46490 = n24019 & ~n25610 ;
  assign n46491 = n46490 ^ n14285 ^ 1'b0 ;
  assign n46489 = ( n19131 & n19991 ) | ( n19131 & ~n28218 ) | ( n19991 & ~n28218 ) ;
  assign n46492 = n46491 ^ n46489 ^ n38294 ;
  assign n46493 = ( n2516 & n7981 ) | ( n2516 & ~n23455 ) | ( n7981 & ~n23455 ) ;
  assign n46494 = n15825 | n28594 ;
  assign n46495 = ( n23072 & n25892 ) | ( n23072 & ~n46494 ) | ( n25892 & ~n46494 ) ;
  assign n46496 = ~n24895 & n46495 ;
  assign n46497 = ( n6691 & n9239 ) | ( n6691 & n46496 ) | ( n9239 & n46496 ) ;
  assign n46498 = n20027 & n33438 ;
  assign n46499 = ~n37572 & n46498 ;
  assign n46500 = n28020 & ~n39258 ;
  assign n46501 = ~n21733 & n46500 ;
  assign n46502 = n14809 ^ n4897 ^ 1'b0 ;
  assign n46503 = n20290 | n40150 ;
  assign n46504 = n46503 ^ n30503 ^ 1'b0 ;
  assign n46505 = n29859 ^ n27950 ^ 1'b0 ;
  assign n46506 = n46505 ^ n28534 ^ n5320 ;
  assign n46507 = ( n18179 & n40555 ) | ( n18179 & n41947 ) | ( n40555 & n41947 ) ;
  assign n46508 = n23357 & n25575 ;
  assign n46509 = n46508 ^ n19076 ^ 1'b0 ;
  assign n46510 = ( ~n11447 & n32624 ) | ( ~n11447 & n46509 ) | ( n32624 & n46509 ) ;
  assign n46511 = ( n1990 & ~n6252 ) | ( n1990 & n9514 ) | ( ~n6252 & n9514 ) ;
  assign n46512 = n46511 ^ n45198 ^ n21997 ;
  assign n46513 = ( ~n8088 & n37480 ) | ( ~n8088 & n46512 ) | ( n37480 & n46512 ) ;
  assign n46514 = ( n659 & n5485 ) | ( n659 & n12260 ) | ( n5485 & n12260 ) ;
  assign n46515 = n15064 ^ n3250 ^ 1'b0 ;
  assign n46516 = n21572 | n46515 ;
  assign n46517 = ( n8122 & ~n32642 ) | ( n8122 & n41986 ) | ( ~n32642 & n41986 ) ;
  assign n46518 = ~n3231 & n46517 ;
  assign n46519 = n26870 & n46518 ;
  assign n46520 = n22140 ^ n1646 ^ 1'b0 ;
  assign n46521 = n22646 & ~n46520 ;
  assign n46522 = ~n14765 & n15815 ;
  assign n46523 = ~n22265 & n46522 ;
  assign n46524 = n46523 ^ n26665 ^ n13578 ;
  assign n46525 = ( n40435 & n46521 ) | ( n40435 & n46524 ) | ( n46521 & n46524 ) ;
  assign n46526 = n17589 & ~n46525 ;
  assign n46527 = n8979 & n46526 ;
  assign n46528 = n21119 ^ n12518 ^ 1'b0 ;
  assign n46529 = n38309 & ~n46528 ;
  assign n46530 = ~n21990 & n46529 ;
  assign n46531 = ( ~n14232 & n31593 ) | ( ~n14232 & n46530 ) | ( n31593 & n46530 ) ;
  assign n46532 = n46531 ^ n1028 ^ 1'b0 ;
  assign n46533 = n43213 ^ n21351 ^ n12946 ;
  assign n46534 = n4171 ^ n4150 ^ 1'b0 ;
  assign n46535 = n16697 & n46534 ;
  assign n46536 = n46535 ^ n26211 ^ 1'b0 ;
  assign n46537 = n46536 ^ n45980 ^ n45526 ;
  assign n46538 = n15352 ^ n15248 ^ n2367 ;
  assign n46539 = n46538 ^ n20103 ^ x14 ;
  assign n46540 = n42036 ^ n41304 ^ n24178 ;
  assign n46541 = n30848 ^ n30037 ^ 1'b0 ;
  assign n46542 = n34750 ^ n23471 ^ n14016 ;
  assign n46543 = n14342 & ~n46542 ;
  assign n46544 = n27179 & n46543 ;
  assign n46545 = n13962 ^ n8745 ^ 1'b0 ;
  assign n46546 = ~n10469 & n46545 ;
  assign n46547 = ~n16702 & n35599 ;
  assign n46548 = n46547 ^ n16744 ^ 1'b0 ;
  assign n46549 = n25739 ^ n25563 ^ n4732 ;
  assign n46550 = n46549 ^ n3793 ^ 1'b0 ;
  assign n46551 = n16951 & n46550 ;
  assign n46552 = n11507 & ~n25846 ;
  assign n46554 = ~n12479 & n29200 ;
  assign n46555 = n46554 ^ n14223 ^ 1'b0 ;
  assign n46553 = ( n5446 & n12863 ) | ( n5446 & n35969 ) | ( n12863 & n35969 ) ;
  assign n46556 = n46555 ^ n46553 ^ 1'b0 ;
  assign n46557 = n18631 | n39313 ;
  assign n46558 = n9621 ^ n9142 ^ 1'b0 ;
  assign n46559 = n16751 & n46558 ;
  assign n46560 = ( ~n610 & n22763 ) | ( ~n610 & n46559 ) | ( n22763 & n46559 ) ;
  assign n46561 = n35368 & n46560 ;
  assign n46562 = n45783 ^ n36045 ^ 1'b0 ;
  assign n46563 = ( n8804 & n13314 ) | ( n8804 & n14046 ) | ( n13314 & n14046 ) ;
  assign n46564 = n46563 ^ n31891 ^ n8308 ;
  assign n46565 = n46400 ^ n19819 ^ n16515 ;
  assign n46566 = ( n7890 & n21829 ) | ( n7890 & ~n46565 ) | ( n21829 & ~n46565 ) ;
  assign n46567 = ( ~n2097 & n20672 ) | ( ~n2097 & n46566 ) | ( n20672 & n46566 ) ;
  assign n46568 = n29206 & n31102 ;
  assign n46569 = ( n622 & ~n14060 ) | ( n622 & n43081 ) | ( ~n14060 & n43081 ) ;
  assign n46570 = n14568 & n21407 ;
  assign n46571 = ~n46569 & n46570 ;
  assign n46572 = ( n8674 & ~n15957 ) | ( n8674 & n17964 ) | ( ~n15957 & n17964 ) ;
  assign n46573 = n658 | n21219 ;
  assign n46574 = n29245 & ~n46573 ;
  assign n46575 = n46574 ^ n37124 ^ n32211 ;
  assign n46576 = ( n11611 & n11827 ) | ( n11611 & ~n12337 ) | ( n11827 & ~n12337 ) ;
  assign n46577 = n46576 ^ n1496 ^ 1'b0 ;
  assign n46578 = n46577 ^ n13069 ^ n7684 ;
  assign n46581 = n5626 & n7699 ;
  assign n46579 = n1996 | n9797 ;
  assign n46580 = n37148 & ~n46579 ;
  assign n46582 = n46581 ^ n46580 ^ n24020 ;
  assign n46583 = ~n21325 & n21754 ;
  assign n46584 = n31559 ^ n19283 ^ n5799 ;
  assign n46585 = n2397 & ~n46584 ;
  assign n46586 = n3374 & ~n4109 ;
  assign n46587 = n46586 ^ n5599 ^ 1'b0 ;
  assign n46588 = ( n16191 & n18072 ) | ( n16191 & n25340 ) | ( n18072 & n25340 ) ;
  assign n46589 = n2706 & n46588 ;
  assign n46590 = ( ~n1242 & n26902 ) | ( ~n1242 & n27598 ) | ( n26902 & n27598 ) ;
  assign n46592 = n31017 ^ n10700 ^ 1'b0 ;
  assign n46591 = ( n16578 & ~n30773 ) | ( n16578 & n33448 ) | ( ~n30773 & n33448 ) ;
  assign n46593 = n46592 ^ n46591 ^ n1155 ;
  assign n46594 = n46593 ^ n11649 ^ 1'b0 ;
  assign n46595 = n46590 & n46594 ;
  assign n46601 = ( n21274 & n30937 ) | ( n21274 & n36281 ) | ( n30937 & n36281 ) ;
  assign n46596 = ( n1805 & ~n17837 ) | ( n1805 & n18152 ) | ( ~n17837 & n18152 ) ;
  assign n46597 = n8932 & n19613 ;
  assign n46598 = n46597 ^ n7727 ^ 1'b0 ;
  assign n46599 = ( ~n9712 & n21248 ) | ( ~n9712 & n39935 ) | ( n21248 & n39935 ) ;
  assign n46600 = ( n46596 & n46598 ) | ( n46596 & n46599 ) | ( n46598 & n46599 ) ;
  assign n46602 = n46601 ^ n46600 ^ n28684 ;
  assign n46603 = n46602 ^ n44750 ^ n43980 ;
  assign n46604 = ( n5711 & n29253 ) | ( n5711 & ~n36030 ) | ( n29253 & ~n36030 ) ;
  assign n46605 = ( ~n18054 & n21061 ) | ( ~n18054 & n34634 ) | ( n21061 & n34634 ) ;
  assign n46606 = ~n45969 & n46605 ;
  assign n46607 = n15626 & ~n16094 ;
  assign n46608 = n46607 ^ n25398 ^ 1'b0 ;
  assign n46609 = n46608 ^ n21051 ^ n3411 ;
  assign n46610 = n19365 ^ n15510 ^ 1'b0 ;
  assign n46611 = n17029 ^ n12017 ^ n7086 ;
  assign n46612 = ( n42921 & n46415 ) | ( n42921 & n46611 ) | ( n46415 & n46611 ) ;
  assign n46613 = ~n8017 & n19299 ;
  assign n46614 = n42528 & n44979 ;
  assign n46615 = n46614 ^ n10082 ^ 1'b0 ;
  assign n46616 = ( n19136 & n22458 ) | ( n19136 & n25396 ) | ( n22458 & n25396 ) ;
  assign n46617 = n20469 & n25402 ;
  assign n46618 = ~n46616 & n46617 ;
  assign n46619 = n21546 ^ n16352 ^ 1'b0 ;
  assign n46620 = n8187 & ~n46619 ;
  assign n46621 = ( n30920 & ~n33260 ) | ( n30920 & n46620 ) | ( ~n33260 & n46620 ) ;
  assign n46622 = n3420 & ~n6394 ;
  assign n46623 = n1887 & n46622 ;
  assign n46624 = n46623 ^ n19946 ^ n10415 ;
  assign n46625 = n38037 ^ n26796 ^ n12910 ;
  assign n46626 = ( n2652 & ~n13508 ) | ( n2652 & n15930 ) | ( ~n13508 & n15930 ) ;
  assign n46627 = ( n10243 & n25486 ) | ( n10243 & ~n33938 ) | ( n25486 & ~n33938 ) ;
  assign n46628 = n29972 ^ x131 ^ 1'b0 ;
  assign n46629 = n9542 | n46628 ;
  assign n46630 = ~n8175 & n36156 ;
  assign n46631 = n46630 ^ n7599 ^ 1'b0 ;
  assign n46632 = n28678 & n46631 ;
  assign n46633 = n46632 ^ n44585 ^ 1'b0 ;
  assign n46634 = ( n2388 & n8510 ) | ( n2388 & ~n46633 ) | ( n8510 & ~n46633 ) ;
  assign n46635 = n16769 ^ n6431 ^ 1'b0 ;
  assign n46636 = n5484 & ~n46635 ;
  assign n46637 = n18693 ^ n1736 ^ 1'b0 ;
  assign n46638 = n12794 & n46637 ;
  assign n46639 = n26355 & n46638 ;
  assign n46642 = n35119 ^ n8168 ^ n1973 ;
  assign n46640 = ( n2190 & n22178 ) | ( n2190 & ~n39759 ) | ( n22178 & ~n39759 ) ;
  assign n46641 = n11485 | n46640 ;
  assign n46643 = n46642 ^ n46641 ^ 1'b0 ;
  assign n46644 = n2749 & ~n9370 ;
  assign n46645 = ~n1227 & n13838 ;
  assign n46646 = n3789 & n46645 ;
  assign n46647 = n15845 | n25483 ;
  assign n46648 = ~n16615 & n30554 ;
  assign n46649 = ~n25452 & n46648 ;
  assign n46650 = ( n46646 & n46647 ) | ( n46646 & ~n46649 ) | ( n46647 & ~n46649 ) ;
  assign n46651 = n40243 ^ n31567 ^ n9393 ;
  assign n46652 = ( n4921 & ~n31110 ) | ( n4921 & n45187 ) | ( ~n31110 & n45187 ) ;
  assign n46653 = ( n20849 & ~n25439 ) | ( n20849 & n31135 ) | ( ~n25439 & n31135 ) ;
  assign n46654 = n46653 ^ n21993 ^ 1'b0 ;
  assign n46655 = n30296 | n35180 ;
  assign n46656 = n46655 ^ n7222 ^ 1'b0 ;
  assign n46657 = ( ~n11060 & n35723 ) | ( ~n11060 & n46656 ) | ( n35723 & n46656 ) ;
  assign n46658 = n24595 ^ n17110 ^ n10587 ;
  assign n46659 = n46658 ^ n26659 ^ 1'b0 ;
  assign n46660 = n1867 & ~n46659 ;
  assign n46661 = n15341 | n26984 ;
  assign n46662 = n38317 | n46661 ;
  assign n46663 = n37103 ^ n34602 ^ n29842 ;
  assign n46664 = n44952 ^ n40119 ^ n38283 ;
  assign n46665 = n46664 ^ n43595 ^ n16985 ;
  assign n46666 = n33403 ^ n20921 ^ n12143 ;
  assign n46667 = ( ~n10238 & n11804 ) | ( ~n10238 & n25569 ) | ( n11804 & n25569 ) ;
  assign n46668 = ( n12810 & ~n19415 ) | ( n12810 & n46667 ) | ( ~n19415 & n46667 ) ;
  assign n46669 = n46668 ^ n20414 ^ n13693 ;
  assign n46670 = n29333 ^ n23961 ^ 1'b0 ;
  assign n46671 = n18808 & ~n44760 ;
  assign n46672 = n23440 ^ n18150 ^ 1'b0 ;
  assign n46673 = n46671 & n46672 ;
  assign n46674 = n12189 ^ n371 ^ 1'b0 ;
  assign n46675 = n1191 | n46674 ;
  assign n46676 = n46675 ^ n8688 ^ n7782 ;
  assign n46677 = ( n22832 & ~n22962 ) | ( n22832 & n46676 ) | ( ~n22962 & n46676 ) ;
  assign n46681 = n30051 ^ n13667 ^ n10699 ;
  assign n46678 = n16864 ^ n5659 ^ 1'b0 ;
  assign n46679 = n461 & ~n46678 ;
  assign n46680 = n12273 & n46679 ;
  assign n46682 = n46681 ^ n46680 ^ 1'b0 ;
  assign n46683 = n46677 & ~n46682 ;
  assign n46684 = n46683 ^ n21897 ^ 1'b0 ;
  assign n46685 = n39465 ^ n16117 ^ n14986 ;
  assign n46686 = n3549 | n37595 ;
  assign n46687 = n45224 ^ n11042 ^ 1'b0 ;
  assign n46688 = n24589 | n46687 ;
  assign n46689 = ( n3432 & ~n46686 ) | ( n3432 & n46688 ) | ( ~n46686 & n46688 ) ;
  assign n46690 = n6894 ^ n2948 ^ n2826 ;
  assign n46691 = ~n3550 & n46690 ;
  assign n46692 = n46691 ^ n26868 ^ n15335 ;
  assign n46693 = n46692 ^ n26816 ^ n3744 ;
  assign n46694 = n26074 | n46693 ;
  assign n46695 = n11878 & n44166 ;
  assign n46696 = ( n8113 & n33283 ) | ( n8113 & ~n46695 ) | ( n33283 & ~n46695 ) ;
  assign n46697 = n43464 ^ n1712 ^ x42 ;
  assign n46698 = n9337 & n16371 ;
  assign n46699 = n1832 & n46698 ;
  assign n46700 = n16828 ^ n13398 ^ 1'b0 ;
  assign n46701 = n28967 | n46700 ;
  assign n46702 = ( n12681 & n46699 ) | ( n12681 & ~n46701 ) | ( n46699 & ~n46701 ) ;
  assign n46703 = n33943 ^ n18521 ^ n4262 ;
  assign n46704 = n46703 ^ n45912 ^ 1'b0 ;
  assign n46705 = n7746 ^ n3859 ^ 1'b0 ;
  assign n46706 = n46704 & n46705 ;
  assign n46707 = n6846 & n29473 ;
  assign n46708 = n3493 ^ n1550 ^ 1'b0 ;
  assign n46709 = ( ~n9540 & n13367 ) | ( ~n9540 & n46708 ) | ( n13367 & n46708 ) ;
  assign n46710 = n46707 | n46709 ;
  assign n46711 = n14675 | n38595 ;
  assign n46713 = n11684 ^ n3933 ^ 1'b0 ;
  assign n46714 = n6964 | n46713 ;
  assign n46715 = ( ~n40972 & n41164 ) | ( ~n40972 & n46714 ) | ( n41164 & n46714 ) ;
  assign n46712 = n18284 ^ n10670 ^ n4475 ;
  assign n46716 = n46715 ^ n46712 ^ n19408 ;
  assign n46717 = ( n4694 & ~n8918 ) | ( n4694 & n9291 ) | ( ~n8918 & n9291 ) ;
  assign n46718 = n16225 & ~n46717 ;
  assign n46725 = n30852 ^ n24620 ^ 1'b0 ;
  assign n46726 = n21580 | n46725 ;
  assign n46719 = ( n2696 & n18077 ) | ( n2696 & n42438 ) | ( n18077 & n42438 ) ;
  assign n46720 = n6136 & ~n46719 ;
  assign n46721 = n30749 & n46720 ;
  assign n46722 = ~n4917 & n14544 ;
  assign n46723 = n46721 & n46722 ;
  assign n46724 = ( n13854 & n31247 ) | ( n13854 & ~n46723 ) | ( n31247 & ~n46723 ) ;
  assign n46727 = n46726 ^ n46724 ^ n32852 ;
  assign n46728 = n8388 & n13942 ;
  assign n46729 = n46728 ^ n40270 ^ 1'b0 ;
  assign n46730 = x208 & n20855 ;
  assign n46731 = n46730 ^ n27288 ^ 1'b0 ;
  assign n46732 = n33513 ^ n24476 ^ 1'b0 ;
  assign n46733 = n17673 | n22179 ;
  assign n46734 = n46732 | n46733 ;
  assign n46735 = x6 & n46649 ;
  assign n46736 = ( ~n2182 & n10433 ) | ( ~n2182 & n21248 ) | ( n10433 & n21248 ) ;
  assign n46737 = ( n21023 & n22358 ) | ( n21023 & ~n46736 ) | ( n22358 & ~n46736 ) ;
  assign n46738 = n36196 ^ n36087 ^ n30154 ;
  assign n46739 = n43398 ^ n42948 ^ n34869 ;
  assign n46740 = n46739 ^ n18064 ^ n702 ;
  assign n46741 = n30894 ^ n19104 ^ n8745 ;
  assign n46742 = n46741 ^ n22646 ^ n2294 ;
  assign n46743 = n39693 ^ n30503 ^ 1'b0 ;
  assign n46748 = n12956 ^ n10606 ^ 1'b0 ;
  assign n46749 = n11055 & n46748 ;
  assign n46744 = n4339 | n8526 ;
  assign n46745 = n46744 ^ n30805 ^ 1'b0 ;
  assign n46746 = n17589 ^ n7254 ^ 1'b0 ;
  assign n46747 = ( ~n9065 & n46745 ) | ( ~n9065 & n46746 ) | ( n46745 & n46746 ) ;
  assign n46750 = n46749 ^ n46747 ^ n3031 ;
  assign n46751 = n21642 ^ n14713 ^ 1'b0 ;
  assign n46752 = n25857 ^ n6465 ^ 1'b0 ;
  assign n46753 = n39184 ^ n18767 ^ n16774 ;
  assign n46754 = n15960 | n44369 ;
  assign n46755 = n46754 ^ n12264 ^ n10230 ;
  assign n46756 = n29113 ^ n25598 ^ 1'b0 ;
  assign n46757 = n17517 | n46756 ;
  assign n46758 = n12476 & ~n25701 ;
  assign n46759 = n46758 ^ n19050 ^ 1'b0 ;
  assign n46760 = n37681 & n46759 ;
  assign n46761 = n46760 ^ n36788 ^ n6878 ;
  assign n46762 = ( n7031 & ~n46757 ) | ( n7031 & n46761 ) | ( ~n46757 & n46761 ) ;
  assign n46763 = n38479 ^ n11218 ^ 1'b0 ;
  assign n46764 = n9408 | n46763 ;
  assign n46765 = n31236 | n46764 ;
  assign n46766 = n3813 & ~n46765 ;
  assign n46767 = ( n8742 & ~n24204 ) | ( n8742 & n46766 ) | ( ~n24204 & n46766 ) ;
  assign n46772 = ~n11194 & n19943 ;
  assign n46768 = n16752 ^ n643 ^ 1'b0 ;
  assign n46769 = n414 | n46768 ;
  assign n46770 = n6386 & ~n46769 ;
  assign n46771 = n46770 ^ n36440 ^ 1'b0 ;
  assign n46773 = n46772 ^ n46771 ^ n33499 ;
  assign n46774 = ( n3048 & ~n20693 ) | ( n3048 & n28501 ) | ( ~n20693 & n28501 ) ;
  assign n46775 = ( ~n2742 & n8620 ) | ( ~n2742 & n33230 ) | ( n8620 & n33230 ) ;
  assign n46776 = ( n30033 & n46774 ) | ( n30033 & ~n46775 ) | ( n46774 & ~n46775 ) ;
  assign n46777 = n30919 ^ n15930 ^ 1'b0 ;
  assign n46778 = n46777 ^ n6365 ^ n3594 ;
  assign n46779 = ( n23090 & ~n46389 ) | ( n23090 & n46778 ) | ( ~n46389 & n46778 ) ;
  assign n46781 = ( ~n13325 & n14579 ) | ( ~n13325 & n19546 ) | ( n14579 & n19546 ) ;
  assign n46780 = ( n5324 & ~n13786 ) | ( n5324 & n21294 ) | ( ~n13786 & n21294 ) ;
  assign n46782 = n46781 ^ n46780 ^ 1'b0 ;
  assign n46785 = ( n10940 & ~n39648 ) | ( n10940 & n43302 ) | ( ~n39648 & n43302 ) ;
  assign n46783 = n1323 & ~n1956 ;
  assign n46784 = ~n17557 & n46783 ;
  assign n46786 = n46785 ^ n46784 ^ n7741 ;
  assign n46787 = ~n3898 & n37273 ;
  assign n46788 = n45577 & n46787 ;
  assign n46789 = n46788 ^ n41118 ^ n4438 ;
  assign n46790 = n5110 & n46789 ;
  assign n46791 = n46790 ^ n44669 ^ 1'b0 ;
  assign n46793 = n42837 ^ n29382 ^ 1'b0 ;
  assign n46794 = n31053 | n46793 ;
  assign n46792 = n12695 & n20049 ;
  assign n46795 = n46794 ^ n46792 ^ 1'b0 ;
  assign n46796 = ~n13017 & n34460 ;
  assign n46797 = n31137 ^ n25518 ^ n13473 ;
  assign n46798 = ~n8519 & n31283 ;
  assign n46799 = n46798 ^ n6498 ^ 1'b0 ;
  assign n46800 = n1122 | n5098 ;
  assign n46801 = n8484 & ~n46800 ;
  assign n46802 = n46801 ^ n36956 ^ n35840 ;
  assign n46803 = ( ~n20458 & n46799 ) | ( ~n20458 & n46802 ) | ( n46799 & n46802 ) ;
  assign n46804 = n43335 ^ n17084 ^ n9783 ;
  assign n46806 = n13794 ^ n13543 ^ 1'b0 ;
  assign n46805 = n40595 ^ n18732 ^ n16122 ;
  assign n46807 = n46806 ^ n46805 ^ 1'b0 ;
  assign n46811 = n6209 ^ x71 ^ 1'b0 ;
  assign n46809 = n17513 ^ n10358 ^ n3351 ;
  assign n46808 = n32208 ^ n19205 ^ n566 ;
  assign n46810 = n46809 ^ n46808 ^ n931 ;
  assign n46812 = n46811 ^ n46810 ^ n24811 ;
  assign n46813 = n23061 ^ n11668 ^ 1'b0 ;
  assign n46814 = n26231 | n46813 ;
  assign n46815 = ( ~n13776 & n24518 ) | ( ~n13776 & n46814 ) | ( n24518 & n46814 ) ;
  assign n46816 = ( n14684 & ~n15333 ) | ( n14684 & n27913 ) | ( ~n15333 & n27913 ) ;
  assign n46817 = n2742 & n46816 ;
  assign n46818 = n29919 ^ n496 ^ 1'b0 ;
  assign n46819 = n46818 ^ n13143 ^ n3502 ;
  assign n46820 = ( n10059 & n33495 ) | ( n10059 & ~n45995 ) | ( n33495 & ~n45995 ) ;
  assign n46821 = n5899 & n46820 ;
  assign n46822 = n46821 ^ n32880 ^ 1'b0 ;
  assign n46823 = n32252 ^ n4243 ^ 1'b0 ;
  assign n46824 = n36027 ^ n2548 ^ 1'b0 ;
  assign n46825 = n12237 & n46824 ;
  assign n46826 = ( ~n5641 & n45863 ) | ( ~n5641 & n46825 ) | ( n45863 & n46825 ) ;
  assign n46827 = n41979 ^ n21603 ^ 1'b0 ;
  assign n46828 = n46827 ^ n23810 ^ n8828 ;
  assign n46829 = n21943 ^ n3342 ^ x193 ;
  assign n46830 = n8525 & n46829 ;
  assign n46831 = n46421 ^ n40352 ^ n25359 ;
  assign n46832 = n28573 ^ n27104 ^ n11756 ;
  assign n46833 = ( n12812 & n22999 ) | ( n12812 & ~n33563 ) | ( n22999 & ~n33563 ) ;
  assign n46834 = ( n14552 & ~n19576 ) | ( n14552 & n46833 ) | ( ~n19576 & n46833 ) ;
  assign n46835 = n15335 & ~n46834 ;
  assign n46836 = n17450 ^ n13403 ^ n4130 ;
  assign n46837 = n7137 & n19746 ;
  assign n46838 = ~n40521 & n46837 ;
  assign n46839 = n46838 ^ n15365 ^ 1'b0 ;
  assign n46840 = n46836 & ~n46839 ;
  assign n46841 = ( n26000 & n29431 ) | ( n26000 & ~n38652 ) | ( n29431 & ~n38652 ) ;
  assign n46842 = ( n21664 & ~n41652 ) | ( n21664 & n46094 ) | ( ~n41652 & n46094 ) ;
  assign n46843 = n15309 ^ n7601 ^ 1'b0 ;
  assign n46844 = n7856 & ~n46843 ;
  assign n46845 = n46844 ^ n9870 ^ n713 ;
  assign n46846 = ( n1309 & ~n27909 ) | ( n1309 & n31139 ) | ( ~n27909 & n31139 ) ;
  assign n46847 = ( ~n20656 & n32865 ) | ( ~n20656 & n46846 ) | ( n32865 & n46846 ) ;
  assign n46848 = n46847 ^ n27550 ^ n5484 ;
  assign n46849 = n31120 ^ n4363 ^ 1'b0 ;
  assign n46850 = ~n1417 & n17398 ;
  assign n46851 = n46850 ^ n21325 ^ 1'b0 ;
  assign n46852 = n21147 | n29792 ;
  assign n46853 = n20030 | n46852 ;
  assign n46854 = n10740 | n12115 ;
  assign n46855 = n46854 ^ n35891 ^ 1'b0 ;
  assign n46856 = n34666 ^ n4319 ^ 1'b0 ;
  assign n46857 = n8939 | n46856 ;
  assign n46858 = n30297 ^ n24995 ^ n24985 ;
  assign n46859 = n17615 ^ n16621 ^ n6567 ;
  assign n46860 = n46859 ^ n13066 ^ n473 ;
  assign n46861 = ~n46858 & n46860 ;
  assign n46862 = ( n6281 & ~n6477 ) | ( n6281 & n13412 ) | ( ~n6477 & n13412 ) ;
  assign n46863 = n46862 ^ n38353 ^ n14257 ;
  assign n46864 = ~n8171 & n23168 ;
  assign n46865 = n42343 ^ n4904 ^ n2254 ;
  assign n46866 = ( n15968 & n46864 ) | ( n15968 & ~n46865 ) | ( n46864 & ~n46865 ) ;
  assign n46867 = n36528 ^ n14252 ^ n9314 ;
  assign n46868 = ( ~n16880 & n39353 ) | ( ~n16880 & n46867 ) | ( n39353 & n46867 ) ;
  assign n46869 = n46868 ^ n37760 ^ n35665 ;
  assign n46872 = ~n299 & n9486 ;
  assign n46873 = n11392 & n46872 ;
  assign n46874 = n10403 & ~n46873 ;
  assign n46870 = n332 & n15170 ;
  assign n46871 = ~n5364 & n46870 ;
  assign n46875 = n46874 ^ n46871 ^ n8726 ;
  assign n46876 = n23229 ^ n22523 ^ n3638 ;
  assign n46877 = n7207 ^ n6915 ^ 1'b0 ;
  assign n46878 = n19262 ^ n13119 ^ n7290 ;
  assign n46879 = n27950 ^ n5488 ^ 1'b0 ;
  assign n46880 = ( ~n46877 & n46878 ) | ( ~n46877 & n46879 ) | ( n46878 & n46879 ) ;
  assign n46881 = ( n28652 & n30002 ) | ( n28652 & ~n46880 ) | ( n30002 & ~n46880 ) ;
  assign n46882 = ( n770 & n13986 ) | ( n770 & ~n32927 ) | ( n13986 & ~n32927 ) ;
  assign n46883 = n46882 ^ n5861 ^ 1'b0 ;
  assign n46884 = n20396 | n46883 ;
  assign n46885 = n3476 ^ n478 ^ 1'b0 ;
  assign n46886 = n46885 ^ n31510 ^ 1'b0 ;
  assign n46887 = n38849 ^ n35700 ^ n12781 ;
  assign n46888 = ( ~n845 & n16559 ) | ( ~n845 & n46887 ) | ( n16559 & n46887 ) ;
  assign n46889 = n46886 & n46888 ;
  assign n46890 = n22211 ^ n16033 ^ n14849 ;
  assign n46891 = n46890 ^ n24521 ^ n1473 ;
  assign n46892 = n11061 ^ n6494 ^ 1'b0 ;
  assign n46893 = n5951 & ~n28157 ;
  assign n46895 = ( n12610 & ~n32642 ) | ( n12610 & n45017 ) | ( ~n32642 & n45017 ) ;
  assign n46894 = n14395 ^ n7224 ^ n2685 ;
  assign n46896 = n46895 ^ n46894 ^ n8097 ;
  assign n46897 = ( n27036 & ~n38844 ) | ( n27036 & n41977 ) | ( ~n38844 & n41977 ) ;
  assign n46898 = n6188 | n11471 ;
  assign n46899 = n24192 & ~n46898 ;
  assign n46900 = n46899 ^ n46882 ^ 1'b0 ;
  assign n46902 = ( n3548 & ~n9047 ) | ( n3548 & n14211 ) | ( ~n9047 & n14211 ) ;
  assign n46903 = n46902 ^ n12059 ^ 1'b0 ;
  assign n46904 = ( n3151 & ~n7950 ) | ( n3151 & n46903 ) | ( ~n7950 & n46903 ) ;
  assign n46901 = n4997 | n12202 ;
  assign n46905 = n46904 ^ n46901 ^ 1'b0 ;
  assign n46906 = ( n2134 & n8390 ) | ( n2134 & ~n9808 ) | ( n8390 & ~n9808 ) ;
  assign n46907 = n44465 ^ n39468 ^ 1'b0 ;
  assign n46908 = n46906 | n46907 ;
  assign n46909 = n26155 ^ n24275 ^ n12796 ;
  assign n46910 = n14438 ^ n11529 ^ n5484 ;
  assign n46911 = n46910 ^ n14772 ^ 1'b0 ;
  assign n46912 = n46909 | n46911 ;
  assign n46913 = n46912 ^ n22337 ^ n17470 ;
  assign n46914 = ( n9727 & n25548 ) | ( n9727 & n40981 ) | ( n25548 & n40981 ) ;
  assign n46915 = ( n12121 & n23498 ) | ( n12121 & ~n43375 ) | ( n23498 & ~n43375 ) ;
  assign n46917 = n5113 & ~n30670 ;
  assign n46916 = n21936 ^ n1202 ^ n966 ;
  assign n46918 = n46917 ^ n46916 ^ n21506 ;
  assign n46919 = n21162 ^ n13207 ^ n6509 ;
  assign n46920 = n23001 | n46919 ;
  assign n46921 = ( ~n14455 & n18773 ) | ( ~n14455 & n46920 ) | ( n18773 & n46920 ) ;
  assign n46922 = n33388 ^ n22240 ^ n14563 ;
  assign n46923 = n5662 & ~n13729 ;
  assign n46924 = n38077 ^ n15640 ^ 1'b0 ;
  assign n46925 = n3522 & ~n22113 ;
  assign n46926 = n46925 ^ n23715 ^ 1'b0 ;
  assign n46927 = ( n16200 & ~n24586 ) | ( n16200 & n29573 ) | ( ~n24586 & n29573 ) ;
  assign n46928 = ( ~n8570 & n25527 ) | ( ~n8570 & n28973 ) | ( n25527 & n28973 ) ;
  assign n46929 = ( n5754 & n12190 ) | ( n5754 & n19588 ) | ( n12190 & n19588 ) ;
  assign n46930 = ( ~n3751 & n5827 ) | ( ~n3751 & n25118 ) | ( n5827 & n25118 ) ;
  assign n46931 = ( n6554 & n19893 ) | ( n6554 & ~n46930 ) | ( n19893 & ~n46930 ) ;
  assign n46932 = n8383 & ~n39384 ;
  assign n46933 = n12035 & n46932 ;
  assign n46936 = ( n6695 & n19983 ) | ( n6695 & n20488 ) | ( n19983 & n20488 ) ;
  assign n46934 = n30326 ^ n7151 ^ 1'b0 ;
  assign n46935 = n22878 & ~n46934 ;
  assign n46937 = n46936 ^ n46935 ^ n21580 ;
  assign n46938 = n4463 | n15093 ;
  assign n46939 = n45083 ^ n25191 ^ 1'b0 ;
  assign n46940 = n17516 & ~n46939 ;
  assign n46941 = n34976 ^ n12376 ^ n4250 ;
  assign n46942 = ( ~n24080 & n46940 ) | ( ~n24080 & n46941 ) | ( n46940 & n46941 ) ;
  assign n46943 = ~n36557 & n41633 ;
  assign n46944 = n44881 ^ n13307 ^ 1'b0 ;
  assign n46945 = ( n7153 & n42861 ) | ( n7153 & ~n46944 ) | ( n42861 & ~n46944 ) ;
  assign n46948 = n2994 & ~n7662 ;
  assign n46949 = ( ~n3697 & n44006 ) | ( ~n3697 & n46948 ) | ( n44006 & n46948 ) ;
  assign n46946 = n9105 & n12260 ;
  assign n46947 = n46946 ^ n10734 ^ n5578 ;
  assign n46950 = n46949 ^ n46947 ^ n27746 ;
  assign n46951 = n10545 & n25130 ;
  assign n46952 = n46951 ^ n20493 ^ n1620 ;
  assign n46953 = ( n6985 & n20013 ) | ( n6985 & n46952 ) | ( n20013 & n46952 ) ;
  assign n46954 = ~n13199 & n46953 ;
  assign n46955 = n46954 ^ n34383 ^ 1'b0 ;
  assign n46956 = n5825 & n41583 ;
  assign n46957 = n46956 ^ n25053 ^ 1'b0 ;
  assign n46958 = ~n17676 & n46957 ;
  assign n46959 = n23532 & n46958 ;
  assign n46960 = n46959 ^ n2185 ^ 1'b0 ;
  assign n46961 = n36754 ^ n14208 ^ 1'b0 ;
  assign n46962 = n44533 ^ n35205 ^ n17951 ;
  assign n46963 = ( n31504 & ~n35184 ) | ( n31504 & n41846 ) | ( ~n35184 & n41846 ) ;
  assign n46964 = ( n8846 & ~n13135 ) | ( n8846 & n46963 ) | ( ~n13135 & n46963 ) ;
  assign n46965 = n39162 ^ n30017 ^ n18386 ;
  assign n46966 = ( ~n2078 & n5937 ) | ( ~n2078 & n12092 ) | ( n5937 & n12092 ) ;
  assign n46967 = n18935 ^ n9951 ^ n2394 ;
  assign n46968 = ( ~n14958 & n46966 ) | ( ~n14958 & n46967 ) | ( n46966 & n46967 ) ;
  assign n46969 = ( ~n34988 & n44206 ) | ( ~n34988 & n46968 ) | ( n44206 & n46968 ) ;
  assign n46970 = ( n1921 & ~n7692 ) | ( n1921 & n9746 ) | ( ~n7692 & n9746 ) ;
  assign n46971 = ( n27812 & n36540 ) | ( n27812 & ~n46970 ) | ( n36540 & ~n46970 ) ;
  assign n46972 = n1873 ^ n1503 ^ 1'b0 ;
  assign n46973 = n4684 & ~n46972 ;
  assign n46974 = n46973 ^ n31218 ^ n27979 ;
  assign n46975 = n46974 ^ n39600 ^ n5255 ;
  assign n46976 = ( n7770 & n46971 ) | ( n7770 & n46975 ) | ( n46971 & n46975 ) ;
  assign n46977 = ( n22314 & n41286 ) | ( n22314 & n41873 ) | ( n41286 & n41873 ) ;
  assign n46978 = n38925 ^ n38130 ^ 1'b0 ;
  assign n46979 = n23500 ^ n23209 ^ n12436 ;
  assign n46980 = n42380 ^ n29945 ^ 1'b0 ;
  assign n46981 = ~n46979 & n46980 ;
  assign n46982 = ~n19849 & n35539 ;
  assign n46983 = n46982 ^ n23276 ^ 1'b0 ;
  assign n46984 = n11792 & n15851 ;
  assign n46985 = n27251 | n33108 ;
  assign n46986 = n41243 | n46985 ;
  assign n46987 = ( n23089 & ~n35458 ) | ( n23089 & n46986 ) | ( ~n35458 & n46986 ) ;
  assign n46988 = n484 | n28263 ;
  assign n46989 = n26293 ^ n24214 ^ n21050 ;
  assign n46990 = ( n23030 & n34583 ) | ( n23030 & ~n46989 ) | ( n34583 & ~n46989 ) ;
  assign n46993 = n5736 & ~n46646 ;
  assign n46994 = n28193 & n46993 ;
  assign n46995 = n46994 ^ n27167 ^ 1'b0 ;
  assign n46991 = n36299 & n37248 ;
  assign n46992 = n46991 ^ n4174 ^ 1'b0 ;
  assign n46996 = n46995 ^ n46992 ^ n32612 ;
  assign n46997 = ( ~n4288 & n5262 ) | ( ~n4288 & n11824 ) | ( n5262 & n11824 ) ;
  assign n46998 = ~n40796 & n46997 ;
  assign n46999 = n6015 & n17265 ;
  assign n47000 = n46999 ^ n10300 ^ 1'b0 ;
  assign n47001 = ( ~n16258 & n21537 ) | ( ~n16258 & n47000 ) | ( n21537 & n47000 ) ;
  assign n47003 = ( ~n18687 & n20420 ) | ( ~n18687 & n23506 ) | ( n20420 & n23506 ) ;
  assign n47002 = n1422 & n19003 ;
  assign n47004 = n47003 ^ n47002 ^ 1'b0 ;
  assign n47005 = n24116 ^ n11924 ^ n10735 ;
  assign n47006 = ( n10254 & n40374 ) | ( n10254 & ~n40656 ) | ( n40374 & ~n40656 ) ;
  assign n47007 = n1951 | n18618 ;
  assign n47008 = n47007 ^ n5938 ^ 1'b0 ;
  assign n47009 = n5478 & ~n47008 ;
  assign n47010 = n47009 ^ n7456 ^ n563 ;
  assign n47011 = n46252 ^ n24898 ^ 1'b0 ;
  assign n47012 = n9596 & ~n47011 ;
  assign n47013 = ( n13832 & n17502 ) | ( n13832 & n47012 ) | ( n17502 & n47012 ) ;
  assign n47014 = ( n8659 & n12069 ) | ( n8659 & n16623 ) | ( n12069 & n16623 ) ;
  assign n47015 = ( n13864 & n22513 ) | ( n13864 & ~n47014 ) | ( n22513 & ~n47014 ) ;
  assign n47016 = ~n740 & n12058 ;
  assign n47017 = ~n34146 & n47016 ;
  assign n47018 = ( n1979 & ~n47015 ) | ( n1979 & n47017 ) | ( ~n47015 & n47017 ) ;
  assign n47019 = n47018 ^ n14633 ^ 1'b0 ;
  assign n47020 = n47019 ^ n6102 ^ n1131 ;
  assign n47021 = ( n956 & ~n6481 ) | ( n956 & n23170 ) | ( ~n6481 & n23170 ) ;
  assign n47022 = n47021 ^ n26130 ^ n13681 ;
  assign n47023 = n18402 & ~n40313 ;
  assign n47024 = n45604 & n47023 ;
  assign n47025 = n7637 & n36789 ;
  assign n47026 = n42122 & n47025 ;
  assign n47027 = n44189 ^ n27829 ^ 1'b0 ;
  assign n47028 = n24809 | n47027 ;
  assign n47030 = ~n16019 & n34411 ;
  assign n47029 = ( n6005 & ~n15051 ) | ( n6005 & n15995 ) | ( ~n15051 & n15995 ) ;
  assign n47031 = n47030 ^ n47029 ^ n2725 ;
  assign n47032 = ( n10612 & ~n15498 ) | ( n10612 & n19143 ) | ( ~n15498 & n19143 ) ;
  assign n47036 = ( ~n13134 & n20102 ) | ( ~n13134 & n40696 ) | ( n20102 & n40696 ) ;
  assign n47033 = n23926 ^ n16455 ^ n10712 ;
  assign n47034 = ( ~x193 & n8357 ) | ( ~x193 & n15576 ) | ( n8357 & n15576 ) ;
  assign n47035 = ( n35153 & ~n47033 ) | ( n35153 & n47034 ) | ( ~n47033 & n47034 ) ;
  assign n47037 = n47036 ^ n47035 ^ x245 ;
  assign n47040 = n29536 ^ n10741 ^ n5418 ;
  assign n47038 = n28356 ^ n6436 ^ n3620 ;
  assign n47039 = n47038 ^ n22012 ^ n8884 ;
  assign n47041 = n47040 ^ n47039 ^ n23129 ;
  assign n47042 = ( n6376 & ~n10805 ) | ( n6376 & n11737 ) | ( ~n10805 & n11737 ) ;
  assign n47043 = ~n15603 & n47042 ;
  assign n47044 = n21238 & n47043 ;
  assign n47045 = ( n3441 & n28341 ) | ( n3441 & n34091 ) | ( n28341 & n34091 ) ;
  assign n47046 = n47045 ^ n21104 ^ 1'b0 ;
  assign n47047 = ~n16275 & n47046 ;
  assign n47048 = n13193 & ~n22202 ;
  assign n47049 = ( n27355 & ~n44120 ) | ( n27355 & n47048 ) | ( ~n44120 & n47048 ) ;
  assign n47050 = n47049 ^ n31306 ^ 1'b0 ;
  assign n47051 = n950 & ~n47050 ;
  assign n47052 = ~n3116 & n19904 ;
  assign n47053 = n47052 ^ n28281 ^ n15959 ;
  assign n47054 = ( ~n6867 & n10583 ) | ( ~n6867 & n20097 ) | ( n10583 & n20097 ) ;
  assign n47055 = n47054 ^ n33475 ^ n2379 ;
  assign n47056 = ( n9198 & ~n30827 ) | ( n9198 & n33924 ) | ( ~n30827 & n33924 ) ;
  assign n47057 = ~n2579 & n15754 ;
  assign n47058 = n5619 & n47057 ;
  assign n47059 = n47058 ^ n1774 ^ 1'b0 ;
  assign n47060 = n43272 ^ n32532 ^ n8495 ;
  assign n47061 = n37379 ^ n36939 ^ 1'b0 ;
  assign n47062 = ( ~n7304 & n7729 ) | ( ~n7304 & n10952 ) | ( n7729 & n10952 ) ;
  assign n47063 = n5593 & n20576 ;
  assign n47064 = n47063 ^ n34220 ^ 1'b0 ;
  assign n47065 = n44366 | n47064 ;
  assign n47066 = n47062 & ~n47065 ;
  assign n47067 = n47066 ^ n17846 ^ 1'b0 ;
  assign n47068 = ~n26779 & n47067 ;
  assign n47069 = n5312 & ~n12126 ;
  assign n47070 = n8834 & ~n30855 ;
  assign n47071 = n47070 ^ n22992 ^ 1'b0 ;
  assign n47072 = n18752 ^ n8982 ^ n1466 ;
  assign n47073 = n46018 | n47072 ;
  assign n47074 = n19175 & n47073 ;
  assign n47075 = n7425 & ~n47074 ;
  assign n47076 = ( ~n1246 & n15471 ) | ( ~n1246 & n31979 ) | ( n15471 & n31979 ) ;
  assign n47077 = n6583 & ~n30171 ;
  assign n47078 = n14209 ^ n4014 ^ x210 ;
  assign n47079 = n16965 | n47078 ;
  assign n47080 = n47079 ^ n21191 ^ n19190 ;
  assign n47085 = n38077 ^ n12087 ^ 1'b0 ;
  assign n47086 = ~n13225 & n47085 ;
  assign n47081 = n20584 ^ n12849 ^ n3137 ;
  assign n47082 = ( ~n15322 & n16707 ) | ( ~n15322 & n34171 ) | ( n16707 & n34171 ) ;
  assign n47083 = n9211 & n47082 ;
  assign n47084 = n47081 & ~n47083 ;
  assign n47087 = n47086 ^ n47084 ^ 1'b0 ;
  assign n47088 = ( n6041 & n14014 ) | ( n6041 & n25396 ) | ( n14014 & n25396 ) ;
  assign n47089 = n32175 ^ n19554 ^ n8222 ;
  assign n47090 = n21955 | n47089 ;
  assign n47091 = ~n47088 & n47090 ;
  assign n47092 = ( n5733 & n6229 ) | ( n5733 & ~n47091 ) | ( n6229 & ~n47091 ) ;
  assign n47093 = ( ~n8335 & n16385 ) | ( ~n8335 & n45808 ) | ( n16385 & n45808 ) ;
  assign n47094 = ~n2341 & n47093 ;
  assign n47095 = n47094 ^ n5234 ^ 1'b0 ;
  assign n47096 = ( ~n10259 & n25957 ) | ( ~n10259 & n47095 ) | ( n25957 & n47095 ) ;
  assign n47097 = n3826 | n13135 ;
  assign n47098 = n8638 | n47097 ;
  assign n47099 = n47098 ^ n13522 ^ 1'b0 ;
  assign n47100 = n42251 ^ n17960 ^ n2557 ;
  assign n47101 = n47100 ^ n42756 ^ n11686 ;
  assign n47102 = n32045 ^ n27873 ^ n22585 ;
  assign n47103 = ( n18528 & ~n19608 ) | ( n18528 & n47102 ) | ( ~n19608 & n47102 ) ;
  assign n47104 = ( n27985 & ~n28331 ) | ( n27985 & n42328 ) | ( ~n28331 & n42328 ) ;
  assign n47105 = n31170 ^ n29155 ^ n22429 ;
  assign n47106 = n47105 ^ n36176 ^ n13130 ;
  assign n47107 = n20801 & ~n45253 ;
  assign n47108 = n15805 ^ n6159 ^ 1'b0 ;
  assign n47109 = n47108 ^ n25167 ^ n10162 ;
  assign n47110 = n24650 & ~n47109 ;
  assign n47111 = n40731 ^ n24560 ^ n624 ;
  assign n47115 = n27918 ^ n23360 ^ 1'b0 ;
  assign n47112 = n20407 ^ n5789 ^ n5122 ;
  assign n47113 = ( n1476 & n45444 ) | ( n1476 & n47112 ) | ( n45444 & n47112 ) ;
  assign n47114 = ~n18947 & n47113 ;
  assign n47116 = n47115 ^ n47114 ^ 1'b0 ;
  assign n47117 = n3819 & ~n14911 ;
  assign n47118 = n47117 ^ n10807 ^ 1'b0 ;
  assign n47119 = ( n5078 & n40521 ) | ( n5078 & n47118 ) | ( n40521 & n47118 ) ;
  assign n47120 = n47119 ^ n28140 ^ n6126 ;
  assign n47121 = n20148 & ~n41775 ;
  assign n47122 = n47121 ^ n12314 ^ 1'b0 ;
  assign n47123 = n20123 & n22259 ;
  assign n47124 = ~n19126 & n35350 ;
  assign n47125 = ( n13042 & n32698 ) | ( n13042 & n35192 ) | ( n32698 & n35192 ) ;
  assign n47126 = n1928 & ~n14413 ;
  assign n47127 = n10338 ^ n1223 ^ 1'b0 ;
  assign n47128 = ( ~n1028 & n4619 ) | ( ~n1028 & n27526 ) | ( n4619 & n27526 ) ;
  assign n47129 = n20341 ^ n5921 ^ n1409 ;
  assign n47130 = n23950 & n47129 ;
  assign n47131 = ( x84 & x163 ) | ( x84 & ~n32420 ) | ( x163 & ~n32420 ) ;
  assign n47132 = ( n34411 & n47130 ) | ( n34411 & n47131 ) | ( n47130 & n47131 ) ;
  assign n47133 = n19749 | n25787 ;
  assign n47134 = n47132 & ~n47133 ;
  assign n47135 = n45406 ^ n26139 ^ n17354 ;
  assign n47136 = ~n7907 & n21776 ;
  assign n47137 = n45793 ^ n44480 ^ n25986 ;
  assign n47138 = n40555 ^ n19227 ^ n9494 ;
  assign n47139 = n42211 & ~n47138 ;
  assign n47140 = ( n5216 & ~n10163 ) | ( n5216 & n19019 ) | ( ~n10163 & n19019 ) ;
  assign n47141 = n3736 ^ n1520 ^ n444 ;
  assign n47142 = n47141 ^ n1060 ^ n442 ;
  assign n47143 = n40175 ^ n36542 ^ n25861 ;
  assign n47144 = ( ~n9728 & n34918 ) | ( ~n9728 & n47143 ) | ( n34918 & n47143 ) ;
  assign n47145 = n21579 & ~n47144 ;
  assign n47146 = n331 & n47145 ;
  assign n47147 = n47142 & ~n47146 ;
  assign n47148 = n22175 & n47147 ;
  assign n47149 = n19480 ^ n7706 ^ 1'b0 ;
  assign n47150 = n15140 & n47149 ;
  assign n47151 = ( n23072 & ~n45145 ) | ( n23072 & n47150 ) | ( ~n45145 & n47150 ) ;
  assign n47152 = n47151 ^ n27084 ^ n12302 ;
  assign n47153 = n1054 & ~n47152 ;
  assign n47154 = n41218 ^ n19848 ^ 1'b0 ;
  assign n47155 = n23922 | n47154 ;
  assign n47156 = n26639 ^ n13672 ^ n10728 ;
  assign n47157 = n47156 ^ n39001 ^ 1'b0 ;
  assign n47158 = n19349 & n47157 ;
  assign n47159 = ( ~n26111 & n38699 ) | ( ~n26111 & n45966 ) | ( n38699 & n45966 ) ;
  assign n47160 = ( n2473 & ~n5953 ) | ( n2473 & n22219 ) | ( ~n5953 & n22219 ) ;
  assign n47161 = ( ~n12105 & n12304 ) | ( ~n12105 & n47160 ) | ( n12304 & n47160 ) ;
  assign n47162 = ( n34218 & ~n41576 ) | ( n34218 & n47161 ) | ( ~n41576 & n47161 ) ;
  assign n47163 = ( ~n8754 & n13131 ) | ( ~n8754 & n30849 ) | ( n13131 & n30849 ) ;
  assign n47164 = n4184 ^ n3876 ^ 1'b0 ;
  assign n47165 = ( n1526 & ~n33896 ) | ( n1526 & n47164 ) | ( ~n33896 & n47164 ) ;
  assign n47166 = n42437 ^ n25862 ^ n5939 ;
  assign n47167 = n40615 & ~n47166 ;
  assign n47168 = n4118 ^ n916 ^ 1'b0 ;
  assign n47169 = n23856 & n47168 ;
  assign n47170 = n8106 | n15075 ;
  assign n47171 = n23449 | n47170 ;
  assign n47172 = ( n11011 & n37036 ) | ( n11011 & ~n47171 ) | ( n37036 & ~n47171 ) ;
  assign n47173 = n45968 ^ n23826 ^ 1'b0 ;
  assign n47174 = ~n47172 & n47173 ;
  assign n47175 = ~n47169 & n47174 ;
  assign n47178 = n38535 ^ n10483 ^ 1'b0 ;
  assign n47176 = n39458 ^ n33003 ^ n6878 ;
  assign n47177 = n45037 | n47176 ;
  assign n47179 = n47178 ^ n47177 ^ 1'b0 ;
  assign n47180 = n34495 & n45617 ;
  assign n47181 = n47180 ^ n45538 ^ 1'b0 ;
  assign n47182 = n8081 & n27531 ;
  assign n47183 = ( n11497 & n41464 ) | ( n11497 & n47182 ) | ( n41464 & n47182 ) ;
  assign n47184 = ( n15738 & n17626 ) | ( n15738 & ~n23460 ) | ( n17626 & ~n23460 ) ;
  assign n47185 = n42682 ^ n38461 ^ n29071 ;
  assign n47186 = n34680 ^ n32676 ^ n6535 ;
  assign n47187 = n18885 & ~n24124 ;
  assign n47188 = n32654 & n47187 ;
  assign n47189 = ( ~n6460 & n13131 ) | ( ~n6460 & n47188 ) | ( n13131 & n47188 ) ;
  assign n47190 = n47189 ^ n41434 ^ n5602 ;
  assign n47192 = n1238 | n12125 ;
  assign n47191 = n1979 & ~n27750 ;
  assign n47193 = n47192 ^ n47191 ^ n42854 ;
  assign n47195 = n4842 & n10294 ;
  assign n47194 = n6388 | n29595 ;
  assign n47196 = n47195 ^ n47194 ^ 1'b0 ;
  assign n47197 = n46029 ^ n6235 ^ 1'b0 ;
  assign n47198 = n47196 | n47197 ;
  assign n47199 = ~n44179 & n47198 ;
  assign n47200 = ( ~n3597 & n47193 ) | ( ~n3597 & n47199 ) | ( n47193 & n47199 ) ;
  assign n47201 = ~n11540 & n21582 ;
  assign n47204 = n3735 | n6761 ;
  assign n47205 = n47204 ^ n16527 ^ 1'b0 ;
  assign n47202 = n22727 ^ n12528 ^ n7110 ;
  assign n47203 = n35433 & ~n47202 ;
  assign n47206 = n47205 ^ n47203 ^ 1'b0 ;
  assign n47207 = ~n8199 & n47206 ;
  assign n47208 = n47207 ^ n7485 ^ 1'b0 ;
  assign n47209 = ~n3800 & n5517 ;
  assign n47210 = n16539 & n47209 ;
  assign n47212 = n25122 ^ n7682 ^ n4397 ;
  assign n47213 = ( n4923 & n6420 ) | ( n4923 & ~n47212 ) | ( n6420 & ~n47212 ) ;
  assign n47211 = n22745 ^ n6806 ^ 1'b0 ;
  assign n47214 = n47213 ^ n47211 ^ n19033 ;
  assign n47215 = ~n27749 & n47214 ;
  assign n47216 = ( x146 & n47210 ) | ( x146 & n47215 ) | ( n47210 & n47215 ) ;
  assign n47219 = n8834 ^ n7782 ^ n4033 ;
  assign n47217 = n43426 ^ n36156 ^ 1'b0 ;
  assign n47218 = ~n27128 & n47217 ;
  assign n47220 = n47219 ^ n47218 ^ n24984 ;
  assign n47221 = n47220 ^ n30306 ^ n1287 ;
  assign n47222 = n14579 & n22599 ;
  assign n47223 = ( n24197 & n44709 ) | ( n24197 & ~n47222 ) | ( n44709 & ~n47222 ) ;
  assign n47224 = n39714 ^ n8308 ^ 1'b0 ;
  assign n47225 = n41719 & n47224 ;
  assign n47226 = n19315 ^ n2433 ^ 1'b0 ;
  assign n47227 = n15625 ^ n10333 ^ n1058 ;
  assign n47228 = ( ~n25252 & n45936 ) | ( ~n25252 & n47227 ) | ( n45936 & n47227 ) ;
  assign n47229 = n31237 ^ n8892 ^ n766 ;
  assign n47230 = ( n5929 & n28462 ) | ( n5929 & ~n47229 ) | ( n28462 & ~n47229 ) ;
  assign n47231 = n47230 ^ n5957 ^ 1'b0 ;
  assign n47232 = n15885 | n47231 ;
  assign n47233 = n14318 ^ n8644 ^ n3534 ;
  assign n47234 = ~n13917 & n47233 ;
  assign n47235 = ~n1801 & n47234 ;
  assign n47236 = n25164 ^ n24385 ^ n2705 ;
  assign n47237 = ( n4279 & n33564 ) | ( n4279 & n47236 ) | ( n33564 & n47236 ) ;
  assign n47238 = ~n21637 & n47237 ;
  assign n47239 = ~n27455 & n47238 ;
  assign n47240 = n47239 ^ n35247 ^ n3780 ;
  assign n47241 = ( n1590 & n2629 ) | ( n1590 & ~n9949 ) | ( n2629 & ~n9949 ) ;
  assign n47242 = n47241 ^ n36727 ^ n28941 ;
  assign n47243 = ( n312 & ~n31928 ) | ( n312 & n34146 ) | ( ~n31928 & n34146 ) ;
  assign n47244 = x133 & ~n3710 ;
  assign n47245 = n47244 ^ n11692 ^ 1'b0 ;
  assign n47246 = n38464 ^ n37075 ^ n10618 ;
  assign n47247 = ( n29685 & ~n47245 ) | ( n29685 & n47246 ) | ( ~n47245 & n47246 ) ;
  assign n47248 = ( ~n25529 & n28711 ) | ( ~n25529 & n33397 ) | ( n28711 & n33397 ) ;
  assign n47249 = ~n463 & n41166 ;
  assign n47250 = ~n12697 & n47249 ;
  assign n47251 = x71 & ~n47250 ;
  assign n47252 = ~n1198 & n47251 ;
  assign n47253 = ( ~n4897 & n11752 ) | ( ~n4897 & n41618 ) | ( n11752 & n41618 ) ;
  assign n47254 = ~n11043 & n35633 ;
  assign n47255 = ~n34258 & n47254 ;
  assign n47256 = ~n47253 & n47255 ;
  assign n47257 = n5525 | n8412 ;
  assign n47258 = n47257 ^ n9318 ^ 1'b0 ;
  assign n47259 = n28250 | n37231 ;
  assign n47260 = n47258 | n47259 ;
  assign n47261 = n23013 & ~n27653 ;
  assign n47262 = n47261 ^ n38241 ^ n12792 ;
  assign n47263 = n11941 & ~n27047 ;
  assign n47264 = n8684 ^ n2866 ^ 1'b0 ;
  assign n47265 = n5911 & ~n24267 ;
  assign n47266 = ( n5811 & ~n15411 ) | ( n5811 & n39706 ) | ( ~n15411 & n39706 ) ;
  assign n47267 = n47266 ^ n47115 ^ n24648 ;
  assign n47268 = ( n10503 & ~n14167 ) | ( n10503 & n41132 ) | ( ~n14167 & n41132 ) ;
  assign n47269 = n10352 | n47268 ;
  assign n47270 = n10347 ^ n6168 ^ 1'b0 ;
  assign n47271 = n555 & ~n5609 ;
  assign n47272 = n40056 & n47271 ;
  assign n47273 = ( n4282 & n4992 ) | ( n4282 & ~n12387 ) | ( n4992 & ~n12387 ) ;
  assign n47274 = ~n47272 & n47273 ;
  assign n47275 = n47274 ^ n1356 ^ 1'b0 ;
  assign n47276 = n12198 & ~n47275 ;
  assign n47277 = n47276 ^ n19457 ^ 1'b0 ;
  assign n47278 = n1324 | n31816 ;
  assign n47279 = n2510 & n42260 ;
  assign n47280 = ~n44881 & n47279 ;
  assign n47281 = ~n29225 & n47280 ;
  assign n47282 = n17919 ^ n8598 ^ n3471 ;
  assign n47283 = n47282 ^ n44482 ^ n21565 ;
  assign n47284 = ~n3505 & n13948 ;
  assign n47285 = ( n7223 & n14968 ) | ( n7223 & n47284 ) | ( n14968 & n47284 ) ;
  assign n47286 = ( n17400 & ~n22362 ) | ( n17400 & n36840 ) | ( ~n22362 & n36840 ) ;
  assign n47287 = ( ~n16628 & n47285 ) | ( ~n16628 & n47286 ) | ( n47285 & n47286 ) ;
  assign n47288 = n40021 ^ n19503 ^ 1'b0 ;
  assign n47289 = n34332 & n47288 ;
  assign n47290 = ~n24983 & n47289 ;
  assign n47291 = ( n1040 & n5368 ) | ( n1040 & n5613 ) | ( n5368 & n5613 ) ;
  assign n47292 = n47291 ^ n3169 ^ x16 ;
  assign n47293 = n37362 ^ n7932 ^ 1'b0 ;
  assign n47294 = n21197 ^ n8668 ^ 1'b0 ;
  assign n47295 = n47294 ^ n36159 ^ n14485 ;
  assign n47296 = n47295 ^ n34596 ^ n6925 ;
  assign n47297 = n1217 | n11446 ;
  assign n47298 = n47297 ^ n29635 ^ 1'b0 ;
  assign n47300 = n16649 & ~n23757 ;
  assign n47299 = n3676 & n22757 ;
  assign n47301 = n47300 ^ n47299 ^ 1'b0 ;
  assign n47304 = ( n6229 & n20221 ) | ( n6229 & n41576 ) | ( n20221 & n41576 ) ;
  assign n47305 = n47304 ^ n35250 ^ n16552 ;
  assign n47302 = n31865 ^ n6619 ^ 1'b0 ;
  assign n47303 = ~n29724 & n47302 ;
  assign n47306 = n47305 ^ n47303 ^ 1'b0 ;
  assign n47307 = n40245 ^ n35812 ^ n33557 ;
  assign n47308 = n7633 ^ n3524 ^ 1'b0 ;
  assign n47309 = n47308 ^ n2878 ^ n2162 ;
  assign n47310 = ( x101 & n20729 ) | ( x101 & ~n44662 ) | ( n20729 & ~n44662 ) ;
  assign n47311 = ( n5700 & n33603 ) | ( n5700 & n41545 ) | ( n33603 & n41545 ) ;
  assign n47312 = n47311 ^ n26296 ^ n18704 ;
  assign n47313 = ( n27103 & ~n47310 ) | ( n27103 & n47312 ) | ( ~n47310 & n47312 ) ;
  assign n47314 = n31824 ^ n19532 ^ 1'b0 ;
  assign n47315 = n1230 & n29703 ;
  assign n47316 = ~n25642 & n47315 ;
  assign n47317 = n47316 ^ n30234 ^ n24463 ;
  assign n47318 = n31363 ^ n27836 ^ n21320 ;
  assign n47319 = n31760 | n44382 ;
  assign n47320 = n47319 ^ n27775 ^ 1'b0 ;
  assign n47321 = n20715 ^ n10128 ^ 1'b0 ;
  assign n47322 = ~n37006 & n47321 ;
  assign n47323 = n13018 ^ n11782 ^ 1'b0 ;
  assign n47324 = n6658 | n47323 ;
  assign n47325 = n47324 ^ n13712 ^ n12953 ;
  assign n47326 = n47325 ^ n39131 ^ n24628 ;
  assign n47327 = ( n11951 & n13828 ) | ( n11951 & n30904 ) | ( n13828 & n30904 ) ;
  assign n47328 = n47327 ^ n41861 ^ n6226 ;
  assign n47329 = n47328 ^ n6994 ^ 1'b0 ;
  assign n47330 = n11858 ^ n11144 ^ n4209 ;
  assign n47331 = ( n12673 & n22142 ) | ( n12673 & ~n47330 ) | ( n22142 & ~n47330 ) ;
  assign n47332 = n23694 ^ n2412 ^ 1'b0 ;
  assign n47333 = n14395 & ~n47332 ;
  assign n47334 = ( ~n3444 & n4346 ) | ( ~n3444 & n47333 ) | ( n4346 & n47333 ) ;
  assign n47335 = n11017 & n13100 ;
  assign n47336 = n24354 & ~n47335 ;
  assign n47337 = n47336 ^ n10642 ^ n711 ;
  assign n47338 = n17136 & ~n44188 ;
  assign n47339 = ( n5329 & n27848 ) | ( n5329 & n47338 ) | ( n27848 & n47338 ) ;
  assign n47340 = n20753 ^ n8285 ^ n4415 ;
  assign n47341 = n47340 ^ n31952 ^ 1'b0 ;
  assign n47342 = ~n47339 & n47341 ;
  assign n47343 = ~n1733 & n2943 ;
  assign n47344 = n47343 ^ n1131 ^ 1'b0 ;
  assign n47345 = n39662 & ~n47344 ;
  assign n47346 = ~n10368 & n17106 ;
  assign n47347 = n14026 & n47346 ;
  assign n47348 = n15822 ^ n13272 ^ n4781 ;
  assign n47349 = n47348 ^ n13452 ^ n7821 ;
  assign n47350 = n47349 ^ n33910 ^ n28206 ;
  assign n47351 = n21943 ^ n17154 ^ n1904 ;
  assign n47352 = n47351 ^ n41150 ^ n29789 ;
  assign n47353 = ( ~n5923 & n23679 ) | ( ~n5923 & n27404 ) | ( n23679 & n27404 ) ;
  assign n47354 = n20516 & n47353 ;
  assign n47355 = ( ~n34823 & n39197 ) | ( ~n34823 & n46558 ) | ( n39197 & n46558 ) ;
  assign n47356 = n21334 ^ n8279 ^ n4272 ;
  assign n47357 = ( n33777 & n38789 ) | ( n33777 & n47356 ) | ( n38789 & n47356 ) ;
  assign n47358 = ( n19102 & n47355 ) | ( n19102 & n47357 ) | ( n47355 & n47357 ) ;
  assign n47359 = n28028 ^ n16624 ^ n8819 ;
  assign n47360 = ( ~n5438 & n11625 ) | ( ~n5438 & n25773 ) | ( n11625 & n25773 ) ;
  assign n47361 = ~n17400 & n39455 ;
  assign n47362 = ~n18222 & n47361 ;
  assign n47363 = n25901 ^ n15521 ^ 1'b0 ;
  assign n47364 = n36513 & n47363 ;
  assign n47366 = n34021 ^ n17368 ^ n16624 ;
  assign n47367 = ( n552 & n19044 ) | ( n552 & ~n47366 ) | ( n19044 & ~n47366 ) ;
  assign n47365 = n21103 | n37179 ;
  assign n47368 = n47367 ^ n47365 ^ 1'b0 ;
  assign n47369 = ~n3581 & n47368 ;
  assign n47370 = n47369 ^ n40502 ^ 1'b0 ;
  assign n47371 = n16013 ^ n10825 ^ 1'b0 ;
  assign n47372 = ( n8302 & n14513 ) | ( n8302 & ~n23671 ) | ( n14513 & ~n23671 ) ;
  assign n47373 = n42294 ^ n25480 ^ n7000 ;
  assign n47374 = ( n10821 & n47372 ) | ( n10821 & ~n47373 ) | ( n47372 & ~n47373 ) ;
  assign n47375 = ( n390 & n8193 ) | ( n390 & n37306 ) | ( n8193 & n37306 ) ;
  assign n47376 = ( n2242 & n9518 ) | ( n2242 & n22981 ) | ( n9518 & n22981 ) ;
  assign n47377 = n24297 ^ n19955 ^ 1'b0 ;
  assign n47378 = ~n1722 & n47377 ;
  assign n47379 = ( ~n13859 & n15143 ) | ( ~n13859 & n47378 ) | ( n15143 & n47378 ) ;
  assign n47380 = n29493 ^ n27669 ^ 1'b0 ;
  assign n47381 = ( ~n15321 & n22450 ) | ( ~n15321 & n47380 ) | ( n22450 & n47380 ) ;
  assign n47382 = n9766 ^ n2202 ^ 1'b0 ;
  assign n47383 = n31919 | n47382 ;
  assign n47384 = ~n16748 & n27368 ;
  assign n47385 = n47384 ^ n2457 ^ 1'b0 ;
  assign n47386 = n28580 ^ n5309 ^ n2903 ;
  assign n47387 = n5453 | n47386 ;
  assign n47388 = n47387 ^ n21583 ^ 1'b0 ;
  assign n47389 = n36621 ^ n13940 ^ n11219 ;
  assign n47390 = n39663 ^ n871 ^ n598 ;
  assign n47391 = ( n35527 & n47389 ) | ( n35527 & ~n47390 ) | ( n47389 & ~n47390 ) ;
  assign n47392 = n42861 ^ n36365 ^ n30666 ;
  assign n47393 = n35485 ^ n23454 ^ n6908 ;
  assign n47394 = n31721 ^ n18751 ^ n7303 ;
  assign n47395 = ( ~n4614 & n44986 ) | ( ~n4614 & n47394 ) | ( n44986 & n47394 ) ;
  assign n47396 = ( ~n24961 & n47393 ) | ( ~n24961 & n47395 ) | ( n47393 & n47395 ) ;
  assign n47397 = n23172 ^ n20180 ^ 1'b0 ;
  assign n47398 = n44991 | n47397 ;
  assign n47399 = n40821 ^ n7367 ^ n1213 ;
  assign n47400 = ( n17601 & n37798 ) | ( n17601 & n47399 ) | ( n37798 & n47399 ) ;
  assign n47401 = n36312 ^ n35710 ^ n5418 ;
  assign n47402 = n11171 & ~n23032 ;
  assign n47403 = n47402 ^ n33327 ^ 1'b0 ;
  assign n47404 = n5645 & ~n40500 ;
  assign n47405 = n47404 ^ n17876 ^ 1'b0 ;
  assign n47406 = n47368 & n47405 ;
  assign n47407 = n47403 & n47406 ;
  assign n47408 = n27638 & n35658 ;
  assign n47409 = ~n30899 & n47408 ;
  assign n47410 = ( n7010 & n14170 ) | ( n7010 & ~n21717 ) | ( n14170 & ~n21717 ) ;
  assign n47411 = n15988 & n17397 ;
  assign n47412 = ( n25355 & n47410 ) | ( n25355 & ~n47411 ) | ( n47410 & ~n47411 ) ;
  assign n47414 = n32266 & ~n42068 ;
  assign n47413 = ~n11117 & n20135 ;
  assign n47415 = n47414 ^ n47413 ^ n36509 ;
  assign n47416 = n47415 ^ n29760 ^ n16611 ;
  assign n47417 = ~n14172 & n41441 ;
  assign n47418 = n2793 & ~n16159 ;
  assign n47419 = ~n3704 & n47418 ;
  assign n47420 = n28838 | n47419 ;
  assign n47421 = n47420 ^ n5107 ^ 1'b0 ;
  assign n47422 = ( n14744 & ~n23955 ) | ( n14744 & n24017 ) | ( ~n23955 & n24017 ) ;
  assign n47423 = ~n30441 & n47422 ;
  assign n47424 = n47421 & n47423 ;
  assign n47425 = n47417 & ~n47424 ;
  assign n47426 = ( ~n2004 & n14226 ) | ( ~n2004 & n18775 ) | ( n14226 & n18775 ) ;
  assign n47427 = n16064 ^ n10352 ^ 1'b0 ;
  assign n47428 = ( n13562 & ~n47426 ) | ( n13562 & n47427 ) | ( ~n47426 & n47427 ) ;
  assign n47429 = ( n4697 & ~n19040 ) | ( n4697 & n29631 ) | ( ~n19040 & n29631 ) ;
  assign n47430 = ~n19362 & n22156 ;
  assign n47431 = n47430 ^ n40415 ^ 1'b0 ;
  assign n47432 = n34139 ^ n25639 ^ n6768 ;
  assign n47433 = n39540 & n47432 ;
  assign n47434 = ~n13348 & n18068 ;
  assign n47435 = n37001 & n47434 ;
  assign n47436 = n12195 ^ n2763 ^ 1'b0 ;
  assign n47437 = ( n1495 & ~n7813 ) | ( n1495 & n34389 ) | ( ~n7813 & n34389 ) ;
  assign n47442 = n26708 ^ n24516 ^ n1808 ;
  assign n47443 = ( n34087 & ~n42138 ) | ( n34087 & n47442 ) | ( ~n42138 & n47442 ) ;
  assign n47438 = n2275 | n7572 ;
  assign n47439 = n47438 ^ n10538 ^ 1'b0 ;
  assign n47440 = ( n4042 & n12296 ) | ( n4042 & ~n47439 ) | ( n12296 & ~n47439 ) ;
  assign n47441 = ( n8903 & n11577 ) | ( n8903 & n47440 ) | ( n11577 & n47440 ) ;
  assign n47444 = n47443 ^ n47441 ^ n23839 ;
  assign n47445 = n2120 & n10378 ;
  assign n47446 = n47445 ^ n33804 ^ 1'b0 ;
  assign n47447 = n26834 | n47446 ;
  assign n47448 = ( n12068 & n15593 ) | ( n12068 & n47447 ) | ( n15593 & n47447 ) ;
  assign n47449 = n47448 ^ n35986 ^ n11241 ;
  assign n47450 = n15009 ^ n10352 ^ 1'b0 ;
  assign n47451 = n6038 & n47450 ;
  assign n47452 = n47451 ^ n38582 ^ n16815 ;
  assign n47453 = ( n2347 & ~n24323 ) | ( n2347 & n28910 ) | ( ~n24323 & n28910 ) ;
  assign n47455 = n24836 ^ n16266 ^ n4823 ;
  assign n47454 = n28451 | n30556 ;
  assign n47456 = n47455 ^ n47454 ^ 1'b0 ;
  assign n47457 = ( x248 & n16759 ) | ( x248 & n45964 ) | ( n16759 & n45964 ) ;
  assign n47458 = ( ~n9176 & n16921 ) | ( ~n9176 & n18188 ) | ( n16921 & n18188 ) ;
  assign n47459 = n47458 ^ n42859 ^ n33941 ;
  assign n47460 = n853 & n15518 ;
  assign n47461 = n8503 & n47460 ;
  assign n47462 = ( n20557 & ~n35382 ) | ( n20557 & n47461 ) | ( ~n35382 & n47461 ) ;
  assign n47463 = n22063 ^ n16733 ^ 1'b0 ;
  assign n47464 = ~n18861 & n47463 ;
  assign n47465 = n1900 & n47464 ;
  assign n47466 = ( ~n1550 & n4957 ) | ( ~n1550 & n9979 ) | ( n4957 & n9979 ) ;
  assign n47467 = ( n5811 & ~n7498 ) | ( n5811 & n47466 ) | ( ~n7498 & n47466 ) ;
  assign n47468 = n43852 ^ n7307 ^ 1'b0 ;
  assign n47469 = ( n10219 & n44704 ) | ( n10219 & ~n47468 ) | ( n44704 & ~n47468 ) ;
  assign n47470 = n47469 ^ n44140 ^ n33587 ;
  assign n47471 = n7863 ^ n6604 ^ n5002 ;
  assign n47472 = n15003 & n47471 ;
  assign n47473 = ( n707 & n22243 ) | ( n707 & n47472 ) | ( n22243 & n47472 ) ;
  assign n47474 = n5962 & ~n47473 ;
  assign n47475 = ( ~n8547 & n26924 ) | ( ~n8547 & n43155 ) | ( n26924 & n43155 ) ;
  assign n47477 = n22856 ^ n14352 ^ n13933 ;
  assign n47476 = ( n10817 & n20822 ) | ( n10817 & ~n31581 ) | ( n20822 & ~n31581 ) ;
  assign n47478 = n47477 ^ n47476 ^ n5894 ;
  assign n47479 = ( ~x42 & n3926 ) | ( ~x42 & n21535 ) | ( n3926 & n21535 ) ;
  assign n47480 = n27491 ^ n2896 ^ 1'b0 ;
  assign n47481 = n28948 & ~n47480 ;
  assign n47482 = n21442 ^ n5045 ^ n1553 ;
  assign n47483 = n22634 & ~n47482 ;
  assign n47484 = n47483 ^ n12744 ^ 1'b0 ;
  assign n47485 = n20310 & ~n37501 ;
  assign n47486 = n4667 & n47485 ;
  assign n47487 = n46979 ^ n28698 ^ n8228 ;
  assign n47488 = n44744 ^ n30683 ^ n15829 ;
  assign n47489 = ( n5696 & n15738 ) | ( n5696 & n31956 ) | ( n15738 & n31956 ) ;
  assign n47490 = ~n8506 & n22420 ;
  assign n47491 = n39998 & n47490 ;
  assign n47492 = n27055 ^ n1410 ^ 1'b0 ;
  assign n47493 = n13802 & ~n47492 ;
  assign n47494 = n44183 & ~n47493 ;
  assign n47495 = n47494 ^ n18038 ^ 1'b0 ;
  assign n47496 = n9348 & ~n41794 ;
  assign n47497 = ~n32238 & n32350 ;
  assign n47498 = ~n21289 & n47497 ;
  assign n47499 = n35917 & n47498 ;
  assign n47500 = ~n5207 & n5232 ;
  assign n47501 = n8539 & n47500 ;
  assign n47502 = ( n2381 & ~n7876 ) | ( n2381 & n47501 ) | ( ~n7876 & n47501 ) ;
  assign n47503 = n47502 ^ n34849 ^ n8184 ;
  assign n47504 = ~n10152 & n12036 ;
  assign n47505 = n22385 & n47504 ;
  assign n47506 = n47505 ^ n12453 ^ 1'b0 ;
  assign n47507 = n16494 & n47506 ;
  assign n47508 = n47507 ^ n37857 ^ n19480 ;
  assign n47509 = ( n15748 & n23914 ) | ( n15748 & n46261 ) | ( n23914 & n46261 ) ;
  assign n47510 = n4911 | n12550 ;
  assign n47511 = n47510 ^ n36027 ^ n28020 ;
  assign n47512 = ~n28019 & n35647 ;
  assign n47513 = n9072 & n47512 ;
  assign n47514 = n12853 & ~n44548 ;
  assign n47515 = ( n1520 & ~n7147 ) | ( n1520 & n11102 ) | ( ~n7147 & n11102 ) ;
  assign n47516 = ( n4527 & n30871 ) | ( n4527 & ~n47515 ) | ( n30871 & ~n47515 ) ;
  assign n47517 = n3574 & ~n38800 ;
  assign n47518 = ~n47516 & n47517 ;
  assign n47521 = n21111 ^ n1194 ^ 1'b0 ;
  assign n47519 = n20899 ^ n11021 ^ 1'b0 ;
  assign n47520 = ( n23460 & ~n23706 ) | ( n23460 & n47519 ) | ( ~n23706 & n47519 ) ;
  assign n47522 = n47521 ^ n47520 ^ n29930 ;
  assign n47523 = ( ~n6882 & n16838 ) | ( ~n6882 & n31079 ) | ( n16838 & n31079 ) ;
  assign n47524 = ~n20041 & n32157 ;
  assign n47525 = n15411 ^ n10523 ^ n2848 ;
  assign n47526 = n10601 & n17972 ;
  assign n47527 = ( n9249 & ~n31936 ) | ( n9249 & n47526 ) | ( ~n31936 & n47526 ) ;
  assign n47528 = ( n3573 & ~n16601 ) | ( n3573 & n47527 ) | ( ~n16601 & n47527 ) ;
  assign n47529 = ( ~n30678 & n40175 ) | ( ~n30678 & n45909 ) | ( n40175 & n45909 ) ;
  assign n47530 = n31908 | n44596 ;
  assign n47531 = n47529 | n47530 ;
  assign n47533 = n5037 ^ n3944 ^ 1'b0 ;
  assign n47532 = n35824 & ~n46264 ;
  assign n47534 = n47533 ^ n47532 ^ 1'b0 ;
  assign n47535 = ~n32438 & n47534 ;
  assign n47536 = n15600 & n47535 ;
  assign n47538 = ( n1762 & n4850 ) | ( n1762 & ~n10676 ) | ( n4850 & ~n10676 ) ;
  assign n47537 = n369 | n6454 ;
  assign n47539 = n47538 ^ n47537 ^ 1'b0 ;
  assign n47540 = ( ~n7883 & n13067 ) | ( ~n7883 & n42184 ) | ( n13067 & n42184 ) ;
  assign n47542 = n23915 ^ n9920 ^ n7322 ;
  assign n47543 = n47542 ^ n26562 ^ n17329 ;
  assign n47541 = n23637 ^ n9295 ^ n4230 ;
  assign n47544 = n47543 ^ n47541 ^ 1'b0 ;
  assign n47545 = n28463 ^ n23564 ^ n7756 ;
  assign n47546 = n25940 & ~n47545 ;
  assign n47547 = n650 & ~n6587 ;
  assign n47548 = n47547 ^ n41737 ^ n15194 ;
  assign n47549 = n42251 ^ n22927 ^ n19369 ;
  assign n47550 = n26281 ^ n6699 ^ 1'b0 ;
  assign n47551 = n2913 & n47550 ;
  assign n47556 = x75 & ~n17386 ;
  assign n47557 = n17386 & n47556 ;
  assign n47555 = ( n766 & n17549 ) | ( n766 & n19528 ) | ( n17549 & n19528 ) ;
  assign n47558 = n47557 ^ n47555 ^ 1'b0 ;
  assign n47552 = n34775 ^ n3337 ^ 1'b0 ;
  assign n47553 = n3948 & n47552 ;
  assign n47554 = ( n266 & ~n17855 ) | ( n266 & n47553 ) | ( ~n17855 & n47553 ) ;
  assign n47559 = n47558 ^ n47554 ^ n25126 ;
  assign n47560 = n18225 & n47559 ;
  assign n47561 = x67 & n30139 ;
  assign n47562 = ~n9349 & n47561 ;
  assign n47563 = n45458 ^ n23067 ^ 1'b0 ;
  assign n47564 = n13200 & n47563 ;
  assign n47565 = n1705 & n39827 ;
  assign n47566 = n8027 | n47565 ;
  assign n47567 = n47566 ^ n1407 ^ 1'b0 ;
  assign n47568 = n47567 ^ n28835 ^ n14964 ;
  assign n47569 = n22625 ^ n12629 ^ n9892 ;
  assign n47570 = ( n264 & n18602 ) | ( n264 & ~n47569 ) | ( n18602 & ~n47569 ) ;
  assign n47571 = n34595 ^ n33680 ^ n28933 ;
  assign n47572 = ( ~n22787 & n47570 ) | ( ~n22787 & n47571 ) | ( n47570 & n47571 ) ;
  assign n47573 = n47572 ^ n22131 ^ 1'b0 ;
  assign n47574 = n18200 & ~n40367 ;
  assign n47575 = ( ~n11621 & n13901 ) | ( ~n11621 & n33452 ) | ( n13901 & n33452 ) ;
  assign n47576 = n47575 ^ n24294 ^ n5721 ;
  assign n47577 = n47576 ^ n42085 ^ n12836 ;
  assign n47578 = n31189 ^ n24370 ^ n22180 ;
  assign n47579 = n47578 ^ n37946 ^ n24765 ;
  assign n47580 = n15986 & ~n22270 ;
  assign n47581 = n8373 & n47580 ;
  assign n47582 = ( n4812 & ~n8571 ) | ( n4812 & n23601 ) | ( ~n8571 & n23601 ) ;
  assign n47583 = ( n2161 & n47581 ) | ( n2161 & n47582 ) | ( n47581 & n47582 ) ;
  assign n47584 = n47583 ^ n3588 ^ 1'b0 ;
  assign n47585 = ~n29101 & n47584 ;
  assign n47586 = n47585 ^ n19648 ^ n19543 ;
  assign n47587 = ( n26823 & n32282 ) | ( n26823 & n47586 ) | ( n32282 & n47586 ) ;
  assign n47588 = n33268 ^ n13494 ^ 1'b0 ;
  assign n47589 = n4986 & ~n38634 ;
  assign n47590 = n2720 & n47589 ;
  assign n47591 = ( ~n1140 & n7942 ) | ( ~n1140 & n16338 ) | ( n7942 & n16338 ) ;
  assign n47592 = n47591 ^ n8303 ^ n2164 ;
  assign n47593 = ~n19818 & n20945 ;
  assign n47594 = n47593 ^ n38538 ^ 1'b0 ;
  assign n47595 = ( n2408 & n17732 ) | ( n2408 & n20972 ) | ( n17732 & n20972 ) ;
  assign n47599 = ( ~n24003 & n24075 ) | ( ~n24003 & n43870 ) | ( n24075 & n43870 ) ;
  assign n47596 = n1758 & ~n2830 ;
  assign n47597 = n47596 ^ n27460 ^ 1'b0 ;
  assign n47598 = ( n15397 & n33575 ) | ( n15397 & ~n47597 ) | ( n33575 & ~n47597 ) ;
  assign n47600 = n47599 ^ n47598 ^ 1'b0 ;
  assign n47602 = n10428 & ~n20121 ;
  assign n47601 = n8173 | n35607 ;
  assign n47603 = n47602 ^ n47601 ^ 1'b0 ;
  assign n47604 = n19917 ^ n15782 ^ 1'b0 ;
  assign n47605 = n29671 | n47604 ;
  assign n47606 = n47605 ^ n27016 ^ 1'b0 ;
  assign n47607 = ( n3795 & n6429 ) | ( n3795 & ~n6646 ) | ( n6429 & ~n6646 ) ;
  assign n47608 = n5172 ^ n1121 ^ 1'b0 ;
  assign n47609 = n5378 & n47608 ;
  assign n47610 = n47609 ^ n41577 ^ n1549 ;
  assign n47611 = ( n19578 & n47607 ) | ( n19578 & n47610 ) | ( n47607 & n47610 ) ;
  assign n47612 = n3633 & ~n11462 ;
  assign n47613 = ( n23574 & n45072 ) | ( n23574 & ~n47612 ) | ( n45072 & ~n47612 ) ;
  assign n47615 = ~n3741 & n15062 ;
  assign n47614 = n30064 ^ n10656 ^ n7225 ;
  assign n47616 = n47615 ^ n47614 ^ n33765 ;
  assign n47617 = n47616 ^ n44456 ^ n11661 ;
  assign n47618 = ( n3310 & n6059 ) | ( n3310 & n30530 ) | ( n6059 & n30530 ) ;
  assign n47619 = ( n8900 & n26867 ) | ( n8900 & n42448 ) | ( n26867 & n42448 ) ;
  assign n47620 = n13045 ^ n8583 ^ n6737 ;
  assign n47621 = n3241 & n45452 ;
  assign n47622 = n47621 ^ n29634 ^ n5097 ;
  assign n47623 = ( n37254 & n40051 ) | ( n37254 & n47622 ) | ( n40051 & n47622 ) ;
  assign n47624 = ( ~n6500 & n28337 ) | ( ~n6500 & n47623 ) | ( n28337 & n47623 ) ;
  assign n47625 = ~n47620 & n47624 ;
  assign n47626 = n13118 & ~n38377 ;
  assign n47627 = n12136 & n47626 ;
  assign n47628 = ( n2125 & ~n17182 ) | ( n2125 & n17281 ) | ( ~n17182 & n17281 ) ;
  assign n47629 = n12471 | n26651 ;
  assign n47630 = n47628 & ~n47629 ;
  assign n47631 = n36339 ^ n18092 ^ n13109 ;
  assign n47635 = n14581 ^ n2427 ^ 1'b0 ;
  assign n47636 = ( ~n6527 & n26554 ) | ( ~n6527 & n47635 ) | ( n26554 & n47635 ) ;
  assign n47632 = n3701 & ~n32598 ;
  assign n47633 = ~x4 & n47632 ;
  assign n47634 = n47633 ^ n20596 ^ n9036 ;
  assign n47637 = n47636 ^ n47634 ^ n29059 ;
  assign n47638 = ( n17870 & n47631 ) | ( n17870 & ~n47637 ) | ( n47631 & ~n47637 ) ;
  assign n47639 = ( n916 & n19517 ) | ( n916 & ~n24196 ) | ( n19517 & ~n24196 ) ;
  assign n47640 = ( n13718 & n19098 ) | ( n13718 & n47639 ) | ( n19098 & n47639 ) ;
  assign n47641 = n47640 ^ n14892 ^ n9202 ;
  assign n47642 = n47641 ^ n15616 ^ 1'b0 ;
  assign n47643 = n37797 ^ n7314 ^ 1'b0 ;
  assign n47644 = n31008 ^ n29062 ^ n1955 ;
  assign n47645 = n3658 ^ n3325 ^ 1'b0 ;
  assign n47646 = ( ~n4166 & n23472 ) | ( ~n4166 & n47645 ) | ( n23472 & n47645 ) ;
  assign n47647 = n44953 ^ n14720 ^ n6841 ;
  assign n47648 = n17121 ^ n6052 ^ n1886 ;
  assign n47649 = n26286 ^ n11716 ^ 1'b0 ;
  assign n47650 = n18111 & ~n47649 ;
  assign n47651 = n1674 & ~n5475 ;
  assign n47652 = ~n8234 & n47651 ;
  assign n47653 = n2188 & n12696 ;
  assign n47654 = n47653 ^ n19814 ^ 1'b0 ;
  assign n47655 = ~n484 & n29281 ;
  assign n47656 = n41843 & n47655 ;
  assign n47657 = ( n3104 & n30863 ) | ( n3104 & ~n47656 ) | ( n30863 & ~n47656 ) ;
  assign n47658 = ( n21968 & n26311 ) | ( n21968 & ~n37111 ) | ( n26311 & ~n37111 ) ;
  assign n47659 = ~n7345 & n9507 ;
  assign n47660 = n47659 ^ n21782 ^ 1'b0 ;
  assign n47661 = n11550 | n19157 ;
  assign n47662 = n47661 ^ n11863 ^ 1'b0 ;
  assign n47663 = ( ~n2135 & n47660 ) | ( ~n2135 & n47662 ) | ( n47660 & n47662 ) ;
  assign n47667 = n32444 ^ n18002 ^ 1'b0 ;
  assign n47668 = n16296 & n47667 ;
  assign n47666 = n1972 | n25962 ;
  assign n47669 = n47668 ^ n47666 ^ 1'b0 ;
  assign n47664 = n29553 & ~n36796 ;
  assign n47665 = ~n45709 & n47664 ;
  assign n47670 = n47669 ^ n47665 ^ n11537 ;
  assign n47671 = n19523 ^ n3111 ^ 1'b0 ;
  assign n47672 = ( ~n13584 & n27110 ) | ( ~n13584 & n37578 ) | ( n27110 & n37578 ) ;
  assign n47673 = ( n5430 & ~n34487 ) | ( n5430 & n37069 ) | ( ~n34487 & n37069 ) ;
  assign n47674 = n9221 & n9642 ;
  assign n47675 = n47674 ^ n24088 ^ 1'b0 ;
  assign n47676 = n27480 ^ n22011 ^ 1'b0 ;
  assign n47677 = ~n11056 & n36019 ;
  assign n47678 = n47677 ^ n3715 ^ 1'b0 ;
  assign n47679 = n28876 ^ n16004 ^ 1'b0 ;
  assign n47680 = n9789 ^ n9571 ^ 1'b0 ;
  assign n47681 = ( n11697 & n45699 ) | ( n11697 & ~n47680 ) | ( n45699 & ~n47680 ) ;
  assign n47682 = n47681 ^ n47157 ^ n11433 ;
  assign n47683 = ( ~n9345 & n10615 ) | ( ~n9345 & n10949 ) | ( n10615 & n10949 ) ;
  assign n47684 = n47683 ^ n9787 ^ 1'b0 ;
  assign n47689 = n19795 ^ n5430 ^ n595 ;
  assign n47686 = n33931 ^ n26084 ^ n6375 ;
  assign n47687 = n45508 ^ n8258 ^ 1'b0 ;
  assign n47688 = n47686 & ~n47687 ;
  assign n47685 = n42106 | n42403 ;
  assign n47690 = n47689 ^ n47688 ^ n47685 ;
  assign n47691 = ( n4792 & n6711 ) | ( n4792 & n22887 ) | ( n6711 & n22887 ) ;
  assign n47692 = ( n3842 & ~n45231 ) | ( n3842 & n47691 ) | ( ~n45231 & n47691 ) ;
  assign n47693 = n47692 ^ n32527 ^ n23997 ;
  assign n47694 = n3284 & n34757 ;
  assign n47695 = n47694 ^ n2730 ^ 1'b0 ;
  assign n47696 = n7911 & n47695 ;
  assign n47697 = n3310 & n18368 ;
  assign n47698 = ~n546 & n47697 ;
  assign n47703 = n5466 | n34820 ;
  assign n47699 = n47112 ^ n25478 ^ n6531 ;
  assign n47700 = n21817 ^ n18972 ^ 1'b0 ;
  assign n47701 = ~n47699 & n47700 ;
  assign n47702 = n32553 & n47701 ;
  assign n47704 = n47703 ^ n47702 ^ 1'b0 ;
  assign n47706 = n22138 ^ n7651 ^ n4832 ;
  assign n47705 = n23591 ^ n9272 ^ n4784 ;
  assign n47707 = n47706 ^ n47705 ^ n20127 ;
  assign n47708 = n27376 ^ n12366 ^ n8499 ;
  assign n47709 = n23134 ^ n15359 ^ 1'b0 ;
  assign n47710 = ( n26933 & n46274 ) | ( n26933 & n47709 ) | ( n46274 & n47709 ) ;
  assign n47711 = ( n3351 & ~n31065 ) | ( n3351 & n47710 ) | ( ~n31065 & n47710 ) ;
  assign n47712 = n28620 ^ n24125 ^ n4666 ;
  assign n47713 = ( n3398 & ~n10700 ) | ( n3398 & n15533 ) | ( ~n10700 & n15533 ) ;
  assign n47714 = n47713 ^ n20789 ^ 1'b0 ;
  assign n47715 = n38480 ^ n17154 ^ 1'b0 ;
  assign n47716 = n37337 ^ n27267 ^ n21246 ;
  assign n47717 = ( n1230 & n14678 ) | ( n1230 & ~n47716 ) | ( n14678 & ~n47716 ) ;
  assign n47718 = n30306 & n47717 ;
  assign n47719 = n9356 & n46677 ;
  assign n47720 = n12521 & n47719 ;
  assign n47721 = n13778 | n39389 ;
  assign n47722 = ( ~x115 & n17812 ) | ( ~x115 & n34953 ) | ( n17812 & n34953 ) ;
  assign n47723 = n28168 ^ n24509 ^ 1'b0 ;
  assign n47724 = ( n28685 & n33328 ) | ( n28685 & ~n37933 ) | ( n33328 & ~n37933 ) ;
  assign n47725 = n47724 ^ n42895 ^ n3376 ;
  assign n47726 = ( n6564 & n7264 ) | ( n6564 & ~n40447 ) | ( n7264 & ~n40447 ) ;
  assign n47727 = n47726 ^ n12695 ^ n11534 ;
  assign n47728 = ( ~n8180 & n46701 ) | ( ~n8180 & n47727 ) | ( n46701 & n47727 ) ;
  assign n47729 = n47054 ^ n18768 ^ n10852 ;
  assign n47730 = n12294 ^ n3717 ^ 1'b0 ;
  assign n47731 = n10259 | n47730 ;
  assign n47732 = n18461 ^ n918 ^ 1'b0 ;
  assign n47733 = n18253 & ~n47732 ;
  assign n47734 = n9421 ^ n3763 ^ 1'b0 ;
  assign n47735 = n18036 ^ n17015 ^ n10943 ;
  assign n47736 = ( ~n3525 & n7973 ) | ( ~n3525 & n47735 ) | ( n7973 & n47735 ) ;
  assign n47737 = n44819 ^ n23004 ^ 1'b0 ;
  assign n47738 = n22189 ^ n14177 ^ n1539 ;
  assign n47739 = n47738 ^ n6986 ^ n5540 ;
  assign n47740 = n24799 ^ n20171 ^ n3654 ;
  assign n47741 = ( n43930 & n47739 ) | ( n43930 & n47740 ) | ( n47739 & n47740 ) ;
  assign n47742 = n12257 ^ n2231 ^ 1'b0 ;
  assign n47743 = n19861 & ~n47742 ;
  assign n47744 = n4034 | n47743 ;
  assign n47745 = n42523 ^ n22853 ^ 1'b0 ;
  assign n47746 = n27490 ^ n2559 ^ 1'b0 ;
  assign n47747 = n32582 | n47746 ;
  assign n47748 = ( n6747 & n12809 ) | ( n6747 & n24032 ) | ( n12809 & n24032 ) ;
  assign n47749 = ( n9452 & n46187 ) | ( n9452 & n47748 ) | ( n46187 & n47748 ) ;
  assign n47750 = n28274 | n47749 ;
  assign n47751 = ( n2612 & n28594 ) | ( n2612 & n47607 ) | ( n28594 & n47607 ) ;
  assign n47752 = ( ~n2781 & n23120 ) | ( ~n2781 & n47751 ) | ( n23120 & n47751 ) ;
  assign n47753 = ~n31769 & n47752 ;
  assign n47754 = ( n7010 & n7104 ) | ( n7010 & n32705 ) | ( n7104 & n32705 ) ;
  assign n47755 = ( n18458 & ~n20263 ) | ( n18458 & n34576 ) | ( ~n20263 & n34576 ) ;
  assign n47756 = n47755 ^ n26959 ^ x196 ;
  assign n47760 = n4970 & ~n29703 ;
  assign n47757 = ( n1372 & n1600 ) | ( n1372 & n17752 ) | ( n1600 & n17752 ) ;
  assign n47758 = n47757 ^ n33826 ^ 1'b0 ;
  assign n47759 = n45215 | n47758 ;
  assign n47761 = n47760 ^ n47759 ^ n27588 ;
  assign n47762 = n4349 & ~n21405 ;
  assign n47763 = ( n17829 & n28458 ) | ( n17829 & n40144 ) | ( n28458 & n40144 ) ;
  assign n47764 = ( n6517 & n17332 ) | ( n6517 & ~n30735 ) | ( n17332 & ~n30735 ) ;
  assign n47765 = n14595 ^ n11102 ^ n4507 ;
  assign n47766 = n47765 ^ n14813 ^ n11795 ;
  assign n47767 = n18351 | n47766 ;
  assign n47768 = n47767 ^ n32610 ^ 1'b0 ;
  assign n47769 = n47768 ^ n9294 ^ x226 ;
  assign n47770 = n6363 & ~n47769 ;
  assign n47771 = ~n36164 & n41114 ;
  assign n47772 = n46485 ^ n30302 ^ n28160 ;
  assign n47773 = n47772 ^ n40859 ^ n6445 ;
  assign n47774 = n11424 & n30255 ;
  assign n47775 = n47773 & n47774 ;
  assign n47776 = n5920 & ~n39215 ;
  assign n47777 = ( ~n4302 & n5329 ) | ( ~n4302 & n14073 ) | ( n5329 & n14073 ) ;
  assign n47778 = n47270 ^ n40754 ^ n15904 ;
  assign n47779 = n33654 ^ n30672 ^ n16147 ;
  assign n47780 = n30219 ^ n23028 ^ 1'b0 ;
  assign n47781 = ~n383 & n23017 ;
  assign n47782 = n8510 | n12600 ;
  assign n47783 = ~n19323 & n36469 ;
  assign n47784 = ~n26476 & n47783 ;
  assign n47785 = n47784 ^ n47685 ^ 1'b0 ;
  assign n47786 = n9574 & n36693 ;
  assign n47787 = n47786 ^ n26756 ^ 1'b0 ;
  assign n47788 = n39342 ^ n36087 ^ 1'b0 ;
  assign n47789 = n47787 & ~n47788 ;
  assign n47790 = ~n21357 & n24063 ;
  assign n47791 = ~n7801 & n47790 ;
  assign n47792 = n4804 & ~n47791 ;
  assign n47793 = ~n24350 & n47792 ;
  assign n47794 = n7863 ^ n7355 ^ 1'b0 ;
  assign n47795 = ( n7856 & n10370 ) | ( n7856 & n47794 ) | ( n10370 & n47794 ) ;
  assign n47796 = ( ~n25200 & n37938 ) | ( ~n25200 & n47795 ) | ( n37938 & n47795 ) ;
  assign n47799 = n2866 | n21017 ;
  assign n47800 = n1678 | n47799 ;
  assign n47797 = n6994 & ~n47681 ;
  assign n47798 = n11143 & n47797 ;
  assign n47801 = n47800 ^ n47798 ^ x176 ;
  assign n47802 = n11314 ^ n7925 ^ 1'b0 ;
  assign n47803 = ~n10422 & n47802 ;
  assign n47804 = n29460 ^ n7942 ^ n7866 ;
  assign n47805 = n47804 ^ n42117 ^ n30914 ;
  assign n47809 = n9904 ^ n9422 ^ 1'b0 ;
  assign n47808 = ( ~n21322 & n22874 ) | ( ~n21322 & n28963 ) | ( n22874 & n28963 ) ;
  assign n47806 = ~n28271 & n28363 ;
  assign n47807 = n47806 ^ n7476 ^ 1'b0 ;
  assign n47810 = n47809 ^ n47808 ^ n47807 ;
  assign n47815 = n12895 | n13539 ;
  assign n47816 = n36416 & ~n47815 ;
  assign n47813 = n41294 ^ n29493 ^ n2694 ;
  assign n47814 = ( n18103 & ~n22336 ) | ( n18103 & n47813 ) | ( ~n22336 & n47813 ) ;
  assign n47817 = n47816 ^ n47814 ^ n18830 ;
  assign n47811 = ( n3898 & ~n6262 ) | ( n3898 & n9228 ) | ( ~n6262 & n9228 ) ;
  assign n47812 = n47811 ^ n3387 ^ 1'b0 ;
  assign n47818 = n47817 ^ n47812 ^ 1'b0 ;
  assign n47819 = n23995 | n28573 ;
  assign n47820 = ( ~n3517 & n19795 ) | ( ~n3517 & n27401 ) | ( n19795 & n27401 ) ;
  assign n47821 = ~n6150 & n47820 ;
  assign n47823 = n42277 ^ n24626 ^ n1313 ;
  assign n47824 = ( n10665 & n29733 ) | ( n10665 & ~n47823 ) | ( n29733 & ~n47823 ) ;
  assign n47822 = n25033 & ~n39671 ;
  assign n47825 = n47824 ^ n47822 ^ 1'b0 ;
  assign n47826 = n14012 | n47825 ;
  assign n47827 = n47826 ^ n4812 ^ 1'b0 ;
  assign n47828 = n25861 ^ n9068 ^ 1'b0 ;
  assign n47829 = ( n38059 & ~n47543 ) | ( n38059 & n47828 ) | ( ~n47543 & n47828 ) ;
  assign n47830 = ( ~n7979 & n8104 ) | ( ~n7979 & n47829 ) | ( n8104 & n47829 ) ;
  assign n47831 = x70 & n11061 ;
  assign n47832 = ( ~n1341 & n4419 ) | ( ~n1341 & n27909 ) | ( n4419 & n27909 ) ;
  assign n47833 = n6518 ^ n3423 ^ 1'b0 ;
  assign n47834 = n28929 | n47833 ;
  assign n47835 = ( ~n3969 & n14284 ) | ( ~n3969 & n27480 ) | ( n14284 & n27480 ) ;
  assign n47836 = ( n5019 & ~n14482 ) | ( n5019 & n47835 ) | ( ~n14482 & n47835 ) ;
  assign n47837 = ( n42438 & n47834 ) | ( n42438 & ~n47836 ) | ( n47834 & ~n47836 ) ;
  assign n47838 = n23640 ^ n9151 ^ n3976 ;
  assign n47839 = n47838 ^ n25036 ^ n5974 ;
  assign n47840 = ( n11709 & n28301 ) | ( n11709 & n40245 ) | ( n28301 & n40245 ) ;
  assign n47843 = ( ~n460 & n1382 ) | ( ~n460 & n7098 ) | ( n1382 & n7098 ) ;
  assign n47844 = ( n6073 & n35616 ) | ( n6073 & ~n47843 ) | ( n35616 & ~n47843 ) ;
  assign n47841 = n29067 ^ n1916 ^ 1'b0 ;
  assign n47842 = n23698 & ~n47841 ;
  assign n47845 = n47844 ^ n47842 ^ n45505 ;
  assign n47846 = n24103 | n25573 ;
  assign n47847 = n28527 & ~n47846 ;
  assign n47848 = ( ~n2151 & n18857 ) | ( ~n2151 & n23768 ) | ( n18857 & n23768 ) ;
  assign n47849 = n31189 ^ n27249 ^ n11233 ;
  assign n47850 = n47652 | n47849 ;
  assign n47851 = n47848 | n47850 ;
  assign n47852 = ( n8337 & ~n11148 ) | ( n8337 & n21685 ) | ( ~n11148 & n21685 ) ;
  assign n47853 = n47852 ^ n16896 ^ 1'b0 ;
  assign n47854 = n31787 | n47853 ;
  assign n47855 = n585 | n25738 ;
  assign n47856 = n13350 & n15869 ;
  assign n47857 = ~n47855 & n47856 ;
  assign n47858 = n37690 ^ n10303 ^ 1'b0 ;
  assign n47859 = ( ~n17923 & n32497 ) | ( ~n17923 & n44367 ) | ( n32497 & n44367 ) ;
  assign n47860 = ( ~x176 & n20054 ) | ( ~x176 & n25465 ) | ( n20054 & n25465 ) ;
  assign n47861 = n45031 ^ n39803 ^ n9877 ;
  assign n47862 = ( n987 & n14433 ) | ( n987 & ~n18285 ) | ( n14433 & ~n18285 ) ;
  assign n47863 = n7553 & ~n14648 ;
  assign n47864 = ~n19443 & n47863 ;
  assign n47865 = n47864 ^ n11048 ^ 1'b0 ;
  assign n47866 = n6760 | n36762 ;
  assign n47867 = n47865 | n47866 ;
  assign n47868 = n482 | n13444 ;
  assign n47869 = n14099 | n47868 ;
  assign n47870 = ( n34047 & ~n43066 ) | ( n34047 & n44184 ) | ( ~n43066 & n44184 ) ;
  assign n47871 = ( n13017 & n20908 ) | ( n13017 & ~n47870 ) | ( n20908 & ~n47870 ) ;
  assign n47872 = n38910 ^ n32404 ^ 1'b0 ;
  assign n47873 = n17410 ^ n10623 ^ 1'b0 ;
  assign n47874 = n9458 | n13800 ;
  assign n47875 = n4456 & n6662 ;
  assign n47876 = n12315 & n47875 ;
  assign n47877 = n47876 ^ n25355 ^ n21249 ;
  assign n47883 = n3255 & n28394 ;
  assign n47884 = ~n9851 & n47883 ;
  assign n47878 = ( n473 & ~n12236 ) | ( n473 & n13597 ) | ( ~n12236 & n13597 ) ;
  assign n47879 = n14808 & ~n28117 ;
  assign n47880 = ~n47878 & n47879 ;
  assign n47881 = n45703 ^ n15419 ^ n787 ;
  assign n47882 = n47880 | n47881 ;
  assign n47885 = n47884 ^ n47882 ^ n17074 ;
  assign n47886 = n23018 ^ n4261 ^ 1'b0 ;
  assign n47887 = n1126 | n32363 ;
  assign n47888 = n47887 ^ n40371 ^ 1'b0 ;
  assign n47889 = n24670 ^ n17770 ^ 1'b0 ;
  assign n47890 = n287 & ~n47889 ;
  assign n47891 = n26697 & n47890 ;
  assign n47892 = ~n1537 & n20307 ;
  assign n47893 = n7233 ^ n4837 ^ 1'b0 ;
  assign n47894 = ( n2156 & n19143 ) | ( n2156 & n35762 ) | ( n19143 & n35762 ) ;
  assign n47895 = ( ~n7515 & n17966 ) | ( ~n7515 & n47894 ) | ( n17966 & n47894 ) ;
  assign n47896 = n44077 & ~n47895 ;
  assign n47897 = n4558 & n8912 ;
  assign n47898 = n47897 ^ n47583 ^ n15893 ;
  assign n47899 = ( ~n24536 & n28491 ) | ( ~n24536 & n35616 ) | ( n28491 & n35616 ) ;
  assign n47901 = n4991 & n14707 ;
  assign n47902 = n5892 & n47901 ;
  assign n47900 = ( n21821 & n24822 ) | ( n21821 & n27163 ) | ( n24822 & n27163 ) ;
  assign n47903 = n47902 ^ n47900 ^ n14525 ;
  assign n47904 = n47903 ^ n45535 ^ 1'b0 ;
  assign n47905 = ( n14299 & ~n19588 ) | ( n14299 & n27501 ) | ( ~n19588 & n27501 ) ;
  assign n47906 = n43524 & n47905 ;
  assign n47907 = ~n37955 & n47906 ;
  assign n47908 = n26889 & n27973 ;
  assign n47909 = ( n13651 & ~n16841 ) | ( n13651 & n41966 ) | ( ~n16841 & n41966 ) ;
  assign n47910 = ( n21194 & ~n47908 ) | ( n21194 & n47909 ) | ( ~n47908 & n47909 ) ;
  assign n47911 = n8184 & n24661 ;
  assign n47912 = ( n310 & n8189 ) | ( n310 & ~n47911 ) | ( n8189 & ~n47911 ) ;
  assign n47913 = ( n1973 & n24209 ) | ( n1973 & ~n41516 ) | ( n24209 & ~n41516 ) ;
  assign n47914 = ( n12176 & n27554 ) | ( n12176 & n29598 ) | ( n27554 & n29598 ) ;
  assign n47915 = n38089 ^ n22273 ^ 1'b0 ;
  assign n47916 = ~n8140 & n44411 ;
  assign n47917 = n29852 & n47916 ;
  assign n47918 = n47917 ^ n21497 ^ n3549 ;
  assign n47919 = ( ~n3432 & n8898 ) | ( ~n3432 & n47918 ) | ( n8898 & n47918 ) ;
  assign n47920 = ( n16976 & n35319 ) | ( n16976 & ~n47919 ) | ( n35319 & ~n47919 ) ;
  assign n47921 = n27838 ^ n24015 ^ 1'b0 ;
  assign n47922 = ~n47565 & n47921 ;
  assign n47923 = n10089 ^ n7539 ^ 1'b0 ;
  assign n47924 = n38386 ^ n26179 ^ 1'b0 ;
  assign n47925 = n30098 ^ n23281 ^ 1'b0 ;
  assign n47926 = ~n47924 & n47925 ;
  assign n47928 = ~n35254 & n46816 ;
  assign n47929 = n22795 & n47928 ;
  assign n47927 = n7009 & n10745 ;
  assign n47930 = n47929 ^ n47927 ^ 1'b0 ;
  assign n47931 = n7503 & ~n42954 ;
  assign n47933 = ~n6403 & n7265 ;
  assign n47932 = ~n8504 & n40971 ;
  assign n47934 = n47933 ^ n47932 ^ n1949 ;
  assign n47935 = n47934 ^ n37233 ^ n8438 ;
  assign n47936 = ( n731 & ~n21088 ) | ( n731 & n39007 ) | ( ~n21088 & n39007 ) ;
  assign n47937 = n46838 ^ n8835 ^ 1'b0 ;
  assign n47938 = n13494 ^ n8102 ^ n5548 ;
  assign n47939 = n866 & ~n47938 ;
  assign n47940 = n3664 & n47939 ;
  assign n47941 = n2659 & ~n24831 ;
  assign n47942 = n47940 & n47941 ;
  assign n47943 = n12930 & ~n20539 ;
  assign n47944 = n29020 & n47943 ;
  assign n47945 = n25548 | n34122 ;
  assign n47946 = n18183 | n47945 ;
  assign n47947 = ~n22078 & n47946 ;
  assign n47948 = n9138 & n9538 ;
  assign n47949 = n47948 ^ n17605 ^ n17215 ;
  assign n47950 = n37961 ^ n20543 ^ n9105 ;
  assign n47951 = n31580 ^ n9353 ^ n8426 ;
  assign n47952 = ( n12379 & n33899 ) | ( n12379 & ~n47951 ) | ( n33899 & ~n47951 ) ;
  assign n47953 = n18680 ^ n16298 ^ n3162 ;
  assign n47954 = ( n1875 & n45835 ) | ( n1875 & ~n47953 ) | ( n45835 & ~n47953 ) ;
  assign n47955 = n8566 | n19499 ;
  assign n47956 = n38108 & ~n47955 ;
  assign n47957 = n16365 ^ n14558 ^ n1003 ;
  assign n47958 = n23297 ^ n10162 ^ 1'b0 ;
  assign n47959 = n47957 & ~n47958 ;
  assign n47960 = n42645 ^ n9029 ^ 1'b0 ;
  assign n47961 = n42837 | n47960 ;
  assign n47963 = n14230 & ~n32833 ;
  assign n47962 = n571 & ~n23853 ;
  assign n47964 = n47963 ^ n47962 ^ n4005 ;
  assign n47967 = n5675 & ~n8443 ;
  assign n47965 = ( n803 & n32993 ) | ( n803 & n45168 ) | ( n32993 & n45168 ) ;
  assign n47966 = ( ~n2737 & n21123 ) | ( ~n2737 & n47965 ) | ( n21123 & n47965 ) ;
  assign n47968 = n47967 ^ n47966 ^ n6351 ;
  assign n47969 = n7478 & ~n35970 ;
  assign n47970 = n42250 ^ n25175 ^ n2203 ;
  assign n47971 = n47970 ^ n36303 ^ n20719 ;
  assign n47972 = n17577 ^ n13831 ^ 1'b0 ;
  assign n47973 = n9870 & n47972 ;
  assign n47974 = n40098 | n43475 ;
  assign n47975 = n47973 | n47974 ;
  assign n47976 = n34742 ^ n12425 ^ 1'b0 ;
  assign n47977 = ( ~n6478 & n21264 ) | ( ~n6478 & n39985 ) | ( n21264 & n39985 ) ;
  assign n47978 = ( ~n11251 & n38645 ) | ( ~n11251 & n47977 ) | ( n38645 & n47977 ) ;
  assign n47979 = n47978 ^ n45348 ^ n10398 ;
  assign n47980 = ( n30075 & n41810 ) | ( n30075 & n42380 ) | ( n41810 & n42380 ) ;
  assign n47981 = ~n8311 & n47980 ;
  assign n47982 = n2252 ^ n983 ^ 1'b0 ;
  assign n47983 = ( ~n20469 & n42540 ) | ( ~n20469 & n47982 ) | ( n42540 & n47982 ) ;
  assign n47984 = ( n6668 & ~n25465 ) | ( n6668 & n33888 ) | ( ~n25465 & n33888 ) ;
  assign n47985 = ( ~n7037 & n9080 ) | ( ~n7037 & n10175 ) | ( n9080 & n10175 ) ;
  assign n47986 = n47985 ^ n26242 ^ n13935 ;
  assign n47987 = ( n3303 & n21632 ) | ( n3303 & ~n47986 ) | ( n21632 & ~n47986 ) ;
  assign n47988 = ( n21074 & n37246 ) | ( n21074 & ~n47987 ) | ( n37246 & ~n47987 ) ;
  assign n47989 = ( n3914 & n9065 ) | ( n3914 & ~n14720 ) | ( n9065 & ~n14720 ) ;
  assign n47990 = n47989 ^ n1538 ^ 1'b0 ;
  assign n47991 = n47990 ^ n34179 ^ n15228 ;
  assign n47992 = ( n28476 & n45636 ) | ( n28476 & ~n47991 ) | ( n45636 & ~n47991 ) ;
  assign n47993 = n47992 ^ n34427 ^ n12551 ;
  assign n47994 = ( n39260 & n47988 ) | ( n39260 & n47993 ) | ( n47988 & n47993 ) ;
  assign n47995 = n2045 & ~n7736 ;
  assign n47996 = ~n10271 & n47995 ;
  assign n47997 = n14058 & n35867 ;
  assign n47998 = ~x67 & n47997 ;
  assign n47999 = ( n21322 & ~n26020 ) | ( n21322 & n39255 ) | ( ~n26020 & n39255 ) ;
  assign n48000 = n17999 | n47120 ;
  assign n48001 = n47999 | n48000 ;
  assign n48002 = ( ~n19535 & n23832 ) | ( ~n19535 & n29307 ) | ( n23832 & n29307 ) ;
  assign n48003 = n41179 & n48002 ;
  assign n48004 = n18802 & ~n26044 ;
  assign n48006 = ( n5603 & n7910 ) | ( n5603 & n8398 ) | ( n7910 & n8398 ) ;
  assign n48005 = ( n24245 & n39149 ) | ( n24245 & n43776 ) | ( n39149 & n43776 ) ;
  assign n48007 = n48006 ^ n48005 ^ n11596 ;
  assign n48008 = ( n15836 & n40095 ) | ( n15836 & ~n48007 ) | ( n40095 & ~n48007 ) ;
  assign n48009 = n17662 & n29123 ;
  assign n48010 = n34182 ^ n27363 ^ 1'b0 ;
  assign n48011 = ( ~n28218 & n33268 ) | ( ~n28218 & n48010 ) | ( n33268 & n48010 ) ;
  assign n48012 = n48011 ^ n23074 ^ 1'b0 ;
  assign n48013 = n3281 & ~n9993 ;
  assign n48014 = ( n13487 & n16345 ) | ( n13487 & n32938 ) | ( n16345 & n32938 ) ;
  assign n48015 = n6327 & ~n23453 ;
  assign n48016 = ~n48014 & n48015 ;
  assign n48017 = n2588 & n36298 ;
  assign n48018 = n48017 ^ n17452 ^ 1'b0 ;
  assign n48019 = ( n16536 & ~n16881 ) | ( n16536 & n31215 ) | ( ~n16881 & n31215 ) ;
  assign n48020 = ~n2014 & n19754 ;
  assign n48021 = ~n20285 & n48020 ;
  assign n48022 = ( n35237 & ~n41940 ) | ( n35237 & n48021 ) | ( ~n41940 & n48021 ) ;
  assign n48023 = ~n17199 & n25420 ;
  assign n48024 = ( n13947 & n32528 ) | ( n13947 & n34406 ) | ( n32528 & n34406 ) ;
  assign n48025 = n14226 ^ n13960 ^ n863 ;
  assign n48026 = n48025 ^ n26873 ^ n7225 ;
  assign n48027 = n48026 ^ n28321 ^ n9756 ;
  assign n48028 = n31194 ^ n3545 ^ 1'b0 ;
  assign n48029 = n31222 ^ n10032 ^ 1'b0 ;
  assign n48030 = n21495 | n48029 ;
  assign n48033 = n15663 & ~n15714 ;
  assign n48031 = n15329 ^ n10171 ^ 1'b0 ;
  assign n48032 = n38959 & ~n48031 ;
  assign n48034 = n48033 ^ n48032 ^ n10249 ;
  assign n48035 = n23399 ^ n20152 ^ n15816 ;
  assign n48036 = n1209 | n32479 ;
  assign n48037 = n25639 ^ n5203 ^ n2813 ;
  assign n48038 = ( x4 & n4750 ) | ( x4 & ~n25891 ) | ( n4750 & ~n25891 ) ;
  assign n48039 = n4884 & n48038 ;
  assign n48040 = ~n48037 & n48039 ;
  assign n48041 = ( n40113 & n48036 ) | ( n40113 & n48040 ) | ( n48036 & n48040 ) ;
  assign n48042 = n42394 ^ n32010 ^ n22398 ;
  assign n48043 = n43853 ^ n36053 ^ n6123 ;
  assign n48044 = n26766 & n48043 ;
  assign n48045 = n290 | n12209 ;
  assign n48046 = n48045 ^ n18491 ^ 1'b0 ;
  assign n48047 = n20690 ^ n9360 ^ n5293 ;
  assign n48048 = n48047 ^ n18365 ^ n6101 ;
  assign n48049 = n48048 ^ n35927 ^ n19120 ;
  assign n48050 = ~n13999 & n19399 ;
  assign n48051 = n21540 & n48050 ;
  assign n48052 = n24049 & ~n48051 ;
  assign n48053 = n48049 & n48052 ;
  assign n48054 = n18933 & ~n37745 ;
  assign n48055 = n48054 ^ n23832 ^ 1'b0 ;
  assign n48056 = ( n29365 & n46553 ) | ( n29365 & n48055 ) | ( n46553 & n48055 ) ;
  assign n48057 = n48056 ^ n37092 ^ n14377 ;
  assign n48058 = n8395 & n36392 ;
  assign n48059 = n15928 & n48058 ;
  assign n48060 = n17811 | n48059 ;
  assign n48061 = n48060 ^ n8388 ^ 1'b0 ;
  assign n48062 = ( n20486 & n27937 ) | ( n20486 & n48061 ) | ( n27937 & n48061 ) ;
  assign n48063 = n19424 ^ n8341 ^ 1'b0 ;
  assign n48064 = n45908 ^ n15123 ^ 1'b0 ;
  assign n48065 = n8913 | n13994 ;
  assign n48066 = n6149 | n48065 ;
  assign n48067 = n48066 ^ n45368 ^ n3938 ;
  assign n48068 = n42522 ^ n10504 ^ 1'b0 ;
  assign n48069 = ~n48067 & n48068 ;
  assign n48070 = n29252 ^ n26639 ^ n14468 ;
  assign n48071 = ( n6399 & ~n21729 ) | ( n6399 & n48070 ) | ( ~n21729 & n48070 ) ;
  assign n48072 = ( n6373 & n40548 ) | ( n6373 & ~n48071 ) | ( n40548 & ~n48071 ) ;
  assign n48073 = n35846 | n48072 ;
  assign n48074 = ~n23538 & n40538 ;
  assign n48075 = n48074 ^ n46559 ^ n20529 ;
  assign n48076 = n31320 ^ n21394 ^ 1'b0 ;
  assign n48077 = n28073 ^ n20150 ^ n3439 ;
  assign n48078 = ( n5907 & n7809 ) | ( n5907 & n48077 ) | ( n7809 & n48077 ) ;
  assign n48079 = ~n13368 & n30882 ;
  assign n48080 = ( ~n22133 & n48078 ) | ( ~n22133 & n48079 ) | ( n48078 & n48079 ) ;
  assign n48081 = ( ~n3144 & n13808 ) | ( ~n3144 & n33217 ) | ( n13808 & n33217 ) ;
  assign n48082 = n25883 ^ n2697 ^ 1'b0 ;
  assign n48083 = n9575 & ~n48082 ;
  assign n48084 = ~n22306 & n48083 ;
  assign n48085 = n16415 & n48084 ;
  assign n48086 = n28198 ^ n20123 ^ n5918 ;
  assign n48087 = n48086 ^ n12578 ^ 1'b0 ;
  assign n48088 = ~n5626 & n34853 ;
  assign n48089 = n48088 ^ n2265 ^ 1'b0 ;
  assign n48090 = ( n5177 & n12764 ) | ( n5177 & ~n34259 ) | ( n12764 & ~n34259 ) ;
  assign n48091 = ( n10245 & ~n36159 ) | ( n10245 & n48090 ) | ( ~n36159 & n48090 ) ;
  assign n48092 = n23700 ^ n20540 ^ 1'b0 ;
  assign n48093 = n16493 ^ n8102 ^ n1597 ;
  assign n48094 = n7855 ^ n5380 ^ n2157 ;
  assign n48095 = n15221 ^ n12554 ^ n4623 ;
  assign n48096 = ( n3397 & n48094 ) | ( n3397 & ~n48095 ) | ( n48094 & ~n48095 ) ;
  assign n48097 = n7487 | n18715 ;
  assign n48098 = n41441 | n48097 ;
  assign n48099 = n31626 ^ n2217 ^ 1'b0 ;
  assign n48100 = n48098 & ~n48099 ;
  assign n48101 = ~n4998 & n30277 ;
  assign n48102 = n48101 ^ n5973 ^ 1'b0 ;
  assign n48103 = n18707 & ~n45714 ;
  assign n48104 = n40157 ^ n23820 ^ n15013 ;
  assign n48105 = ~n39771 & n48104 ;
  assign n48106 = n48105 ^ n3085 ^ 1'b0 ;
  assign n48107 = n23088 ^ n21323 ^ n3402 ;
  assign n48108 = n24760 ^ n10043 ^ 1'b0 ;
  assign n48109 = ( n7062 & n7856 ) | ( n7062 & n48108 ) | ( n7856 & n48108 ) ;
  assign n48110 = n48109 ^ n13466 ^ n562 ;
  assign n48111 = n48110 ^ n4826 ^ 1'b0 ;
  assign n48112 = ( n36575 & n37088 ) | ( n36575 & ~n48111 ) | ( n37088 & ~n48111 ) ;
  assign n48113 = ( ~n4022 & n16803 ) | ( ~n4022 & n22730 ) | ( n16803 & n22730 ) ;
  assign n48114 = n45093 ^ n10314 ^ n300 ;
  assign n48115 = n8762 & n48114 ;
  assign n48116 = n29096 ^ n16454 ^ 1'b0 ;
  assign n48117 = n7326 & ~n29609 ;
  assign n48118 = ~n27122 & n48117 ;
  assign n48119 = n48118 ^ n7498 ^ 1'b0 ;
  assign n48120 = n20067 & ~n24257 ;
  assign n48121 = ( ~n30257 & n33013 ) | ( ~n30257 & n48120 ) | ( n33013 & n48120 ) ;
  assign n48122 = ~n9907 & n11214 ;
  assign n48123 = n2054 | n9478 ;
  assign n48124 = n48123 ^ n11461 ^ 1'b0 ;
  assign n48125 = ( n1005 & n2789 ) | ( n1005 & ~n32510 ) | ( n2789 & ~n32510 ) ;
  assign n48126 = n48125 ^ n24239 ^ n7938 ;
  assign n48127 = n14161 | n48126 ;
  assign n48128 = n48127 ^ n22693 ^ 1'b0 ;
  assign n48129 = n48128 ^ n33827 ^ 1'b0 ;
  assign n48131 = n45940 ^ n25350 ^ n12136 ;
  assign n48130 = n40665 ^ n19294 ^ n982 ;
  assign n48132 = n48131 ^ n48130 ^ n41370 ;
  assign n48133 = n22697 & n40485 ;
  assign n48135 = ( ~n4042 & n6742 ) | ( ~n4042 & n38950 ) | ( n6742 & n38950 ) ;
  assign n48136 = ~n2306 & n48135 ;
  assign n48134 = ( ~n6309 & n10007 ) | ( ~n6309 & n21810 ) | ( n10007 & n21810 ) ;
  assign n48137 = n48136 ^ n48134 ^ n1679 ;
  assign n48138 = ( n1519 & n6142 ) | ( n1519 & n8092 ) | ( n6142 & n8092 ) ;
  assign n48139 = n43839 ^ n22121 ^ 1'b0 ;
  assign n48140 = n48138 | n48139 ;
  assign n48141 = n6109 & ~n42684 ;
  assign n48142 = ~n18576 & n48141 ;
  assign n48143 = ( ~n817 & n13393 ) | ( ~n817 & n19486 ) | ( n13393 & n19486 ) ;
  assign n48144 = n16770 | n48143 ;
  assign n48145 = n6161 | n48144 ;
  assign n48146 = n8021 & ~n28847 ;
  assign n48147 = n48146 ^ n8011 ^ 1'b0 ;
  assign n48148 = n48147 ^ n38767 ^ n12320 ;
  assign n48149 = n21761 ^ n8813 ^ n7596 ;
  assign n48150 = ( n38259 & ~n40998 ) | ( n38259 & n48149 ) | ( ~n40998 & n48149 ) ;
  assign n48152 = ( n4549 & n15774 ) | ( n4549 & n22969 ) | ( n15774 & n22969 ) ;
  assign n48151 = n38666 & ~n38765 ;
  assign n48153 = n48152 ^ n48151 ^ n25080 ;
  assign n48154 = ( n10731 & n31616 ) | ( n10731 & n43645 ) | ( n31616 & n43645 ) ;
  assign n48155 = n48154 ^ n46867 ^ n16565 ;
  assign n48156 = n17386 | n18493 ;
  assign n48157 = n19453 & ~n48156 ;
  assign n48158 = n48157 ^ n15544 ^ n5434 ;
  assign n48159 = ~n3379 & n11567 ;
  assign n48160 = n48159 ^ n18919 ^ 1'b0 ;
  assign n48161 = n48160 ^ n523 ^ 1'b0 ;
  assign n48162 = n35471 ^ n9892 ^ n7104 ;
  assign n48163 = n47012 ^ n23069 ^ 1'b0 ;
  assign n48164 = ~n39311 & n48163 ;
  assign n48165 = n46878 ^ n10455 ^ 1'b0 ;
  assign n48166 = n45964 & n48165 ;
  assign n48167 = n23028 ^ n16955 ^ n12561 ;
  assign n48168 = ( n3383 & n10841 ) | ( n3383 & n48167 ) | ( n10841 & n48167 ) ;
  assign n48169 = n1026 | n48168 ;
  assign n48170 = n21426 & ~n48169 ;
  assign n48171 = n48170 ^ n15134 ^ n9737 ;
  assign n48172 = n21798 ^ n12133 ^ 1'b0 ;
  assign n48173 = ~n24520 & n48172 ;
  assign n48174 = n18751 ^ n14262 ^ n8641 ;
  assign n48175 = n18400 & n24261 ;
  assign n48176 = n48175 ^ n7259 ^ 1'b0 ;
  assign n48177 = n48176 ^ n5502 ^ 1'b0 ;
  assign n48178 = n42789 ^ n29663 ^ n9078 ;
  assign n48179 = n48178 ^ n29689 ^ n21489 ;
  assign n48180 = n19210 ^ n1813 ^ x88 ;
  assign n48181 = n48180 ^ n11684 ^ 1'b0 ;
  assign n48182 = n45323 & ~n48181 ;
  assign n48183 = ( n4623 & ~n18288 ) | ( n4623 & n26976 ) | ( ~n18288 & n26976 ) ;
  assign n48184 = n15975 & ~n48183 ;
  assign n48191 = n22494 ^ n22484 ^ n7348 ;
  assign n48189 = n47441 ^ n23667 ^ 1'b0 ;
  assign n48190 = n6780 | n48189 ;
  assign n48185 = n34205 | n39515 ;
  assign n48186 = n11631 & ~n48185 ;
  assign n48187 = n29417 ^ n16300 ^ n6638 ;
  assign n48188 = ( n18464 & ~n48186 ) | ( n18464 & n48187 ) | ( ~n48186 & n48187 ) ;
  assign n48192 = n48191 ^ n48190 ^ n48188 ;
  assign n48193 = n6936 & ~n11942 ;
  assign n48194 = n10151 | n25629 ;
  assign n48195 = n48194 ^ n3126 ^ 1'b0 ;
  assign n48196 = ( ~n310 & n12726 ) | ( ~n310 & n48195 ) | ( n12726 & n48195 ) ;
  assign n48197 = n15382 ^ n12249 ^ 1'b0 ;
  assign n48198 = n1101 & n34907 ;
  assign n48199 = n48198 ^ n12465 ^ 1'b0 ;
  assign n48200 = ( n33563 & n48197 ) | ( n33563 & ~n48199 ) | ( n48197 & ~n48199 ) ;
  assign n48201 = n22629 & n43853 ;
  assign n48204 = n18416 ^ n10500 ^ 1'b0 ;
  assign n48205 = n26104 & ~n48204 ;
  assign n48203 = n9546 ^ n3305 ^ 1'b0 ;
  assign n48206 = n48205 ^ n48203 ^ n30413 ;
  assign n48202 = n41126 ^ n26959 ^ n3838 ;
  assign n48207 = n48206 ^ n48202 ^ n12547 ;
  assign n48208 = n25195 | n48207 ;
  assign n48209 = n48201 & ~n48208 ;
  assign n48210 = n46721 ^ n20883 ^ n12852 ;
  assign n48211 = n35674 & ~n48210 ;
  assign n48212 = ( n31811 & ~n41164 ) | ( n31811 & n44831 ) | ( ~n41164 & n44831 ) ;
  assign n48213 = n29247 ^ n16018 ^ n4676 ;
  assign n48214 = n42379 ^ n3947 ^ 1'b0 ;
  assign n48215 = n24149 ^ n11285 ^ 1'b0 ;
  assign n48216 = ~n6430 & n26296 ;
  assign n48217 = n48216 ^ n11006 ^ 1'b0 ;
  assign n48218 = ( n21319 & n48215 ) | ( n21319 & ~n48217 ) | ( n48215 & ~n48217 ) ;
  assign n48219 = n25558 ^ n2870 ^ 1'b0 ;
  assign n48220 = n7886 | n8819 ;
  assign n48221 = n48220 ^ n25375 ^ 1'b0 ;
  assign n48222 = ( ~n4353 & n12932 ) | ( ~n4353 & n48221 ) | ( n12932 & n48221 ) ;
  assign n48223 = n2659 & n17917 ;
  assign n48224 = n48222 & n48223 ;
  assign n48225 = ( n14933 & ~n48219 ) | ( n14933 & n48224 ) | ( ~n48219 & n48224 ) ;
  assign n48226 = n8375 & n43051 ;
  assign n48227 = ( n18906 & ~n23982 ) | ( n18906 & n44324 ) | ( ~n23982 & n44324 ) ;
  assign n48228 = n20952 ^ n15751 ^ n1356 ;
  assign n48229 = n42788 | n48228 ;
  assign n48230 = n48227 & ~n48229 ;
  assign n48231 = n15684 ^ n9148 ^ n7601 ;
  assign n48232 = n2295 | n19197 ;
  assign n48233 = n48231 & ~n48232 ;
  assign n48234 = ~n7679 & n23607 ;
  assign n48235 = ~n44880 & n48234 ;
  assign n48236 = n24175 & n40902 ;
  assign n48237 = ~n9870 & n48236 ;
  assign n48238 = n48237 ^ n14046 ^ n11126 ;
  assign n48239 = n10598 & n48238 ;
  assign n48240 = n41527 ^ n38648 ^ n2203 ;
  assign n48244 = n19064 ^ n12786 ^ n7169 ;
  assign n48241 = n28121 ^ n1261 ^ 1'b0 ;
  assign n48242 = n48241 ^ n3327 ^ 1'b0 ;
  assign n48243 = n14834 & n48242 ;
  assign n48245 = n48244 ^ n48243 ^ n24448 ;
  assign n48246 = n26518 ^ n18565 ^ n8814 ;
  assign n48247 = n26651 & ~n48246 ;
  assign n48248 = n6024 | n24717 ;
  assign n48249 = ( n13277 & ~n21731 ) | ( n13277 & n33263 ) | ( ~n21731 & n33263 ) ;
  assign n48250 = ~n1716 & n20956 ;
  assign n48251 = ~n28188 & n32564 ;
  assign n48252 = n48251 ^ n1955 ^ 1'b0 ;
  assign n48253 = n2385 & ~n15157 ;
  assign n48254 = n48253 ^ n46070 ^ 1'b0 ;
  assign n48255 = n7293 & ~n14513 ;
  assign n48256 = n47565 ^ n39131 ^ n22030 ;
  assign n48257 = n7181 | n14581 ;
  assign n48258 = n11757 | n48257 ;
  assign n48259 = n2657 & ~n48258 ;
  assign n48260 = ( ~n1464 & n7860 ) | ( ~n1464 & n48259 ) | ( n7860 & n48259 ) ;
  assign n48261 = n48260 ^ n45116 ^ n9107 ;
  assign n48262 = n35057 ^ n28201 ^ n15900 ;
  assign n48263 = n28437 ^ n13605 ^ 1'b0 ;
  assign n48264 = n36577 ^ n4229 ^ 1'b0 ;
  assign n48265 = n48263 & n48264 ;
  assign n48266 = x38 & ~n1833 ;
  assign n48267 = n30450 & n48266 ;
  assign n48268 = ( n24380 & ~n32659 ) | ( n24380 & n36787 ) | ( ~n32659 & n36787 ) ;
  assign n48269 = n4225 & n7980 ;
  assign n48270 = n18554 & n48269 ;
  assign n48271 = ( ~n12454 & n13397 ) | ( ~n12454 & n21675 ) | ( n13397 & n21675 ) ;
  assign n48272 = n48271 ^ n22141 ^ n1681 ;
  assign n48273 = n48272 ^ n22372 ^ n9929 ;
  assign n48274 = ( n11414 & ~n13187 ) | ( n11414 & n17120 ) | ( ~n13187 & n17120 ) ;
  assign n48275 = ~n4406 & n48274 ;
  assign n48276 = ~n48273 & n48275 ;
  assign n48277 = ( n11207 & ~n48270 ) | ( n11207 & n48276 ) | ( ~n48270 & n48276 ) ;
  assign n48278 = n48277 ^ n18403 ^ n10213 ;
  assign n48279 = n35960 ^ n29377 ^ n13340 ;
  assign n48284 = n13268 ^ n3452 ^ n1498 ;
  assign n48280 = ~n18898 & n25864 ;
  assign n48281 = n48280 ^ n7316 ^ 1'b0 ;
  assign n48282 = ( n16612 & n21982 ) | ( n16612 & n48281 ) | ( n21982 & n48281 ) ;
  assign n48283 = n48282 ^ n36550 ^ n30669 ;
  assign n48285 = n48284 ^ n48283 ^ n31824 ;
  assign n48286 = ( ~n21596 & n33870 ) | ( ~n21596 & n34645 ) | ( n33870 & n34645 ) ;
  assign n48287 = ( ~n5248 & n12470 ) | ( ~n5248 & n15647 ) | ( n12470 & n15647 ) ;
  assign n48288 = ( ~n23722 & n43038 ) | ( ~n23722 & n48287 ) | ( n43038 & n48287 ) ;
  assign n48289 = ( n8859 & ~n20958 ) | ( n8859 & n46676 ) | ( ~n20958 & n46676 ) ;
  assign n48290 = n11905 ^ n9805 ^ 1'b0 ;
  assign n48291 = n814 & ~n48290 ;
  assign n48292 = ( n39509 & n48289 ) | ( n39509 & ~n48291 ) | ( n48289 & ~n48291 ) ;
  assign n48293 = n1752 & n48292 ;
  assign n48294 = n13501 & n48293 ;
  assign n48295 = ( n3879 & n14789 ) | ( n3879 & ~n41349 ) | ( n14789 & ~n41349 ) ;
  assign n48296 = ~n29359 & n48295 ;
  assign n48297 = n48296 ^ n24727 ^ 1'b0 ;
  assign n48298 = n2859 | n48297 ;
  assign n48299 = n29635 & ~n48298 ;
  assign n48300 = n22275 & ~n24462 ;
  assign n48301 = ~n44846 & n48300 ;
  assign n48302 = n1077 & n13821 ;
  assign n48303 = ( n2257 & n6338 ) | ( n2257 & n14874 ) | ( n6338 & n14874 ) ;
  assign n48304 = n23860 ^ n22372 ^ 1'b0 ;
  assign n48305 = ~n13969 & n45269 ;
  assign n48306 = n25101 & n48305 ;
  assign n48307 = n48306 ^ n29049 ^ n17913 ;
  assign n48308 = ( n7447 & ~n23942 ) | ( n7447 & n48307 ) | ( ~n23942 & n48307 ) ;
  assign n48309 = ( ~n32308 & n36540 ) | ( ~n32308 & n40058 ) | ( n36540 & n40058 ) ;
  assign n48311 = ( n14311 & n16071 ) | ( n14311 & n43458 ) | ( n16071 & n43458 ) ;
  assign n48310 = n23718 & ~n24111 ;
  assign n48312 = n48311 ^ n48310 ^ 1'b0 ;
  assign n48313 = ( n2348 & n35930 ) | ( n2348 & ~n48312 ) | ( n35930 & ~n48312 ) ;
  assign n48314 = n18461 ^ n11089 ^ 1'b0 ;
  assign n48315 = n48313 | n48314 ;
  assign n48316 = n2717 & n10062 ;
  assign n48317 = n42111 ^ n41094 ^ n28684 ;
  assign n48318 = n48317 ^ n11242 ^ n7277 ;
  assign n48319 = n20744 ^ n647 ^ 1'b0 ;
  assign n48320 = n18258 | n48319 ;
  assign n48321 = n48320 ^ n17110 ^ n1924 ;
  assign n48322 = n15552 ^ n12843 ^ 1'b0 ;
  assign n48323 = ( n10644 & n27404 ) | ( n10644 & ~n29687 ) | ( n27404 & ~n29687 ) ;
  assign n48324 = n48322 & n48323 ;
  assign n48325 = n32515 ^ n3385 ^ n1196 ;
  assign n48326 = ( n15227 & n25993 ) | ( n15227 & ~n36459 ) | ( n25993 & ~n36459 ) ;
  assign n48327 = n28331 & ~n30804 ;
  assign n48328 = n30922 ^ n17849 ^ n1870 ;
  assign n48329 = ( n11192 & ~n48327 ) | ( n11192 & n48328 ) | ( ~n48327 & n48328 ) ;
  assign n48330 = n9480 ^ n1096 ^ 1'b0 ;
  assign n48331 = n4572 & ~n48330 ;
  assign n48332 = n3654 | n6279 ;
  assign n48333 = n48331 | n48332 ;
  assign n48334 = n48333 ^ n9366 ^ 1'b0 ;
  assign n48335 = ( n2736 & n6605 ) | ( n2736 & n39570 ) | ( n6605 & n39570 ) ;
  assign n48336 = ~n7171 & n27275 ;
  assign n48337 = n48336 ^ n39222 ^ 1'b0 ;
  assign n48338 = ~n48335 & n48337 ;
  assign n48339 = ( n4138 & n10047 ) | ( n4138 & n29354 ) | ( n10047 & n29354 ) ;
  assign n48340 = n5071 & n39651 ;
  assign n48341 = n48340 ^ n8954 ^ 1'b0 ;
  assign n48342 = n34144 & ~n48341 ;
  assign n48343 = ~n3670 & n16018 ;
  assign n48344 = n48343 ^ n20058 ^ n12339 ;
  assign n48345 = n17549 ^ n9828 ^ n9807 ;
  assign n48346 = ( n4192 & n36155 ) | ( n4192 & ~n48345 ) | ( n36155 & ~n48345 ) ;
  assign n48347 = n44939 ^ n44812 ^ n44087 ;
  assign n48348 = n48347 ^ n40213 ^ 1'b0 ;
  assign n48349 = n24559 & ~n48348 ;
  assign n48350 = n11448 ^ n3940 ^ 1'b0 ;
  assign n48351 = ~n19474 & n48350 ;
  assign n48352 = n9362 & ~n26928 ;
  assign n48353 = n5863 & n48352 ;
  assign n48354 = n48353 ^ n23759 ^ 1'b0 ;
  assign n48355 = n21404 & ~n27778 ;
  assign n48356 = n48355 ^ n44852 ^ 1'b0 ;
  assign n48357 = n27959 ^ n22290 ^ n16931 ;
  assign n48358 = n12328 & ~n35395 ;
  assign n48359 = n48358 ^ n18958 ^ 1'b0 ;
  assign n48360 = ~n8030 & n48359 ;
  assign n48361 = n22175 ^ n12946 ^ n12295 ;
  assign n48362 = n48361 ^ n41446 ^ n20708 ;
  assign n48363 = ( n18618 & ~n30811 ) | ( n18618 & n31553 ) | ( ~n30811 & n31553 ) ;
  assign n48365 = ( n988 & n12750 ) | ( n988 & ~n24241 ) | ( n12750 & ~n24241 ) ;
  assign n48364 = ( n3808 & n27956 ) | ( n3808 & n45868 ) | ( n27956 & n45868 ) ;
  assign n48366 = n48365 ^ n48364 ^ n12739 ;
  assign n48367 = n48366 ^ n34452 ^ n16955 ;
  assign n48368 = n43306 ^ n16558 ^ 1'b0 ;
  assign n48369 = ~n12257 & n35839 ;
  assign n48370 = n48369 ^ n33382 ^ 1'b0 ;
  assign n48371 = ~n25282 & n37401 ;
  assign n48372 = ( n27341 & n32342 ) | ( n27341 & n48371 ) | ( n32342 & n48371 ) ;
  assign n48373 = ( n655 & n12625 ) | ( n655 & n27033 ) | ( n12625 & n27033 ) ;
  assign n48374 = ( n2626 & ~n8410 ) | ( n2626 & n13619 ) | ( ~n8410 & n13619 ) ;
  assign n48375 = n48374 ^ n22571 ^ 1'b0 ;
  assign n48376 = n3689 & ~n27480 ;
  assign n48377 = n8315 ^ n2926 ^ 1'b0 ;
  assign n48378 = n37371 ^ n5970 ^ n1449 ;
  assign n48379 = n15703 & ~n46999 ;
  assign n48380 = n30788 & ~n48379 ;
  assign n48381 = n48378 & n48380 ;
  assign n48382 = ( ~x81 & n48377 ) | ( ~x81 & n48381 ) | ( n48377 & n48381 ) ;
  assign n48383 = ( n8301 & n17838 ) | ( n8301 & ~n22879 ) | ( n17838 & ~n22879 ) ;
  assign n48391 = ( n502 & n2927 ) | ( n502 & ~n5261 ) | ( n2927 & ~n5261 ) ;
  assign n48392 = n48391 ^ n13793 ^ n8873 ;
  assign n48389 = n3644 & n17419 ;
  assign n48390 = n48389 ^ n14336 ^ 1'b0 ;
  assign n48393 = n48392 ^ n48390 ^ n7702 ;
  assign n48388 = n36722 ^ n24109 ^ n3894 ;
  assign n48384 = ( n1080 & n25860 ) | ( n1080 & n26100 ) | ( n25860 & n26100 ) ;
  assign n48385 = n7859 | n19441 ;
  assign n48386 = n48385 ^ n29494 ^ 1'b0 ;
  assign n48387 = ( n36692 & n48384 ) | ( n36692 & ~n48386 ) | ( n48384 & ~n48386 ) ;
  assign n48394 = n48393 ^ n48388 ^ n48387 ;
  assign n48395 = ~n1564 & n7151 ;
  assign n48396 = n48395 ^ n30547 ^ 1'b0 ;
  assign n48397 = n28829 ^ n8138 ^ 1'b0 ;
  assign n48398 = ~n31961 & n48397 ;
  assign n48399 = n47794 ^ n431 ^ 1'b0 ;
  assign n48400 = n23571 & n30116 ;
  assign n48401 = n39567 ^ n17743 ^ n4523 ;
  assign n48402 = ( n1225 & n9107 ) | ( n1225 & ~n40854 ) | ( n9107 & ~n40854 ) ;
  assign n48403 = n7640 ^ n6788 ^ 1'b0 ;
  assign n48404 = n48403 ^ n3990 ^ n2818 ;
  assign n48405 = n48404 ^ n36068 ^ n31008 ;
  assign n48406 = n13082 | n16940 ;
  assign n48407 = n28594 & ~n46675 ;
  assign n48408 = ( n5829 & n8958 ) | ( n5829 & ~n31651 ) | ( n8958 & ~n31651 ) ;
  assign n48409 = ( n22802 & n32642 ) | ( n22802 & ~n48408 ) | ( n32642 & ~n48408 ) ;
  assign n48410 = n11400 & n12107 ;
  assign n48411 = ~n12275 & n48410 ;
  assign n48412 = n9516 & ~n45188 ;
  assign n48413 = n22012 ^ n21707 ^ n738 ;
  assign n48414 = n48413 ^ n27933 ^ n20106 ;
  assign n48415 = ( n32131 & n39498 ) | ( n32131 & n43178 ) | ( n39498 & n43178 ) ;
  assign n48418 = ( n12509 & n13436 ) | ( n12509 & ~n37911 ) | ( n13436 & ~n37911 ) ;
  assign n48419 = n48418 ^ n7766 ^ 1'b0 ;
  assign n48416 = n25601 | n28026 ;
  assign n48417 = n10277 & n48416 ;
  assign n48420 = n48419 ^ n48417 ^ 1'b0 ;
  assign n48421 = n7805 | n27746 ;
  assign n48422 = n48421 ^ n5992 ^ 1'b0 ;
  assign n48424 = n4410 | n13146 ;
  assign n48423 = ~n14821 & n26902 ;
  assign n48425 = n48424 ^ n48423 ^ n22356 ;
  assign n48426 = n29648 | n48425 ;
  assign n48427 = n48422 & ~n48426 ;
  assign n48428 = n39381 ^ n6144 ^ 1'b0 ;
  assign n48429 = n39731 ^ n13759 ^ n13634 ;
  assign n48430 = ( x251 & n7363 ) | ( x251 & ~n19110 ) | ( n7363 & ~n19110 ) ;
  assign n48431 = ( n21681 & n22937 ) | ( n21681 & n48430 ) | ( n22937 & n48430 ) ;
  assign n48432 = n42102 ^ n38742 ^ n37486 ;
  assign n48433 = ( n7558 & ~n40406 ) | ( n7558 & n48374 ) | ( ~n40406 & n48374 ) ;
  assign n48434 = n35866 ^ n27374 ^ n11300 ;
  assign n48435 = n12539 | n21707 ;
  assign n48436 = n10488 & ~n48435 ;
  assign n48437 = n47970 & n48436 ;
  assign n48438 = n30627 ^ n15997 ^ n10863 ;
  assign n48439 = n30887 ^ n8951 ^ n7249 ;
  assign n48440 = n41170 & n48439 ;
  assign n48444 = n5449 | n26817 ;
  assign n48445 = n13802 | n48444 ;
  assign n48446 = n48445 ^ n18056 ^ n8950 ;
  assign n48441 = ~n6676 & n31254 ;
  assign n48442 = n47973 ^ n9205 ^ 1'b0 ;
  assign n48443 = n48441 & n48442 ;
  assign n48447 = n48446 ^ n48443 ^ n14438 ;
  assign n48449 = n8776 ^ n1567 ^ 1'b0 ;
  assign n48450 = ~n10228 & n48449 ;
  assign n48448 = n30770 ^ n20596 ^ n6450 ;
  assign n48451 = n48450 ^ n48448 ^ n31382 ;
  assign n48452 = ( n5918 & ~n21318 ) | ( n5918 & n48451 ) | ( ~n21318 & n48451 ) ;
  assign n48453 = n33210 ^ n8193 ^ n1099 ;
  assign n48454 = n48453 ^ n9758 ^ n8727 ;
  assign n48455 = ( n7223 & n11367 ) | ( n7223 & ~n26912 ) | ( n11367 & ~n26912 ) ;
  assign n48456 = ( ~n3274 & n23734 ) | ( ~n3274 & n24315 ) | ( n23734 & n24315 ) ;
  assign n48457 = ( n5234 & n48455 ) | ( n5234 & ~n48456 ) | ( n48455 & ~n48456 ) ;
  assign n48458 = n34738 ^ n19479 ^ n14657 ;
  assign n48459 = n48458 ^ n6189 ^ 1'b0 ;
  assign n48460 = ~n23715 & n48459 ;
  assign n48461 = ( n19372 & n39212 ) | ( n19372 & ~n46469 ) | ( n39212 & ~n46469 ) ;
  assign n48465 = n43563 ^ n5594 ^ 1'b0 ;
  assign n48466 = n48465 ^ n45378 ^ n22585 ;
  assign n48462 = n26891 ^ n4703 ^ 1'b0 ;
  assign n48463 = ( ~x30 & n30469 ) | ( ~x30 & n34319 ) | ( n30469 & n34319 ) ;
  assign n48464 = ( n24075 & n48462 ) | ( n24075 & n48463 ) | ( n48462 & n48463 ) ;
  assign n48467 = n48466 ^ n48464 ^ n27759 ;
  assign n48468 = ( ~n10137 & n12047 ) | ( ~n10137 & n31260 ) | ( n12047 & n31260 ) ;
  assign n48469 = ( ~n20485 & n33955 ) | ( ~n20485 & n35289 ) | ( n33955 & n35289 ) ;
  assign n48470 = n14823 | n47205 ;
  assign n48471 = n23798 | n48470 ;
  assign n48472 = n24327 ^ n20513 ^ 1'b0 ;
  assign n48473 = ( n4482 & n34037 ) | ( n4482 & n48472 ) | ( n34037 & n48472 ) ;
  assign n48474 = ( ~n19575 & n38383 ) | ( ~n19575 & n41555 ) | ( n38383 & n41555 ) ;
  assign n48475 = n3520 & ~n14805 ;
  assign n48476 = n48475 ^ n6677 ^ 1'b0 ;
  assign n48477 = n414 & ~n25596 ;
  assign n48478 = n48477 ^ n10549 ^ 1'b0 ;
  assign n48479 = ( n3390 & ~n8864 ) | ( n3390 & n48478 ) | ( ~n8864 & n48478 ) ;
  assign n48480 = n26195 ^ n18362 ^ n13712 ;
  assign n48481 = n48480 ^ n5628 ^ 1'b0 ;
  assign n48482 = n1257 & ~n48481 ;
  assign n48483 = ( n431 & ~n7766 ) | ( n431 & n26778 ) | ( ~n7766 & n26778 ) ;
  assign n48484 = n28073 & n43543 ;
  assign n48485 = ( n21115 & n23886 ) | ( n21115 & n48484 ) | ( n23886 & n48484 ) ;
  assign n48486 = ( n10360 & n10446 ) | ( n10360 & ~n13277 ) | ( n10446 & ~n13277 ) ;
  assign n48487 = ( ~n30815 & n37924 ) | ( ~n30815 & n48486 ) | ( n37924 & n48486 ) ;
  assign n48488 = n28717 & ~n47424 ;
  assign n48489 = n48488 ^ n18092 ^ 1'b0 ;
  assign n48490 = n48489 ^ n3663 ^ n2800 ;
  assign n48491 = n37797 ^ n887 ^ 1'b0 ;
  assign n48492 = n41270 & n48491 ;
  assign n48493 = ( n8289 & ~n30437 ) | ( n8289 & n42157 ) | ( ~n30437 & n42157 ) ;
  assign n48494 = n24750 ^ n18219 ^ 1'b0 ;
  assign n48495 = ~n37364 & n48494 ;
  assign n48496 = ( n4154 & n48493 ) | ( n4154 & ~n48495 ) | ( n48493 & ~n48495 ) ;
  assign n48497 = n20392 ^ n7525 ^ n1246 ;
  assign n48498 = n48497 ^ n38298 ^ n7577 ;
  assign n48499 = n7870 & n29867 ;
  assign n48500 = n40933 & n48499 ;
  assign n48501 = ( n343 & n29946 ) | ( n343 & ~n48500 ) | ( n29946 & ~n48500 ) ;
  assign n48502 = n48501 ^ n4397 ^ n2797 ;
  assign n48503 = n34175 ^ n30320 ^ n26651 ;
  assign n48504 = ( n31872 & n33119 ) | ( n31872 & ~n41717 ) | ( n33119 & ~n41717 ) ;
  assign n48505 = n48504 ^ n5863 ^ n5405 ;
  assign n48506 = n16791 ^ n5635 ^ n2621 ;
  assign n48507 = n37631 ^ n22248 ^ 1'b0 ;
  assign n48508 = n40351 | n48507 ;
  assign n48509 = n42103 ^ n5524 ^ n2069 ;
  assign n48510 = n48509 ^ n30171 ^ 1'b0 ;
  assign n48511 = x79 & n48510 ;
  assign n48512 = ( n700 & n9426 ) | ( n700 & n33017 ) | ( n9426 & n33017 ) ;
  assign n48513 = n17552 ^ n16511 ^ 1'b0 ;
  assign n48514 = ( n9400 & ~n27810 ) | ( n9400 & n48513 ) | ( ~n27810 & n48513 ) ;
  assign n48515 = n6148 ^ n3089 ^ n1463 ;
  assign n48516 = n48515 ^ n30565 ^ n2001 ;
  assign n48517 = n1142 & ~n7805 ;
  assign n48518 = ~n42096 & n48517 ;
  assign n48519 = n48518 ^ n18409 ^ 1'b0 ;
  assign n48520 = ( n2240 & n22501 ) | ( n2240 & n26629 ) | ( n22501 & n26629 ) ;
  assign n48521 = ( n749 & n6299 ) | ( n749 & n15933 ) | ( n6299 & n15933 ) ;
  assign n48522 = n48521 ^ n16897 ^ n5697 ;
  assign n48523 = ( n17732 & n35980 ) | ( n17732 & n48522 ) | ( n35980 & n48522 ) ;
  assign n48526 = ( n2408 & n16359 ) | ( n2408 & n18321 ) | ( n16359 & n18321 ) ;
  assign n48524 = ~n9918 & n10019 ;
  assign n48525 = ~n5409 & n48524 ;
  assign n48527 = n48526 ^ n48525 ^ n872 ;
  assign n48528 = n28609 & n38362 ;
  assign n48529 = n48528 ^ n3217 ^ 1'b0 ;
  assign n48530 = ( n8338 & ~n39548 ) | ( n8338 & n43820 ) | ( ~n39548 & n43820 ) ;
  assign n48531 = n17533 | n48530 ;
  assign n48532 = ~n4046 & n8652 ;
  assign n48533 = n48532 ^ n35582 ^ 1'b0 ;
  assign n48534 = n48533 ^ n33297 ^ n11357 ;
  assign n48535 = n38130 ^ n1942 ^ n1689 ;
  assign n48536 = ( n6355 & ~n11195 ) | ( n6355 & n48535 ) | ( ~n11195 & n48535 ) ;
  assign n48537 = n37614 ^ n28715 ^ n20750 ;
  assign n48538 = n27709 ^ n9200 ^ n3180 ;
  assign n48539 = n24026 ^ n19203 ^ n3044 ;
  assign n48540 = ( n33810 & ~n37096 ) | ( n33810 & n44220 ) | ( ~n37096 & n44220 ) ;
  assign n48541 = n2872 | n37994 ;
  assign n48542 = n44690 ^ n17026 ^ 1'b0 ;
  assign n48543 = ~n47726 & n48542 ;
  assign n48546 = n5581 ^ n2955 ^ 1'b0 ;
  assign n48544 = n3679 & n34047 ;
  assign n48545 = ~n1752 & n48544 ;
  assign n48547 = n48546 ^ n48545 ^ 1'b0 ;
  assign n48548 = n48547 ^ n30859 ^ n19893 ;
  assign n48549 = n15939 & n48548 ;
  assign n48550 = n31399 & n48549 ;
  assign n48554 = ( n1805 & ~n17833 ) | ( n1805 & n20998 ) | ( ~n17833 & n20998 ) ;
  assign n48552 = ( ~n14373 & n16303 ) | ( ~n14373 & n38321 ) | ( n16303 & n38321 ) ;
  assign n48551 = n41935 ^ n35510 ^ n702 ;
  assign n48553 = n48552 ^ n48551 ^ n38145 ;
  assign n48555 = n48554 ^ n48553 ^ n3766 ;
  assign n48556 = n22381 ^ n11976 ^ 1'b0 ;
  assign n48557 = n38227 | n48556 ;
  assign n48558 = n48557 ^ n24691 ^ 1'b0 ;
  assign n48559 = n23772 ^ n18601 ^ n5307 ;
  assign n48560 = n28538 & ~n48559 ;
  assign n48561 = n47825 ^ n33632 ^ n17608 ;
  assign n48562 = n4438 | n37727 ;
  assign n48563 = ~n11641 & n48562 ;
  assign n48564 = n48563 ^ n25901 ^ 1'b0 ;
  assign n48565 = ( n15687 & n34093 ) | ( n15687 & ~n48564 ) | ( n34093 & ~n48564 ) ;
  assign n48566 = n28322 ^ n19090 ^ n18439 ;
  assign n48567 = ( n12432 & n43923 ) | ( n12432 & n48566 ) | ( n43923 & n48566 ) ;
  assign n48568 = n22877 ^ n16712 ^ n7023 ;
  assign n48569 = ( ~n17762 & n27297 ) | ( ~n17762 & n29362 ) | ( n27297 & n29362 ) ;
  assign n48570 = ( n9247 & n27237 ) | ( n9247 & ~n34821 ) | ( n27237 & ~n34821 ) ;
  assign n48571 = n48570 ^ n24840 ^ 1'b0 ;
  assign n48572 = n8241 | n38871 ;
  assign n48573 = n48572 ^ n16007 ^ 1'b0 ;
  assign n48574 = n11430 & n48573 ;
  assign n48575 = n10216 ^ n1280 ^ 1'b0 ;
  assign n48576 = n26179 & ~n48575 ;
  assign n48577 = n23613 & n48576 ;
  assign n48578 = n41144 & ~n48577 ;
  assign n48579 = ~n4844 & n48578 ;
  assign n48580 = n8451 ^ n6139 ^ n5211 ;
  assign n48581 = ( n24500 & ~n42900 ) | ( n24500 & n43027 ) | ( ~n42900 & n43027 ) ;
  assign n48582 = ( n3979 & n8279 ) | ( n3979 & ~n35206 ) | ( n8279 & ~n35206 ) ;
  assign n48583 = ( ~n26121 & n35633 ) | ( ~n26121 & n37088 ) | ( n35633 & n37088 ) ;
  assign n48584 = n30003 ^ n869 ^ 1'b0 ;
  assign n48585 = n14034 & n48584 ;
  assign n48586 = n30711 | n43856 ;
  assign n48587 = n17784 ^ n15651 ^ n2296 ;
  assign n48588 = n48587 ^ n30232 ^ n17727 ;
  assign n48589 = ( n4978 & n37802 ) | ( n4978 & n48078 ) | ( n37802 & n48078 ) ;
  assign n48590 = n48589 ^ n26649 ^ n17418 ;
  assign n48591 = ( n20858 & n23451 ) | ( n20858 & ~n29719 ) | ( n23451 & ~n29719 ) ;
  assign n48592 = n48591 ^ n9136 ^ 1'b0 ;
  assign n48593 = ~n13057 & n48592 ;
  assign n48594 = ~n31359 & n48593 ;
  assign n48595 = n17583 ^ n9851 ^ n2889 ;
  assign n48596 = n8027 | n20564 ;
  assign n48597 = n48596 ^ n16606 ^ n12270 ;
  assign n48598 = n13301 ^ n5038 ^ 1'b0 ;
  assign n48599 = n9632 & ~n48598 ;
  assign n48600 = ( n12694 & n30274 ) | ( n12694 & n46260 ) | ( n30274 & n46260 ) ;
  assign n48601 = n33685 | n48600 ;
  assign n48602 = n48601 ^ n15602 ^ 1'b0 ;
  assign n48603 = ~n16817 & n34317 ;
  assign n48604 = ( n39155 & n45904 ) | ( n39155 & ~n48603 ) | ( n45904 & ~n48603 ) ;
  assign n48605 = n19382 ^ n17485 ^ n8688 ;
  assign n48606 = n37727 ^ n23415 ^ n2751 ;
  assign n48607 = n48606 ^ n33328 ^ n5448 ;
  assign n48608 = n37480 ^ n15696 ^ n14158 ;
  assign n48609 = ( n6306 & ~n9804 ) | ( n6306 & n26568 ) | ( ~n9804 & n26568 ) ;
  assign n48610 = n3592 | n48609 ;
  assign n48611 = ~n21177 & n48610 ;
  assign n48612 = ( n3074 & ~n12847 ) | ( n3074 & n23363 ) | ( ~n12847 & n23363 ) ;
  assign n48613 = n5657 | n48612 ;
  assign n48614 = n48613 ^ n10691 ^ 1'b0 ;
  assign n48615 = n19321 & ~n26870 ;
  assign n48616 = n48615 ^ n2408 ^ 1'b0 ;
  assign n48617 = n9033 ^ n7897 ^ n5911 ;
  assign n48618 = n48617 ^ n18906 ^ n8726 ;
  assign n48619 = n27043 ^ n20160 ^ n15997 ;
  assign n48620 = n41010 ^ n33856 ^ n10100 ;
  assign n48621 = ( n48618 & ~n48619 ) | ( n48618 & n48620 ) | ( ~n48619 & n48620 ) ;
  assign n48622 = n11048 ^ n6424 ^ 1'b0 ;
  assign n48623 = ( n15099 & n41941 ) | ( n15099 & n48622 ) | ( n41941 & n48622 ) ;
  assign n48624 = n7655 | n22597 ;
  assign n48625 = ~n21587 & n48624 ;
  assign n48626 = ( n5237 & ~n7924 ) | ( n5237 & n37817 ) | ( ~n7924 & n37817 ) ;
  assign n48627 = ~n3845 & n17669 ;
  assign n48628 = n48627 ^ n9416 ^ n3776 ;
  assign n48629 = n5043 & n22676 ;
  assign n48630 = n48629 ^ n25929 ^ 1'b0 ;
  assign n48631 = ( n3461 & n31363 ) | ( n3461 & ~n48630 ) | ( n31363 & ~n48630 ) ;
  assign n48635 = ( n744 & n26566 ) | ( n744 & ~n37461 ) | ( n26566 & ~n37461 ) ;
  assign n48632 = n22930 ^ n5018 ^ 1'b0 ;
  assign n48633 = n31042 & ~n48632 ;
  assign n48634 = ~n11912 & n48633 ;
  assign n48636 = n48635 ^ n48634 ^ 1'b0 ;
  assign n48637 = x17 & ~n9670 ;
  assign n48638 = ( n18691 & n48313 ) | ( n18691 & n48637 ) | ( n48313 & n48637 ) ;
  assign n48639 = n2070 & ~n20899 ;
  assign n48640 = ( n5553 & ~n27832 ) | ( n5553 & n48639 ) | ( ~n27832 & n48639 ) ;
  assign n48641 = n48640 ^ n47353 ^ n20131 ;
  assign n48642 = n21062 ^ n9608 ^ n302 ;
  assign n48643 = n35073 ^ n8462 ^ 1'b0 ;
  assign n48644 = ~n48642 & n48643 ;
  assign n48645 = ~n2143 & n40687 ;
  assign n48646 = n48645 ^ n2976 ^ 1'b0 ;
  assign n48647 = ( ~n1997 & n24322 ) | ( ~n1997 & n48646 ) | ( n24322 & n48646 ) ;
  assign n48648 = ( ~n14308 & n48644 ) | ( ~n14308 & n48647 ) | ( n48644 & n48647 ) ;
  assign n48649 = n31237 ^ n7325 ^ 1'b0 ;
  assign n48650 = n48649 ^ n14267 ^ 1'b0 ;
  assign n48651 = ( n2591 & n37323 ) | ( n2591 & ~n48650 ) | ( n37323 & ~n48650 ) ;
  assign n48652 = n48651 ^ n15466 ^ 1'b0 ;
  assign n48653 = ~n38211 & n48652 ;
  assign n48654 = n24565 ^ n16597 ^ n7891 ;
  assign n48655 = n3254 & n4182 ;
  assign n48659 = n5598 & ~n17897 ;
  assign n48656 = n8503 ^ n7452 ^ x57 ;
  assign n48657 = n48656 ^ n13629 ^ 1'b0 ;
  assign n48658 = n13385 & n48657 ;
  assign n48660 = n48659 ^ n48658 ^ n8001 ;
  assign n48661 = ( ~n10639 & n11367 ) | ( ~n10639 & n48660 ) | ( n11367 & n48660 ) ;
  assign n48662 = n14247 | n21573 ;
  assign n48663 = ( ~n1806 & n32743 ) | ( ~n1806 & n41040 ) | ( n32743 & n41040 ) ;
  assign n48664 = n11608 | n16874 ;
  assign n48665 = n48664 ^ n20318 ^ n5058 ;
  assign n48666 = n48665 ^ n5260 ^ 1'b0 ;
  assign n48667 = ~n48663 & n48666 ;
  assign n48668 = n14653 ^ n14244 ^ n2720 ;
  assign n48669 = n48668 ^ n7404 ^ n6988 ;
  assign n48670 = n37424 ^ n31000 ^ n18870 ;
  assign n48671 = n36946 ^ n19662 ^ n19471 ;
  assign n48672 = ( n8877 & ~n36914 ) | ( n8877 & n48671 ) | ( ~n36914 & n48671 ) ;
  assign n48676 = ( n13042 & n33153 ) | ( n13042 & n39249 ) | ( n33153 & n39249 ) ;
  assign n48673 = n22408 ^ n3904 ^ n499 ;
  assign n48674 = n44222 ^ n17208 ^ 1'b0 ;
  assign n48675 = n48673 & ~n48674 ;
  assign n48677 = n48676 ^ n48675 ^ n30667 ;
  assign n48678 = ~n3855 & n7635 ;
  assign n48679 = n5771 & n48678 ;
  assign n48680 = ( ~n21334 & n29775 ) | ( ~n21334 & n48679 ) | ( n29775 & n48679 ) ;
  assign n48681 = ( n501 & ~n4758 ) | ( n501 & n20890 ) | ( ~n4758 & n20890 ) ;
  assign n48682 = n48681 ^ n18067 ^ n2426 ;
  assign n48683 = ( n23072 & n25778 ) | ( n23072 & ~n48682 ) | ( n25778 & ~n48682 ) ;
  assign n48684 = ( n45468 & ~n48680 ) | ( n45468 & n48683 ) | ( ~n48680 & n48683 ) ;
  assign n48685 = n492 & n26791 ;
  assign n48686 = n11443 & ~n43737 ;
  assign n48687 = n37734 & n48686 ;
  assign n48688 = n4100 & n7009 ;
  assign n48689 = ~n1519 & n48688 ;
  assign n48690 = n48689 ^ n11327 ^ 1'b0 ;
  assign n48691 = n28844 & ~n48690 ;
  assign n48692 = n37011 ^ n25673 ^ n4493 ;
  assign n48693 = n18958 ^ n13406 ^ n1925 ;
  assign n48694 = ( n40197 & n48692 ) | ( n40197 & ~n48693 ) | ( n48692 & ~n48693 ) ;
  assign n48696 = n23815 ^ n5667 ^ 1'b0 ;
  assign n48697 = n7996 & n48696 ;
  assign n48698 = n48697 ^ n22727 ^ n1313 ;
  assign n48695 = n4212 & n37092 ;
  assign n48699 = n48698 ^ n48695 ^ 1'b0 ;
  assign n48700 = n48699 ^ n7476 ^ n6801 ;
  assign n48703 = n34855 ^ n34150 ^ 1'b0 ;
  assign n48704 = n8552 | n48703 ;
  assign n48701 = ( n636 & ~n10394 ) | ( n636 & n16256 ) | ( ~n10394 & n16256 ) ;
  assign n48702 = n48701 ^ n29162 ^ 1'b0 ;
  assign n48705 = n48704 ^ n48702 ^ n45269 ;
  assign n48706 = n5919 | n13562 ;
  assign n48707 = n48706 ^ n24483 ^ 1'b0 ;
  assign n48708 = n48707 ^ n9756 ^ n2308 ;
  assign n48709 = n3791 & ~n12404 ;
  assign n48710 = n48709 ^ n23673 ^ 1'b0 ;
  assign n48711 = n48710 ^ n46458 ^ n12746 ;
  assign n48712 = ( n22549 & n22600 ) | ( n22549 & ~n48711 ) | ( n22600 & ~n48711 ) ;
  assign n48713 = ( n2665 & n12111 ) | ( n2665 & ~n15588 ) | ( n12111 & ~n15588 ) ;
  assign n48714 = n48713 ^ n13600 ^ n977 ;
  assign n48715 = n48714 ^ n27323 ^ n21497 ;
  assign n48716 = n41897 ^ n39001 ^ n25624 ;
  assign n48717 = ( n27389 & n42671 ) | ( n27389 & n48716 ) | ( n42671 & n48716 ) ;
  assign n48718 = ( n25312 & ~n39705 ) | ( n25312 & n48717 ) | ( ~n39705 & n48717 ) ;
  assign n48719 = n31941 | n36924 ;
  assign n48720 = n36080 | n48719 ;
  assign n48721 = n44189 ^ n9782 ^ 1'b0 ;
  assign n48722 = n7927 & n11359 ;
  assign n48723 = n48722 ^ n38101 ^ 1'b0 ;
  assign n48724 = ( n12656 & n41464 ) | ( n12656 & n47948 ) | ( n41464 & n47948 ) ;
  assign n48725 = ( n1184 & n1475 ) | ( n1184 & n7326 ) | ( n1475 & n7326 ) ;
  assign n48726 = n48725 ^ n11656 ^ n4466 ;
  assign n48727 = n48726 ^ n39768 ^ n14056 ;
  assign n48728 = n48727 ^ n27385 ^ n4586 ;
  assign n48729 = ( n16542 & n22393 ) | ( n16542 & n41677 ) | ( n22393 & n41677 ) ;
  assign n48730 = n43336 ^ n22200 ^ n10257 ;
  assign n48732 = ~n18347 & n39621 ;
  assign n48733 = n47411 & n48732 ;
  assign n48731 = ~n1486 & n40033 ;
  assign n48734 = n48733 ^ n48731 ^ n39650 ;
  assign n48735 = n3923 | n6609 ;
  assign n48736 = n13555 ^ n11198 ^ n1848 ;
  assign n48739 = ( n1862 & n11211 ) | ( n1862 & n25833 ) | ( n11211 & n25833 ) ;
  assign n48737 = ~n8067 & n36049 ;
  assign n48738 = n46530 & n48737 ;
  assign n48740 = n48739 ^ n48738 ^ n15475 ;
  assign n48741 = ( n9174 & ~n22415 ) | ( n9174 & n48270 ) | ( ~n22415 & n48270 ) ;
  assign n48742 = n28052 & ~n28292 ;
  assign n48743 = n48742 ^ n11046 ^ 1'b0 ;
  assign n48744 = ( n4472 & n5492 ) | ( n4472 & ~n48743 ) | ( n5492 & ~n48743 ) ;
  assign n48745 = n16702 ^ n15386 ^ n8911 ;
  assign n48746 = n48744 & ~n48745 ;
  assign n48747 = n5567 ^ n3390 ^ 1'b0 ;
  assign n48748 = ~n16332 & n48747 ;
  assign n48749 = ( n11684 & ~n33559 ) | ( n11684 & n48748 ) | ( ~n33559 & n48748 ) ;
  assign n48750 = n6232 ^ n5352 ^ n4741 ;
  assign n48751 = n48750 ^ n15777 ^ n14042 ;
  assign n48752 = n48751 ^ n33441 ^ n23026 ;
  assign n48753 = n41458 ^ n22884 ^ 1'b0 ;
  assign n48754 = n48753 ^ n13091 ^ 1'b0 ;
  assign n48755 = n6289 ^ n959 ^ 1'b0 ;
  assign n48756 = ( n2258 & n17726 ) | ( n2258 & n39837 ) | ( n17726 & n39837 ) ;
  assign n48757 = ( n1789 & ~n48755 ) | ( n1789 & n48756 ) | ( ~n48755 & n48756 ) ;
  assign n48758 = n48757 ^ n34755 ^ 1'b0 ;
  assign n48759 = n7160 & ~n48758 ;
  assign n48760 = n3045 & n5442 ;
  assign n48763 = n48125 ^ n42834 ^ n25130 ;
  assign n48761 = n1647 | n15770 ;
  assign n48762 = n48761 ^ n18664 ^ n16125 ;
  assign n48764 = n48763 ^ n48762 ^ n19406 ;
  assign n48765 = n33005 | n48764 ;
  assign n48766 = ( ~n13546 & n37192 ) | ( ~n13546 & n48765 ) | ( n37192 & n48765 ) ;
  assign n48767 = n12632 & ~n44815 ;
  assign n48768 = ( n29530 & n40315 ) | ( n29530 & n41867 ) | ( n40315 & n41867 ) ;
  assign n48769 = ~n14606 & n22714 ;
  assign n48770 = n48769 ^ n682 ^ 1'b0 ;
  assign n48771 = n5766 & n20525 ;
  assign n48772 = ( ~n8986 & n30875 ) | ( ~n8986 & n48771 ) | ( n30875 & n48771 ) ;
  assign n48773 = n45571 ^ n19394 ^ n7337 ;
  assign n48774 = n48773 ^ n20453 ^ 1'b0 ;
  assign n48775 = n48772 | n48774 ;
  assign n48776 = ( n4030 & n9134 ) | ( n4030 & n17838 ) | ( n9134 & n17838 ) ;
  assign n48777 = n48776 ^ n27894 ^ n13111 ;
  assign n48778 = ( n48770 & n48775 ) | ( n48770 & n48777 ) | ( n48775 & n48777 ) ;
  assign n48779 = ( ~n20103 & n38933 ) | ( ~n20103 & n43832 ) | ( n38933 & n43832 ) ;
  assign n48780 = ( n724 & ~n21220 ) | ( n724 & n27106 ) | ( ~n21220 & n27106 ) ;
  assign n48782 = n42759 ^ n12293 ^ n2525 ;
  assign n48781 = n29472 ^ n24659 ^ 1'b0 ;
  assign n48783 = n48782 ^ n48781 ^ n25025 ;
  assign n48784 = ~n22861 & n46269 ;
  assign n48785 = n8454 & n48784 ;
  assign n48786 = n35515 ^ n25899 ^ 1'b0 ;
  assign n48787 = ~n12438 & n48786 ;
  assign n48788 = n13032 ^ n9589 ^ n2254 ;
  assign n48789 = ( ~n668 & n26152 ) | ( ~n668 & n48788 ) | ( n26152 & n48788 ) ;
  assign n48790 = ( n5827 & n21737 ) | ( n5827 & ~n48789 ) | ( n21737 & ~n48789 ) ;
  assign n48791 = n5471 & n30717 ;
  assign n48792 = n48791 ^ n37122 ^ n16967 ;
  assign n48793 = ( n290 & n19999 ) | ( n290 & ~n25359 ) | ( n19999 & ~n25359 ) ;
  assign n48794 = n48793 ^ n13292 ^ n9093 ;
  assign n48795 = ( n11997 & ~n12334 ) | ( n11997 & n22176 ) | ( ~n12334 & n22176 ) ;
  assign n48796 = ( n13597 & ~n48794 ) | ( n13597 & n48795 ) | ( ~n48794 & n48795 ) ;
  assign n48797 = ~n3441 & n6162 ;
  assign n48798 = ~n3154 & n9799 ;
  assign n48799 = n48798 ^ n15310 ^ 1'b0 ;
  assign n48800 = ~n34963 & n48799 ;
  assign n48801 = ( ~n3545 & n13028 ) | ( ~n3545 & n26743 ) | ( n13028 & n26743 ) ;
  assign n48802 = n48801 ^ n39661 ^ 1'b0 ;
  assign n48803 = n23452 ^ n12685 ^ n7467 ;
  assign n48804 = n17762 & n21479 ;
  assign n48805 = n48804 ^ n8855 ^ n5398 ;
  assign n48806 = n48803 | n48805 ;
  assign n48807 = n2077 & n11444 ;
  assign n48808 = n17515 & n29330 ;
  assign n48809 = n48808 ^ n14324 ^ 1'b0 ;
  assign n48810 = n48809 ^ n24223 ^ 1'b0 ;
  assign n48811 = ( n17276 & n28527 ) | ( n17276 & ~n48810 ) | ( n28527 & ~n48810 ) ;
  assign n48812 = n10594 | n18018 ;
  assign n48813 = ( n14753 & n24914 ) | ( n14753 & n36519 ) | ( n24914 & n36519 ) ;
  assign n48814 = ( n9486 & n20990 ) | ( n9486 & n24650 ) | ( n20990 & n24650 ) ;
  assign n48815 = n20877 & ~n30915 ;
  assign n48816 = n48815 ^ n13744 ^ 1'b0 ;
  assign n48817 = n48816 ^ n27159 ^ 1'b0 ;
  assign n48818 = ~n17751 & n39201 ;
  assign n48819 = n48818 ^ n9930 ^ 1'b0 ;
  assign n48820 = n21219 & ~n48819 ;
  assign n48823 = n16836 & n31549 ;
  assign n48824 = n48823 ^ n13349 ^ 1'b0 ;
  assign n48821 = ~n545 & n9218 ;
  assign n48822 = n48821 ^ n22096 ^ 1'b0 ;
  assign n48825 = n48824 ^ n48822 ^ 1'b0 ;
  assign n48826 = n37325 & n48825 ;
  assign n48827 = n17798 ^ n5513 ^ 1'b0 ;
  assign n48828 = n40792 | n44891 ;
  assign n48829 = n48589 | n48828 ;
  assign n48830 = n40886 ^ n991 ^ 1'b0 ;
  assign n48831 = n19646 ^ n16356 ^ n5723 ;
  assign n48832 = ( ~n8047 & n8759 ) | ( ~n8047 & n48831 ) | ( n8759 & n48831 ) ;
  assign n48834 = n2399 & n22506 ;
  assign n48833 = ( n1996 & n2039 ) | ( n1996 & n44116 ) | ( n2039 & n44116 ) ;
  assign n48835 = n48834 ^ n48833 ^ n33955 ;
  assign n48836 = x241 & n24103 ;
  assign n48837 = ( ~n23390 & n42488 ) | ( ~n23390 & n48836 ) | ( n42488 & n48836 ) ;
  assign n48838 = n48837 ^ n23637 ^ n14589 ;
  assign n48839 = n48835 & ~n48838 ;
  assign n48840 = n15231 ^ n2488 ^ n599 ;
  assign n48841 = n31490 ^ n11862 ^ n1288 ;
  assign n48842 = n21622 ^ n16248 ^ n11476 ;
  assign n48843 = n16288 & n41907 ;
  assign n48844 = n26815 & n48843 ;
  assign n48845 = n19725 ^ n8400 ^ 1'b0 ;
  assign n48846 = n1465 & ~n48845 ;
  assign n48847 = n45503 & n48846 ;
  assign n48848 = n8004 | n41755 ;
  assign n48849 = n25374 ^ n8967 ^ n3450 ;
  assign n48850 = n48849 ^ n30311 ^ n16400 ;
  assign n48851 = ( n9358 & ~n24507 ) | ( n9358 & n25939 ) | ( ~n24507 & n25939 ) ;
  assign n48852 = n48851 ^ n33698 ^ 1'b0 ;
  assign n48853 = n24892 ^ n3510 ^ 1'b0 ;
  assign n48854 = n12023 ^ n6114 ^ 1'b0 ;
  assign n48855 = ~n284 & n48854 ;
  assign n48856 = n48855 ^ n1124 ^ 1'b0 ;
  assign n48857 = n4949 & ~n48856 ;
  assign n48858 = ~n5504 & n17437 ;
  assign n48859 = n24016 ^ n14033 ^ n13412 ;
  assign n48860 = n8022 & n33640 ;
  assign n48861 = ( n36999 & n48859 ) | ( n36999 & ~n48860 ) | ( n48859 & ~n48860 ) ;
  assign n48862 = ( n41458 & n45064 ) | ( n41458 & ~n48861 ) | ( n45064 & ~n48861 ) ;
  assign n48863 = ( n4700 & n48858 ) | ( n4700 & ~n48862 ) | ( n48858 & ~n48862 ) ;
  assign n48864 = n6484 | n27955 ;
  assign n48865 = n5666 | n48864 ;
  assign n48868 = n8744 ^ n8743 ^ n5963 ;
  assign n48866 = ( n1490 & n11480 ) | ( n1490 & n34036 ) | ( n11480 & n34036 ) ;
  assign n48867 = n39853 & ~n48866 ;
  assign n48869 = n48868 ^ n48867 ^ n14866 ;
  assign n48871 = n41787 | n45455 ;
  assign n48870 = n45718 ^ n36316 ^ n21159 ;
  assign n48872 = n48871 ^ n48870 ^ n14482 ;
  assign n48873 = ( ~n5894 & n16659 ) | ( ~n5894 & n21440 ) | ( n16659 & n21440 ) ;
  assign n48874 = n30027 ^ n9249 ^ 1'b0 ;
  assign n48875 = n48873 & n48874 ;
  assign n48876 = n48875 ^ n44847 ^ n17344 ;
  assign n48877 = n10248 & n42080 ;
  assign n48878 = n18517 & n29040 ;
  assign n48879 = n48878 ^ n5552 ^ 1'b0 ;
  assign n48880 = n48879 ^ n46838 ^ n9605 ;
  assign n48883 = ( n11131 & n12264 ) | ( n11131 & n24100 ) | ( n12264 & n24100 ) ;
  assign n48881 = ~n40175 & n46521 ;
  assign n48882 = n44513 & n48881 ;
  assign n48884 = n48883 ^ n48882 ^ n33466 ;
  assign n48885 = ( n18094 & ~n28658 ) | ( n18094 & n28953 ) | ( ~n28658 & n28953 ) ;
  assign n48886 = n5986 | n9698 ;
  assign n48887 = n7455 & ~n43007 ;
  assign n48888 = n48887 ^ n22686 ^ 1'b0 ;
  assign n48889 = n38328 ^ n35300 ^ 1'b0 ;
  assign n48890 = n28917 | n48889 ;
  assign n48891 = ( ~n31157 & n32881 ) | ( ~n31157 & n48890 ) | ( n32881 & n48890 ) ;
  assign n48892 = ( n3014 & ~n10033 ) | ( n3014 & n29340 ) | ( ~n10033 & n29340 ) ;
  assign n48893 = ( n12271 & n13123 ) | ( n12271 & n40453 ) | ( n13123 & n40453 ) ;
  assign n48894 = ( n5786 & n25468 ) | ( n5786 & n48893 ) | ( n25468 & n48893 ) ;
  assign n48897 = n7585 & ~n37932 ;
  assign n48896 = ( ~x190 & n16578 ) | ( ~x190 & n18935 ) | ( n16578 & n18935 ) ;
  assign n48895 = n34325 ^ n13689 ^ n9565 ;
  assign n48898 = n48897 ^ n48896 ^ n48895 ;
  assign n48899 = ( n7177 & n23850 ) | ( n7177 & n48898 ) | ( n23850 & n48898 ) ;
  assign n48900 = ( n5723 & n27305 ) | ( n5723 & n33207 ) | ( n27305 & n33207 ) ;
  assign n48901 = ( ~n15172 & n35227 ) | ( ~n15172 & n48900 ) | ( n35227 & n48900 ) ;
  assign n48902 = n42386 & n48901 ;
  assign n48903 = n8697 & n48902 ;
  assign n48904 = n48259 ^ n11546 ^ 1'b0 ;
  assign n48905 = ( n1649 & ~n4438 ) | ( n1649 & n25674 ) | ( ~n4438 & n25674 ) ;
  assign n48906 = n9007 & ~n48905 ;
  assign n48907 = ( n19134 & ~n33724 ) | ( n19134 & n38915 ) | ( ~n33724 & n38915 ) ;
  assign n48908 = n31170 & ~n48907 ;
  assign n48909 = n38244 ^ n1549 ^ 1'b0 ;
  assign n48910 = ~n48908 & n48909 ;
  assign n48911 = n26062 ^ n2866 ^ 1'b0 ;
  assign n48912 = n37706 ^ n21023 ^ n8155 ;
  assign n48914 = n14649 | n14760 ;
  assign n48915 = n48914 ^ n26406 ^ 1'b0 ;
  assign n48916 = n48915 ^ n36469 ^ n32927 ;
  assign n48913 = n48273 ^ n21816 ^ n2795 ;
  assign n48917 = n48916 ^ n48913 ^ n8389 ;
  assign n48918 = n12215 | n12634 ;
  assign n48919 = ( n12045 & n20532 ) | ( n12045 & n34058 ) | ( n20532 & n34058 ) ;
  assign n48920 = ( n11406 & n36320 ) | ( n11406 & ~n48919 ) | ( n36320 & ~n48919 ) ;
  assign n48921 = ( ~n1334 & n1973 ) | ( ~n1334 & n12371 ) | ( n1973 & n12371 ) ;
  assign n48922 = n14203 & n29689 ;
  assign n48923 = n7778 & n48922 ;
  assign n48924 = n12074 ^ n7456 ^ n6208 ;
  assign n48925 = n6102 & n48924 ;
  assign n48926 = n14698 | n47072 ;
  assign n48927 = n41548 ^ n10101 ^ 1'b0 ;
  assign n48928 = n13775 & n27974 ;
  assign n48929 = n48928 ^ n36126 ^ 1'b0 ;
  assign n48930 = n48929 ^ n22010 ^ 1'b0 ;
  assign n48931 = n9785 & n36557 ;
  assign n48932 = n14822 ^ n5396 ^ n1855 ;
  assign n48933 = n48932 ^ n38061 ^ n16596 ;
  assign n48934 = n5844 | n48933 ;
  assign n48935 = n5686 ^ n3542 ^ 1'b0 ;
  assign n48936 = ( n2060 & n11345 ) | ( n2060 & ~n48935 ) | ( n11345 & ~n48935 ) ;
  assign n48937 = n23234 ^ n21414 ^ 1'b0 ;
  assign n48938 = n6008 & n48937 ;
  assign n48939 = n48938 ^ n20558 ^ 1'b0 ;
  assign n48940 = n5622 & ~n30156 ;
  assign n48941 = n6576 & n39581 ;
  assign n48942 = ~n399 & n48941 ;
  assign n48943 = n48942 ^ n32896 ^ n5417 ;
  assign n48944 = n45741 ^ n14048 ^ n6056 ;
  assign n48945 = n29730 ^ n25702 ^ 1'b0 ;
  assign n48946 = ~n34087 & n48945 ;
  assign n48947 = n46337 ^ n10421 ^ n1137 ;
  assign n48948 = n11331 ^ n9775 ^ n8067 ;
  assign n48949 = ~n14439 & n48948 ;
  assign n48950 = n22553 ^ n18405 ^ n7150 ;
  assign n48951 = n5491 & ~n48950 ;
  assign n48952 = n14808 & n25299 ;
  assign n48953 = n47325 & n48952 ;
  assign n48954 = n28837 & n33636 ;
  assign n48955 = ~n21101 & n48954 ;
  assign n48956 = n9416 ^ n2142 ^ 1'b0 ;
  assign n48957 = ~n18583 & n48956 ;
  assign n48958 = n21862 ^ n3015 ^ 1'b0 ;
  assign n48959 = n12986 & ~n31797 ;
  assign n48960 = n48959 ^ n39407 ^ 1'b0 ;
  assign n48961 = n35239 | n44381 ;
  assign n48962 = n48960 | n48961 ;
  assign n48963 = ( n26311 & n48958 ) | ( n26311 & n48962 ) | ( n48958 & n48962 ) ;
  assign n48965 = ( n3287 & n3822 ) | ( n3287 & ~n5261 ) | ( n3822 & ~n5261 ) ;
  assign n48966 = n48965 ^ n16451 ^ n13675 ;
  assign n48964 = n11256 & ~n32288 ;
  assign n48967 = n48966 ^ n48964 ^ n16904 ;
  assign n48968 = n5040 & ~n37150 ;
  assign n48969 = ( n2862 & n7322 ) | ( n2862 & ~n22780 ) | ( n7322 & ~n22780 ) ;
  assign n48970 = n48969 ^ n45992 ^ n983 ;
  assign n48971 = n46217 ^ n15987 ^ n2125 ;
  assign n48972 = n23018 | n39735 ;
  assign n48973 = n48972 ^ n3728 ^ 1'b0 ;
  assign n48974 = ( n1096 & n10101 ) | ( n1096 & n23745 ) | ( n10101 & n23745 ) ;
  assign n48975 = n7244 & n48974 ;
  assign n48976 = ~n4728 & n18097 ;
  assign n48977 = n48976 ^ n29548 ^ 1'b0 ;
  assign n48978 = n45090 ^ n21624 ^ n21371 ;
  assign n48979 = n48978 ^ n12360 ^ n2762 ;
  assign n48980 = n32465 ^ n14952 ^ n9366 ;
  assign n48981 = n38851 ^ n20448 ^ n5719 ;
  assign n48982 = ( n17123 & ~n27363 ) | ( n17123 & n48981 ) | ( ~n27363 & n48981 ) ;
  assign n48983 = ( ~n903 & n37716 ) | ( ~n903 & n48982 ) | ( n37716 & n48982 ) ;
  assign n48984 = n2244 & n6477 ;
  assign n48985 = ( n10398 & ~n22904 ) | ( n10398 & n35973 ) | ( ~n22904 & n35973 ) ;
  assign n48986 = ( ~n15947 & n48984 ) | ( ~n15947 & n48985 ) | ( n48984 & n48985 ) ;
  assign n48987 = n31242 ^ n25788 ^ 1'b0 ;
  assign n48988 = ( ~n12815 & n28812 ) | ( ~n12815 & n31401 ) | ( n28812 & n31401 ) ;
  assign n48989 = ~n3721 & n16788 ;
  assign n48990 = ( n12593 & n15437 ) | ( n12593 & ~n48989 ) | ( n15437 & ~n48989 ) ;
  assign n48991 = ~n34018 & n48990 ;
  assign n48992 = n4163 ^ n3782 ^ 1'b0 ;
  assign n48993 = n6109 & ~n48992 ;
  assign n48994 = n41294 ^ n33584 ^ n7247 ;
  assign n48995 = n15819 & ~n19209 ;
  assign n48996 = n48995 ^ n8397 ^ 1'b0 ;
  assign n48998 = n16343 & n19604 ;
  assign n48999 = n48998 ^ n15737 ^ 1'b0 ;
  assign n48997 = n33173 & n43099 ;
  assign n49000 = n48999 ^ n48997 ^ 1'b0 ;
  assign n49001 = ~n24035 & n33065 ;
  assign n49002 = n49001 ^ n1538 ^ 1'b0 ;
  assign n49003 = ( n48996 & n49000 ) | ( n48996 & n49002 ) | ( n49000 & n49002 ) ;
  assign n49004 = n44327 ^ n32825 ^ 1'b0 ;
  assign n49005 = n17350 | n20119 ;
  assign n49006 = n45537 ^ n35861 ^ n31053 ;
  assign n49007 = n49006 ^ n19900 ^ 1'b0 ;
  assign n49008 = n49005 & n49007 ;
  assign n49009 = ~n10877 & n49008 ;
  assign n49010 = n8412 & n49009 ;
  assign n49011 = n49010 ^ n18645 ^ n11880 ;
  assign n49012 = n30553 ^ n9631 ^ n4692 ;
  assign n49013 = n49012 ^ n40527 ^ n38449 ;
  assign n49015 = ( n1173 & n27033 ) | ( n1173 & ~n30695 ) | ( n27033 & ~n30695 ) ;
  assign n49016 = ( n12409 & n32373 ) | ( n12409 & n49015 ) | ( n32373 & n49015 ) ;
  assign n49014 = ~n29656 & n45396 ;
  assign n49017 = n49016 ^ n49014 ^ 1'b0 ;
  assign n49018 = n1555 & n24505 ;
  assign n49019 = n49018 ^ n4397 ^ 1'b0 ;
  assign n49020 = n49019 ^ n7636 ^ 1'b0 ;
  assign n49021 = n28568 ^ n16227 ^ n10725 ;
  assign n49022 = n47206 ^ n35916 ^ n18029 ;
  assign n49023 = n25297 ^ n8423 ^ 1'b0 ;
  assign n49025 = ( n1686 & n24424 ) | ( n1686 & n25861 ) | ( n24424 & n25861 ) ;
  assign n49024 = ( n7890 & ~n28151 ) | ( n7890 & n37947 ) | ( ~n28151 & n37947 ) ;
  assign n49026 = n49025 ^ n49024 ^ n9214 ;
  assign n49027 = ( n22317 & n24850 ) | ( n22317 & ~n47275 ) | ( n24850 & ~n47275 ) ;
  assign n49028 = n28680 ^ n16514 ^ n9888 ;
  assign n49029 = ( n30414 & ~n39507 ) | ( n30414 & n40910 ) | ( ~n39507 & n40910 ) ;
  assign n49030 = ~n15647 & n17009 ;
  assign n49031 = n18663 & n49030 ;
  assign n49032 = n37414 ^ n23048 ^ n9997 ;
  assign n49033 = n49032 ^ n32624 ^ 1'b0 ;
  assign n49034 = n24854 ^ n24409 ^ n5319 ;
  assign n49035 = ~n35553 & n49034 ;
  assign n49036 = ~n44657 & n49035 ;
  assign n49037 = ( n273 & n11795 ) | ( n273 & n31649 ) | ( n11795 & n31649 ) ;
  assign n49038 = n3330 | n49037 ;
  assign n49039 = n28805 & ~n49038 ;
  assign n49040 = ( n12776 & n20528 ) | ( n12776 & ~n25338 ) | ( n20528 & ~n25338 ) ;
  assign n49041 = ~n545 & n6529 ;
  assign n49042 = ~n7168 & n49041 ;
  assign n49043 = ~n4493 & n49042 ;
  assign n49044 = n6596 & ~n49043 ;
  assign n49045 = n13090 & n49044 ;
  assign n49046 = n49045 ^ n35670 ^ n2281 ;
  assign n49047 = n19261 & n21106 ;
  assign n49048 = n44397 ^ n19742 ^ n273 ;
  assign n49049 = n25275 & n44769 ;
  assign n49050 = n25834 ^ n6999 ^ n3288 ;
  assign n49051 = n12234 ^ n2939 ^ n1394 ;
  assign n49052 = n6587 | n49051 ;
  assign n49053 = n49052 ^ n44663 ^ 1'b0 ;
  assign n49054 = n10249 ^ n8290 ^ n2174 ;
  assign n49055 = n49054 ^ n31811 ^ 1'b0 ;
  assign n49056 = n49053 & ~n49055 ;
  assign n49057 = n43490 ^ n30961 ^ 1'b0 ;
  assign n49058 = n34554 ^ n24228 ^ n7665 ;
  assign n49059 = ( n3638 & n26293 ) | ( n3638 & ~n45869 ) | ( n26293 & ~n45869 ) ;
  assign n49060 = n49059 ^ n42756 ^ 1'b0 ;
  assign n49061 = ( n9153 & n36053 ) | ( n9153 & n39133 ) | ( n36053 & n39133 ) ;
  assign n49062 = ( ~n13083 & n17732 ) | ( ~n13083 & n34218 ) | ( n17732 & n34218 ) ;
  assign n49063 = ( n38902 & n49061 ) | ( n38902 & n49062 ) | ( n49061 & n49062 ) ;
  assign n49064 = n22913 ^ n16600 ^ n6923 ;
  assign n49065 = ~n10020 & n49064 ;
  assign n49066 = n42602 & ~n49065 ;
  assign n49067 = n2062 ^ n698 ^ 1'b0 ;
  assign n49068 = ( n7197 & n49066 ) | ( n7197 & n49067 ) | ( n49066 & n49067 ) ;
  assign n49072 = ( n3227 & ~n10830 ) | ( n3227 & n22420 ) | ( ~n10830 & n22420 ) ;
  assign n49069 = ( ~n3502 & n8470 ) | ( ~n3502 & n10765 ) | ( n8470 & n10765 ) ;
  assign n49070 = ( n704 & n1420 ) | ( n704 & n27468 ) | ( n1420 & n27468 ) ;
  assign n49071 = ( n40479 & n49069 ) | ( n40479 & ~n49070 ) | ( n49069 & ~n49070 ) ;
  assign n49073 = n49072 ^ n49071 ^ n46959 ;
  assign n49074 = n29560 ^ n14641 ^ 1'b0 ;
  assign n49075 = n49074 ^ n28781 ^ n18424 ;
  assign n49076 = n49075 ^ n44642 ^ n32073 ;
  assign n49077 = ~n23490 & n26059 ;
  assign n49078 = n26334 & ~n49077 ;
  assign n49080 = ( n2697 & n17589 ) | ( n2697 & ~n25996 ) | ( n17589 & ~n25996 ) ;
  assign n49079 = n6191 | n21682 ;
  assign n49081 = n49080 ^ n49079 ^ 1'b0 ;
  assign n49082 = ( n7013 & ~n11044 ) | ( n7013 & n29864 ) | ( ~n11044 & n29864 ) ;
  assign n49083 = ~n2981 & n22424 ;
  assign n49084 = n12038 | n16130 ;
  assign n49085 = n22132 & ~n49084 ;
  assign n49086 = n49085 ^ n33986 ^ n19867 ;
  assign n49087 = n27864 ^ n15436 ^ 1'b0 ;
  assign n49088 = ( ~n21934 & n49086 ) | ( ~n21934 & n49087 ) | ( n49086 & n49087 ) ;
  assign n49089 = n8456 & ~n37482 ;
  assign n49090 = n3402 | n3501 ;
  assign n49091 = n49090 ^ n9096 ^ 1'b0 ;
  assign n49092 = ~n26976 & n49091 ;
  assign n49094 = n13762 ^ n10945 ^ 1'b0 ;
  assign n49095 = ~n46392 & n49094 ;
  assign n49093 = ( n7609 & n16753 ) | ( n7609 & ~n38341 ) | ( n16753 & ~n38341 ) ;
  assign n49096 = n49095 ^ n49093 ^ 1'b0 ;
  assign n49097 = n42499 ^ n29844 ^ 1'b0 ;
  assign n49098 = n37386 & n49097 ;
  assign n49099 = n32527 ^ n15912 ^ 1'b0 ;
  assign n49100 = n18388 & ~n47110 ;
  assign n49101 = ~n21988 & n49100 ;
  assign n49102 = n28106 ^ n2825 ^ 1'b0 ;
  assign n49103 = n44334 ^ n24456 ^ n7635 ;
  assign n49104 = n4995 ^ n2139 ^ x128 ;
  assign n49105 = n49104 ^ n18032 ^ n15400 ;
  assign n49106 = ( n3716 & ~n16684 ) | ( n3716 & n34903 ) | ( ~n16684 & n34903 ) ;
  assign n49107 = n34484 ^ n15515 ^ n3111 ;
  assign n49108 = ( n17343 & ~n49106 ) | ( n17343 & n49107 ) | ( ~n49106 & n49107 ) ;
  assign n49109 = n31736 ^ n22080 ^ n8463 ;
  assign n49110 = n29680 ^ n14507 ^ 1'b0 ;
  assign n49111 = ( x16 & n13374 ) | ( x16 & ~n49110 ) | ( n13374 & ~n49110 ) ;
  assign n49113 = n26084 ^ n13883 ^ 1'b0 ;
  assign n49112 = n29079 | n30574 ;
  assign n49114 = n49113 ^ n49112 ^ n3713 ;
  assign n49115 = ( n21038 & ~n29067 ) | ( n21038 & n49114 ) | ( ~n29067 & n49114 ) ;
  assign n49116 = n24965 ^ n3999 ^ 1'b0 ;
  assign n49117 = n8310 & n28938 ;
  assign n49118 = n6556 & n49117 ;
  assign n49119 = ( n31433 & n49116 ) | ( n31433 & ~n49118 ) | ( n49116 & ~n49118 ) ;
  assign n49121 = n6252 & ~n6886 ;
  assign n49122 = n49121 ^ n19262 ^ 1'b0 ;
  assign n49120 = n10870 & n31302 ;
  assign n49123 = n49122 ^ n49120 ^ 1'b0 ;
  assign n49124 = ~n23527 & n37737 ;
  assign n49125 = n49124 ^ n31191 ^ 1'b0 ;
  assign n49127 = ( n8000 & n15352 ) | ( n8000 & ~n22197 ) | ( n15352 & ~n22197 ) ;
  assign n49126 = ( n819 & n10970 ) | ( n819 & ~n31300 ) | ( n10970 & ~n31300 ) ;
  assign n49128 = n49127 ^ n49126 ^ n35412 ;
  assign n49129 = n48152 ^ n25593 ^ n1133 ;
  assign n49130 = n27570 ^ n21126 ^ n13540 ;
  assign n49131 = ( n3026 & ~n7627 ) | ( n3026 & n33461 ) | ( ~n7627 & n33461 ) ;
  assign n49132 = ( n5396 & ~n26281 ) | ( n5396 & n45426 ) | ( ~n26281 & n45426 ) ;
  assign n49133 = ( n36097 & ~n49131 ) | ( n36097 & n49132 ) | ( ~n49131 & n49132 ) ;
  assign n49134 = ( n4066 & n4368 ) | ( n4066 & ~n27864 ) | ( n4368 & ~n27864 ) ;
  assign n49135 = n49134 ^ n26198 ^ n15600 ;
  assign n49136 = ( n11293 & n20244 ) | ( n11293 & ~n49135 ) | ( n20244 & ~n49135 ) ;
  assign n49137 = n49136 ^ n40376 ^ n35033 ;
  assign n49138 = ( n5064 & n18473 ) | ( n5064 & n21327 ) | ( n18473 & n21327 ) ;
  assign n49139 = ( n1610 & n36549 ) | ( n1610 & ~n49138 ) | ( n36549 & ~n49138 ) ;
  assign n49140 = n46605 ^ n18637 ^ n12781 ;
  assign n49141 = n34144 & ~n49140 ;
  assign n49142 = n49141 ^ n21051 ^ 1'b0 ;
  assign n49143 = n21823 | n49142 ;
  assign n49145 = n36924 ^ n31401 ^ n25711 ;
  assign n49144 = ~n16564 & n44599 ;
  assign n49146 = n49145 ^ n49144 ^ 1'b0 ;
  assign n49147 = n1743 | n49146 ;
  assign n49148 = n49147 ^ n27614 ^ 1'b0 ;
  assign n49149 = n5597 & n45615 ;
  assign n49150 = n10514 & n49149 ;
  assign n49151 = ~n28355 & n37670 ;
  assign n49152 = n42556 & n49151 ;
  assign n49153 = n43813 ^ n27438 ^ n7013 ;
  assign n49154 = n49153 ^ n31052 ^ n20175 ;
  assign n49155 = n35524 ^ n29783 ^ n18162 ;
  assign n49156 = n49155 ^ x62 ^ 1'b0 ;
  assign n49157 = n45808 ^ n34596 ^ 1'b0 ;
  assign n49158 = ( ~n18932 & n44850 ) | ( ~n18932 & n49157 ) | ( n44850 & n49157 ) ;
  assign n49159 = n26883 ^ n17910 ^ n4000 ;
  assign n49160 = ( n26907 & n41596 ) | ( n26907 & n42612 ) | ( n41596 & n42612 ) ;
  assign n49161 = n25117 & ~n43072 ;
  assign n49162 = n27988 & n49161 ;
  assign n49163 = n19640 ^ n7859 ^ 1'b0 ;
  assign n49164 = ~n12842 & n49163 ;
  assign n49165 = ( n11063 & n34684 ) | ( n11063 & ~n37256 ) | ( n34684 & ~n37256 ) ;
  assign n49166 = ( n5750 & ~n9908 ) | ( n5750 & n19674 ) | ( ~n9908 & n19674 ) ;
  assign n49167 = ( ~n9466 & n35247 ) | ( ~n9466 & n49166 ) | ( n35247 & n49166 ) ;
  assign n49169 = n21143 ^ n20099 ^ n7950 ;
  assign n49168 = n16984 & ~n42099 ;
  assign n49170 = n49169 ^ n49168 ^ 1'b0 ;
  assign n49171 = ( ~n14372 & n49167 ) | ( ~n14372 & n49170 ) | ( n49167 & n49170 ) ;
  assign n49172 = n16540 | n22830 ;
  assign n49173 = ( n9176 & n40435 ) | ( n9176 & n49172 ) | ( n40435 & n49172 ) ;
  assign n49174 = n49173 ^ n21629 ^ n14172 ;
  assign n49175 = n43914 ^ n8410 ^ n602 ;
  assign n49176 = ( ~n13080 & n26454 ) | ( ~n13080 & n36370 ) | ( n26454 & n36370 ) ;
  assign n49177 = ( n7279 & ~n49175 ) | ( n7279 & n49176 ) | ( ~n49175 & n49176 ) ;
  assign n49178 = n35205 ^ n26952 ^ n14310 ;
  assign n49179 = ( ~n5370 & n18917 ) | ( ~n5370 & n45619 ) | ( n18917 & n45619 ) ;
  assign n49180 = n31345 ^ n22713 ^ 1'b0 ;
  assign n49181 = n36679 ^ n16999 ^ 1'b0 ;
  assign n49182 = n30551 & ~n49181 ;
  assign n49183 = ( n14468 & n28094 ) | ( n14468 & n33334 ) | ( n28094 & n33334 ) ;
  assign n49184 = n6351 & n49183 ;
  assign n49185 = n48559 & n49184 ;
  assign n49186 = n14897 & ~n41439 ;
  assign n49187 = n43537 & n49186 ;
  assign n49188 = ( n8356 & n20873 ) | ( n8356 & n37806 ) | ( n20873 & n37806 ) ;
  assign n49189 = n42488 ^ n12646 ^ 1'b0 ;
  assign n49190 = n43656 ^ n23653 ^ n7922 ;
  assign n49191 = ( n14976 & n18431 ) | ( n14976 & ~n42751 ) | ( n18431 & ~n42751 ) ;
  assign n49192 = n7531 & n23129 ;
  assign n49193 = ( n19511 & ~n34480 ) | ( n19511 & n49192 ) | ( ~n34480 & n49192 ) ;
  assign n49194 = n23562 ^ n3912 ^ 1'b0 ;
  assign n49195 = n582 & n49194 ;
  assign n49196 = ( n2568 & ~n5876 ) | ( n2568 & n49195 ) | ( ~n5876 & n49195 ) ;
  assign n49197 = n535 | n4397 ;
  assign n49198 = n14203 | n49197 ;
  assign n49199 = ( n10257 & ~n17993 ) | ( n10257 & n29431 ) | ( ~n17993 & n29431 ) ;
  assign n49200 = n49199 ^ n3758 ^ 1'b0 ;
  assign n49201 = ~n31380 & n49200 ;
  assign n49202 = ~n1819 & n49201 ;
  assign n49203 = ( n14010 & n49198 ) | ( n14010 & ~n49202 ) | ( n49198 & ~n49202 ) ;
  assign n49204 = n15775 & ~n29752 ;
  assign n49205 = ~n49203 & n49204 ;
  assign n49206 = n29702 ^ n1031 ^ 1'b0 ;
  assign n49207 = n15846 & ~n49206 ;
  assign n49208 = ~n4279 & n14771 ;
  assign n49209 = n40256 & n49208 ;
  assign n49210 = n21271 ^ n8804 ^ 1'b0 ;
  assign n49211 = ( n5521 & ~n33479 ) | ( n5521 & n49210 ) | ( ~n33479 & n49210 ) ;
  assign n49212 = ( ~n4736 & n20567 ) | ( ~n4736 & n49211 ) | ( n20567 & n49211 ) ;
  assign n49213 = n46736 ^ n28999 ^ n2039 ;
  assign n49214 = n39061 ^ n12806 ^ 1'b0 ;
  assign n49215 = n49214 ^ n7224 ^ n275 ;
  assign n49216 = n44162 ^ n35435 ^ n1188 ;
  assign n49217 = n26322 ^ n3444 ^ 1'b0 ;
  assign n49218 = ( n34613 & n42172 ) | ( n34613 & ~n47852 ) | ( n42172 & ~n47852 ) ;
  assign n49219 = ( n22172 & n25845 ) | ( n22172 & ~n39118 ) | ( n25845 & ~n39118 ) ;
  assign n49220 = n49219 ^ n2903 ^ 1'b0 ;
  assign n49221 = n6298 & ~n16956 ;
  assign n49222 = ~n16267 & n49221 ;
  assign n49225 = n9408 ^ n7824 ^ n4399 ;
  assign n49223 = n40759 ^ n35575 ^ n12086 ;
  assign n49224 = n11405 & ~n49223 ;
  assign n49226 = n49225 ^ n49224 ^ 1'b0 ;
  assign n49227 = ( n14771 & n17619 ) | ( n14771 & n26642 ) | ( n17619 & n26642 ) ;
  assign n49228 = n49227 ^ n37467 ^ 1'b0 ;
  assign n49229 = n48048 | n49228 ;
  assign n49230 = n8383 ^ n5881 ^ 1'b0 ;
  assign n49231 = n46373 & ~n49230 ;
  assign n49232 = n35644 ^ n35518 ^ n14203 ;
  assign n49233 = ( ~n3387 & n4160 ) | ( ~n3387 & n9974 ) | ( n4160 & n9974 ) ;
  assign n49234 = ( n9542 & ~n13710 ) | ( n9542 & n25983 ) | ( ~n13710 & n25983 ) ;
  assign n49235 = x227 & n1146 ;
  assign n49236 = ( n3216 & n8405 ) | ( n3216 & ~n49235 ) | ( n8405 & ~n49235 ) ;
  assign n49237 = n26834 ^ n2465 ^ 1'b0 ;
  assign n49238 = ( n7865 & ~n13935 ) | ( n7865 & n49237 ) | ( ~n13935 & n49237 ) ;
  assign n49239 = n30627 ^ n21325 ^ n13757 ;
  assign n49240 = ( n11916 & n35776 ) | ( n11916 & ~n37296 ) | ( n35776 & ~n37296 ) ;
  assign n49241 = ( n1603 & ~n49239 ) | ( n1603 & n49240 ) | ( ~n49239 & n49240 ) ;
  assign n49242 = n48160 ^ n36152 ^ n33201 ;
  assign n49243 = n33509 ^ n2528 ^ 1'b0 ;
  assign n49244 = ( n2091 & n4537 ) | ( n2091 & n27045 ) | ( n4537 & n27045 ) ;
  assign n49245 = n38617 | n49244 ;
  assign n49246 = ( ~n8062 & n36159 ) | ( ~n8062 & n38415 ) | ( n36159 & n38415 ) ;
  assign n49247 = n49246 ^ n15552 ^ n7010 ;
  assign n49248 = n7735 & ~n34838 ;
  assign n49249 = ( ~n36699 & n49247 ) | ( ~n36699 & n49248 ) | ( n49247 & n49248 ) ;
  assign n49250 = n20715 ^ n11475 ^ n3905 ;
  assign n49251 = ~n27416 & n33739 ;
  assign n49252 = n28916 | n44156 ;
  assign n49253 = n49252 ^ n18681 ^ n17408 ;
  assign n49254 = ( n1855 & n2519 ) | ( n1855 & n49253 ) | ( n2519 & n49253 ) ;
  assign n49255 = n12639 ^ n4788 ^ 1'b0 ;
  assign n49256 = n5948 & ~n49255 ;
  assign n49257 = ~n2417 & n10455 ;
  assign n49258 = n9117 & n49257 ;
  assign n49259 = n49258 ^ n28252 ^ n6365 ;
  assign n49260 = ( n8418 & ~n8904 ) | ( n8418 & n16834 ) | ( ~n8904 & n16834 ) ;
  assign n49261 = n49260 ^ n42513 ^ n23049 ;
  assign n49262 = n9778 ^ n9144 ^ n1583 ;
  assign n49263 = n4405 & n22344 ;
  assign n49264 = ( n15388 & n19603 ) | ( n15388 & n49263 ) | ( n19603 & n49263 ) ;
  assign n49267 = x195 & n10778 ;
  assign n49268 = n29935 & n49267 ;
  assign n49265 = ( n8033 & ~n8712 ) | ( n8033 & n12328 ) | ( ~n8712 & n12328 ) ;
  assign n49266 = x78 & ~n49265 ;
  assign n49269 = n49268 ^ n49266 ^ n3157 ;
  assign n49270 = ( n49262 & n49264 ) | ( n49262 & ~n49269 ) | ( n49264 & ~n49269 ) ;
  assign n49271 = ( n20433 & n24717 ) | ( n20433 & n25646 ) | ( n24717 & n25646 ) ;
  assign n49272 = n49271 ^ n43936 ^ n16368 ;
  assign n49273 = n48464 ^ n38753 ^ n31248 ;
  assign n49276 = ~n639 & n8799 ;
  assign n49277 = n49276 ^ n4554 ^ 1'b0 ;
  assign n49274 = ( n11051 & n29139 ) | ( n11051 & ~n43991 ) | ( n29139 & ~n43991 ) ;
  assign n49275 = n49274 ^ n12736 ^ 1'b0 ;
  assign n49278 = n49277 ^ n49275 ^ n11734 ;
  assign n49279 = n46970 ^ n15490 ^ 1'b0 ;
  assign n49280 = n16961 | n49279 ;
  assign n49281 = n49280 ^ n37355 ^ 1'b0 ;
  assign n49282 = n9655 & n25020 ;
  assign n49283 = ~n24026 & n49282 ;
  assign n49284 = n8923 ^ n4530 ^ 1'b0 ;
  assign n49285 = ~n21993 & n49284 ;
  assign n49286 = ( n2098 & n41436 ) | ( n2098 & n49285 ) | ( n41436 & n49285 ) ;
  assign n49287 = n11558 ^ n7437 ^ n4726 ;
  assign n49288 = n6732 ^ n1391 ^ n1152 ;
  assign n49289 = ( n18592 & ~n49287 ) | ( n18592 & n49288 ) | ( ~n49287 & n49288 ) ;
  assign n49290 = n30348 ^ n29362 ^ n5385 ;
  assign n49291 = n3729 & ~n33294 ;
  assign n49292 = x222 & ~n28466 ;
  assign n49293 = ~n43483 & n49292 ;
  assign n49294 = n49293 ^ n38845 ^ n16845 ;
  assign n49295 = ( n26015 & n46428 ) | ( n26015 & n49294 ) | ( n46428 & n49294 ) ;
  assign n49297 = ( n9940 & ~n27636 ) | ( n9940 & n29428 ) | ( ~n27636 & n29428 ) ;
  assign n49296 = n12209 ^ n3754 ^ 1'b0 ;
  assign n49298 = n49297 ^ n49296 ^ n35509 ;
  assign n49299 = n24920 ^ n19119 ^ n19083 ;
  assign n49300 = n5032 | n49299 ;
  assign n49301 = n16720 & ~n49300 ;
  assign n49302 = n22198 & n40851 ;
  assign n49303 = ~n19139 & n49302 ;
  assign n49304 = n33138 ^ n24835 ^ 1'b0 ;
  assign n49305 = n41912 | n49304 ;
  assign n49306 = n49305 ^ n37048 ^ 1'b0 ;
  assign n49307 = ( n37349 & ~n41788 ) | ( n37349 & n49306 ) | ( ~n41788 & n49306 ) ;
  assign n49308 = ( n31065 & n48500 ) | ( n31065 & n49307 ) | ( n48500 & n49307 ) ;
  assign n49309 = ( ~n8726 & n13675 ) | ( ~n8726 & n21402 ) | ( n13675 & n21402 ) ;
  assign n49310 = n7641 ^ n2484 ^ 1'b0 ;
  assign n49311 = n6544 & n49310 ;
  assign n49313 = ~n14141 & n27589 ;
  assign n49314 = n49313 ^ n41136 ^ 1'b0 ;
  assign n49315 = ( n9151 & n31110 ) | ( n9151 & n49314 ) | ( n31110 & n49314 ) ;
  assign n49312 = n18829 & n22942 ;
  assign n49316 = n49315 ^ n49312 ^ 1'b0 ;
  assign n49317 = ( n5625 & ~n21875 ) | ( n5625 & n49316 ) | ( ~n21875 & n49316 ) ;
  assign n49318 = n10991 ^ n7254 ^ 1'b0 ;
  assign n49319 = n9361 | n49318 ;
  assign n49320 = n16002 & ~n49319 ;
  assign n49321 = n49320 ^ n43662 ^ 1'b0 ;
  assign n49322 = ~n11935 & n49321 ;
  assign n49323 = n21569 | n43481 ;
  assign n49324 = n2234 | n12741 ;
  assign n49325 = n4478 & ~n49324 ;
  assign n49326 = n26793 ^ n14231 ^ 1'b0 ;
  assign n49327 = n41485 | n49326 ;
  assign n49328 = ( n468 & n5146 ) | ( n468 & ~n31723 ) | ( n5146 & ~n31723 ) ;
  assign n49329 = x239 & ~n11330 ;
  assign n49330 = n49329 ^ n37401 ^ 1'b0 ;
  assign n49331 = n49330 ^ n49275 ^ n43569 ;
  assign n49332 = n8653 & ~n16250 ;
  assign n49333 = ~n9687 & n49332 ;
  assign n49334 = n49333 ^ n27350 ^ n9983 ;
  assign n49335 = ( n728 & n9383 ) | ( n728 & n21756 ) | ( n9383 & n21756 ) ;
  assign n49336 = n42179 & ~n49335 ;
  assign n49337 = ( n21541 & ~n49334 ) | ( n21541 & n49336 ) | ( ~n49334 & n49336 ) ;
  assign n49338 = ( n4707 & ~n12000 ) | ( n4707 & n17057 ) | ( ~n12000 & n17057 ) ;
  assign n49339 = n49338 ^ n10880 ^ n5983 ;
  assign n49340 = n43592 ^ n26122 ^ n18094 ;
  assign n49341 = n49340 ^ n41861 ^ n2181 ;
  assign n49342 = n39581 ^ n36951 ^ 1'b0 ;
  assign n49343 = n5737 & n49342 ;
  assign n49344 = n49343 ^ n27110 ^ n23429 ;
  assign n49345 = ( n6774 & n27520 ) | ( n6774 & ~n30659 ) | ( n27520 & ~n30659 ) ;
  assign n49346 = ( n1869 & ~n28786 ) | ( n1869 & n49345 ) | ( ~n28786 & n49345 ) ;
  assign n49347 = n34186 ^ n12095 ^ n6030 ;
  assign n49348 = n20481 & ~n49347 ;
  assign n49349 = ~n10853 & n49348 ;
  assign n49350 = n49349 ^ n47448 ^ n18769 ;
  assign n49351 = n440 & n2198 ;
  assign n49352 = n49351 ^ n11936 ^ 1'b0 ;
  assign n49353 = n39493 ^ n22869 ^ 1'b0 ;
  assign n49354 = n5844 & n49353 ;
  assign n49355 = ~n3315 & n49354 ;
  assign n49356 = n48187 & n49355 ;
  assign n49357 = n39797 & ~n49356 ;
  assign n49358 = ( ~n14934 & n17574 ) | ( ~n14934 & n23474 ) | ( n17574 & n23474 ) ;
  assign n49359 = n31223 ^ n10721 ^ n2934 ;
  assign n49360 = n49358 | n49359 ;
  assign n49361 = ( n13811 & ~n36681 ) | ( n13811 & n49024 ) | ( ~n36681 & n49024 ) ;
  assign n49364 = ( n13180 & ~n16758 ) | ( n13180 & n45018 ) | ( ~n16758 & n45018 ) ;
  assign n49362 = x158 & n3162 ;
  assign n49363 = n49362 ^ n42786 ^ n35361 ;
  assign n49365 = n49364 ^ n49363 ^ n9674 ;
  assign n49366 = n20408 & n39253 ;
  assign n49367 = ~n38615 & n49366 ;
  assign n49368 = ( n1637 & ~n16150 ) | ( n1637 & n23498 ) | ( ~n16150 & n23498 ) ;
  assign n49369 = ~n25573 & n37220 ;
  assign n49370 = ~n49368 & n49369 ;
  assign n49371 = n1519 & ~n5638 ;
  assign n49372 = ~n8216 & n49371 ;
  assign n49373 = ( n8284 & n10074 ) | ( n8284 & ~n49372 ) | ( n10074 & ~n49372 ) ;
  assign n49374 = n42504 & n49373 ;
  assign n49375 = n47211 & n49374 ;
  assign n49376 = n6379 ^ n1550 ^ 1'b0 ;
  assign n49377 = n49375 | n49376 ;
  assign n49378 = ( n12939 & n15140 ) | ( n12939 & n28356 ) | ( n15140 & n28356 ) ;
  assign n49379 = n37808 ^ n11775 ^ n10919 ;
  assign n49380 = ( n4627 & ~n21983 ) | ( n4627 & n49379 ) | ( ~n21983 & n49379 ) ;
  assign n49381 = n49380 ^ n16201 ^ x153 ;
  assign n49382 = ( n3980 & n5504 ) | ( n3980 & ~n19621 ) | ( n5504 & ~n19621 ) ;
  assign n49383 = n49382 ^ n47373 ^ n36470 ;
  assign n49384 = n26347 ^ n8659 ^ n2770 ;
  assign n49385 = ( n34842 & n46381 ) | ( n34842 & n49384 ) | ( n46381 & n49384 ) ;
  assign n49386 = ( ~n1602 & n2565 ) | ( ~n1602 & n9854 ) | ( n2565 & n9854 ) ;
  assign n49387 = n40532 | n49386 ;
  assign n49388 = n49387 ^ n44552 ^ 1'b0 ;
  assign n49389 = n33770 & n34762 ;
  assign n49390 = n49388 & n49389 ;
  assign n49391 = n49390 ^ n43870 ^ n7925 ;
  assign n49392 = n39366 ^ n27950 ^ n21289 ;
  assign n49393 = ( n13285 & ~n23018 ) | ( n13285 & n31892 ) | ( ~n23018 & n31892 ) ;
  assign n49394 = n49392 & ~n49393 ;
  assign n49395 = x102 & ~n21330 ;
  assign n49396 = n49395 ^ n12216 ^ 1'b0 ;
  assign n49397 = n3312 ^ n3303 ^ 1'b0 ;
  assign n49398 = n38652 | n49397 ;
  assign n49399 = n49398 ^ n26735 ^ n16359 ;
  assign n49400 = ( n8684 & n12940 ) | ( n8684 & n18041 ) | ( n12940 & n18041 ) ;
  assign n49401 = n49400 ^ n18452 ^ n6802 ;
  assign n49402 = n49401 ^ n48435 ^ n28593 ;
  assign n49403 = ( ~n21733 & n37421 ) | ( ~n21733 & n37568 ) | ( n37421 & n37568 ) ;
  assign n49404 = n49403 ^ n24536 ^ n17998 ;
  assign n49405 = ( n19370 & ~n46616 ) | ( n19370 & n49404 ) | ( ~n46616 & n49404 ) ;
  assign n49406 = ( ~n15036 & n47048 ) | ( ~n15036 & n49405 ) | ( n47048 & n49405 ) ;
  assign n49407 = ( ~n982 & n15537 ) | ( ~n982 & n16558 ) | ( n15537 & n16558 ) ;
  assign n49412 = n14007 ^ n13671 ^ n9369 ;
  assign n49408 = n49277 ^ n16701 ^ n786 ;
  assign n49409 = n49408 ^ n1561 ^ 1'b0 ;
  assign n49410 = n5887 | n49409 ;
  assign n49411 = n49410 ^ n26333 ^ 1'b0 ;
  assign n49413 = n49412 ^ n49411 ^ 1'b0 ;
  assign n49414 = ( n21772 & n24646 ) | ( n21772 & ~n39831 ) | ( n24646 & ~n39831 ) ;
  assign n49415 = n11324 ^ n10316 ^ n8909 ;
  assign n49416 = ( n5739 & ~n11004 ) | ( n5739 & n49415 ) | ( ~n11004 & n49415 ) ;
  assign n49417 = ~n18388 & n49416 ;
  assign n49418 = n3906 ^ n3515 ^ n2150 ;
  assign n49419 = n49418 ^ n31395 ^ 1'b0 ;
  assign n49420 = ~n16200 & n49419 ;
  assign n49421 = ~n49417 & n49420 ;
  assign n49422 = n45771 ^ n1471 ^ 1'b0 ;
  assign n49423 = n34666 ^ n8916 ^ 1'b0 ;
  assign n49424 = n15530 ^ n14365 ^ n13879 ;
  assign n49425 = n20421 | n49424 ;
  assign n49426 = n37419 ^ n12048 ^ 1'b0 ;
  assign n49427 = ~n9839 & n49426 ;
  assign n49428 = ( n7940 & ~n26610 ) | ( n7940 & n49427 ) | ( ~n26610 & n49427 ) ;
  assign n49429 = n48776 ^ n37566 ^ 1'b0 ;
  assign n49434 = n27243 ^ n3262 ^ n368 ;
  assign n49435 = ( n5815 & n16314 ) | ( n5815 & n49434 ) | ( n16314 & n49434 ) ;
  assign n49432 = ( n20565 & n34395 ) | ( n20565 & ~n38094 ) | ( n34395 & ~n38094 ) ;
  assign n49433 = n32705 | n49432 ;
  assign n49436 = n49435 ^ n49433 ^ 1'b0 ;
  assign n49430 = n15217 | n36818 ;
  assign n49431 = n49430 ^ n13217 ^ 1'b0 ;
  assign n49437 = n49436 ^ n49431 ^ n38187 ;
  assign n49438 = n48702 ^ n26748 ^ n20492 ;
  assign n49439 = n36356 ^ n14580 ^ 1'b0 ;
  assign n49440 = n37031 & n49439 ;
  assign n49441 = n49440 ^ n32674 ^ n25071 ;
  assign n49442 = ~n21605 & n44935 ;
  assign n49443 = n49442 ^ n33940 ^ 1'b0 ;
  assign n49444 = ( n11715 & n18840 ) | ( n11715 & ~n33525 ) | ( n18840 & ~n33525 ) ;
  assign n49445 = ~n28930 & n49444 ;
  assign n49446 = n49445 ^ n25158 ^ 1'b0 ;
  assign n49452 = ( n16559 & ~n24160 ) | ( n16559 & n43662 ) | ( ~n24160 & n43662 ) ;
  assign n49449 = ( ~n9069 & n28443 ) | ( ~n9069 & n38786 ) | ( n28443 & n38786 ) ;
  assign n49450 = n49449 ^ n37691 ^ n24187 ;
  assign n49448 = n20998 ^ n4539 ^ n4381 ;
  assign n49451 = n49450 ^ n49448 ^ n20762 ;
  assign n49447 = n33646 ^ n7115 ^ n5726 ;
  assign n49453 = n49452 ^ n49451 ^ n49447 ;
  assign n49454 = ( n13751 & n27671 ) | ( n13751 & n40464 ) | ( n27671 & n40464 ) ;
  assign n49455 = n19222 | n44310 ;
  assign n49456 = n14045 | n26896 ;
  assign n49457 = ( n12795 & ~n38466 ) | ( n12795 & n49456 ) | ( ~n38466 & n49456 ) ;
  assign n49462 = n3745 ^ n3441 ^ n1365 ;
  assign n49463 = ( n1192 & n31455 ) | ( n1192 & n49462 ) | ( n31455 & n49462 ) ;
  assign n49459 = n29086 ^ n13335 ^ n7182 ;
  assign n49460 = ( ~n2964 & n6314 ) | ( ~n2964 & n49459 ) | ( n6314 & n49459 ) ;
  assign n49458 = ( n13564 & ~n22035 ) | ( n13564 & n22467 ) | ( ~n22035 & n22467 ) ;
  assign n49461 = n49460 ^ n49458 ^ n4487 ;
  assign n49464 = n49463 ^ n49461 ^ 1'b0 ;
  assign n49465 = ~n21756 & n35755 ;
  assign n49466 = n49465 ^ n48794 ^ n36425 ;
  assign n49468 = n6398 & n42895 ;
  assign n49469 = n10154 & n49468 ;
  assign n49467 = ( n10431 & n32664 ) | ( n10431 & ~n41809 ) | ( n32664 & ~n41809 ) ;
  assign n49470 = n49469 ^ n49467 ^ n42260 ;
  assign n49471 = n4567 | n24546 ;
  assign n49472 = ~n3454 & n13736 ;
  assign n49473 = n49471 & n49472 ;
  assign n49474 = n35595 ^ n13236 ^ 1'b0 ;
  assign n49475 = ~n22556 & n49474 ;
  assign n49476 = n6239 & n14339 ;
  assign n49477 = n37969 & n49476 ;
  assign n49478 = n42453 ^ n27240 ^ 1'b0 ;
  assign n49479 = n22824 & ~n49478 ;
  assign n49480 = ( ~n7629 & n30742 ) | ( ~n7629 & n49479 ) | ( n30742 & n49479 ) ;
  assign n49481 = n32072 ^ n5887 ^ 1'b0 ;
  assign n49482 = n49480 | n49481 ;
  assign n49483 = ( ~n1491 & n19833 ) | ( ~n1491 & n26171 ) | ( n19833 & n26171 ) ;
  assign n49484 = n28941 & ~n49483 ;
  assign n49485 = n49484 ^ n446 ^ 1'b0 ;
  assign n49486 = n49485 ^ n22198 ^ n7286 ;
  assign n49487 = n2863 & n18186 ;
  assign n49488 = n49487 ^ n6243 ^ 1'b0 ;
  assign n49489 = n12292 ^ n8552 ^ n6512 ;
  assign n49490 = ( ~n24232 & n49488 ) | ( ~n24232 & n49489 ) | ( n49488 & n49489 ) ;
  assign n49494 = n48896 ^ n21572 ^ n17853 ;
  assign n49492 = n23926 ^ n3043 ^ 1'b0 ;
  assign n49493 = n21957 | n49492 ;
  assign n49491 = n3308 & n34686 ;
  assign n49495 = n49494 ^ n49493 ^ n49491 ;
  assign n49496 = n32367 ^ n30328 ^ n12666 ;
  assign n49497 = n3498 & n49496 ;
  assign n49498 = ( n2203 & n14016 ) | ( n2203 & n40933 ) | ( n14016 & n40933 ) ;
  assign n49499 = n9276 ^ n8174 ^ 1'b0 ;
  assign n49500 = n3522 & n49499 ;
  assign n49501 = n49500 ^ n39515 ^ n6422 ;
  assign n49502 = n5231 ^ n1312 ^ 1'b0 ;
  assign n49503 = n16834 & n37009 ;
  assign n49504 = n49503 ^ n42213 ^ 1'b0 ;
  assign n49509 = n37616 ^ n27862 ^ 1'b0 ;
  assign n49510 = n4835 | n49509 ;
  assign n49505 = ( n555 & n2920 ) | ( n555 & n5110 ) | ( n2920 & n5110 ) ;
  assign n49506 = n21149 ^ n12689 ^ n12181 ;
  assign n49507 = n49506 ^ n16291 ^ 1'b0 ;
  assign n49508 = n49505 & n49507 ;
  assign n49511 = n49510 ^ n49508 ^ n42609 ;
  assign n49512 = ( n9571 & n10030 ) | ( n9571 & n14779 ) | ( n10030 & n14779 ) ;
  assign n49513 = n32010 ^ n23679 ^ n14195 ;
  assign n49514 = ( n30012 & n49512 ) | ( n30012 & ~n49513 ) | ( n49512 & ~n49513 ) ;
  assign n49515 = n8265 ^ x148 ^ x99 ;
  assign n49516 = ~n47483 & n49515 ;
  assign n49517 = ( n12551 & n16897 ) | ( n12551 & n19321 ) | ( n16897 & n19321 ) ;
  assign n49518 = ( n9963 & n47620 ) | ( n9963 & n49517 ) | ( n47620 & n49517 ) ;
  assign n49522 = ( n8455 & n31957 ) | ( n8455 & ~n35092 ) | ( n31957 & ~n35092 ) ;
  assign n49519 = x142 & n568 ;
  assign n49520 = n49519 ^ n1631 ^ 1'b0 ;
  assign n49521 = n49520 ^ n29806 ^ n18126 ;
  assign n49523 = n49522 ^ n49521 ^ n17307 ;
  assign n49524 = n47064 ^ n28025 ^ n8728 ;
  assign n49526 = ( n13991 & n17276 ) | ( n13991 & ~n27553 ) | ( n17276 & ~n27553 ) ;
  assign n49525 = n15663 & ~n17519 ;
  assign n49527 = n49526 ^ n49525 ^ 1'b0 ;
  assign n49528 = n42531 & ~n45025 ;
  assign n49529 = n49528 ^ n7270 ^ 1'b0 ;
  assign n49530 = n7780 & ~n35283 ;
  assign n49531 = n38025 ^ n19064 ^ n4531 ;
  assign n49532 = ( n27764 & ~n47405 ) | ( n27764 & n49531 ) | ( ~n47405 & n49531 ) ;
  assign n49533 = ( n21325 & n29596 ) | ( n21325 & n44735 ) | ( n29596 & n44735 ) ;
  assign n49534 = n32084 ^ n8679 ^ n6947 ;
  assign n49535 = n31930 ^ n13438 ^ n10925 ;
  assign n49536 = n2438 & ~n35938 ;
  assign n49537 = n49536 ^ n20283 ^ 1'b0 ;
  assign n49538 = n49537 ^ n26751 ^ 1'b0 ;
  assign n49539 = n10174 & n20753 ;
  assign n49540 = n49539 ^ n40687 ^ 1'b0 ;
  assign n49541 = n4557 | n6441 ;
  assign n49542 = n49541 ^ n16598 ^ 1'b0 ;
  assign n49543 = n13466 ^ n9649 ^ 1'b0 ;
  assign n49544 = n5920 & ~n49543 ;
  assign n49545 = ( n2964 & n21007 ) | ( n2964 & n36682 ) | ( n21007 & n36682 ) ;
  assign n49546 = ( ~n14707 & n19005 ) | ( ~n14707 & n35973 ) | ( n19005 & n35973 ) ;
  assign n49547 = n49546 ^ n44535 ^ n43216 ;
  assign n49548 = n6765 | n12833 ;
  assign n49549 = n680 & ~n49548 ;
  assign n49550 = n49549 ^ n25536 ^ n11250 ;
  assign n49551 = ( n2926 & n4630 ) | ( n2926 & n22630 ) | ( n4630 & n22630 ) ;
  assign n49552 = n49551 ^ n32729 ^ 1'b0 ;
  assign n49553 = ( n16251 & n34205 ) | ( n16251 & n49552 ) | ( n34205 & n49552 ) ;
  assign n49554 = n30383 ^ n23479 ^ n10059 ;
  assign n49555 = n49554 ^ n26936 ^ n8584 ;
  assign n49556 = ( n6373 & n25897 ) | ( n6373 & n49555 ) | ( n25897 & n49555 ) ;
  assign n49557 = n35927 ^ n32264 ^ n17697 ;
  assign n49558 = ( ~n11934 & n27133 ) | ( ~n11934 & n49557 ) | ( n27133 & n49557 ) ;
  assign n49559 = ( ~n2160 & n20113 ) | ( ~n2160 & n24070 ) | ( n20113 & n24070 ) ;
  assign n49560 = ( n2192 & n17409 ) | ( n2192 & ~n49559 ) | ( n17409 & ~n49559 ) ;
  assign n49561 = ( n20428 & n29426 ) | ( n20428 & ~n48984 ) | ( n29426 & ~n48984 ) ;
  assign n49562 = n30105 & ~n49561 ;
  assign n49563 = n49562 ^ n7888 ^ 1'b0 ;
  assign n49564 = n1677 & ~n9634 ;
  assign n49565 = n26695 & n49564 ;
  assign n49566 = ( n2976 & ~n20444 ) | ( n2976 & n36066 ) | ( ~n20444 & n36066 ) ;
  assign n49567 = ( ~n27750 & n49565 ) | ( ~n27750 & n49566 ) | ( n49565 & n49566 ) ;
  assign n49568 = n28387 & n49567 ;
  assign n49569 = n49568 ^ n18837 ^ 1'b0 ;
  assign n49570 = n45455 ^ n29356 ^ n17955 ;
  assign n49572 = n37644 ^ n21389 ^ n10807 ;
  assign n49571 = ( n2800 & ~n7493 ) | ( n2800 & n31097 ) | ( ~n7493 & n31097 ) ;
  assign n49573 = n49572 ^ n49571 ^ n11065 ;
  assign n49574 = n3017 & n10985 ;
  assign n49575 = ( ~n8963 & n18685 ) | ( ~n8963 & n49505 ) | ( n18685 & n49505 ) ;
  assign n49576 = ~n49574 & n49575 ;
  assign n49577 = n49576 ^ n2993 ^ 1'b0 ;
  assign n49578 = ( ~n12416 & n26745 ) | ( ~n12416 & n49577 ) | ( n26745 & n49577 ) ;
  assign n49579 = n49578 ^ n29271 ^ n2613 ;
  assign n49580 = n2234 & n4260 ;
  assign n49581 = n49580 ^ n17936 ^ n15808 ;
  assign n49582 = n16759 | n35659 ;
  assign n49583 = ( n13787 & n18921 ) | ( n13787 & ~n49582 ) | ( n18921 & ~n49582 ) ;
  assign n49587 = n18661 ^ n10211 ^ 1'b0 ;
  assign n49588 = n9771 & n49587 ;
  assign n49589 = n49588 ^ n15300 ^ n12898 ;
  assign n49590 = n49589 ^ n29436 ^ n3430 ;
  assign n49584 = ( ~n4627 & n22402 ) | ( ~n4627 & n26856 ) | ( n22402 & n26856 ) ;
  assign n49585 = n15184 & n49584 ;
  assign n49586 = ~n21950 & n49585 ;
  assign n49591 = n49590 ^ n49586 ^ n17680 ;
  assign n49592 = ~n7479 & n12968 ;
  assign n49593 = ~x28 & n49592 ;
  assign n49594 = n1198 & ~n2701 ;
  assign n49595 = n49594 ^ n24333 ^ 1'b0 ;
  assign n49599 = n33365 ^ n9820 ^ 1'b0 ;
  assign n49600 = n13362 & n49599 ;
  assign n49596 = n32978 ^ n12481 ^ n5403 ;
  assign n49597 = n49596 ^ n14545 ^ n8625 ;
  assign n49598 = n49597 ^ n44916 ^ n8275 ;
  assign n49601 = n49600 ^ n49598 ^ n13077 ;
  assign n49602 = ~n32299 & n49601 ;
  assign n49603 = n45389 & n49602 ;
  assign n49604 = n47421 ^ n43635 ^ n37088 ;
  assign n49605 = n10309 & n20408 ;
  assign n49606 = ~n8760 & n49605 ;
  assign n49607 = n47772 ^ n35956 ^ 1'b0 ;
  assign n49608 = n49607 ^ n33834 ^ n28691 ;
  assign n49609 = n49606 | n49608 ;
  assign n49610 = n6675 ^ n6523 ^ n1315 ;
  assign n49611 = ( n382 & n43086 ) | ( n382 & n49610 ) | ( n43086 & n49610 ) ;
  assign n49612 = n49611 ^ n38864 ^ n23295 ;
  assign n49613 = n12243 ^ n8037 ^ n1998 ;
  assign n49614 = ( n1756 & n38536 ) | ( n1756 & n49613 ) | ( n38536 & n49613 ) ;
  assign n49615 = ( n26447 & n28129 ) | ( n26447 & ~n46935 ) | ( n28129 & ~n46935 ) ;
  assign n49616 = ~n8673 & n10527 ;
  assign n49617 = ( n19109 & n25772 ) | ( n19109 & ~n33690 ) | ( n25772 & ~n33690 ) ;
  assign n49618 = n44710 ^ n15194 ^ 1'b0 ;
  assign n49619 = ~n49617 & n49618 ;
  assign n49620 = n41154 ^ n25867 ^ 1'b0 ;
  assign n49621 = ( n21855 & ~n29248 ) | ( n21855 & n46105 ) | ( ~n29248 & n46105 ) ;
  assign n49622 = n45245 ^ n30874 ^ n8469 ;
  assign n49623 = n28837 ^ n14552 ^ 1'b0 ;
  assign n49624 = ( n5542 & ~n37249 ) | ( n5542 & n40930 ) | ( ~n37249 & n40930 ) ;
  assign n49625 = n49624 ^ n29901 ^ n6548 ;
  assign n49626 = ( n1116 & ~n32743 ) | ( n1116 & n38211 ) | ( ~n32743 & n38211 ) ;
  assign n49627 = n14800 & n22178 ;
  assign n49628 = n23541 & n49627 ;
  assign n49629 = n49628 ^ n1129 ^ 1'b0 ;
  assign n49630 = n12141 | n23783 ;
  assign n49631 = ~n538 & n18374 ;
  assign n49632 = ( n904 & ~n13522 ) | ( n904 & n45716 ) | ( ~n13522 & n45716 ) ;
  assign n49633 = ( n2841 & ~n14304 ) | ( n2841 & n14749 ) | ( ~n14304 & n14749 ) ;
  assign n49634 = n14914 & ~n49633 ;
  assign n49635 = n49632 & n49634 ;
  assign n49636 = n24199 ^ n15171 ^ n12486 ;
  assign n49637 = n49636 ^ n3943 ^ 1'b0 ;
  assign n49638 = n45668 | n49637 ;
  assign n49639 = n21825 & ~n49638 ;
  assign n49640 = n42581 ^ n34188 ^ n15678 ;
  assign n49641 = ( ~n19036 & n34884 ) | ( ~n19036 & n49640 ) | ( n34884 & n49640 ) ;
  assign n49642 = n13150 | n43009 ;
  assign n49643 = n19869 ^ n8351 ^ 1'b0 ;
  assign n49644 = n20276 ^ n13664 ^ n3039 ;
  assign n49645 = ( ~n4855 & n33017 ) | ( ~n4855 & n49644 ) | ( n33017 & n49644 ) ;
  assign n49646 = n8929 ^ n1915 ^ 1'b0 ;
  assign n49647 = n8799 | n49646 ;
  assign n49648 = n34474 ^ n14595 ^ n456 ;
  assign n49649 = ( n9293 & n10403 ) | ( n9293 & ~n13536 ) | ( n10403 & ~n13536 ) ;
  assign n49650 = n49649 ^ n37042 ^ n17867 ;
  assign n49651 = n49650 ^ n11687 ^ 1'b0 ;
  assign n49652 = n15664 ^ n9972 ^ 1'b0 ;
  assign n49653 = n49652 ^ n1130 ^ 1'b0 ;
  assign n49654 = ( ~n16372 & n23293 ) | ( ~n16372 & n49653 ) | ( n23293 & n49653 ) ;
  assign n49655 = n12848 ^ n6509 ^ 1'b0 ;
  assign n49656 = n49655 ^ n14275 ^ n2955 ;
  assign n49657 = n4713 & ~n6031 ;
  assign n49658 = ~n24573 & n49657 ;
  assign n49659 = ( n10735 & n40760 ) | ( n10735 & ~n49658 ) | ( n40760 & ~n49658 ) ;
  assign n49660 = n49659 ^ n2105 ^ 1'b0 ;
  assign n49661 = n7429 | n16595 ;
  assign n49662 = ( n10861 & n24572 ) | ( n10861 & ~n49661 ) | ( n24572 & ~n49661 ) ;
  assign n49663 = ( ~n2022 & n3777 ) | ( ~n2022 & n49662 ) | ( n3777 & n49662 ) ;
  assign n49665 = n3748 | n20641 ;
  assign n49664 = ( n10800 & ~n12401 ) | ( n10800 & n19402 ) | ( ~n12401 & n19402 ) ;
  assign n49666 = n49665 ^ n49664 ^ 1'b0 ;
  assign n49670 = ( n9082 & ~n10711 ) | ( n9082 & n29958 ) | ( ~n10711 & n29958 ) ;
  assign n49667 = n47142 ^ n41969 ^ n12071 ;
  assign n49668 = n12617 ^ n3353 ^ 1'b0 ;
  assign n49669 = n49667 | n49668 ;
  assign n49671 = n49670 ^ n49669 ^ n48932 ;
  assign n49672 = ( n3676 & ~n25756 ) | ( n3676 & n41195 ) | ( ~n25756 & n41195 ) ;
  assign n49673 = n49672 ^ n9533 ^ n7687 ;
  assign n49674 = n31261 ^ n1257 ^ 1'b0 ;
  assign n49675 = n13762 & ~n49674 ;
  assign n49676 = ( n16714 & n22785 ) | ( n16714 & n36369 ) | ( n22785 & n36369 ) ;
  assign n49677 = n49676 ^ n20135 ^ n19654 ;
  assign n49678 = n38762 ^ n32679 ^ n26241 ;
  assign n49679 = n49677 & n49678 ;
  assign n49680 = ( n21458 & n36919 ) | ( n21458 & ~n39648 ) | ( n36919 & ~n39648 ) ;
  assign n49681 = n16709 ^ n12764 ^ 1'b0 ;
  assign n49682 = n49680 & n49681 ;
  assign n49686 = n14702 ^ n14098 ^ n11660 ;
  assign n49683 = n28037 ^ n3361 ^ 1'b0 ;
  assign n49684 = n16681 & n49683 ;
  assign n49685 = ( n31512 & n33804 ) | ( n31512 & n49684 ) | ( n33804 & n49684 ) ;
  assign n49687 = n49686 ^ n49685 ^ n23301 ;
  assign n49689 = n41823 ^ n8745 ^ n3697 ;
  assign n49690 = n49689 ^ n37661 ^ 1'b0 ;
  assign n49688 = ( n17430 & ~n20322 ) | ( n17430 & n34545 ) | ( ~n20322 & n34545 ) ;
  assign n49691 = n49690 ^ n49688 ^ n41378 ;
  assign n49692 = ~n39116 & n49691 ;
  assign n49693 = ( ~n20899 & n49687 ) | ( ~n20899 & n49692 ) | ( n49687 & n49692 ) ;
  assign n49694 = n13573 & n32079 ;
  assign n49695 = ( n10007 & ~n17154 ) | ( n10007 & n32235 ) | ( ~n17154 & n32235 ) ;
  assign n49697 = n16976 ^ n16722 ^ 1'b0 ;
  assign n49696 = n2268 & n14183 ;
  assign n49698 = n49697 ^ n49696 ^ 1'b0 ;
  assign n49699 = n49698 ^ n40581 ^ n9589 ;
  assign n49700 = n2638 & ~n49699 ;
  assign n49701 = ( n4230 & n32001 ) | ( n4230 & ~n49700 ) | ( n32001 & ~n49700 ) ;
  assign n49702 = n22724 ^ n9866 ^ 1'b0 ;
  assign n49703 = ( n19303 & ~n42497 ) | ( n19303 & n49702 ) | ( ~n42497 & n49702 ) ;
  assign n49704 = n49703 ^ n33896 ^ n21137 ;
  assign n49705 = n49704 ^ n25936 ^ n3753 ;
  assign n49706 = n37607 ^ n31049 ^ n26034 ;
  assign n49707 = n2144 & n14291 ;
  assign n49708 = ~n13452 & n49707 ;
  assign n49709 = n49708 ^ n27855 ^ 1'b0 ;
  assign n49710 = n27614 ^ n7429 ^ n5346 ;
  assign n49711 = ~n1562 & n27926 ;
  assign n49712 = n49710 & n49711 ;
  assign n49713 = n49712 ^ n19938 ^ 1'b0 ;
  assign n49714 = ( n17682 & ~n23124 ) | ( n17682 & n28857 ) | ( ~n23124 & n28857 ) ;
  assign n49715 = n49714 ^ n41740 ^ 1'b0 ;
  assign n49716 = n49713 & ~n49715 ;
  assign n49717 = ~n29820 & n39253 ;
  assign n49718 = n2058 & n49717 ;
  assign n49719 = n29165 & n37123 ;
  assign n49720 = n49719 ^ n39066 ^ 1'b0 ;
  assign n49721 = ( ~n29858 & n42583 ) | ( ~n29858 & n49720 ) | ( n42583 & n49720 ) ;
  assign n49722 = n11688 ^ n9857 ^ 1'b0 ;
  assign n49723 = ~n5295 & n49722 ;
  assign n49724 = n49723 ^ n47417 ^ 1'b0 ;
  assign n49725 = n28465 & n45212 ;
  assign n49726 = n34642 | n35563 ;
  assign n49727 = n23197 | n49726 ;
  assign n49728 = n49727 ^ n26132 ^ 1'b0 ;
  assign n49729 = n33001 ^ n8558 ^ n7116 ;
  assign n49730 = x144 & ~n12191 ;
  assign n49731 = n49730 ^ n11120 ^ 1'b0 ;
  assign n49732 = ( n2379 & n2413 ) | ( n2379 & ~n23183 ) | ( n2413 & ~n23183 ) ;
  assign n49733 = n49732 ^ n27175 ^ n13518 ;
  assign n49734 = n49733 ^ n28494 ^ n16694 ;
  assign n49735 = n49734 ^ n31510 ^ n22673 ;
  assign n49736 = n8806 & ~n49735 ;
  assign n49737 = n40786 ^ n29214 ^ n3120 ;
  assign n49738 = ( ~n22448 & n33758 ) | ( ~n22448 & n37624 ) | ( n33758 & n37624 ) ;
  assign n49739 = ~n22509 & n39196 ;
  assign n49740 = ~n8675 & n27279 ;
  assign n49741 = n32138 ^ n30003 ^ 1'b0 ;
  assign n49742 = n28580 & ~n49741 ;
  assign n49743 = n49742 ^ n24346 ^ n19108 ;
  assign n49744 = n12718 & n17490 ;
  assign n49745 = n19563 ^ n11072 ^ n7760 ;
  assign n49746 = ( ~n3784 & n8344 ) | ( ~n3784 & n24483 ) | ( n8344 & n24483 ) ;
  assign n49747 = n18875 | n49746 ;
  assign n49748 = ( n9716 & n15343 ) | ( n9716 & n49747 ) | ( n15343 & n49747 ) ;
  assign n49749 = ( n27099 & n49745 ) | ( n27099 & ~n49748 ) | ( n49745 & ~n49748 ) ;
  assign n49750 = n7760 | n24267 ;
  assign n49751 = n49134 ^ n25394 ^ 1'b0 ;
  assign n49752 = n49750 | n49751 ;
  assign n49753 = n42789 ^ n7050 ^ n1466 ;
  assign n49754 = n1402 | n18390 ;
  assign n49755 = n49753 & ~n49754 ;
  assign n49756 = n45085 ^ n3609 ^ 1'b0 ;
  assign n49757 = ~n48381 & n49756 ;
  assign n49758 = n38326 ^ n20603 ^ n6511 ;
  assign n49759 = n48671 ^ n15278 ^ n14561 ;
  assign n49760 = ( n5910 & n35184 ) | ( n5910 & n37587 ) | ( n35184 & n37587 ) ;
  assign n49761 = ( n36371 & ~n45020 ) | ( n36371 & n49760 ) | ( ~n45020 & n49760 ) ;
  assign n49763 = n40198 ^ n9247 ^ 1'b0 ;
  assign n49764 = ~n13631 & n49763 ;
  assign n49765 = ~n22162 & n49764 ;
  assign n49762 = n29756 ^ n27945 ^ n13711 ;
  assign n49766 = n49765 ^ n49762 ^ n38490 ;
  assign n49767 = n19867 & ~n21532 ;
  assign n49768 = n49767 ^ n29086 ^ 1'b0 ;
  assign n49769 = ( n22536 & n24665 ) | ( n22536 & n36946 ) | ( n24665 & n36946 ) ;
  assign n49770 = n8897 | n49769 ;
  assign n49771 = n49768 | n49770 ;
  assign n49773 = n41605 | n42072 ;
  assign n49774 = n28403 | n49773 ;
  assign n49775 = ~n29631 & n49774 ;
  assign n49772 = n20409 & n35880 ;
  assign n49776 = n49775 ^ n49772 ^ 1'b0 ;
  assign n49777 = ~n11317 & n16640 ;
  assign n49778 = ~n6244 & n49777 ;
  assign n49779 = n15321 & n49778 ;
  assign n49780 = n49779 ^ n1408 ^ 1'b0 ;
  assign n49781 = n7338 | n31396 ;
  assign n49782 = n31602 | n49781 ;
  assign n49783 = n24779 ^ n15905 ^ n5689 ;
  assign n49784 = ( n11269 & ~n49782 ) | ( n11269 & n49783 ) | ( ~n49782 & n49783 ) ;
  assign n49785 = n45050 ^ n13923 ^ n6364 ;
  assign n49786 = n49785 ^ n25192 ^ 1'b0 ;
  assign n49787 = n35561 ^ n4824 ^ 1'b0 ;
  assign n49788 = n5575 | n10831 ;
  assign n49789 = ( n21872 & ~n29319 ) | ( n21872 & n30378 ) | ( ~n29319 & n30378 ) ;
  assign n49790 = ~n28039 & n49789 ;
  assign n49791 = n47918 ^ n29872 ^ n6609 ;
  assign n49792 = n49791 ^ n49246 ^ n13136 ;
  assign n49793 = n27099 ^ n10662 ^ 1'b0 ;
  assign n49794 = n20663 | n49793 ;
  assign n49795 = n49794 ^ n30249 ^ 1'b0 ;
  assign n49796 = ( n14349 & ~n20132 ) | ( n14349 & n49795 ) | ( ~n20132 & n49795 ) ;
  assign n49797 = n15376 & ~n27463 ;
  assign n49798 = n47144 ^ n45963 ^ 1'b0 ;
  assign n49799 = n10611 | n13554 ;
  assign n49800 = n20006 ^ n3143 ^ 1'b0 ;
  assign n49801 = ( n17727 & n49799 ) | ( n17727 & ~n49800 ) | ( n49799 & ~n49800 ) ;
  assign n49802 = ~n8739 & n15893 ;
  assign n49803 = n34121 ^ n31400 ^ n5873 ;
  assign n49805 = n19979 ^ n11833 ^ n3200 ;
  assign n49804 = n40066 | n42143 ;
  assign n49806 = n49805 ^ n49804 ^ 1'b0 ;
  assign n49807 = n3291 | n22012 ;
  assign n49808 = n11933 ^ n6114 ^ 1'b0 ;
  assign n49809 = n18677 ^ n12728 ^ 1'b0 ;
  assign n49810 = n32232 | n49809 ;
  assign n49812 = ( n9582 & n12190 ) | ( n9582 & ~n26219 ) | ( n12190 & ~n26219 ) ;
  assign n49811 = n16270 & n29846 ;
  assign n49813 = n49812 ^ n49811 ^ 1'b0 ;
  assign n49814 = n21162 ^ n9261 ^ n631 ;
  assign n49815 = n49814 ^ n2373 ^ 1'b0 ;
  assign n49816 = ~n19828 & n49815 ;
  assign n49817 = n49816 ^ n9930 ^ n7339 ;
  assign n49818 = n36840 ^ n25459 ^ n22687 ;
  assign n49822 = ( n1561 & n7366 ) | ( n1561 & n38455 ) | ( n7366 & n38455 ) ;
  assign n49819 = n5663 | n36454 ;
  assign n49820 = n25483 ^ n8870 ^ 1'b0 ;
  assign n49821 = n49819 & n49820 ;
  assign n49823 = n49822 ^ n49821 ^ n5599 ;
  assign n49824 = n45114 & ~n49823 ;
  assign n49826 = n5774 ^ n5214 ^ 1'b0 ;
  assign n49825 = n8717 & ~n37686 ;
  assign n49827 = n49826 ^ n49825 ^ 1'b0 ;
  assign n49828 = n28729 ^ n12132 ^ n6019 ;
  assign n49829 = n39688 ^ n37212 ^ n28997 ;
  assign n49830 = n21974 & ~n49829 ;
  assign n49831 = ( n8134 & n23409 ) | ( n8134 & ~n49830 ) | ( n23409 & ~n49830 ) ;
  assign n49832 = ( n25960 & n27951 ) | ( n25960 & ~n34369 ) | ( n27951 & ~n34369 ) ;
  assign n49834 = n18155 | n42788 ;
  assign n49833 = ~n13517 & n18166 ;
  assign n49835 = n49834 ^ n49833 ^ 1'b0 ;
  assign n49836 = ~n16110 & n18280 ;
  assign n49837 = n16527 | n17465 ;
  assign n49838 = n43051 & ~n49837 ;
  assign n49839 = ( n23051 & n49836 ) | ( n23051 & ~n49838 ) | ( n49836 & ~n49838 ) ;
  assign n49840 = n43670 & ~n49839 ;
  assign n49841 = n49840 ^ n3557 ^ 1'b0 ;
  assign n49842 = ( ~n22348 & n24666 ) | ( ~n22348 & n27924 ) | ( n24666 & n27924 ) ;
  assign n49843 = n31839 ^ n15112 ^ n1809 ;
  assign n49844 = n15309 ^ n2367 ^ n1596 ;
  assign n49845 = n49844 ^ n21233 ^ n16252 ;
  assign n49846 = ~n49843 & n49845 ;
  assign n49847 = n29373 & ~n45677 ;
  assign n49848 = n23636 & n49847 ;
  assign n49849 = n49848 ^ n36444 ^ 1'b0 ;
  assign n49850 = n16954 ^ n1605 ^ 1'b0 ;
  assign n49851 = n22125 & ~n49850 ;
  assign n49852 = n49851 ^ n15502 ^ n10344 ;
  assign n49853 = ~n525 & n18395 ;
  assign n49854 = n7889 & ~n25488 ;
  assign n49855 = ( n10387 & ~n27378 ) | ( n10387 & n35483 ) | ( ~n27378 & n35483 ) ;
  assign n49856 = n7345 | n12486 ;
  assign n49857 = n49856 ^ n22296 ^ 1'b0 ;
  assign n49858 = n39144 ^ n9486 ^ n4983 ;
  assign n49859 = ( ~n15979 & n18752 ) | ( ~n15979 & n49858 ) | ( n18752 & n49858 ) ;
  assign n49860 = n49859 ^ n17776 ^ n9616 ;
  assign n49861 = n15022 | n19617 ;
  assign n49862 = n49860 & ~n49861 ;
  assign n49864 = n36871 ^ n13104 ^ n1130 ;
  assign n49863 = n26249 | n34669 ;
  assign n49865 = n49864 ^ n49863 ^ 1'b0 ;
  assign n49866 = n31071 | n33605 ;
  assign n49867 = n17878 & ~n49866 ;
  assign n49869 = n28707 ^ n7665 ^ 1'b0 ;
  assign n49870 = ~n24502 & n49869 ;
  assign n49868 = n825 & ~n47917 ;
  assign n49871 = n49870 ^ n49868 ^ 1'b0 ;
  assign n49872 = ( n19425 & n33619 ) | ( n19425 & n49871 ) | ( n33619 & n49871 ) ;
  assign n49873 = ~n20789 & n22012 ;
  assign n49874 = n49873 ^ n16782 ^ 1'b0 ;
  assign n49875 = n49874 ^ n26349 ^ n24086 ;
  assign n49876 = n3251 & n18643 ;
  assign n49877 = ~n11816 & n49876 ;
  assign n49878 = n49877 ^ n5406 ^ 1'b0 ;
  assign n49880 = ~n1504 & n30775 ;
  assign n49879 = n24903 ^ n14589 ^ 1'b0 ;
  assign n49881 = n49880 ^ n49879 ^ n13635 ;
  assign n49882 = n49881 ^ n36934 ^ n30654 ;
  assign n49883 = n5712 | n27996 ;
  assign n49884 = n49883 ^ n16733 ^ 1'b0 ;
  assign n49885 = ( n6724 & n28478 ) | ( n6724 & ~n49884 ) | ( n28478 & ~n49884 ) ;
  assign n49886 = n18269 & ~n43213 ;
  assign n49887 = ~n2764 & n49886 ;
  assign n49888 = n653 & ~n3111 ;
  assign n49889 = n44336 & n49888 ;
  assign n49890 = n38664 ^ n17486 ^ 1'b0 ;
  assign n49891 = ( n13048 & ~n14834 ) | ( n13048 & n30535 ) | ( ~n14834 & n30535 ) ;
  assign n49892 = n5232 & ~n41746 ;
  assign n49893 = ( n42607 & n49891 ) | ( n42607 & n49892 ) | ( n49891 & n49892 ) ;
  assign n49894 = n2620 & n12358 ;
  assign n49895 = ~n40615 & n49894 ;
  assign n49896 = n49895 ^ n33799 ^ n26097 ;
  assign n49897 = n31643 ^ n15992 ^ n12249 ;
  assign n49898 = ( n13811 & ~n30602 ) | ( n13811 & n49897 ) | ( ~n30602 & n49897 ) ;
  assign n49899 = n21281 ^ n18237 ^ n15049 ;
  assign n49900 = ( n27799 & n27954 ) | ( n27799 & ~n49899 ) | ( n27954 & ~n49899 ) ;
  assign n49901 = ~n18633 & n24716 ;
  assign n49902 = n49901 ^ n9252 ^ 1'b0 ;
  assign n49903 = n28022 & n49902 ;
  assign n49904 = n17978 & n18467 ;
  assign n49905 = ~n20435 & n49904 ;
  assign n49906 = n9785 ^ n1223 ^ 1'b0 ;
  assign n49907 = n9389 & ~n49906 ;
  assign n49908 = n12166 ^ n8438 ^ n6063 ;
  assign n49909 = n49908 ^ n41282 ^ n11065 ;
  assign n49910 = n49909 ^ n17570 ^ n16474 ;
  assign n49911 = n11558 & n38626 ;
  assign n49912 = n49911 ^ n16371 ^ 1'b0 ;
  assign n49913 = ( n18565 & n49821 ) | ( n18565 & ~n49912 ) | ( n49821 & ~n49912 ) ;
  assign n49914 = n12569 & ~n44262 ;
  assign n49915 = n30616 & n49914 ;
  assign n49916 = ( ~n42255 & n49913 ) | ( ~n42255 & n49915 ) | ( n49913 & n49915 ) ;
  assign n49920 = ( n14314 & ~n14455 ) | ( n14314 & n18511 ) | ( ~n14455 & n18511 ) ;
  assign n49921 = n49920 ^ n22023 ^ n16818 ;
  assign n49917 = n20026 ^ n14077 ^ 1'b0 ;
  assign n49918 = x103 & n49917 ;
  assign n49919 = ( ~n22264 & n28005 ) | ( ~n22264 & n49918 ) | ( n28005 & n49918 ) ;
  assign n49922 = n49921 ^ n49919 ^ n1527 ;
  assign n49923 = ~n44781 & n46944 ;
  assign n49924 = n33651 & ~n48221 ;
  assign n49925 = n7251 & n49924 ;
  assign n49926 = n49925 ^ n36442 ^ n14324 ;
  assign n49927 = n49926 ^ n40812 ^ 1'b0 ;
  assign n49928 = n49927 ^ n17035 ^ n15429 ;
  assign n49929 = n2710 | n29842 ;
  assign n49930 = n49929 ^ n11597 ^ 1'b0 ;
  assign n49931 = ( n27251 & n33276 ) | ( n27251 & n49930 ) | ( n33276 & n49930 ) ;
  assign n49932 = n30477 ^ n883 ^ 1'b0 ;
  assign n49933 = n29655 ^ n18529 ^ 1'b0 ;
  assign n49934 = n37579 ^ n18134 ^ 1'b0 ;
  assign n49935 = n22752 | n49934 ;
  assign n49936 = n6281 & n40293 ;
  assign n49937 = n36593 ^ n16381 ^ n8580 ;
  assign n49938 = n3731 | n8034 ;
  assign n49939 = ( n15379 & n24668 ) | ( n15379 & n49938 ) | ( n24668 & n49938 ) ;
  assign n49940 = n4441 | n11724 ;
  assign n49941 = ( n19261 & ~n25558 ) | ( n19261 & n49940 ) | ( ~n25558 & n49940 ) ;
  assign n49942 = n24416 ^ n12263 ^ n5514 ;
  assign n49943 = n37275 ^ n29431 ^ n28614 ;
  assign n49944 = ( ~x69 & n49942 ) | ( ~x69 & n49943 ) | ( n49942 & n49943 ) ;
  assign n49945 = n49944 ^ n18972 ^ 1'b0 ;
  assign n49946 = n49945 ^ n29869 ^ n25667 ;
  assign n49947 = ( n615 & ~n9224 ) | ( n615 & n31988 ) | ( ~n9224 & n31988 ) ;
  assign n49948 = n3391 & ~n5720 ;
  assign n49949 = ~n8659 & n49948 ;
  assign n49950 = n49949 ^ n3752 ^ 1'b0 ;
  assign n49951 = n28317 & n49950 ;
  assign n49952 = n49951 ^ n17388 ^ 1'b0 ;
  assign n49953 = ( n1307 & n3462 ) | ( n1307 & ~n30355 ) | ( n3462 & ~n30355 ) ;
  assign n49954 = n49953 ^ n9131 ^ n8781 ;
  assign n49955 = n7986 & n49954 ;
  assign n49956 = ~n49952 & n49955 ;
  assign n49957 = n26080 ^ n11364 ^ n5795 ;
  assign n49958 = n2032 ^ n645 ^ 1'b0 ;
  assign n49959 = ( n24371 & n31915 ) | ( n24371 & n49958 ) | ( n31915 & n49958 ) ;
  assign n49960 = n49959 ^ n46517 ^ 1'b0 ;
  assign n49961 = ~n49957 & n49960 ;
  assign n49962 = ( n1905 & ~n11727 ) | ( n1905 & n29773 ) | ( ~n11727 & n29773 ) ;
  assign n49963 = n49962 ^ n1561 ^ 1'b0 ;
  assign n49964 = n8615 & ~n49963 ;
  assign n49965 = n7949 ^ n2477 ^ 1'b0 ;
  assign n49966 = n49964 & n49965 ;
  assign n49967 = ~n8119 & n49966 ;
  assign n49968 = n40835 & n49967 ;
  assign n49969 = n28359 ^ n23419 ^ 1'b0 ;
  assign n49970 = n49880 ^ n25303 ^ n21274 ;
  assign n49971 = ( n26522 & ~n33640 ) | ( n26522 & n36057 ) | ( ~n33640 & n36057 ) ;
  assign n49972 = n6731 & ~n13149 ;
  assign n49973 = ~n3980 & n49972 ;
  assign n49974 = n49973 ^ n33174 ^ n5054 ;
  assign n49975 = n37605 ^ n20202 ^ 1'b0 ;
  assign n49976 = n27145 & ~n36855 ;
  assign n49977 = n11325 & ~n21948 ;
  assign n49978 = n8909 & n49108 ;
  assign n49979 = n49977 & n49978 ;
  assign n49980 = n27914 ^ n12084 ^ 1'b0 ;
  assign n49981 = n28113 ^ n27074 ^ n6407 ;
  assign n49982 = n27478 & n49981 ;
  assign n49983 = n47836 ^ n35078 ^ 1'b0 ;
  assign n49984 = n31847 ^ n16883 ^ n7241 ;
  assign n49985 = ~n16881 & n22002 ;
  assign n49986 = ( x122 & n10345 ) | ( x122 & ~n18906 ) | ( n10345 & ~n18906 ) ;
  assign n49987 = ( n3979 & n7562 ) | ( n3979 & ~n36132 ) | ( n7562 & ~n36132 ) ;
  assign n49988 = n49987 ^ n2070 ^ 1'b0 ;
  assign n49989 = n49988 ^ n28591 ^ n1329 ;
  assign n49990 = n23376 | n42169 ;
  assign n49992 = n6157 & n31232 ;
  assign n49993 = n49992 ^ n19655 ^ x49 ;
  assign n49991 = ~n37224 & n37861 ;
  assign n49994 = n49993 ^ n49991 ^ 1'b0 ;
  assign n49995 = n38239 ^ n32899 ^ n31925 ;
  assign n49996 = n7089 & n34184 ;
  assign n49997 = ~n49995 & n49996 ;
  assign n49998 = n4667 | n49997 ;
  assign n49999 = n580 | n49998 ;
  assign n50000 = x154 & n5697 ;
  assign n50001 = n50000 ^ n19822 ^ 1'b0 ;
  assign n50002 = ( n3974 & ~n27954 ) | ( n3974 & n50001 ) | ( ~n27954 & n50001 ) ;
  assign n50003 = ~n23943 & n50002 ;
  assign n50004 = ~n14350 & n50003 ;
  assign n50005 = n34922 ^ n7689 ^ 1'b0 ;
  assign n50006 = n50005 ^ n30710 ^ n17153 ;
  assign n50007 = n9164 & ~n41348 ;
  assign n50008 = ( n40228 & n50006 ) | ( n40228 & n50007 ) | ( n50006 & n50007 ) ;
  assign n50009 = n47150 ^ n21200 ^ n3691 ;
  assign n50010 = ( n15225 & n16373 ) | ( n15225 & ~n21771 ) | ( n16373 & ~n21771 ) ;
  assign n50011 = n50010 ^ n14616 ^ n6307 ;
  assign n50014 = n21648 & ~n23685 ;
  assign n50012 = ( n27542 & ~n27811 ) | ( n27542 & n27937 ) | ( ~n27811 & n27937 ) ;
  assign n50013 = ~n12444 & n50012 ;
  assign n50015 = n50014 ^ n50013 ^ n49000 ;
  assign n50017 = n22334 & ~n30206 ;
  assign n50016 = n2228 & n8424 ;
  assign n50018 = n50017 ^ n50016 ^ 1'b0 ;
  assign n50019 = n50018 ^ n29855 ^ n3609 ;
  assign n50020 = n50019 ^ n29115 ^ n12709 ;
  assign n50021 = n42220 ^ n32415 ^ n27389 ;
  assign n50022 = n5374 | n25019 ;
  assign n50023 = n25466 & ~n50022 ;
  assign n50024 = n2741 & ~n10151 ;
  assign n50025 = n36337 & n50024 ;
  assign n50026 = n2300 | n19611 ;
  assign n50027 = ( n6470 & n36171 ) | ( n6470 & ~n50026 ) | ( n36171 & ~n50026 ) ;
  assign n50028 = n38921 ^ n16838 ^ n6314 ;
  assign n50029 = n6736 ^ n4760 ^ 1'b0 ;
  assign n50030 = n10403 & n50029 ;
  assign n50031 = ( n1298 & ~n7577 ) | ( n1298 & n13058 ) | ( ~n7577 & n13058 ) ;
  assign n50032 = n12975 ^ n4849 ^ n665 ;
  assign n50033 = ( n23241 & n34877 ) | ( n23241 & n50032 ) | ( n34877 & n50032 ) ;
  assign n50034 = n50033 ^ n3305 ^ 1'b0 ;
  assign n50035 = n50031 | n50034 ;
  assign n50036 = n39011 ^ n32084 ^ n13202 ;
  assign n50037 = ( n17418 & n22767 ) | ( n17418 & ~n38037 ) | ( n22767 & ~n38037 ) ;
  assign n50040 = n12016 | n28837 ;
  assign n50041 = n30082 ^ n27522 ^ n16418 ;
  assign n50042 = n50041 ^ n45275 ^ 1'b0 ;
  assign n50043 = n50040 & n50042 ;
  assign n50038 = n11734 ^ n6300 ^ n2188 ;
  assign n50039 = ( n2535 & n27729 ) | ( n2535 & ~n50038 ) | ( n27729 & ~n50038 ) ;
  assign n50044 = n50043 ^ n50039 ^ n17001 ;
  assign n50045 = n26624 ^ n5277 ^ n1001 ;
  assign n50046 = ( n9982 & ~n12040 ) | ( n9982 & n50045 ) | ( ~n12040 & n50045 ) ;
  assign n50047 = n50046 ^ n19773 ^ n12841 ;
  assign n50048 = ~n2451 & n32218 ;
  assign n50049 = n11241 & n50048 ;
  assign n50050 = ( n8582 & ~n28798 ) | ( n8582 & n50049 ) | ( ~n28798 & n50049 ) ;
  assign n50051 = ~n50047 & n50050 ;
  assign n50052 = n898 & ~n15888 ;
  assign n50053 = n40439 ^ n35617 ^ n15851 ;
  assign n50054 = n23500 ^ n22697 ^ n14627 ;
  assign n50055 = n50054 ^ n27476 ^ n16414 ;
  assign n50056 = ( n31102 & ~n50053 ) | ( n31102 & n50055 ) | ( ~n50053 & n50055 ) ;
  assign n50057 = n14638 ^ n5313 ^ 1'b0 ;
  assign n50058 = n10656 | n50057 ;
  assign n50059 = n50058 ^ n27546 ^ n22034 ;
  assign n50060 = n33887 ^ n2151 ^ 1'b0 ;
  assign n50061 = n10827 | n50060 ;
  assign n50062 = n50061 ^ n27673 ^ n3781 ;
  assign n50064 = n48331 ^ n23727 ^ n8068 ;
  assign n50063 = ( ~n7139 & n20807 ) | ( ~n7139 & n34356 ) | ( n20807 & n34356 ) ;
  assign n50065 = n50064 ^ n50063 ^ n7056 ;
  assign n50066 = n39898 ^ n22801 ^ n11762 ;
  assign n50067 = n42348 & ~n42743 ;
  assign n50068 = n45817 & n50067 ;
  assign n50069 = n50068 ^ n7465 ^ n4081 ;
  assign n50070 = n16281 ^ n3872 ^ 1'b0 ;
  assign n50071 = ~n4524 & n34123 ;
  assign n50072 = n50071 ^ n40361 ^ 1'b0 ;
  assign n50073 = n45145 ^ n13586 ^ 1'b0 ;
  assign n50074 = n48966 ^ n17822 ^ n2038 ;
  assign n50075 = ( n6141 & n15616 ) | ( n6141 & n50074 ) | ( n15616 & n50074 ) ;
  assign n50076 = n41385 ^ n25900 ^ n12423 ;
  assign n50077 = ( ~x236 & n8819 ) | ( ~x236 & n50076 ) | ( n8819 & n50076 ) ;
  assign n50078 = n50077 ^ n43464 ^ 1'b0 ;
  assign n50079 = n7957 & ~n50078 ;
  assign n50080 = n50079 ^ n21030 ^ n12467 ;
  assign n50081 = ( n7954 & n18688 ) | ( n7954 & ~n41228 ) | ( n18688 & ~n41228 ) ;
  assign n50082 = n10625 & ~n42220 ;
  assign n50083 = ~x52 & n50082 ;
  assign n50084 = n50083 ^ n14634 ^ n8089 ;
  assign n50085 = ( n17533 & ~n20512 ) | ( n17533 & n50084 ) | ( ~n20512 & n50084 ) ;
  assign n50086 = n15811 | n50085 ;
  assign n50087 = ( ~n24351 & n36116 ) | ( ~n24351 & n50086 ) | ( n36116 & n50086 ) ;
  assign n50088 = ( n8958 & n10444 ) | ( n8958 & n18453 ) | ( n10444 & n18453 ) ;
  assign n50089 = n50088 ^ n48134 ^ n46811 ;
  assign n50090 = ( n15732 & n33119 ) | ( n15732 & n50089 ) | ( n33119 & n50089 ) ;
  assign n50091 = ( n3639 & n14112 ) | ( n3639 & n21862 ) | ( n14112 & n21862 ) ;
  assign n50092 = n938 & n3483 ;
  assign n50093 = n39526 ^ n25021 ^ n5684 ;
  assign n50094 = ~n45847 & n50093 ;
  assign n50095 = n37640 ^ n19373 ^ n15550 ;
  assign n50096 = n50095 ^ n13897 ^ 1'b0 ;
  assign n50097 = ~n2302 & n50096 ;
  assign n50098 = n20498 ^ n5777 ^ 1'b0 ;
  assign n50099 = ( ~n2066 & n41720 ) | ( ~n2066 & n50098 ) | ( n41720 & n50098 ) ;
  assign n50100 = n50099 ^ n35011 ^ n12340 ;
  assign n50101 = n9458 & n31187 ;
  assign n50102 = ( ~n3096 & n30496 ) | ( ~n3096 & n38915 ) | ( n30496 & n38915 ) ;
  assign n50103 = n50102 ^ n38330 ^ n22719 ;
  assign n50104 = ~n39868 & n50103 ;
  assign n50105 = ( n1084 & n11273 ) | ( n1084 & ~n12406 ) | ( n11273 & ~n12406 ) ;
  assign n50106 = n4681 | n50105 ;
  assign n50107 = n50106 ^ n7375 ^ 1'b0 ;
  assign n50108 = ( n4049 & n12415 ) | ( n4049 & n50107 ) | ( n12415 & n50107 ) ;
  assign n50109 = ~n8335 & n20031 ;
  assign n50110 = n39595 ^ n33217 ^ n12340 ;
  assign n50111 = ~n9212 & n37521 ;
  assign n50112 = ( n15100 & ~n18280 ) | ( n15100 & n20421 ) | ( ~n18280 & n20421 ) ;
  assign n50113 = ~n23164 & n50112 ;
  assign n50114 = n50113 ^ n26957 ^ 1'b0 ;
  assign n50115 = n44801 & n50114 ;
  assign n50116 = ~n1983 & n50115 ;
  assign n50117 = n12418 | n50116 ;
  assign n50118 = n50117 ^ n1406 ^ 1'b0 ;
  assign n50119 = ~n2752 & n33273 ;
  assign n50120 = n18343 & ~n26788 ;
  assign n50121 = ( ~n5467 & n7089 ) | ( ~n5467 & n50120 ) | ( n7089 & n50120 ) ;
  assign n50122 = n47081 ^ n20221 ^ n2635 ;
  assign n50123 = ~x99 & n3081 ;
  assign n50124 = n17329 ^ n12546 ^ 1'b0 ;
  assign n50125 = n14173 & ~n50124 ;
  assign n50126 = ( ~n22513 & n50123 ) | ( ~n22513 & n50125 ) | ( n50123 & n50125 ) ;
  assign n50127 = n47986 ^ n40409 ^ 1'b0 ;
  assign n50128 = n50127 ^ n49733 ^ n4510 ;
  assign n50130 = n2239 & n10951 ;
  assign n50129 = n13235 | n31039 ;
  assign n50131 = n50130 ^ n50129 ^ 1'b0 ;
  assign n50132 = n46269 ^ n31155 ^ n5811 ;
  assign n50133 = n10292 ^ n5111 ^ n593 ;
  assign n50139 = ~n715 & n13309 ;
  assign n50140 = n2912 & n50139 ;
  assign n50135 = ( n10315 & n11332 ) | ( n10315 & n33996 ) | ( n11332 & n33996 ) ;
  assign n50136 = n38094 ^ n278 ^ 1'b0 ;
  assign n50137 = n50135 | n50136 ;
  assign n50134 = n5409 & ~n40035 ;
  assign n50138 = n50137 ^ n50134 ^ n30025 ;
  assign n50141 = n50140 ^ n50138 ^ n45593 ;
  assign n50142 = ( n5386 & n32240 ) | ( n5386 & n38000 ) | ( n32240 & n38000 ) ;
  assign n50143 = ( n32107 & ~n40355 ) | ( n32107 & n49054 ) | ( ~n40355 & n49054 ) ;
  assign n50144 = ( ~n5628 & n12371 ) | ( ~n5628 & n50143 ) | ( n12371 & n50143 ) ;
  assign n50145 = n44837 ^ n21126 ^ 1'b0 ;
  assign n50146 = n50145 ^ n22101 ^ n10553 ;
  assign n50147 = n16897 ^ n15398 ^ 1'b0 ;
  assign n50148 = n4680 & ~n50147 ;
  assign n50149 = n23882 ^ n13273 ^ n4572 ;
  assign n50150 = n42954 | n49054 ;
  assign n50151 = n14604 & ~n50150 ;
  assign n50152 = n50151 ^ n33984 ^ 1'b0 ;
  assign n50153 = n50152 ^ n14000 ^ 1'b0 ;
  assign n50154 = n50149 & n50153 ;
  assign n50155 = ( n29399 & n35310 ) | ( n29399 & n37552 ) | ( n35310 & n37552 ) ;
  assign n50156 = ( n17373 & ~n21252 ) | ( n17373 & n27669 ) | ( ~n21252 & n27669 ) ;
  assign n50157 = n14227 | n17460 ;
  assign n50158 = ( n1578 & ~n18638 ) | ( n1578 & n45603 ) | ( ~n18638 & n45603 ) ;
  assign n50159 = ( n17291 & n27685 ) | ( n17291 & n46373 ) | ( n27685 & n46373 ) ;
  assign n50161 = n23319 | n30990 ;
  assign n50160 = n35458 & n49966 ;
  assign n50162 = n50161 ^ n50160 ^ 1'b0 ;
  assign n50163 = ( n1144 & n8480 ) | ( n1144 & n34880 ) | ( n8480 & n34880 ) ;
  assign n50164 = n50163 ^ n44363 ^ n8632 ;
  assign n50165 = n11238 | n25674 ;
  assign n50166 = n36802 ^ n5067 ^ 1'b0 ;
  assign n50167 = n48343 ^ n3376 ^ 1'b0 ;
  assign n50171 = n29826 ^ n22615 ^ n9997 ;
  assign n50170 = ( ~n9323 & n21456 ) | ( ~n9323 & n33216 ) | ( n21456 & n33216 ) ;
  assign n50172 = n50171 ^ n50170 ^ n27128 ;
  assign n50168 = n32527 ^ n28837 ^ 1'b0 ;
  assign n50169 = n30057 & n50168 ;
  assign n50173 = n50172 ^ n50169 ^ n23455 ;
  assign n50174 = n9120 | n50173 ;
  assign n50175 = n50174 ^ n10343 ^ 1'b0 ;
  assign n50176 = ( n2613 & n50167 ) | ( n2613 & ~n50175 ) | ( n50167 & ~n50175 ) ;
  assign n50177 = n24976 | n35115 ;
  assign n50178 = n50177 ^ n26327 ^ n23332 ;
  assign n50181 = ( ~n8167 & n8408 ) | ( ~n8167 & n45507 ) | ( n8408 & n45507 ) ;
  assign n50182 = n50181 ^ n30775 ^ n2892 ;
  assign n50179 = n24961 ^ n10623 ^ n2659 ;
  assign n50180 = n50179 ^ n21556 ^ n10773 ;
  assign n50183 = n50182 ^ n50180 ^ n32547 ;
  assign n50184 = ( ~n20320 & n32444 ) | ( ~n20320 & n50183 ) | ( n32444 & n50183 ) ;
  assign n50185 = ( n6296 & n8245 ) | ( n6296 & ~n15650 ) | ( n8245 & ~n15650 ) ;
  assign n50186 = n26519 ^ n24653 ^ 1'b0 ;
  assign n50187 = n36363 ^ n25380 ^ 1'b0 ;
  assign n50188 = n50186 | n50187 ;
  assign n50189 = ~n3518 & n7439 ;
  assign n50190 = n50189 ^ n25713 ^ 1'b0 ;
  assign n50191 = n5037 & n50190 ;
  assign n50192 = ~n31002 & n50191 ;
  assign n50193 = n50192 ^ n50094 ^ 1'b0 ;
  assign n50194 = ~n31936 & n50193 ;
  assign n50195 = n36799 ^ n26767 ^ 1'b0 ;
  assign n50196 = n27730 ^ n19662 ^ n17940 ;
  assign n50197 = n17096 | n28835 ;
  assign n50198 = n50197 ^ n10336 ^ 1'b0 ;
  assign n50199 = n2624 & ~n50198 ;
  assign n50200 = n13420 & n50199 ;
  assign n50201 = n50200 ^ n32620 ^ 1'b0 ;
  assign n50202 = ( n14359 & n38614 ) | ( n14359 & ~n39539 ) | ( n38614 & ~n39539 ) ;
  assign n50203 = n469 | n50202 ;
  assign n50204 = n29079 ^ n24367 ^ n14544 ;
  assign n50205 = n33713 & ~n50204 ;
  assign n50206 = n16064 ^ n11764 ^ 1'b0 ;
  assign n50207 = ~n45090 & n50206 ;
  assign n50208 = n21019 | n47636 ;
  assign n50209 = n50208 ^ n42509 ^ 1'b0 ;
  assign n50210 = n12035 | n28809 ;
  assign n50211 = n50210 ^ n3897 ^ 1'b0 ;
  assign n50212 = ( n25221 & ~n27119 ) | ( n25221 & n45668 ) | ( ~n27119 & n45668 ) ;
  assign n50213 = ( n11166 & n21570 ) | ( n11166 & n23170 ) | ( n21570 & n23170 ) ;
  assign n50214 = n50213 ^ n18226 ^ 1'b0 ;
  assign n50215 = n50212 & n50214 ;
  assign n50216 = ( n18293 & n22537 ) | ( n18293 & n37667 ) | ( n22537 & n37667 ) ;
  assign n50217 = n11590 ^ n460 ^ 1'b0 ;
  assign n50218 = ~n28638 & n50217 ;
  assign n50219 = n50218 ^ n7324 ^ 1'b0 ;
  assign n50220 = ( n9815 & ~n50216 ) | ( n9815 & n50219 ) | ( ~n50216 & n50219 ) ;
  assign n50221 = n12807 & ~n29104 ;
  assign n50222 = n2299 & n50221 ;
  assign n50223 = n23547 ^ n7100 ^ 1'b0 ;
  assign n50224 = n16301 & n17613 ;
  assign n50225 = n50224 ^ n16508 ^ 1'b0 ;
  assign n50226 = ( ~n50222 & n50223 ) | ( ~n50222 & n50225 ) | ( n50223 & n50225 ) ;
  assign n50227 = n43749 ^ n13909 ^ n9480 ;
  assign n50228 = n22250 ^ n19296 ^ 1'b0 ;
  assign n50229 = n50228 ^ n20236 ^ n7714 ;
  assign n50230 = n48731 ^ n27044 ^ n17130 ;
  assign n50231 = n50230 ^ n12635 ^ n6607 ;
  assign n50232 = ( n3456 & ~n27916 ) | ( n3456 & n50231 ) | ( ~n27916 & n50231 ) ;
  assign n50233 = n16990 ^ n1840 ^ 1'b0 ;
  assign n50234 = ~n35092 & n50233 ;
  assign n50235 = ( ~n28988 & n48377 ) | ( ~n28988 & n50234 ) | ( n48377 & n50234 ) ;
  assign n50236 = ( n10737 & n13270 ) | ( n10737 & n31782 ) | ( n13270 & n31782 ) ;
  assign n50237 = ( n28945 & n44852 ) | ( n28945 & ~n50236 ) | ( n44852 & ~n50236 ) ;
  assign n50238 = n29115 & n50085 ;
  assign n50240 = n2325 & ~n11293 ;
  assign n50241 = ~n36023 & n50240 ;
  assign n50239 = x17 & n42907 ;
  assign n50242 = n50241 ^ n50239 ^ 1'b0 ;
  assign n50243 = n25899 | n31639 ;
  assign n50244 = n50243 ^ n5119 ^ 1'b0 ;
  assign n50245 = ( n10767 & n15912 ) | ( n10767 & ~n17577 ) | ( n15912 & ~n17577 ) ;
  assign n50246 = n46070 ^ n3366 ^ n1235 ;
  assign n50247 = n18972 | n46611 ;
  assign n50248 = n33490 ^ n31007 ^ n1461 ;
  assign n50249 = ~n363 & n10723 ;
  assign n50250 = n50249 ^ n9722 ^ 1'b0 ;
  assign n50251 = n50250 ^ n48711 ^ n5285 ;
  assign n50252 = ( n7440 & ~n18496 ) | ( n7440 & n28048 ) | ( ~n18496 & n28048 ) ;
  assign n50253 = ( n15847 & n32386 ) | ( n15847 & n50252 ) | ( n32386 & n50252 ) ;
  assign n50254 = n8068 & ~n31603 ;
  assign n50255 = ~n11847 & n50254 ;
  assign n50256 = ~n8096 & n50255 ;
  assign n50257 = n18774 | n50256 ;
  assign n50258 = n50257 ^ n20817 ^ 1'b0 ;
  assign n50259 = n44220 ^ n22217 ^ n617 ;
  assign n50260 = n8223 & n19961 ;
  assign n50261 = n50260 ^ n20679 ^ 1'b0 ;
  assign n50262 = n28279 ^ n24026 ^ n4389 ;
  assign n50263 = n50262 ^ n39186 ^ 1'b0 ;
  assign n50264 = n18412 ^ n8985 ^ n2054 ;
  assign n50265 = ( n10467 & n29128 ) | ( n10467 & n50264 ) | ( n29128 & n50264 ) ;
  assign n50266 = n35233 ^ n7703 ^ n5682 ;
  assign n50267 = n10349 & n16266 ;
  assign n50268 = n50267 ^ n8182 ^ 1'b0 ;
  assign n50269 = n50268 ^ n18518 ^ n4735 ;
  assign n50270 = n34480 ^ n25327 ^ 1'b0 ;
  assign n50271 = x112 & ~n50270 ;
  assign n50272 = ~n6913 & n13324 ;
  assign n50273 = ~n14603 & n50272 ;
  assign n50274 = n14431 | n50273 ;
  assign n50275 = n5119 | n50274 ;
  assign n50276 = n22103 ^ n15410 ^ n4618 ;
  assign n50277 = n50276 ^ n35418 ^ 1'b0 ;
  assign n50278 = n28054 & ~n50277 ;
  assign n50279 = n29268 ^ n26769 ^ n23478 ;
  assign n50280 = ( n10632 & n11114 ) | ( n10632 & n50279 ) | ( n11114 & n50279 ) ;
  assign n50281 = n4698 & ~n50280 ;
  assign n50282 = n50281 ^ n25663 ^ 1'b0 ;
  assign n50283 = ~n8072 & n50282 ;
  assign n50284 = ~n50278 & n50283 ;
  assign n50285 = n5237 | n13969 ;
  assign n50286 = n15379 ^ n12079 ^ 1'b0 ;
  assign n50287 = n18138 ^ n14838 ^ n3987 ;
  assign n50288 = n50287 ^ n18349 ^ n4866 ;
  assign n50289 = n37538 ^ n13748 ^ 1'b0 ;
  assign n50295 = ( ~n3500 & n11206 ) | ( ~n3500 & n13190 ) | ( n11206 & n13190 ) ;
  assign n50291 = ( ~n2223 & n8160 ) | ( ~n2223 & n9122 ) | ( n8160 & n9122 ) ;
  assign n50292 = n50291 ^ n1813 ^ 1'b0 ;
  assign n50293 = n50292 ^ n30973 ^ 1'b0 ;
  assign n50294 = ~n26297 & n50293 ;
  assign n50290 = n30877 ^ n27373 ^ n2818 ;
  assign n50296 = n50295 ^ n50294 ^ n50290 ;
  assign n50297 = n20178 ^ n7783 ^ 1'b0 ;
  assign n50298 = n21945 | n50297 ;
  assign n50301 = n1548 & ~n5957 ;
  assign n50302 = n50301 ^ n4688 ^ 1'b0 ;
  assign n50299 = ( n12524 & n19888 ) | ( n12524 & ~n45269 ) | ( n19888 & ~n45269 ) ;
  assign n50300 = n13048 & n50299 ;
  assign n50303 = n50302 ^ n50300 ^ 1'b0 ;
  assign n50305 = n11412 ^ n2390 ^ n390 ;
  assign n50304 = ~n19882 & n41117 ;
  assign n50306 = n50305 ^ n50304 ^ 1'b0 ;
  assign n50307 = ( ~n14836 & n41284 ) | ( ~n14836 & n50306 ) | ( n41284 & n50306 ) ;
  assign n50308 = n40890 ^ n19115 ^ 1'b0 ;
  assign n50309 = n50308 ^ n41040 ^ n3808 ;
  assign n50310 = n3536 ^ n467 ^ 1'b0 ;
  assign n50311 = n15825 & n50310 ;
  assign n50312 = n50311 ^ n47757 ^ n41706 ;
  assign n50314 = n19233 ^ n13438 ^ n11855 ;
  assign n50313 = ( ~n6615 & n13674 ) | ( ~n6615 & n26081 ) | ( n13674 & n26081 ) ;
  assign n50315 = n50314 ^ n50313 ^ n2032 ;
  assign n50316 = ( n5617 & n7862 ) | ( n5617 & ~n24428 ) | ( n7862 & ~n24428 ) ;
  assign n50317 = n50316 ^ n28356 ^ n4272 ;
  assign n50318 = n50317 ^ n17075 ^ n11481 ;
  assign n50319 = n37514 ^ n27072 ^ n9695 ;
  assign n50320 = ( n7224 & n16433 ) | ( n7224 & ~n41180 ) | ( n16433 & ~n41180 ) ;
  assign n50321 = n3553 & n15869 ;
  assign n50322 = n50321 ^ n29438 ^ 1'b0 ;
  assign n50323 = n19141 ^ n8044 ^ x23 ;
  assign n50324 = ( n4337 & n47166 ) | ( n4337 & ~n50323 ) | ( n47166 & ~n50323 ) ;
  assign n50325 = ~n42044 & n50324 ;
  assign n50326 = ( n9188 & n10751 ) | ( n9188 & ~n40323 ) | ( n10751 & ~n40323 ) ;
  assign n50327 = n490 & n50326 ;
  assign n50328 = n50325 & n50327 ;
  assign n50329 = n10582 & ~n15265 ;
  assign n50330 = ~n2586 & n50329 ;
  assign n50332 = ( n27617 & ~n28129 ) | ( n27617 & n37827 ) | ( ~n28129 & n37827 ) ;
  assign n50331 = n6253 & ~n16527 ;
  assign n50333 = n50332 ^ n50331 ^ 1'b0 ;
  assign n50334 = ( ~n19091 & n50330 ) | ( ~n19091 & n50333 ) | ( n50330 & n50333 ) ;
  assign n50335 = n46491 | n50334 ;
  assign n50336 = n50328 & ~n50335 ;
  assign n50337 = n49314 ^ n36459 ^ n22778 ;
  assign n50338 = n19901 & ~n47212 ;
  assign n50339 = ( n7467 & n30267 ) | ( n7467 & ~n50338 ) | ( n30267 & ~n50338 ) ;
  assign n50340 = n46775 ^ n33260 ^ 1'b0 ;
  assign n50341 = n36356 ^ n16756 ^ 1'b0 ;
  assign n50342 = n27316 & n50341 ;
  assign n50343 = n8794 | n24705 ;
  assign n50344 = n50343 ^ n24621 ^ 1'b0 ;
  assign n50345 = ( ~n5674 & n37082 ) | ( ~n5674 & n50344 ) | ( n37082 & n50344 ) ;
  assign n50346 = n50345 ^ n49065 ^ 1'b0 ;
  assign n50347 = ~n1560 & n23726 ;
  assign n50348 = n50347 ^ n45187 ^ 1'b0 ;
  assign n50349 = n28754 ^ n12111 ^ 1'b0 ;
  assign n50350 = n49529 ^ n2888 ^ 1'b0 ;
  assign n50351 = n15976 & ~n50350 ;
  assign n50352 = ( n489 & ~n6599 ) | ( n489 & n35817 ) | ( ~n6599 & n35817 ) ;
  assign n50353 = n48005 ^ n23614 ^ 1'b0 ;
  assign n50354 = n28379 ^ n24856 ^ n13512 ;
  assign n50355 = n50354 ^ n33962 ^ n8793 ;
  assign n50356 = n34573 ^ n16212 ^ n10444 ;
  assign n50357 = n50356 ^ n46046 ^ n41320 ;
  assign n50358 = ( n4083 & n10949 ) | ( n4083 & n32295 ) | ( n10949 & n32295 ) ;
  assign n50359 = ~n8967 & n42926 ;
  assign n50360 = n49392 ^ n47074 ^ n42143 ;
  assign n50361 = n48443 ^ n28816 ^ 1'b0 ;
  assign n50362 = ~n44806 & n50361 ;
  assign n50363 = ~n10641 & n50362 ;
  assign n50364 = n6801 ^ n1090 ^ 1'b0 ;
  assign n50365 = n20687 | n50364 ;
  assign n50366 = n13285 & ~n36320 ;
  assign n50367 = n34556 & n50366 ;
  assign n50368 = n26264 ^ n1842 ^ 1'b0 ;
  assign n50369 = n49452 & n50368 ;
  assign n50370 = n17870 & ~n35343 ;
  assign n50371 = n50370 ^ n21229 ^ n10600 ;
  assign n50372 = n29563 ^ n13390 ^ 1'b0 ;
  assign n50373 = ( n834 & n11236 ) | ( n834 & n21533 ) | ( n11236 & n21533 ) ;
  assign n50376 = n802 ^ x195 ^ 1'b0 ;
  assign n50377 = n6191 | n50376 ;
  assign n50374 = ~n38845 & n42213 ;
  assign n50375 = n50374 ^ n31074 ^ 1'b0 ;
  assign n50378 = n50377 ^ n50375 ^ n24672 ;
  assign n50379 = n39569 ^ n23175 ^ n1436 ;
  assign n50381 = n34976 ^ n20656 ^ n20506 ;
  assign n50380 = n9148 | n40518 ;
  assign n50382 = n50381 ^ n50380 ^ 1'b0 ;
  assign n50383 = ( x129 & ~n10456 ) | ( x129 & n19219 ) | ( ~n10456 & n19219 ) ;
  assign n50384 = n3007 & n12831 ;
  assign n50385 = ~n50383 & n50384 ;
  assign n50386 = n3144 & ~n18793 ;
  assign n50387 = ~n5818 & n50386 ;
  assign n50388 = n1893 & n50361 ;
  assign n50389 = n6478 | n34011 ;
  assign n50390 = ( n1119 & ~n48143 ) | ( n1119 & n50389 ) | ( ~n48143 & n50389 ) ;
  assign n50392 = n6873 & ~n40975 ;
  assign n50393 = n50392 ^ n22733 ^ 1'b0 ;
  assign n50391 = n29903 ^ n25327 ^ n11205 ;
  assign n50394 = n50393 ^ n50391 ^ n15712 ;
  assign n50397 = n17032 ^ n14593 ^ n11799 ;
  assign n50395 = n3890 & ~n19494 ;
  assign n50396 = n4939 & n50395 ;
  assign n50398 = n50397 ^ n50396 ^ 1'b0 ;
  assign n50399 = n25069 ^ n18128 ^ 1'b0 ;
  assign n50400 = n21249 & n50399 ;
  assign n50401 = ( n19683 & n21937 ) | ( n19683 & n50400 ) | ( n21937 & n50400 ) ;
  assign n50402 = n50401 ^ n8056 ^ n656 ;
  assign n50403 = ( n10569 & n22912 ) | ( n10569 & n43769 ) | ( n22912 & n43769 ) ;
  assign n50404 = n14897 ^ n10746 ^ n6242 ;
  assign n50405 = n2268 & ~n26010 ;
  assign n50406 = ~n15697 & n50405 ;
  assign n50407 = n16866 & n17587 ;
  assign n50408 = ( n4731 & n15250 ) | ( n4731 & n28017 ) | ( n15250 & n28017 ) ;
  assign n50409 = n13295 & n50408 ;
  assign n50410 = ~n3195 & n20132 ;
  assign n50411 = n50409 & n50410 ;
  assign n50412 = n50411 ^ n10047 ^ 1'b0 ;
  assign n50413 = n41933 & n46771 ;
  assign n50414 = n50413 ^ n46148 ^ 1'b0 ;
  assign n50415 = n3512 | n24521 ;
  assign n50416 = n50415 ^ n7445 ^ 1'b0 ;
  assign n50417 = ( ~n3214 & n13700 ) | ( ~n3214 & n50416 ) | ( n13700 & n50416 ) ;
  assign n50418 = ( n809 & ~n7311 ) | ( n809 & n34694 ) | ( ~n7311 & n34694 ) ;
  assign n50419 = ( x117 & n12287 ) | ( x117 & n50418 ) | ( n12287 & n50418 ) ;
  assign n50420 = n21729 ^ n9314 ^ 1'b0 ;
  assign n50421 = n34040 ^ n34039 ^ n25896 ;
  assign n50422 = ~n33036 & n50421 ;
  assign n50423 = ~n46681 & n50422 ;
  assign n50424 = n50423 ^ n14428 ^ n3868 ;
  assign n50425 = n19552 ^ n16598 ^ n5588 ;
  assign n50426 = n43458 ^ n42866 ^ 1'b0 ;
  assign n50427 = ( n15962 & ~n50425 ) | ( n15962 & n50426 ) | ( ~n50425 & n50426 ) ;
  assign n50428 = ( n3249 & ~n4558 ) | ( n3249 & n35510 ) | ( ~n4558 & n35510 ) ;
  assign n50429 = ( ~n5085 & n8790 ) | ( ~n5085 & n20950 ) | ( n8790 & n20950 ) ;
  assign n50430 = n14004 ^ n2719 ^ 1'b0 ;
  assign n50431 = ~n39914 & n50430 ;
  assign n50432 = ( n496 & n50429 ) | ( n496 & n50431 ) | ( n50429 & n50431 ) ;
  assign n50433 = ~n958 & n2451 ;
  assign n50434 = ~n2649 & n41229 ;
  assign n50435 = ~n14364 & n50434 ;
  assign n50438 = ~n19783 & n29928 ;
  assign n50439 = n50438 ^ n43554 ^ 1'b0 ;
  assign n50436 = ( n3574 & n9485 ) | ( n3574 & ~n9951 ) | ( n9485 & ~n9951 ) ;
  assign n50437 = ~n7373 & n50436 ;
  assign n50440 = n50439 ^ n50437 ^ 1'b0 ;
  assign n50441 = n12310 | n40683 ;
  assign n50442 = n50441 ^ n12209 ^ n4539 ;
  assign n50443 = ( n10538 & n32054 ) | ( n10538 & n50442 ) | ( n32054 & n50442 ) ;
  assign n50444 = n10879 & ~n15306 ;
  assign n50445 = n50444 ^ n25967 ^ 1'b0 ;
  assign n50446 = n50445 ^ n41740 ^ n10790 ;
  assign n50447 = n30590 ^ n8675 ^ 1'b0 ;
  assign n50448 = n38400 ^ n13190 ^ 1'b0 ;
  assign n50449 = ( n22261 & n47083 ) | ( n22261 & n47582 ) | ( n47083 & n47582 ) ;
  assign n50450 = ( n5270 & ~n12010 ) | ( n5270 & n27753 ) | ( ~n12010 & n27753 ) ;
  assign n50451 = n50450 ^ n46758 ^ n16779 ;
  assign n50452 = n50451 ^ n7815 ^ 1'b0 ;
  assign n50453 = n50452 ^ n45683 ^ n32825 ;
  assign n50454 = ~n12694 & n50453 ;
  assign n50455 = n22619 ^ n17105 ^ 1'b0 ;
  assign n50456 = n35907 & n50455 ;
  assign n50457 = ~n12895 & n22230 ;
  assign n50458 = n50457 ^ n25447 ^ 1'b0 ;
  assign n50459 = n50458 ^ n34186 ^ n25234 ;
  assign n50460 = ( n1743 & ~n8344 ) | ( n1743 & n12125 ) | ( ~n8344 & n12125 ) ;
  assign n50461 = n3291 | n50460 ;
  assign n50462 = n39201 & ~n50461 ;
  assign n50463 = ( ~n26568 & n45359 ) | ( ~n26568 & n50462 ) | ( n45359 & n50462 ) ;
  assign n50464 = n20422 ^ n5367 ^ n3181 ;
  assign n50465 = n6955 | n34686 ;
  assign n50466 = n48418 | n50465 ;
  assign n50467 = ( n48086 & n50464 ) | ( n48086 & n50466 ) | ( n50464 & n50466 ) ;
  assign n50471 = n10067 ^ n8259 ^ n7151 ;
  assign n50468 = n14733 | n30082 ;
  assign n50469 = n44054 & ~n50468 ;
  assign n50470 = n50469 ^ n41821 ^ n9639 ;
  assign n50472 = n50471 ^ n50470 ^ n17126 ;
  assign n50473 = ( n3838 & n36761 ) | ( n3838 & n50472 ) | ( n36761 & n50472 ) ;
  assign n50474 = ( n1892 & n20855 ) | ( n1892 & n28565 ) | ( n20855 & n28565 ) ;
  assign n50475 = ( ~n7947 & n31549 ) | ( ~n7947 & n45084 ) | ( n31549 & n45084 ) ;
  assign n50476 = n47543 & n50475 ;
  assign n50477 = n20728 ^ n16628 ^ 1'b0 ;
  assign n50478 = n17892 ^ n12674 ^ 1'b0 ;
  assign n50479 = n36323 ^ n7440 ^ 1'b0 ;
  assign n50480 = n18728 ^ n13172 ^ 1'b0 ;
  assign n50481 = n50479 & n50480 ;
  assign n50482 = n9096 | n20495 ;
  assign n50483 = n48259 ^ n28137 ^ n8651 ;
  assign n50484 = n50483 ^ n36727 ^ 1'b0 ;
  assign n50485 = ( n17970 & n48413 ) | ( n17970 & ~n50484 ) | ( n48413 & ~n50484 ) ;
  assign n50486 = ( ~n9335 & n12433 ) | ( ~n9335 & n33566 ) | ( n12433 & n33566 ) ;
  assign n50487 = n20035 & n43512 ;
  assign n50488 = ( x198 & n3138 ) | ( x198 & ~n50487 ) | ( n3138 & ~n50487 ) ;
  assign n50489 = ~n50486 & n50488 ;
  assign n50490 = n50489 ^ n36621 ^ n9870 ;
  assign n50493 = ( n11089 & n14338 ) | ( n11089 & n27592 ) | ( n14338 & n27592 ) ;
  assign n50491 = n745 & n6855 ;
  assign n50492 = n50491 ^ n32362 ^ 1'b0 ;
  assign n50494 = n50493 ^ n50492 ^ n29159 ;
  assign n50495 = n50494 ^ n8907 ^ n8405 ;
  assign n50496 = ( n3257 & ~n14319 ) | ( n3257 & n35173 ) | ( ~n14319 & n35173 ) ;
  assign n50497 = ( n13202 & n18131 ) | ( n13202 & ~n23150 ) | ( n18131 & ~n23150 ) ;
  assign n50498 = ( ~n41575 & n50496 ) | ( ~n41575 & n50497 ) | ( n50496 & n50497 ) ;
  assign n50499 = ( ~n5000 & n50495 ) | ( ~n5000 & n50498 ) | ( n50495 & n50498 ) ;
  assign n50500 = n44908 ^ n7977 ^ 1'b0 ;
  assign n50501 = ( n22494 & n25539 ) | ( n22494 & ~n33376 ) | ( n25539 & ~n33376 ) ;
  assign n50502 = n14691 ^ n12120 ^ n1072 ;
  assign n50503 = n13350 & n50502 ;
  assign n50504 = n50503 ^ n3752 ^ 1'b0 ;
  assign n50505 = n17409 & n50504 ;
  assign n50506 = n10808 & n50505 ;
  assign n50507 = n4090 & ~n8219 ;
  assign n50508 = n23564 ^ n18096 ^ 1'b0 ;
  assign n50509 = ~n10936 & n50508 ;
  assign n50510 = n14078 ^ n2942 ^ n1535 ;
  assign n50511 = n37583 ^ n27425 ^ n9974 ;
  assign n50512 = n13104 ^ n4601 ^ 1'b0 ;
  assign n50513 = ( n9299 & ~n30488 ) | ( n9299 & n50512 ) | ( ~n30488 & n50512 ) ;
  assign n50514 = ( n14318 & ~n22631 ) | ( n14318 & n41872 ) | ( ~n22631 & n41872 ) ;
  assign n50515 = n43732 ^ n40779 ^ n6241 ;
  assign n50516 = n21450 | n49384 ;
  assign n50517 = n9029 & n29226 ;
  assign n50518 = ( n8938 & ~n29330 ) | ( n8938 & n50517 ) | ( ~n29330 & n50517 ) ;
  assign n50519 = ( n27086 & ~n50516 ) | ( n27086 & n50518 ) | ( ~n50516 & n50518 ) ;
  assign n50520 = n49006 ^ n45265 ^ n1949 ;
  assign n50521 = ~n8190 & n9494 ;
  assign n50522 = n50521 ^ n4182 ^ 1'b0 ;
  assign n50523 = n1577 & ~n50522 ;
  assign n50524 = n30392 & n50523 ;
  assign n50525 = n6708 & ~n10359 ;
  assign n50526 = n50525 ^ n37978 ^ 1'b0 ;
  assign n50527 = n50526 ^ n42823 ^ 1'b0 ;
  assign n50528 = n13536 & ~n50527 ;
  assign n50529 = n45866 ^ n4440 ^ 1'b0 ;
  assign n50530 = n7489 & n17435 ;
  assign n50531 = ~n883 & n50530 ;
  assign n50532 = n43709 ^ n15397 ^ 1'b0 ;
  assign n50533 = ( n18626 & n20175 ) | ( n18626 & n50532 ) | ( n20175 & n50532 ) ;
  assign n50534 = ~n3789 & n6039 ;
  assign n50535 = n46192 ^ n19828 ^ n637 ;
  assign n50536 = n50535 ^ n42031 ^ 1'b0 ;
  assign n50537 = ( n10279 & n41944 ) | ( n10279 & ~n43082 ) | ( n41944 & ~n43082 ) ;
  assign n50538 = n50537 ^ n41843 ^ 1'b0 ;
  assign n50539 = n17307 ^ n13671 ^ 1'b0 ;
  assign n50540 = n26171 ^ n13034 ^ 1'b0 ;
  assign n50541 = ( n2577 & n29225 ) | ( n2577 & ~n50540 ) | ( n29225 & ~n50540 ) ;
  assign n50542 = ( n15050 & n20570 ) | ( n15050 & n32976 ) | ( n20570 & n32976 ) ;
  assign n50543 = ~n19576 & n30134 ;
  assign n50544 = ( n2750 & ~n15051 ) | ( n2750 & n44442 ) | ( ~n15051 & n44442 ) ;
  assign n50545 = ( n25060 & n27789 ) | ( n25060 & ~n40170 ) | ( n27789 & ~n40170 ) ;
  assign n50546 = n41837 ^ n24119 ^ 1'b0 ;
  assign n50547 = n47609 ^ n6375 ^ 1'b0 ;
  assign n50548 = n12985 & n50547 ;
  assign n50550 = n26001 ^ n12608 ^ n12601 ;
  assign n50551 = ( n10235 & ~n11110 ) | ( n10235 & n50550 ) | ( ~n11110 & n50550 ) ;
  assign n50549 = ( ~n22648 & n23579 ) | ( ~n22648 & n40739 ) | ( n23579 & n40739 ) ;
  assign n50552 = n50551 ^ n50549 ^ n19095 ;
  assign n50553 = n2738 & n50552 ;
  assign n50554 = n23365 & n50553 ;
  assign n50555 = n32097 ^ n26008 ^ 1'b0 ;
  assign n50556 = ( n7196 & n12207 ) | ( n7196 & ~n31124 ) | ( n12207 & ~n31124 ) ;
  assign n50558 = ( ~n9288 & n13203 ) | ( ~n9288 & n32504 ) | ( n13203 & n32504 ) ;
  assign n50557 = n38020 ^ n3132 ^ 1'b0 ;
  assign n50559 = n50558 ^ n50557 ^ 1'b0 ;
  assign n50560 = n15899 ^ n9951 ^ n6459 ;
  assign n50561 = ( n24383 & n40874 ) | ( n24383 & ~n50560 ) | ( n40874 & ~n50560 ) ;
  assign n50562 = ( n14670 & ~n19903 ) | ( n14670 & n22769 ) | ( ~n19903 & n22769 ) ;
  assign n50563 = n47640 ^ n46785 ^ n15669 ;
  assign n50564 = n50563 ^ n13657 ^ 1'b0 ;
  assign n50565 = n50564 ^ n7106 ^ 1'b0 ;
  assign n50566 = n34251 ^ n9000 ^ n7155 ;
  assign n50571 = n1756 & n32373 ;
  assign n50567 = n10649 & ~n43301 ;
  assign n50568 = n50567 ^ n25187 ^ 1'b0 ;
  assign n50569 = n50568 ^ n21239 ^ n755 ;
  assign n50570 = ( ~n21852 & n34191 ) | ( ~n21852 & n50569 ) | ( n34191 & n50569 ) ;
  assign n50572 = n50571 ^ n50570 ^ n17150 ;
  assign n50573 = n28970 | n37943 ;
  assign n50574 = n50573 ^ n19752 ^ 1'b0 ;
  assign n50575 = n28301 | n50574 ;
  assign n50576 = n50575 ^ n38839 ^ 1'b0 ;
  assign n50577 = n10825 | n39735 ;
  assign n50578 = n50577 ^ n13511 ^ 1'b0 ;
  assign n50579 = ~n8340 & n22631 ;
  assign n50580 = n33885 ^ n10206 ^ 1'b0 ;
  assign n50581 = ( n14699 & n18097 ) | ( n14699 & n22174 ) | ( n18097 & n22174 ) ;
  assign n50582 = n33343 & n50581 ;
  assign n50583 = n49628 ^ n28893 ^ n4902 ;
  assign n50584 = n45706 ^ n32093 ^ 1'b0 ;
  assign n50585 = n50583 & ~n50584 ;
  assign n50586 = ( n326 & n3589 ) | ( n326 & ~n19081 ) | ( n3589 & ~n19081 ) ;
  assign n50587 = n50586 ^ n24981 ^ n24213 ;
  assign n50588 = ( n41310 & n46128 ) | ( n41310 & n50587 ) | ( n46128 & n50587 ) ;
  assign n50589 = ~n25195 & n30594 ;
  assign n50590 = n6972 & n50589 ;
  assign n50591 = ( ~n28324 & n46664 ) | ( ~n28324 & n50590 ) | ( n46664 & n50590 ) ;
  assign n50592 = n42587 ^ n7498 ^ 1'b0 ;
  assign n50594 = ( n6624 & n11205 ) | ( n6624 & n40615 ) | ( n11205 & n40615 ) ;
  assign n50593 = ( n15283 & n15352 ) | ( n15283 & ~n31345 ) | ( n15352 & ~n31345 ) ;
  assign n50595 = n50594 ^ n50593 ^ n46999 ;
  assign n50596 = n16683 & ~n50423 ;
  assign n50597 = n50596 ^ n8714 ^ 1'b0 ;
  assign n50598 = ~n8053 & n24941 ;
  assign n50599 = ~n34733 & n50598 ;
  assign n50600 = ( n1074 & n18030 ) | ( n1074 & ~n22614 ) | ( n18030 & ~n22614 ) ;
  assign n50601 = n13647 & ~n30507 ;
  assign n50602 = n50601 ^ n33207 ^ n21209 ;
  assign n50603 = n43954 ^ n28250 ^ n9011 ;
  assign n50604 = n39743 ^ n32312 ^ n26634 ;
  assign n50605 = ~n14543 & n50604 ;
  assign n50606 = n44182 ^ n19212 ^ 1'b0 ;
  assign n50607 = ( n18433 & n28206 ) | ( n18433 & n28498 ) | ( n28206 & n28498 ) ;
  assign n50608 = n23685 ^ n14198 ^ n2753 ;
  assign n50609 = ( n4137 & ~n9740 ) | ( n4137 & n13560 ) | ( ~n9740 & n13560 ) ;
  assign n50610 = n50609 ^ n15907 ^ 1'b0 ;
  assign n50611 = n50608 & n50610 ;
  assign n50612 = n11386 & n11989 ;
  assign n50613 = n50612 ^ n14316 ^ 1'b0 ;
  assign n50614 = n24347 & n50613 ;
  assign n50615 = ~n4100 & n50614 ;
  assign n50616 = n15090 ^ n9373 ^ 1'b0 ;
  assign n50617 = n9663 | n50616 ;
  assign n50618 = ( n3103 & n5406 ) | ( n3103 & ~n22519 ) | ( n5406 & ~n22519 ) ;
  assign n50619 = n8495 & ~n50618 ;
  assign n50620 = n50619 ^ n10820 ^ 1'b0 ;
  assign n50623 = n12469 ^ n9920 ^ 1'b0 ;
  assign n50621 = n10060 ^ n10043 ^ n5920 ;
  assign n50622 = ( n4094 & n9609 ) | ( n4094 & ~n50621 ) | ( n9609 & ~n50621 ) ;
  assign n50624 = n50623 ^ n50622 ^ n6381 ;
  assign n50625 = n32555 ^ n26902 ^ n8577 ;
  assign n50626 = ( n475 & n4225 ) | ( n475 & n5745 ) | ( n4225 & n5745 ) ;
  assign n50627 = n33933 ^ n8570 ^ n4931 ;
  assign n50628 = ( n37065 & ~n50626 ) | ( n37065 & n50627 ) | ( ~n50626 & n50627 ) ;
  assign n50629 = n50628 ^ n11831 ^ n5344 ;
  assign n50630 = n3951 | n19200 ;
  assign n50631 = n33669 | n41575 ;
  assign n50632 = n39432 | n50631 ;
  assign n50633 = n50632 ^ n26179 ^ n10980 ;
  assign n50634 = n50633 ^ n40801 ^ 1'b0 ;
  assign n50635 = n4029 ^ n2605 ^ 1'b0 ;
  assign n50636 = n38464 & n50635 ;
  assign n50637 = ( n32393 & ~n39928 ) | ( n32393 & n50636 ) | ( ~n39928 & n50636 ) ;
  assign n50638 = n50637 ^ n17536 ^ n16500 ;
  assign n50639 = n45231 & n46415 ;
  assign n50640 = n11586 ^ n8915 ^ n751 ;
  assign n50641 = n50640 ^ n13807 ^ 1'b0 ;
  assign n50642 = n50639 & ~n50641 ;
  assign n50643 = n4448 & ~n14161 ;
  assign n50644 = n11493 & n50643 ;
  assign n50645 = n16768 ^ n9107 ^ 1'b0 ;
  assign n50646 = n25825 ^ n8537 ^ 1'b0 ;
  assign n50647 = n50646 ^ n26941 ^ n7132 ;
  assign n50648 = ( ~n6834 & n17074 ) | ( ~n6834 & n47029 ) | ( n17074 & n47029 ) ;
  assign n50649 = n21622 ^ n5924 ^ n2186 ;
  assign n50650 = n31490 ^ n29836 ^ 1'b0 ;
  assign n50651 = n2802 & n50650 ;
  assign n50652 = n50651 ^ n9230 ^ 1'b0 ;
  assign n50653 = n50652 ^ n29790 ^ n7306 ;
  assign n50654 = n42718 ^ n3009 ^ 1'b0 ;
  assign n50655 = ~n30553 & n50654 ;
  assign n50656 = n585 & ~n5502 ;
  assign n50657 = n2818 & n12592 ;
  assign n50658 = n50657 ^ n5056 ^ 1'b0 ;
  assign n50659 = n50658 ^ n28149 ^ n27584 ;
  assign n50660 = ( n38995 & ~n39081 ) | ( n38995 & n50659 ) | ( ~n39081 & n50659 ) ;
  assign n50663 = n8910 ^ n747 ^ 1'b0 ;
  assign n50664 = n23395 & ~n50663 ;
  assign n50662 = ( n5725 & ~n11359 ) | ( n5725 & n34290 ) | ( ~n11359 & n34290 ) ;
  assign n50661 = n40578 ^ n24723 ^ x70 ;
  assign n50665 = n50664 ^ n50662 ^ n50661 ;
  assign n50666 = n50665 ^ n12386 ^ n9148 ;
  assign n50667 = ( ~n6405 & n15884 ) | ( ~n6405 & n20311 ) | ( n15884 & n20311 ) ;
  assign n50668 = ( n17245 & n25556 ) | ( n17245 & ~n50667 ) | ( n25556 & ~n50667 ) ;
  assign n50669 = ( n1722 & ~n7236 ) | ( n1722 & n13838 ) | ( ~n7236 & n13838 ) ;
  assign n50670 = n50669 ^ n21232 ^ n13314 ;
  assign n50671 = ( ~n3296 & n16326 ) | ( ~n3296 & n48435 ) | ( n16326 & n48435 ) ;
  assign n50672 = n50671 ^ n19679 ^ n14017 ;
  assign n50674 = ( n10742 & n11895 ) | ( n10742 & ~n12695 ) | ( n11895 & ~n12695 ) ;
  assign n50673 = n17369 ^ n16780 ^ 1'b0 ;
  assign n50675 = n50674 ^ n50673 ^ n40057 ;
  assign n50676 = n4890 & n13106 ;
  assign n50677 = n8238 & n30988 ;
  assign n50678 = n50677 ^ n326 ^ 1'b0 ;
  assign n50679 = n36491 ^ n13631 ^ n5604 ;
  assign n50682 = n4282 & ~n9509 ;
  assign n50683 = n50682 ^ n30877 ^ 1'b0 ;
  assign n50680 = n42049 ^ n1774 ^ 1'b0 ;
  assign n50681 = n2336 & ~n50680 ;
  assign n50684 = n50683 ^ n50681 ^ 1'b0 ;
  assign n50685 = n50679 & ~n50684 ;
  assign n50686 = ~n14418 & n42381 ;
  assign n50687 = ( n7211 & n12473 ) | ( n7211 & n22881 ) | ( n12473 & n22881 ) ;
  assign n50688 = n40141 | n50687 ;
  assign n50689 = n50688 ^ n9247 ^ 1'b0 ;
  assign n50690 = n40835 & ~n50689 ;
  assign n50691 = n16252 | n50690 ;
  assign n50692 = ( n8886 & ~n14343 ) | ( n8886 & n23085 ) | ( ~n14343 & n23085 ) ;
  assign n50693 = ( n4850 & n6290 ) | ( n4850 & ~n50692 ) | ( n6290 & ~n50692 ) ;
  assign n50694 = ( n18069 & n42306 ) | ( n18069 & ~n50693 ) | ( n42306 & ~n50693 ) ;
  assign n50695 = ( n5435 & n6060 ) | ( n5435 & n22048 ) | ( n6060 & n22048 ) ;
  assign n50696 = n48805 ^ n39737 ^ n39442 ;
  assign n50697 = n36025 & ~n50696 ;
  assign n50698 = n4600 ^ n2206 ^ 1'b0 ;
  assign n50699 = ~n40739 & n50698 ;
  assign n50700 = n50699 ^ n42355 ^ n12307 ;
  assign n50701 = n35471 ^ n16172 ^ 1'b0 ;
  assign n50702 = n14145 & ~n50701 ;
  assign n50703 = n50702 ^ n16064 ^ 1'b0 ;
  assign n50704 = n41179 ^ n33846 ^ n5997 ;
  assign n50705 = ~n27562 & n50704 ;
  assign n50706 = n50705 ^ n22949 ^ 1'b0 ;
  assign n50707 = n42793 ^ n30401 ^ n14508 ;
  assign n50708 = ~n3657 & n27771 ;
  assign n50709 = n2435 & n50708 ;
  assign n50710 = n50707 & n50709 ;
  assign n50711 = n3304 ^ x99 ^ 1'b0 ;
  assign n50712 = ( ~n6871 & n7228 ) | ( ~n6871 & n50711 ) | ( n7228 & n50711 ) ;
  assign n50713 = ( ~n12206 & n23883 ) | ( ~n12206 & n50712 ) | ( n23883 & n50712 ) ;
  assign n50715 = n32676 ^ n21236 ^ n1265 ;
  assign n50714 = n22169 ^ n3138 ^ 1'b0 ;
  assign n50716 = n50715 ^ n50714 ^ n48135 ;
  assign n50718 = n4469 | n12781 ;
  assign n50719 = n50718 ^ n3948 ^ 1'b0 ;
  assign n50717 = n34480 ^ n18471 ^ n326 ;
  assign n50720 = n50719 ^ n50717 ^ n19197 ;
  assign n50721 = n46049 ^ n8253 ^ 1'b0 ;
  assign n50722 = n5966 & ~n8426 ;
  assign n50723 = n50722 ^ n30054 ^ n12220 ;
  assign n50724 = n2046 ^ n692 ^ 1'b0 ;
  assign n50725 = ~n42743 & n50724 ;
  assign n50726 = n50725 ^ n30735 ^ n1337 ;
  assign n50727 = ( ~n5561 & n6537 ) | ( ~n5561 & n18131 ) | ( n6537 & n18131 ) ;
  assign n50728 = n50727 ^ n15677 ^ n8651 ;
  assign n50729 = n50728 ^ n28187 ^ n19937 ;
  assign n50730 = n10620 & ~n44781 ;
  assign n50731 = n50730 ^ n47324 ^ 1'b0 ;
  assign n50732 = ( ~n26502 & n39439 ) | ( ~n26502 & n50731 ) | ( n39439 & n50731 ) ;
  assign n50733 = ~n38811 & n50732 ;
  assign n50734 = ~n28713 & n50733 ;
  assign n50737 = n6239 ^ n3281 ^ n2822 ;
  assign n50735 = n41670 ^ n40544 ^ 1'b0 ;
  assign n50736 = n43791 | n50735 ;
  assign n50738 = n50737 ^ n50736 ^ 1'b0 ;
  assign n50739 = n24239 ^ n16097 ^ n2670 ;
  assign n50740 = ( n2528 & n32504 ) | ( n2528 & n35659 ) | ( n32504 & n35659 ) ;
  assign n50741 = n5447 ^ n4651 ^ 1'b0 ;
  assign n50742 = ( ~n8301 & n25543 ) | ( ~n8301 & n35741 ) | ( n25543 & n35741 ) ;
  assign n50743 = ( n10951 & n50741 ) | ( n10951 & n50742 ) | ( n50741 & n50742 ) ;
  assign n50744 = ( ~n22539 & n30334 ) | ( ~n22539 & n39993 ) | ( n30334 & n39993 ) ;
  assign n50745 = ( n5290 & ~n7007 ) | ( n5290 & n43802 ) | ( ~n7007 & n43802 ) ;
  assign n50746 = n45269 ^ n25305 ^ n7181 ;
  assign n50747 = n50746 ^ n49918 ^ n9479 ;
  assign n50748 = n20043 | n44294 ;
  assign n50749 = n32414 & ~n50748 ;
  assign n50750 = n18681 ^ n13268 ^ 1'b0 ;
  assign n50751 = n868 & n30191 ;
  assign n50752 = n50751 ^ n8570 ^ 1'b0 ;
  assign n50753 = n20293 & n30981 ;
  assign n50754 = n20554 ^ n10531 ^ 1'b0 ;
  assign n50755 = n50754 ^ n14377 ^ n4539 ;
  assign n50756 = n24685 ^ n8750 ^ n5693 ;
  assign n50757 = ( n2777 & n32556 ) | ( n2777 & n50756 ) | ( n32556 & n50756 ) ;
  assign n50758 = n37787 & ~n49390 ;
  assign n50759 = n48111 ^ n16897 ^ n8113 ;
  assign n50760 = n50759 ^ n12016 ^ n933 ;
  assign n50761 = n50760 ^ n19212 ^ n16490 ;
  assign n50762 = n12025 & n43569 ;
  assign n50763 = ~n39191 & n50762 ;
  assign n50764 = ( n643 & n1345 ) | ( n643 & ~n26412 ) | ( n1345 & ~n26412 ) ;
  assign n50765 = ~n4070 & n50764 ;
  assign n50766 = ( n2408 & n50763 ) | ( n2408 & n50765 ) | ( n50763 & n50765 ) ;
  assign n50767 = n31813 ^ n3035 ^ 1'b0 ;
  assign n50768 = ( n1383 & n31740 ) | ( n1383 & ~n50767 ) | ( n31740 & ~n50767 ) ;
  assign n50769 = ~n4068 & n21994 ;
  assign n50770 = n50769 ^ n25509 ^ n5823 ;
  assign n50771 = n50770 ^ n33142 ^ n9570 ;
  assign n50772 = x214 & ~n33681 ;
  assign n50773 = n2427 | n26770 ;
  assign n50774 = n17127 | n26590 ;
  assign n50775 = n14011 & ~n50774 ;
  assign n50776 = n2512 & ~n26608 ;
  assign n50777 = n50776 ^ n15421 ^ 1'b0 ;
  assign n50778 = ( n8874 & n15148 ) | ( n8874 & n44172 ) | ( n15148 & n44172 ) ;
  assign n50779 = n34916 ^ n23325 ^ 1'b0 ;
  assign n50780 = n38655 ^ n36304 ^ n33371 ;
  assign n50785 = n1044 & ~n11443 ;
  assign n50783 = n24190 ^ n16037 ^ n10933 ;
  assign n50781 = ( n7615 & ~n14436 ) | ( n7615 & n50460 ) | ( ~n14436 & n50460 ) ;
  assign n50782 = n50781 ^ n32469 ^ n21015 ;
  assign n50784 = n50783 ^ n50782 ^ n33610 ;
  assign n50786 = n50785 ^ n50784 ^ n38648 ;
  assign n50787 = ( x233 & ~n4606 ) | ( x233 & n4832 ) | ( ~n4606 & n4832 ) ;
  assign n50788 = ( n312 & ~n4680 ) | ( n312 & n23594 ) | ( ~n4680 & n23594 ) ;
  assign n50789 = n50788 ^ n3620 ^ 1'b0 ;
  assign n50791 = n41220 ^ n30158 ^ n23082 ;
  assign n50792 = n1067 & n50791 ;
  assign n50793 = n50792 ^ n17350 ^ 1'b0 ;
  assign n50790 = n9271 | n37509 ;
  assign n50794 = n50793 ^ n50790 ^ 1'b0 ;
  assign n50795 = ~n10230 & n13526 ;
  assign n50796 = n45211 & n50795 ;
  assign n50797 = n27767 ^ n20280 ^ 1'b0 ;
  assign n50798 = n44334 & n50797 ;
  assign n50799 = n45861 ^ n25635 ^ n6743 ;
  assign n50800 = n36629 ^ n11236 ^ 1'b0 ;
  assign n50801 = ~n1457 & n50800 ;
  assign n50802 = ( n10442 & n17591 ) | ( n10442 & ~n50801 ) | ( n17591 & ~n50801 ) ;
  assign n50803 = ~n2289 & n43168 ;
  assign n50804 = ~n2021 & n50803 ;
  assign n50805 = ( ~n40532 & n46764 ) | ( ~n40532 & n50804 ) | ( n46764 & n50804 ) ;
  assign n50806 = n49223 ^ n4614 ^ 1'b0 ;
  assign n50807 = n22402 & ~n50806 ;
  assign n50808 = ( n17363 & ~n50173 ) | ( n17363 & n50807 ) | ( ~n50173 & n50807 ) ;
  assign n50810 = n14290 ^ n6067 ^ n4520 ;
  assign n50809 = ( n12614 & ~n37953 ) | ( n12614 & n49010 ) | ( ~n37953 & n49010 ) ;
  assign n50811 = n50810 ^ n50809 ^ n17437 ;
  assign n50814 = ~n3164 & n9163 ;
  assign n50812 = n18944 ^ n1405 ^ 1'b0 ;
  assign n50813 = n15961 & n50812 ;
  assign n50815 = n50814 ^ n50813 ^ 1'b0 ;
  assign n50816 = n50815 ^ n42326 ^ n25950 ;
  assign n50817 = n30952 ^ n13150 ^ n9135 ;
  assign n50818 = ~n35469 & n50817 ;
  assign n50819 = n45184 ^ n12237 ^ 1'b0 ;
  assign n50820 = n50818 | n50819 ;
  assign n50821 = n5574 | n5670 ;
  assign n50822 = n36023 | n50821 ;
  assign n50823 = ( ~n2296 & n17609 ) | ( ~n2296 & n39670 ) | ( n17609 & n39670 ) ;
  assign n50824 = ( n393 & ~n35533 ) | ( n393 & n45177 ) | ( ~n35533 & n45177 ) ;
  assign n50825 = ~n13771 & n20416 ;
  assign n50826 = n41324 & ~n50825 ;
  assign n50827 = n41804 ^ n12843 ^ n7140 ;
  assign n50828 = n16782 ^ n12945 ^ x140 ;
  assign n50829 = ( n15558 & n46909 ) | ( n15558 & ~n50828 ) | ( n46909 & ~n50828 ) ;
  assign n50830 = ~n4333 & n6144 ;
  assign n50831 = ~n20536 & n50830 ;
  assign n50832 = n50831 ^ n19712 ^ 1'b0 ;
  assign n50833 = ~n2779 & n15898 ;
  assign n50834 = n50833 ^ n7553 ^ 1'b0 ;
  assign n50835 = n6391 & n30456 ;
  assign n50836 = ~n15898 & n50835 ;
  assign n50837 = ( n1461 & n15776 ) | ( n1461 & n33957 ) | ( n15776 & n33957 ) ;
  assign n50838 = n45607 ^ n35582 ^ 1'b0 ;
  assign n50839 = n8977 & ~n50838 ;
  assign n50840 = ( n22401 & n50837 ) | ( n22401 & ~n50839 ) | ( n50837 & ~n50839 ) ;
  assign n50841 = ( n20927 & n22246 ) | ( n20927 & n22589 ) | ( n22246 & n22589 ) ;
  assign n50842 = n3767 ^ n1091 ^ 1'b0 ;
  assign n50843 = n11424 & n50842 ;
  assign n50844 = n48026 & n50843 ;
  assign n50845 = ( n14967 & n30295 ) | ( n14967 & ~n32702 ) | ( n30295 & ~n32702 ) ;
  assign n50846 = n18372 | n50845 ;
  assign n50847 = n46930 ^ n37355 ^ 1'b0 ;
  assign n50848 = ~n1848 & n50847 ;
  assign n50849 = n50848 ^ n50338 ^ n16568 ;
  assign n50850 = ~n6907 & n10325 ;
  assign n50851 = ( n4381 & n47668 ) | ( n4381 & ~n50850 ) | ( n47668 & ~n50850 ) ;
  assign n50852 = n9534 | n13502 ;
  assign n50853 = ( n6768 & ~n13577 ) | ( n6768 & n50852 ) | ( ~n13577 & n50852 ) ;
  assign n50854 = n41324 ^ n29810 ^ n7510 ;
  assign n50855 = n50854 ^ n26511 ^ n21719 ;
  assign n50856 = ( n12103 & n19748 ) | ( n12103 & ~n38549 ) | ( n19748 & ~n38549 ) ;
  assign n50857 = n40572 ^ n31869 ^ n2703 ;
  assign n50859 = n34757 ^ n15149 ^ 1'b0 ;
  assign n50858 = ~n45590 & n45649 ;
  assign n50860 = n50859 ^ n50858 ^ n8592 ;
  assign n50861 = n16762 ^ n9334 ^ 1'b0 ;
  assign n50862 = n2846 & n50861 ;
  assign n50863 = n48048 ^ n22450 ^ 1'b0 ;
  assign n50864 = n11684 | n50863 ;
  assign n50865 = ( n37811 & n50862 ) | ( n37811 & n50864 ) | ( n50862 & n50864 ) ;
  assign n50866 = ~n4633 & n25423 ;
  assign n50867 = ~n37841 & n50866 ;
  assign n50868 = n14699 ^ n3999 ^ 1'b0 ;
  assign n50869 = n24361 & ~n50868 ;
  assign n50871 = n5846 | n27822 ;
  assign n50872 = ~n21042 & n50871 ;
  assign n50870 = n47971 | n48676 ;
  assign n50873 = n50872 ^ n50870 ^ 1'b0 ;
  assign n50874 = n27572 ^ n24232 ^ 1'b0 ;
  assign n50875 = n50874 ^ n35532 ^ n380 ;
  assign n50876 = n15851 ^ n8468 ^ n7141 ;
  assign n50877 = ( n22614 & n50875 ) | ( n22614 & n50876 ) | ( n50875 & n50876 ) ;
  assign n50878 = n50877 ^ n8171 ^ 1'b0 ;
  assign n50879 = n23322 | n50878 ;
  assign n50880 = ( n961 & ~n28565 ) | ( n961 & n44801 ) | ( ~n28565 & n44801 ) ;
  assign n50881 = n50880 ^ n46284 ^ n36184 ;
  assign n50882 = ( n8099 & n48383 ) | ( n8099 & ~n50881 ) | ( n48383 & ~n50881 ) ;
  assign n50883 = ~n27676 & n42581 ;
  assign n50884 = ( n375 & n33984 ) | ( n375 & ~n50883 ) | ( n33984 & ~n50883 ) ;
  assign n50885 = n48551 ^ n20737 ^ n16621 ;
  assign n50891 = ~n5463 & n25806 ;
  assign n50886 = x203 & ~n6048 ;
  assign n50887 = ~n10202 & n11055 ;
  assign n50888 = n17787 & ~n50887 ;
  assign n50889 = n50888 ^ n8603 ^ 1'b0 ;
  assign n50890 = ( n31705 & n50886 ) | ( n31705 & n50889 ) | ( n50886 & n50889 ) ;
  assign n50892 = n50891 ^ n50890 ^ n42659 ;
  assign n50893 = ( x220 & ~n11016 ) | ( x220 & n37226 ) | ( ~n11016 & n37226 ) ;
  assign n50894 = ( n2666 & n30665 ) | ( n2666 & ~n50893 ) | ( n30665 & ~n50893 ) ;
  assign n50895 = n26902 ^ n16704 ^ 1'b0 ;
  assign n50896 = ( n10747 & n19891 ) | ( n10747 & n48010 ) | ( n19891 & n48010 ) ;
  assign n50897 = n44272 ^ n12616 ^ 1'b0 ;
  assign n50898 = n35307 | n50897 ;
  assign n50899 = ( n16416 & n28265 ) | ( n16416 & ~n36559 ) | ( n28265 & ~n36559 ) ;
  assign n50900 = ( ~n2408 & n22648 ) | ( ~n2408 & n50899 ) | ( n22648 & n50899 ) ;
  assign n50901 = n50900 ^ n44980 ^ 1'b0 ;
  assign n50902 = n46772 | n50901 ;
  assign n50903 = n9247 ^ n4982 ^ 1'b0 ;
  assign n50904 = n25583 ^ n2420 ^ 1'b0 ;
  assign n50905 = n50904 ^ n50396 ^ n15990 ;
  assign n50906 = ( n8539 & n34302 ) | ( n8539 & n42820 ) | ( n34302 & n42820 ) ;
  assign n50907 = n46453 ^ n29315 ^ n6053 ;
  assign n50908 = ( n6016 & n15396 ) | ( n6016 & ~n50907 ) | ( n15396 & ~n50907 ) ;
  assign n50909 = n12685 ^ n11526 ^ 1'b0 ;
  assign n50911 = ( ~n1891 & n12489 ) | ( ~n1891 & n22422 ) | ( n12489 & n22422 ) ;
  assign n50910 = ( n7747 & ~n22396 ) | ( n7747 & n27650 ) | ( ~n22396 & n27650 ) ;
  assign n50912 = n50911 ^ n50910 ^ n33822 ;
  assign n50913 = ( n20599 & n48576 ) | ( n20599 & n50912 ) | ( n48576 & n50912 ) ;
  assign n50914 = n12920 ^ n2728 ^ x172 ;
  assign n50915 = ( n7649 & ~n28889 ) | ( n7649 & n50914 ) | ( ~n28889 & n50914 ) ;
  assign n50916 = n50915 ^ n4800 ^ n831 ;
  assign n50917 = n17793 | n42055 ;
  assign n50921 = n39153 ^ n9496 ^ n4299 ;
  assign n50918 = n26451 ^ n18452 ^ 1'b0 ;
  assign n50919 = n5240 & n50918 ;
  assign n50920 = ~n11855 & n50919 ;
  assign n50922 = n50921 ^ n50920 ^ 1'b0 ;
  assign n50923 = n50922 ^ n15161 ^ 1'b0 ;
  assign n50924 = n48653 ^ n19136 ^ 1'b0 ;
  assign n50925 = n20672 ^ n15729 ^ 1'b0 ;
  assign n50926 = ~n16087 & n50925 ;
  assign n50927 = n27079 ^ n9518 ^ n8169 ;
  assign n50928 = n48011 ^ n12258 ^ 1'b0 ;
  assign n50929 = n23818 ^ n2011 ^ 1'b0 ;
  assign n50931 = ( n4057 & n17015 ) | ( n4057 & ~n46151 ) | ( n17015 & ~n46151 ) ;
  assign n50930 = ~n2931 & n26430 ;
  assign n50932 = n50931 ^ n50930 ^ 1'b0 ;
  assign n50933 = n50932 ^ n2455 ^ 1'b0 ;
  assign n50934 = n13661 & n50933 ;
  assign n50942 = n47533 ^ n7088 ^ n2282 ;
  assign n50937 = n35776 ^ n22949 ^ 1'b0 ;
  assign n50938 = n21638 | n50937 ;
  assign n50939 = ( ~n3510 & n15042 ) | ( ~n3510 & n50938 ) | ( n15042 & n50938 ) ;
  assign n50940 = n50939 ^ n43342 ^ n8190 ;
  assign n50935 = n16881 ^ n12135 ^ n3505 ;
  assign n50936 = ( n23539 & n41963 ) | ( n23539 & n50935 ) | ( n41963 & n50935 ) ;
  assign n50941 = n50940 ^ n50936 ^ 1'b0 ;
  assign n50943 = n50942 ^ n50941 ^ n40166 ;
  assign n50944 = n35134 ^ n34191 ^ n13243 ;
  assign n50945 = n50944 ^ n6392 ^ n5305 ;
  assign n50946 = n44567 ^ n1417 ^ x220 ;
  assign n50947 = ( n12391 & n25082 ) | ( n12391 & n50946 ) | ( n25082 & n50946 ) ;
  assign n50948 = n50947 ^ n23896 ^ 1'b0 ;
  assign n50949 = n17265 ^ n3892 ^ 1'b0 ;
  assign n50950 = n7342 | n50949 ;
  assign n50951 = n7495 & ~n21654 ;
  assign n50952 = n50951 ^ n7599 ^ 1'b0 ;
  assign n50953 = n13666 | n50952 ;
  assign n50954 = n8212 ^ n1321 ^ 1'b0 ;
  assign n50955 = ( n20291 & ~n23909 ) | ( n20291 & n39547 ) | ( ~n23909 & n39547 ) ;
  assign n50956 = n50955 ^ n44079 ^ 1'b0 ;
  assign n50957 = ( n3185 & ~n4181 ) | ( n3185 & n25620 ) | ( ~n4181 & n25620 ) ;
  assign n50958 = ( ~n7708 & n23968 ) | ( ~n7708 & n50957 ) | ( n23968 & n50957 ) ;
  assign n50959 = n23829 ^ n21976 ^ n12188 ;
  assign n50960 = ( n26473 & ~n42836 ) | ( n26473 & n50959 ) | ( ~n42836 & n50959 ) ;
  assign n50961 = ( ~n12040 & n28621 ) | ( ~n12040 & n38625 ) | ( n28621 & n38625 ) ;
  assign n50962 = ( n4326 & ~n6528 ) | ( n4326 & n38135 ) | ( ~n6528 & n38135 ) ;
  assign n50963 = ( n9505 & n11782 ) | ( n9505 & n13251 ) | ( n11782 & n13251 ) ;
  assign n50964 = n6018 ^ x6 ^ 1'b0 ;
  assign n50965 = n8684 & n50964 ;
  assign n50966 = n50965 ^ n6159 ^ 1'b0 ;
  assign n50967 = ( n773 & ~n6676 ) | ( n773 & n28959 ) | ( ~n6676 & n28959 ) ;
  assign n50968 = ( n12211 & n13038 ) | ( n12211 & n50967 ) | ( n13038 & n50967 ) ;
  assign n50969 = ( n1860 & ~n32312 ) | ( n1860 & n38293 ) | ( ~n32312 & n38293 ) ;
  assign n50970 = ( n50966 & ~n50968 ) | ( n50966 & n50969 ) | ( ~n50968 & n50969 ) ;
  assign n50971 = n16673 & n19983 ;
  assign n50972 = n50971 ^ n13512 ^ 1'b0 ;
  assign n50974 = n9888 ^ n5814 ^ n5425 ;
  assign n50975 = n50974 ^ n17521 ^ n696 ;
  assign n50976 = ( n5770 & n19981 ) | ( n5770 & n50975 ) | ( n19981 & n50975 ) ;
  assign n50973 = n1967 & n2531 ;
  assign n50977 = n50976 ^ n50973 ^ 1'b0 ;
  assign n50978 = ( n1911 & n9239 ) | ( n1911 & n44210 ) | ( n9239 & n44210 ) ;
  assign n50979 = n6760 ^ n2158 ^ 1'b0 ;
  assign n50980 = n860 & ~n50979 ;
  assign n50981 = n50980 ^ n32013 ^ n6911 ;
  assign n50982 = ( ~n36759 & n50978 ) | ( ~n36759 & n50981 ) | ( n50978 & n50981 ) ;
  assign n50983 = n1437 | n9515 ;
  assign n50984 = n24186 | n50983 ;
  assign n50985 = ( n26824 & ~n46993 ) | ( n26824 & n50984 ) | ( ~n46993 & n50984 ) ;
  assign n50986 = ( n2438 & n9177 ) | ( n2438 & n28277 ) | ( n9177 & n28277 ) ;
  assign n50987 = n50986 ^ n27705 ^ 1'b0 ;
  assign n50988 = ( n544 & ~n5678 ) | ( n544 & n13118 ) | ( ~n5678 & n13118 ) ;
  assign n50989 = n21570 ^ n4579 ^ 1'b0 ;
  assign n50990 = n50988 & ~n50989 ;
  assign n50991 = ( n5761 & n16189 ) | ( n5761 & n30734 ) | ( n16189 & n30734 ) ;
  assign n50992 = n48463 ^ n29852 ^ 1'b0 ;
  assign n50993 = ( n4486 & n50991 ) | ( n4486 & ~n50992 ) | ( n50991 & ~n50992 ) ;
  assign n50994 = n50993 ^ n45721 ^ n14688 ;
  assign n50995 = n26889 ^ n12192 ^ 1'b0 ;
  assign n50996 = n50995 ^ n41324 ^ n25527 ;
  assign n50997 = n14685 | n50623 ;
  assign n50998 = n1680 & ~n50997 ;
  assign n50999 = n50998 ^ n41982 ^ 1'b0 ;
  assign n51000 = n39934 ^ n13961 ^ n12954 ;
  assign n51001 = n22747 | n51000 ;
  assign n51002 = n5429 & ~n51001 ;
  assign n51003 = n18593 ^ n1883 ^ 1'b0 ;
  assign n51004 = ( n15191 & n18067 ) | ( n15191 & n51003 ) | ( n18067 & n51003 ) ;
  assign n51007 = ( ~n2364 & n3883 ) | ( ~n2364 & n7819 ) | ( n3883 & n7819 ) ;
  assign n51005 = ~n10469 & n33529 ;
  assign n51006 = n41031 & n51005 ;
  assign n51008 = n51007 ^ n51006 ^ 1'b0 ;
  assign n51009 = ( n10310 & n11064 ) | ( n10310 & ~n46966 ) | ( n11064 & ~n46966 ) ;
  assign n51010 = ( ~n8075 & n48238 ) | ( ~n8075 & n51009 ) | ( n48238 & n51009 ) ;
  assign n51011 = n20047 ^ n3006 ^ n2570 ;
  assign n51012 = n51011 ^ n15464 ^ n5562 ;
  assign n51013 = n32912 ^ n30348 ^ n4126 ;
  assign n51015 = n20058 | n23835 ;
  assign n51014 = n44920 ^ n19780 ^ n13058 ;
  assign n51016 = n51015 ^ n51014 ^ n49950 ;
  assign n51017 = n4116 | n43988 ;
  assign n51018 = n51017 ^ n30922 ^ n14376 ;
  assign n51019 = n20378 | n31226 ;
  assign n51020 = n51019 ^ n40082 ^ 1'b0 ;
  assign n51021 = n20206 ^ n13226 ^ n5811 ;
  assign n51022 = ( n5189 & n9041 ) | ( n5189 & n51021 ) | ( n9041 & n51021 ) ;
  assign n51023 = n51022 ^ n41351 ^ 1'b0 ;
  assign n51024 = n51023 ^ n2869 ^ 1'b0 ;
  assign n51025 = x99 & ~n51024 ;
  assign n51026 = n13737 | n17858 ;
  assign n51027 = n1839 & ~n51026 ;
  assign n51028 = n51027 ^ n43242 ^ n2432 ;
  assign n51029 = ( n11817 & n36369 ) | ( n11817 & n51028 ) | ( n36369 & n51028 ) ;
  assign n51030 = ( ~n21723 & n21883 ) | ( ~n21723 & n40456 ) | ( n21883 & n40456 ) ;
  assign n51031 = n51030 ^ n27604 ^ 1'b0 ;
  assign n51032 = ( n7525 & n10178 ) | ( n7525 & ~n23573 ) | ( n10178 & ~n23573 ) ;
  assign n51033 = n44956 ^ n23152 ^ n7623 ;
  assign n51034 = ( n5141 & n14420 ) | ( n5141 & n17614 ) | ( n14420 & n17614 ) ;
  assign n51035 = ~n875 & n21458 ;
  assign n51036 = n51034 & n51035 ;
  assign n51037 = n51036 ^ n29356 ^ 1'b0 ;
  assign n51038 = n9840 ^ n7995 ^ n575 ;
  assign n51039 = n853 & ~n5074 ;
  assign n51040 = n4808 & n51039 ;
  assign n51041 = n51040 ^ n41633 ^ n14311 ;
  assign n51042 = ( n6024 & ~n8747 ) | ( n6024 & n27762 ) | ( ~n8747 & n27762 ) ;
  assign n51043 = n39572 ^ n17850 ^ 1'b0 ;
  assign n51044 = ~n20580 & n51043 ;
  assign n51045 = ( n51041 & n51042 ) | ( n51041 & ~n51044 ) | ( n51042 & ~n51044 ) ;
  assign n51046 = n2905 | n51045 ;
  assign n51047 = n24692 & ~n51046 ;
  assign n51048 = n14900 & ~n30893 ;
  assign n51049 = n40133 ^ n801 ^ 1'b0 ;
  assign n51050 = ( n21367 & n50914 ) | ( n21367 & ~n51049 ) | ( n50914 & ~n51049 ) ;
  assign n51051 = n29125 ^ n23082 ^ n14654 ;
  assign n51052 = n754 & n23538 ;
  assign n51053 = ~n7237 & n51052 ;
  assign n51054 = n51053 ^ n21606 ^ 1'b0 ;
  assign n51055 = ( n3963 & n51051 ) | ( n3963 & n51054 ) | ( n51051 & n51054 ) ;
  assign n51056 = n34762 ^ n12443 ^ 1'b0 ;
  assign n51057 = ( ~n31559 & n40294 ) | ( ~n31559 & n48493 ) | ( n40294 & n48493 ) ;
  assign n51058 = n11434 ^ n8087 ^ n5261 ;
  assign n51059 = ( n3851 & n4815 ) | ( n3851 & ~n51058 ) | ( n4815 & ~n51058 ) ;
  assign n51060 = ~n5459 & n47598 ;
  assign n51061 = n3018 & n51060 ;
  assign n51062 = n31211 ^ n1472 ^ 1'b0 ;
  assign n51063 = n5431 | n7878 ;
  assign n51067 = n16609 & n48441 ;
  assign n51065 = ( ~n1822 & n2593 ) | ( ~n1822 & n19352 ) | ( n2593 & n19352 ) ;
  assign n51064 = n29612 ^ n15658 ^ n8156 ;
  assign n51066 = n51065 ^ n51064 ^ n15084 ;
  assign n51068 = n51067 ^ n51066 ^ n724 ;
  assign n51069 = n26009 | n42964 ;
  assign n51070 = ( n1976 & ~n2283 ) | ( n1976 & n15674 ) | ( ~n2283 & n15674 ) ;
  assign n51071 = ( n9050 & n51069 ) | ( n9050 & n51070 ) | ( n51069 & n51070 ) ;
  assign n51072 = n15866 ^ n5074 ^ 1'b0 ;
  assign n51073 = ~n9145 & n51072 ;
  assign n51074 = n51073 ^ n47169 ^ 1'b0 ;
  assign n51075 = n51074 ^ n47339 ^ n15773 ;
  assign n51076 = ( n3206 & ~n12207 ) | ( n3206 & n27761 ) | ( ~n12207 & n27761 ) ;
  assign n51077 = ( n3077 & n24194 ) | ( n3077 & n51076 ) | ( n24194 & n51076 ) ;
  assign n51078 = n2116 | n43508 ;
  assign n51079 = ( n9737 & ~n51077 ) | ( n9737 & n51078 ) | ( ~n51077 & n51078 ) ;
  assign n51080 = ( n12855 & n16019 ) | ( n12855 & n22835 ) | ( n16019 & n22835 ) ;
  assign n51081 = ~n13083 & n51080 ;
  assign n51082 = n51081 ^ n44994 ^ 1'b0 ;
  assign n51083 = n6947 & n32841 ;
  assign n51084 = n51083 ^ n25636 ^ 1'b0 ;
  assign n51085 = n24878 ^ n23058 ^ 1'b0 ;
  assign n51086 = n46300 ^ n30595 ^ 1'b0 ;
  assign n51087 = ~n46623 & n51086 ;
  assign n51088 = ( n3557 & ~n28544 ) | ( n3557 & n43187 ) | ( ~n28544 & n43187 ) ;
  assign n51089 = ( n13035 & n15895 ) | ( n13035 & n41340 ) | ( n15895 & n41340 ) ;
  assign n51090 = n12040 & ~n46902 ;
  assign n51091 = ~n51089 & n51090 ;
  assign n51092 = n51091 ^ n37042 ^ n33564 ;
  assign n51093 = n25889 ^ n13250 ^ n7871 ;
  assign n51094 = n51093 ^ n27746 ^ n17107 ;
  assign n51095 = n51094 ^ n33426 ^ n25064 ;
  assign n51096 = n5378 & n12870 ;
  assign n51097 = ~n3557 & n51096 ;
  assign n51098 = n41085 ^ n15182 ^ n6060 ;
  assign n51099 = ~n8852 & n28166 ;
  assign n51100 = n51099 ^ n32243 ^ 1'b0 ;
  assign n51102 = n5916 ^ n3614 ^ 1'b0 ;
  assign n51101 = n21305 ^ n14763 ^ n911 ;
  assign n51103 = n51102 ^ n51101 ^ n34109 ;
  assign n51104 = ~n30456 & n51103 ;
  assign n51105 = ( n14419 & n25130 ) | ( n14419 & n40656 ) | ( n25130 & n40656 ) ;
  assign n51106 = n34776 ^ n5164 ^ n4557 ;
  assign n51107 = n5847 ^ n959 ^ 1'b0 ;
  assign n51108 = n51107 ^ n26188 ^ n23151 ;
  assign n51110 = ( n1358 & n15452 ) | ( n1358 & ~n34665 ) | ( n15452 & ~n34665 ) ;
  assign n51109 = n44641 ^ n20876 ^ 1'b0 ;
  assign n51111 = n51110 ^ n51109 ^ n23488 ;
  assign n51112 = ( n51106 & n51108 ) | ( n51106 & ~n51111 ) | ( n51108 & ~n51111 ) ;
  assign n51113 = n51112 ^ n34272 ^ 1'b0 ;
  assign n51114 = n51105 & ~n51113 ;
  assign n51115 = n18150 ^ n8434 ^ 1'b0 ;
  assign n51116 = ( n5124 & ~n14160 ) | ( n5124 & n25570 ) | ( ~n14160 & n25570 ) ;
  assign n51117 = n40274 ^ n18687 ^ n2851 ;
  assign n51118 = ( n4824 & n6766 ) | ( n4824 & ~n19014 ) | ( n6766 & ~n19014 ) ;
  assign n51119 = n51118 ^ n18774 ^ 1'b0 ;
  assign n51120 = n51119 ^ n36277 ^ n16567 ;
  assign n51121 = ~n50280 & n51120 ;
  assign n51122 = ( n15313 & n16669 ) | ( n15313 & n39639 ) | ( n16669 & n39639 ) ;
  assign n51123 = n22745 ^ n16083 ^ 1'b0 ;
  assign n51124 = ( ~n12307 & n13639 ) | ( ~n12307 & n20606 ) | ( n13639 & n20606 ) ;
  assign n51125 = ( n3484 & n35206 ) | ( n3484 & n40023 ) | ( n35206 & n40023 ) ;
  assign n51126 = n24818 ^ n16683 ^ 1'b0 ;
  assign n51127 = n51126 ^ n10497 ^ n4913 ;
  assign n51128 = n15035 ^ n1428 ^ 1'b0 ;
  assign n51129 = n11072 & n51128 ;
  assign n51130 = n23745 & n51129 ;
  assign n51131 = ~n51127 & n51130 ;
  assign n51132 = n23310 & ~n32231 ;
  assign n51133 = n17095 & ~n51132 ;
  assign n51134 = ~n34620 & n51133 ;
  assign n51140 = n4553 & n25256 ;
  assign n51141 = n51140 ^ n12956 ^ 1'b0 ;
  assign n51142 = n51141 ^ n3185 ^ 1'b0 ;
  assign n51135 = n1446 ^ x135 ^ 1'b0 ;
  assign n51136 = n51135 ^ n37852 ^ n23914 ;
  assign n51137 = ~n49077 & n51136 ;
  assign n51138 = n10546 & n51137 ;
  assign n51139 = n51138 ^ n39095 ^ 1'b0 ;
  assign n51143 = n51142 ^ n51139 ^ n7097 ;
  assign n51144 = n44999 | n51143 ;
  assign n51145 = n51144 ^ n4531 ^ 1'b0 ;
  assign n51146 = n36870 | n51145 ;
  assign n51147 = n2041 & ~n30767 ;
  assign n51148 = ~n51146 & n51147 ;
  assign n51149 = n34035 ^ n20300 ^ 1'b0 ;
  assign n51150 = n25479 ^ n14197 ^ n2318 ;
  assign n51151 = n3262 | n48948 ;
  assign n51152 = n51151 ^ n10775 ^ n1009 ;
  assign n51153 = n7878 | n28557 ;
  assign n51154 = n51152 | n51153 ;
  assign n51155 = n12887 & n36215 ;
  assign n51156 = n51154 & ~n51155 ;
  assign n51160 = n20871 ^ n16505 ^ 1'b0 ;
  assign n51157 = x37 & n3286 ;
  assign n51158 = ~n7999 & n51157 ;
  assign n51159 = n51158 ^ n10411 ^ 1'b0 ;
  assign n51161 = n51160 ^ n51159 ^ n36238 ;
  assign n51162 = ( n7051 & n37872 ) | ( n7051 & n38277 ) | ( n37872 & n38277 ) ;
  assign n51163 = n26705 ^ n12003 ^ n7070 ;
  assign n51164 = n51163 ^ n45885 ^ n17142 ;
  assign n51165 = n1688 | n51164 ;
  assign n51166 = n25519 ^ n24447 ^ n5704 ;
  assign n51167 = n44015 ^ n16756 ^ n15303 ;
  assign n51168 = ~n3877 & n5761 ;
  assign n51169 = n51168 ^ n24541 ^ 1'b0 ;
  assign n51170 = n36442 ^ n16140 ^ 1'b0 ;
  assign n51171 = ~n10303 & n14826 ;
  assign n51172 = n29325 ^ n16568 ^ 1'b0 ;
  assign n51173 = ( ~n14681 & n23686 ) | ( ~n14681 & n51172 ) | ( n23686 & n51172 ) ;
  assign n51174 = ( n906 & n1567 ) | ( n906 & ~n14611 ) | ( n1567 & ~n14611 ) ;
  assign n51175 = n51174 ^ n23685 ^ n10229 ;
  assign n51176 = ( x136 & n632 ) | ( x136 & n32982 ) | ( n632 & n32982 ) ;
  assign n51177 = ( n43392 & n44508 ) | ( n43392 & ~n51176 ) | ( n44508 & ~n51176 ) ;
  assign n51178 = ~x33 & n47325 ;
  assign n51180 = n34188 ^ n14285 ^ n6111 ;
  assign n51179 = ( n6920 & n13170 ) | ( n6920 & ~n50077 ) | ( n13170 & ~n50077 ) ;
  assign n51181 = n51180 ^ n51179 ^ n10092 ;
  assign n51182 = n18667 & n46161 ;
  assign n51183 = ~n4494 & n38394 ;
  assign n51184 = n51183 ^ n4688 ^ 1'b0 ;
  assign n51185 = ~n25816 & n27754 ;
  assign n51186 = n1657 & n51185 ;
  assign n51187 = n1828 & ~n8319 ;
  assign n51188 = n12993 & n51187 ;
  assign n51189 = n30083 ^ n11284 ^ 1'b0 ;
  assign n51190 = ( n1196 & n1308 ) | ( n1196 & n20993 ) | ( n1308 & n20993 ) ;
  assign n51191 = n32668 ^ n8441 ^ 1'b0 ;
  assign n51192 = n40454 ^ n8295 ^ 1'b0 ;
  assign n51193 = ( ~n11781 & n32843 ) | ( ~n11781 & n51192 ) | ( n32843 & n51192 ) ;
  assign n51194 = ( n13782 & n37658 ) | ( n13782 & n51193 ) | ( n37658 & n51193 ) ;
  assign n51195 = n35753 ^ n21204 ^ n11000 ;
  assign n51198 = n37641 ^ n27695 ^ n10243 ;
  assign n51196 = ( n1550 & n4255 ) | ( n1550 & ~n8307 ) | ( n4255 & ~n8307 ) ;
  assign n51197 = n51196 ^ n35562 ^ n13875 ;
  assign n51199 = n51198 ^ n51197 ^ n32889 ;
  assign n51200 = ( n6576 & ~n18539 ) | ( n6576 & n23753 ) | ( ~n18539 & n23753 ) ;
  assign n51201 = n51200 ^ n25643 ^ n20471 ;
  assign n51202 = n51201 ^ n16921 ^ 1'b0 ;
  assign n51203 = ~n5958 & n21889 ;
  assign n51204 = n2872 & n51203 ;
  assign n51206 = n18452 ^ n6663 ^ 1'b0 ;
  assign n51205 = n39256 & ~n45686 ;
  assign n51207 = n51206 ^ n51205 ^ 1'b0 ;
  assign n51208 = n18854 ^ n16833 ^ 1'b0 ;
  assign n51209 = n18601 & n30430 ;
  assign n51210 = n51209 ^ n42585 ^ n22015 ;
  assign n51211 = n33800 ^ n25931 ^ 1'b0 ;
  assign n51212 = n51211 ^ n10865 ^ n3038 ;
  assign n51213 = n40138 ^ n39497 ^ n15880 ;
  assign n51214 = n13692 | n51213 ;
  assign n51215 = n8224 ^ n3932 ^ 1'b0 ;
  assign n51216 = ( n27848 & n51214 ) | ( n27848 & ~n51215 ) | ( n51214 & ~n51215 ) ;
  assign n51217 = n46458 ^ n41673 ^ 1'b0 ;
  assign n51218 = n36277 & ~n51217 ;
  assign n51219 = ( n3144 & n32079 ) | ( n3144 & ~n51218 ) | ( n32079 & ~n51218 ) ;
  assign n51220 = n32157 ^ n18246 ^ n4538 ;
  assign n51221 = ( n8065 & n19114 ) | ( n8065 & n51220 ) | ( n19114 & n51220 ) ;
  assign n51222 = ( n3372 & n8026 ) | ( n3372 & ~n22865 ) | ( n8026 & ~n22865 ) ;
  assign n51223 = n51222 ^ n21775 ^ n7377 ;
  assign n51224 = n33887 ^ n22128 ^ n6765 ;
  assign n51225 = ( n51221 & n51223 ) | ( n51221 & n51224 ) | ( n51223 & n51224 ) ;
  assign n51226 = n49735 ^ n40432 ^ n26956 ;
  assign n51227 = n12519 ^ n1446 ^ x239 ;
  assign n51228 = n51227 ^ n25101 ^ 1'b0 ;
  assign n51229 = n44615 ^ n4494 ^ 1'b0 ;
  assign n51230 = n11450 & n51229 ;
  assign n51231 = n38730 ^ n22635 ^ n9299 ;
  assign n51232 = n51231 ^ n43619 ^ 1'b0 ;
  assign n51233 = ( n18976 & n24420 ) | ( n18976 & ~n45923 ) | ( n24420 & ~n45923 ) ;
  assign n51234 = ( ~n8373 & n26751 ) | ( ~n8373 & n51233 ) | ( n26751 & n51233 ) ;
  assign n51235 = n50123 ^ n35643 ^ n9502 ;
  assign n51236 = ( n4230 & ~n22545 ) | ( n4230 & n27358 ) | ( ~n22545 & n27358 ) ;
  assign n51237 = ( n4883 & n24571 ) | ( n4883 & n25801 ) | ( n24571 & n25801 ) ;
  assign n51238 = ( n6279 & ~n7571 ) | ( n6279 & n44080 ) | ( ~n7571 & n44080 ) ;
  assign n51239 = n19194 & ~n42784 ;
  assign n51240 = ( n1679 & ~n7675 ) | ( n1679 & n20587 ) | ( ~n7675 & n20587 ) ;
  assign n51241 = ~n28273 & n51240 ;
  assign n51242 = n48021 & n51241 ;
  assign n51243 = n3415 ^ n3176 ^ 1'b0 ;
  assign n51244 = n27296 & n51243 ;
  assign n51245 = n2512 | n34177 ;
  assign n51246 = n51245 ^ n33771 ^ 1'b0 ;
  assign n51248 = ( ~n19445 & n45817 ) | ( ~n19445 & n46071 ) | ( n45817 & n46071 ) ;
  assign n51247 = ~n13983 & n22810 ;
  assign n51249 = n51248 ^ n51247 ^ 1'b0 ;
  assign n51254 = n12284 ^ n1877 ^ 1'b0 ;
  assign n51250 = ( n3363 & n3686 ) | ( n3363 & n25879 ) | ( n3686 & n25879 ) ;
  assign n51251 = n51250 ^ n7977 ^ 1'b0 ;
  assign n51252 = n8189 & ~n51251 ;
  assign n51253 = ( n3871 & n50955 ) | ( n3871 & n51252 ) | ( n50955 & n51252 ) ;
  assign n51255 = n51254 ^ n51253 ^ n34495 ;
  assign n51256 = n16909 ^ n6213 ^ n2964 ;
  assign n51257 = n2841 & n51256 ;
  assign n51258 = ~n51255 & n51257 ;
  assign n51259 = ( n3227 & n28621 ) | ( n3227 & n51258 ) | ( n28621 & n51258 ) ;
  assign n51260 = n27314 ^ n23761 ^ n5594 ;
  assign n51261 = n51260 ^ n29159 ^ n8178 ;
  assign n51262 = n15431 & ~n18673 ;
  assign n51263 = n1873 | n10527 ;
  assign n51264 = n3241 | n11858 ;
  assign n51265 = n51264 ^ n16288 ^ 1'b0 ;
  assign n51266 = ( n6464 & n51263 ) | ( n6464 & n51265 ) | ( n51263 & n51265 ) ;
  assign n51267 = n11293 ^ n4141 ^ 1'b0 ;
  assign n51268 = ( ~n1397 & n46577 ) | ( ~n1397 & n51267 ) | ( n46577 & n51267 ) ;
  assign n51269 = n22964 ^ n7197 ^ n438 ;
  assign n51270 = n13642 ^ n10852 ^ 1'b0 ;
  assign n51271 = ( n14143 & ~n35954 ) | ( n14143 & n51270 ) | ( ~n35954 & n51270 ) ;
  assign n51272 = n9153 & ~n45577 ;
  assign n51273 = n51272 ^ n19091 ^ 1'b0 ;
  assign n51274 = n23730 ^ n10719 ^ 1'b0 ;
  assign n51275 = n28821 & n51274 ;
  assign n51276 = n17595 ^ n15354 ^ n9979 ;
  assign n51277 = ~n24918 & n51276 ;
  assign n51278 = n10059 & n27532 ;
  assign n51279 = n10132 ^ n3937 ^ x4 ;
  assign n51280 = ( ~n2715 & n3309 ) | ( ~n2715 & n51279 ) | ( n3309 & n51279 ) ;
  assign n51281 = n51280 ^ n10801 ^ n6584 ;
  assign n51282 = ( ~n12701 & n38950 ) | ( ~n12701 & n51281 ) | ( n38950 & n51281 ) ;
  assign n51283 = n51282 ^ n27196 ^ n5693 ;
  assign n51284 = n48221 ^ n30375 ^ n26492 ;
  assign n51285 = ( n19076 & n32956 ) | ( n19076 & ~n51284 ) | ( n32956 & ~n51284 ) ;
  assign n51286 = ( n21549 & n25816 ) | ( n21549 & n44353 ) | ( n25816 & n44353 ) ;
  assign n51287 = ~n18237 & n51286 ;
  assign n51288 = ( ~n658 & n26301 ) | ( ~n658 & n46345 ) | ( n26301 & n46345 ) ;
  assign n51289 = n418 & n51288 ;
  assign n51290 = ( n1222 & n40127 ) | ( n1222 & ~n51289 ) | ( n40127 & ~n51289 ) ;
  assign n51291 = n12677 ^ n3212 ^ n3120 ;
  assign n51292 = n51291 ^ n48416 ^ n7567 ;
  assign n51293 = n24106 ^ n6168 ^ 1'b0 ;
  assign n51294 = n4594 & ~n51293 ;
  assign n51296 = n21096 ^ n8910 ^ n1996 ;
  assign n51295 = n1029 & ~n34660 ;
  assign n51297 = n51296 ^ n51295 ^ 1'b0 ;
  assign n51298 = n23510 & ~n30687 ;
  assign n51299 = n30171 & n51298 ;
  assign n51300 = ( ~n7468 & n24042 ) | ( ~n7468 & n40589 ) | ( n24042 & n40589 ) ;
  assign n51301 = n41338 ^ n18595 ^ n8157 ;
  assign n51302 = ~n16293 & n51301 ;
  assign n51303 = n51302 ^ n41844 ^ n30624 ;
  assign n51304 = n51300 & n51303 ;
  assign n51305 = ( n11056 & ~n21725 ) | ( n11056 & n49610 ) | ( ~n21725 & n49610 ) ;
  assign n51306 = ( n10789 & ~n27697 ) | ( n10789 & n30220 ) | ( ~n27697 & n30220 ) ;
  assign n51307 = ( ~n17844 & n51305 ) | ( ~n17844 & n51306 ) | ( n51305 & n51306 ) ;
  assign n51308 = n16967 | n19726 ;
  assign n51309 = n14597 | n51308 ;
  assign n51310 = n51309 ^ n40960 ^ n23530 ;
  assign n51312 = ( n11342 & n26327 ) | ( n11342 & n30238 ) | ( n26327 & n30238 ) ;
  assign n51311 = ( n3973 & n4035 ) | ( n3973 & n39574 ) | ( n4035 & n39574 ) ;
  assign n51313 = n51312 ^ n51311 ^ n50932 ;
  assign n51314 = n9008 ^ n3509 ^ 1'b0 ;
  assign n51315 = ~n9067 & n51314 ;
  assign n51316 = n28836 | n34199 ;
  assign n51317 = n51316 ^ n48311 ^ n10217 ;
  assign n51318 = n5186 & ~n51317 ;
  assign n51319 = ~n16146 & n51318 ;
  assign n51320 = n43898 ^ n12968 ^ n10092 ;
  assign n51321 = ( ~n7898 & n14257 ) | ( ~n7898 & n26349 ) | ( n14257 & n26349 ) ;
  assign n51322 = n6643 ^ n6448 ^ 1'b0 ;
  assign n51323 = ( n8510 & n13847 ) | ( n8510 & ~n33910 ) | ( n13847 & ~n33910 ) ;
  assign n51324 = ( n23036 & n51322 ) | ( n23036 & ~n51323 ) | ( n51322 & ~n51323 ) ;
  assign n51326 = n9312 | n21088 ;
  assign n51325 = ~n25741 & n50626 ;
  assign n51327 = n51326 ^ n51325 ^ n27734 ;
  assign n51328 = ( n6590 & ~n8729 ) | ( n6590 & n24160 ) | ( ~n8729 & n24160 ) ;
  assign n51329 = n51328 ^ n43442 ^ n23702 ;
  assign n51330 = n51329 ^ n47842 ^ n2686 ;
  assign n51331 = n4411 | n5293 ;
  assign n51332 = n51331 ^ n2070 ^ 1'b0 ;
  assign n51333 = n51332 ^ n46559 ^ n3128 ;
  assign n51334 = n16522 ^ n11813 ^ x238 ;
  assign n51335 = ( ~n20228 & n51333 ) | ( ~n20228 & n51334 ) | ( n51333 & n51334 ) ;
  assign n51336 = n26849 ^ n22640 ^ n13486 ;
  assign n51337 = ( ~n1754 & n2243 ) | ( ~n1754 & n51336 ) | ( n2243 & n51336 ) ;
  assign n51338 = n2722 & n33973 ;
  assign n51339 = ~n39965 & n49131 ;
  assign n51340 = n51338 & n51339 ;
  assign n51343 = ( n3761 & n4132 ) | ( n3761 & ~n14649 ) | ( n4132 & ~n14649 ) ;
  assign n51344 = n51343 ^ n48525 ^ n3294 ;
  assign n51341 = n26587 ^ n807 ^ 1'b0 ;
  assign n51342 = n51341 ^ n18684 ^ n17557 ;
  assign n51345 = n51344 ^ n51342 ^ n6488 ;
  assign n51346 = ~n1204 & n51345 ;
  assign n51347 = n51346 ^ n7420 ^ 1'b0 ;
  assign n51348 = n40594 & ~n46461 ;
  assign n51349 = n40131 ^ n10298 ^ n4921 ;
  assign n51350 = n51349 ^ n8379 ^ n5564 ;
  assign n51351 = n51350 ^ n49909 ^ n1516 ;
  assign n51352 = n25871 ^ n13596 ^ n1796 ;
  assign n51353 = n37543 ^ n28647 ^ n3599 ;
  assign n51354 = n45727 ^ n21554 ^ 1'b0 ;
  assign n51355 = n35762 | n51354 ;
  assign n51356 = n51355 ^ n21281 ^ n5387 ;
  assign n51357 = n10606 | n51356 ;
  assign n51360 = n17312 ^ n9582 ^ n3138 ;
  assign n51358 = n2152 & ~n26608 ;
  assign n51359 = n14720 & n51358 ;
  assign n51361 = n51360 ^ n51359 ^ n13050 ;
  assign n51362 = n43568 ^ n10739 ^ 1'b0 ;
  assign n51363 = ~n47576 & n51362 ;
  assign n51364 = n16495 ^ n9844 ^ 1'b0 ;
  assign n51365 = ~n11301 & n16445 ;
  assign n51366 = n51365 ^ n12973 ^ 1'b0 ;
  assign n51367 = ( n15914 & n18506 ) | ( n15914 & ~n51366 ) | ( n18506 & ~n51366 ) ;
  assign n51368 = n30081 ^ n6264 ^ 1'b0 ;
  assign n51369 = n9669 & n51368 ;
  assign n51370 = n27520 & n51369 ;
  assign n51371 = n13948 & ~n35556 ;
  assign n51372 = n51371 ^ n29659 ^ 1'b0 ;
  assign n51373 = n7532 ^ n5767 ^ 1'b0 ;
  assign n51374 = ~n606 & n51373 ;
  assign n51375 = n12066 | n51374 ;
  assign n51376 = ( ~n16216 & n26682 ) | ( ~n16216 & n51375 ) | ( n26682 & n51375 ) ;
  assign n51377 = ( ~n9694 & n10267 ) | ( ~n9694 & n17739 ) | ( n10267 & n17739 ) ;
  assign n51379 = ( n21829 & n34836 ) | ( n21829 & ~n35361 ) | ( n34836 & ~n35361 ) ;
  assign n51378 = n5994 & n18843 ;
  assign n51380 = n51379 ^ n51378 ^ 1'b0 ;
  assign n51381 = ( ~n49912 & n51377 ) | ( ~n49912 & n51380 ) | ( n51377 & n51380 ) ;
  assign n51382 = ( n12828 & n14284 ) | ( n12828 & n22236 ) | ( n14284 & n22236 ) ;
  assign n51383 = n45033 ^ n10243 ^ 1'b0 ;
  assign n51384 = n49299 ^ n30675 ^ 1'b0 ;
  assign n51385 = n17913 | n40600 ;
  assign n51386 = n24267 ^ n690 ^ 1'b0 ;
  assign n51387 = n8047 & ~n19411 ;
  assign n51388 = n51387 ^ n47585 ^ 1'b0 ;
  assign n51389 = n51388 ^ n24359 ^ n14165 ;
  assign n51390 = n8107 ^ n6376 ^ 1'b0 ;
  assign n51391 = n51390 ^ n26501 ^ n13640 ;
  assign n51392 = ( n1656 & n2250 ) | ( n1656 & ~n27540 ) | ( n2250 & ~n27540 ) ;
  assign n51393 = n13798 & n48276 ;
  assign n51394 = n51393 ^ n44565 ^ n8549 ;
  assign n51395 = ( ~n6223 & n29911 ) | ( ~n6223 & n40819 ) | ( n29911 & n40819 ) ;
  assign n51396 = n40513 ^ n36320 ^ 1'b0 ;
  assign n51397 = ( n26018 & ~n47193 ) | ( n26018 & n51396 ) | ( ~n47193 & n51396 ) ;
  assign n51398 = n37293 ^ n25392 ^ n10154 ;
  assign n51399 = n24460 ^ n12315 ^ n9576 ;
  assign n51400 = n51398 & n51399 ;
  assign n51401 = n32986 ^ n22568 ^ n13548 ;
  assign n51402 = n51401 ^ n36088 ^ n8369 ;
  assign n51403 = n5748 | n19656 ;
  assign n51404 = n51403 ^ n14232 ^ 1'b0 ;
  assign n51405 = ( ~n6699 & n51402 ) | ( ~n6699 & n51404 ) | ( n51402 & n51404 ) ;
  assign n51406 = n35723 | n51405 ;
  assign n51407 = n51406 ^ n32820 ^ 1'b0 ;
  assign n51408 = n46948 ^ n10156 ^ 1'b0 ;
  assign n51409 = n23881 | n51408 ;
  assign n51410 = n51409 ^ n24585 ^ n13225 ;
  assign n51411 = n23732 | n51410 ;
  assign n51413 = n31000 ^ n14887 ^ 1'b0 ;
  assign n51412 = n8675 & n40438 ;
  assign n51414 = n51413 ^ n51412 ^ 1'b0 ;
  assign n51415 = ( n30039 & n30378 ) | ( n30039 & n32490 ) | ( n30378 & n32490 ) ;
  assign n51416 = n12640 | n51415 ;
  assign n51417 = n1039 & ~n51416 ;
  assign n51418 = n51417 ^ n3633 ^ n1970 ;
  assign n51419 = n16411 ^ n5812 ^ n4342 ;
  assign n51420 = n10367 | n51419 ;
  assign n51421 = n20864 ^ n16921 ^ n7302 ;
  assign n51422 = n51421 ^ n40866 ^ n4792 ;
  assign n51423 = n51422 ^ n12931 ^ n9085 ;
  assign n51424 = ( x241 & ~n4754 ) | ( x241 & n17991 ) | ( ~n4754 & n17991 ) ;
  assign n51425 = ( n13548 & n36234 ) | ( n13548 & n51424 ) | ( n36234 & n51424 ) ;
  assign n51426 = n42515 & ~n51425 ;
  assign n51427 = n11446 ^ n8842 ^ n2849 ;
  assign n51428 = ~n17785 & n51427 ;
  assign n51429 = n14843 | n31030 ;
  assign n51430 = ( n6778 & ~n29225 ) | ( n6778 & n51429 ) | ( ~n29225 & n51429 ) ;
  assign n51431 = ~n5062 & n42086 ;
  assign n51432 = ~n51430 & n51431 ;
  assign n51433 = n44868 ^ n13972 ^ 1'b0 ;
  assign n51434 = n13910 ^ n10548 ^ n2146 ;
  assign n51435 = n51434 ^ n22389 ^ 1'b0 ;
  assign n51436 = n4225 & n51435 ;
  assign n51437 = n2892 & n14094 ;
  assign n51438 = n22540 & ~n51437 ;
  assign n51440 = ( ~n5671 & n19325 ) | ( ~n5671 & n40594 ) | ( n19325 & n40594 ) ;
  assign n51439 = n25486 ^ n17141 ^ n6554 ;
  assign n51441 = n51440 ^ n51439 ^ n462 ;
  assign n51442 = n16186 ^ n8590 ^ n834 ;
  assign n51443 = n5552 & n19550 ;
  assign n51445 = ( n18648 & n20528 ) | ( n18648 & ~n35321 ) | ( n20528 & ~n35321 ) ;
  assign n51444 = n30607 ^ n13627 ^ n887 ;
  assign n51446 = n51445 ^ n51444 ^ n21070 ;
  assign n51450 = n27425 ^ n23266 ^ n2247 ;
  assign n51448 = n25364 ^ n5846 ^ n3498 ;
  assign n51447 = ~n10049 & n51139 ;
  assign n51449 = n51448 ^ n51447 ^ 1'b0 ;
  assign n51451 = n51450 ^ n51449 ^ n10894 ;
  assign n51452 = ~n24613 & n40548 ;
  assign n51453 = n7715 & n51452 ;
  assign n51454 = n51453 ^ n48717 ^ n7449 ;
  assign n51455 = n32046 ^ n19784 ^ n7521 ;
  assign n51456 = n8347 | n25610 ;
  assign n51457 = n51455 & ~n51456 ;
  assign n51458 = n21431 & n39411 ;
  assign n51459 = n51458 ^ n31194 ^ 1'b0 ;
  assign n51460 = n41586 ^ n37052 ^ n28051 ;
  assign n51461 = n51460 ^ n42255 ^ n3977 ;
  assign n51462 = ~n25938 & n51461 ;
  assign n51463 = n26236 ^ n10736 ^ 1'b0 ;
  assign n51464 = n24818 ^ n16003 ^ n3794 ;
  assign n51465 = ( n433 & n12413 ) | ( n433 & ~n23532 ) | ( n12413 & ~n23532 ) ;
  assign n51466 = ( n51309 & ~n51464 ) | ( n51309 & n51465 ) | ( ~n51464 & n51465 ) ;
  assign n51467 = ( n8914 & ~n20013 ) | ( n8914 & n46089 ) | ( ~n20013 & n46089 ) ;
  assign n51468 = n37598 ^ n25459 ^ n7679 ;
  assign n51469 = ~n7944 & n13506 ;
  assign n51470 = n51469 ^ n408 ^ 1'b0 ;
  assign n51471 = n51470 ^ n25822 ^ n11819 ;
  assign n51472 = n51069 ^ n13775 ^ n8059 ;
  assign n51473 = ( n1899 & ~n51471 ) | ( n1899 & n51472 ) | ( ~n51471 & n51472 ) ;
  assign n51474 = n33368 ^ n33328 ^ n32444 ;
  assign n51475 = n4454 & ~n10490 ;
  assign n51476 = n19967 & n51475 ;
  assign n51477 = n45822 ^ n34618 ^ n3644 ;
  assign n51478 = n51477 ^ n4142 ^ 1'b0 ;
  assign n51479 = n48589 & n51478 ;
  assign n51480 = n39768 ^ n26622 ^ n8085 ;
  assign n51481 = ( n7696 & n9283 ) | ( n7696 & ~n51480 ) | ( n9283 & ~n51480 ) ;
  assign n51482 = n51481 ^ n7177 ^ 1'b0 ;
  assign n51483 = ~n17029 & n51482 ;
  assign n51484 = n51483 ^ n11590 ^ 1'b0 ;
  assign n51485 = n26356 & n51484 ;
  assign n51486 = n15270 | n20354 ;
  assign n51487 = n51486 ^ n3975 ^ 1'b0 ;
  assign n51488 = ~n25596 & n51487 ;
  assign n51489 = n48523 & n51488 ;
  assign n51490 = ~n1064 & n51489 ;
  assign n51491 = n25039 ^ n12167 ^ n9473 ;
  assign n51492 = n24315 ^ n11447 ^ 1'b0 ;
  assign n51493 = n23535 & n51492 ;
  assign n51494 = ( n9782 & n48974 ) | ( n9782 & ~n51493 ) | ( n48974 & ~n51493 ) ;
  assign n51495 = ( n5280 & ~n27595 ) | ( n5280 & n42270 ) | ( ~n27595 & n42270 ) ;
  assign n51496 = ( n8896 & n9795 ) | ( n8896 & ~n19396 ) | ( n9795 & ~n19396 ) ;
  assign n51497 = n51496 ^ n50659 ^ n13941 ;
  assign n51500 = ( n3234 & ~n14187 ) | ( n3234 & n20985 ) | ( ~n14187 & n20985 ) ;
  assign n51498 = ( n6342 & ~n9302 ) | ( n6342 & n44623 ) | ( ~n9302 & n44623 ) ;
  assign n51499 = ( ~n40294 & n44815 ) | ( ~n40294 & n51498 ) | ( n44815 & n51498 ) ;
  assign n51501 = n51500 ^ n51499 ^ 1'b0 ;
  assign n51502 = ( n14836 & ~n27010 ) | ( n14836 & n35105 ) | ( ~n27010 & n35105 ) ;
  assign n51503 = n11710 & n28093 ;
  assign n51504 = ~n9245 & n51503 ;
  assign n51505 = n7547 & n38525 ;
  assign n51506 = n51505 ^ n39700 ^ 1'b0 ;
  assign n51507 = ~n32295 & n44676 ;
  assign n51508 = n51507 ^ n44640 ^ 1'b0 ;
  assign n51509 = ~n15667 & n19398 ;
  assign n51510 = n23164 | n47405 ;
  assign n51511 = n51510 ^ n14636 ^ 1'b0 ;
  assign n51512 = n51509 & ~n51511 ;
  assign n51513 = n23074 ^ n1931 ^ 1'b0 ;
  assign n51514 = n47003 ^ n32436 ^ n11078 ;
  assign n51515 = ( n42904 & n49950 ) | ( n42904 & n51514 ) | ( n49950 & n51514 ) ;
  assign n51516 = n17411 & ~n23248 ;
  assign n51517 = ( n3280 & ~n6930 ) | ( n3280 & n15947 ) | ( ~n6930 & n15947 ) ;
  assign n51518 = ( n11481 & n51516 ) | ( n11481 & n51517 ) | ( n51516 & n51517 ) ;
  assign n51519 = n32411 ^ n23940 ^ n6222 ;
  assign n51520 = n40165 ^ n28478 ^ n16032 ;
  assign n51521 = ( n2146 & ~n4226 ) | ( n2146 & n42382 ) | ( ~n4226 & n42382 ) ;
  assign n51522 = n16111 & n46844 ;
  assign n51523 = n51522 ^ n7910 ^ 1'b0 ;
  assign n51524 = n11901 | n44084 ;
  assign n51525 = n46917 | n51524 ;
  assign n51526 = n23576 ^ n11367 ^ n5347 ;
  assign n51527 = n51526 ^ n7859 ^ 1'b0 ;
  assign n51528 = n51527 ^ n22890 ^ 1'b0 ;
  assign n51529 = ( n12374 & ~n22992 ) | ( n12374 & n50425 ) | ( ~n22992 & n50425 ) ;
  assign n51530 = ( n4957 & n46749 ) | ( n4957 & n51529 ) | ( n46749 & n51529 ) ;
  assign n51531 = n48470 ^ n14180 ^ n13358 ;
  assign n51532 = n51531 ^ n39637 ^ n2011 ;
  assign n51533 = n51532 ^ n50804 ^ n9252 ;
  assign n51534 = n1482 | n16880 ;
  assign n51535 = n51534 ^ n17125 ^ 1'b0 ;
  assign n51536 = n51535 ^ n3178 ^ 1'b0 ;
  assign n51537 = ( n14717 & n25835 ) | ( n14717 & n26146 ) | ( n25835 & n26146 ) ;
  assign n51538 = ( ~n20779 & n34385 ) | ( ~n20779 & n42235 ) | ( n34385 & n42235 ) ;
  assign n51539 = ( ~n1676 & n3182 ) | ( ~n1676 & n27089 ) | ( n3182 & n27089 ) ;
  assign n51540 = n51539 ^ n38926 ^ n28846 ;
  assign n51541 = ~n2318 & n21520 ;
  assign n51542 = n34090 ^ n7095 ^ 1'b0 ;
  assign n51543 = ~n12954 & n51542 ;
  assign n51544 = ~n19655 & n51543 ;
  assign n51545 = n3549 ^ n3242 ^ 1'b0 ;
  assign n51546 = n27697 & n51545 ;
  assign n51547 = n51546 ^ n39637 ^ 1'b0 ;
  assign n51548 = n27610 | n51547 ;
  assign n51549 = n24443 ^ n5567 ^ 1'b0 ;
  assign n51550 = n34534 & n51549 ;
  assign n51551 = n24035 ^ n12599 ^ 1'b0 ;
  assign n51552 = n5203 & ~n51551 ;
  assign n51553 = n51552 ^ n16140 ^ n14628 ;
  assign n51554 = ( n39458 & n46483 ) | ( n39458 & n51553 ) | ( n46483 & n51553 ) ;
  assign n51555 = n51554 ^ n50815 ^ n31984 ;
  assign n51556 = ~n10503 & n16139 ;
  assign n51557 = n12413 & n51556 ;
  assign n51558 = ( n11614 & ~n22389 ) | ( n11614 & n51557 ) | ( ~n22389 & n51557 ) ;
  assign n51559 = ( ~n1028 & n11933 ) | ( ~n1028 & n51558 ) | ( n11933 & n51558 ) ;
  assign n51560 = n9610 | n33738 ;
  assign n51561 = ( n7785 & n33283 ) | ( n7785 & n44783 ) | ( n33283 & n44783 ) ;
  assign n51562 = n51561 ^ n2318 ^ 1'b0 ;
  assign n51563 = n41145 ^ n13909 ^ n4150 ;
  assign n51564 = n32423 ^ n32002 ^ n18033 ;
  assign n51565 = ~n4358 & n43665 ;
  assign n51566 = n51565 ^ n23452 ^ 1'b0 ;
  assign n51567 = n1795 & ~n28796 ;
  assign n51568 = n7315 & n51567 ;
  assign n51569 = n17159 & ~n51568 ;
  assign n51570 = ~n12681 & n51569 ;
  assign n51571 = n15290 ^ n466 ^ 1'b0 ;
  assign n51572 = n13959 ^ n8873 ^ 1'b0 ;
  assign n51573 = n37669 ^ n29904 ^ n4819 ;
  assign n51574 = ~n51572 & n51573 ;
  assign n51575 = n51574 ^ n26823 ^ 1'b0 ;
  assign n51576 = ~n16989 & n51575 ;
  assign n51577 = ( ~n4283 & n12690 ) | ( ~n4283 & n26763 ) | ( n12690 & n26763 ) ;
  assign n51578 = ( ~n33981 & n39373 ) | ( ~n33981 & n47889 ) | ( n39373 & n47889 ) ;
  assign n51579 = n39754 ^ n31347 ^ n27906 ;
  assign n51580 = ~n1532 & n1855 ;
  assign n51581 = ( n800 & n8886 ) | ( n800 & ~n33943 ) | ( n8886 & ~n33943 ) ;
  assign n51582 = n4512 & n19945 ;
  assign n51583 = n35492 ^ n25719 ^ n24306 ;
  assign n51584 = ( n40082 & n51582 ) | ( n40082 & ~n51583 ) | ( n51582 & ~n51583 ) ;
  assign n51585 = n17302 ^ n10937 ^ n6658 ;
  assign n51586 = ( n43290 & n45598 ) | ( n43290 & ~n51585 ) | ( n45598 & ~n51585 ) ;
  assign n51588 = n6868 & n12102 ;
  assign n51589 = n5216 & n51588 ;
  assign n51590 = n51589 ^ n44023 ^ n34493 ;
  assign n51587 = ~n1492 & n19120 ;
  assign n51591 = n51590 ^ n51587 ^ 1'b0 ;
  assign n51592 = n51591 ^ n45241 ^ n21473 ;
  assign n51593 = n1182 & ~n51592 ;
  assign n51594 = ~n14433 & n22425 ;
  assign n51595 = ~n32110 & n51594 ;
  assign n51596 = n26731 ^ n7735 ^ n5501 ;
  assign n51597 = ~n6210 & n51596 ;
  assign n51598 = n49814 & n51597 ;
  assign n51599 = ( n8824 & n21745 ) | ( n8824 & ~n49293 ) | ( n21745 & ~n49293 ) ;
  assign n51600 = n30985 ^ n17909 ^ n10552 ;
  assign n51601 = n45956 ^ n31993 ^ 1'b0 ;
  assign n51602 = n49727 & ~n51601 ;
  assign n51603 = ~n5969 & n24979 ;
  assign n51604 = n51603 ^ n46957 ^ 1'b0 ;
  assign n51605 = ( n51174 & n51602 ) | ( n51174 & ~n51604 ) | ( n51602 & ~n51604 ) ;
  assign n51606 = ( ~n28101 & n30846 ) | ( ~n28101 & n42481 ) | ( n30846 & n42481 ) ;
  assign n51611 = n30223 ^ n8649 ^ n3585 ;
  assign n51612 = ( n14510 & n19778 ) | ( n14510 & ~n51611 ) | ( n19778 & ~n51611 ) ;
  assign n51608 = n11198 | n24624 ;
  assign n51609 = n8486 | n37734 ;
  assign n51610 = n51608 | n51609 ;
  assign n51607 = n25820 ^ n4414 ^ 1'b0 ;
  assign n51613 = n51612 ^ n51610 ^ n51607 ;
  assign n51614 = n5021 ^ n4241 ^ n3184 ;
  assign n51615 = n21104 ^ n9943 ^ n747 ;
  assign n51616 = n25697 & ~n51615 ;
  assign n51617 = ( n8184 & n51614 ) | ( n8184 & n51616 ) | ( n51614 & n51616 ) ;
  assign n51618 = ( ~n7213 & n14447 ) | ( ~n7213 & n51617 ) | ( n14447 & n51617 ) ;
  assign n51619 = n51618 ^ n36351 ^ n3747 ;
  assign n51620 = ~n29913 & n51619 ;
  assign n51621 = n24593 & n51620 ;
  assign n51622 = n31060 | n45231 ;
  assign n51623 = n30176 | n32019 ;
  assign n51624 = n47419 & ~n51623 ;
  assign n51625 = ( n18850 & n26838 ) | ( n18850 & ~n51624 ) | ( n26838 & ~n51624 ) ;
  assign n51626 = n45263 ^ n27218 ^ 1'b0 ;
  assign n51627 = n36822 ^ n34049 ^ 1'b0 ;
  assign n51628 = n17936 & ~n51627 ;
  assign n51629 = ( n6722 & n11328 ) | ( n6722 & ~n25064 ) | ( n11328 & ~n25064 ) ;
  assign n51630 = n51628 & n51629 ;
  assign n51631 = n51630 ^ n34877 ^ 1'b0 ;
  assign n51632 = ( n9490 & ~n15483 ) | ( n9490 & n51631 ) | ( ~n15483 & n51631 ) ;
  assign n51633 = n10321 | n44911 ;
  assign n51634 = n39411 ^ n27385 ^ 1'b0 ;
  assign n51635 = n9844 & ~n51634 ;
  assign n51636 = n39797 ^ n22878 ^ 1'b0 ;
  assign n51637 = n51635 & ~n51636 ;
  assign n51638 = ( ~n14356 & n49086 ) | ( ~n14356 & n51637 ) | ( n49086 & n51637 ) ;
  assign n51639 = n37212 ^ n31298 ^ n29021 ;
  assign n51640 = n26431 ^ n22833 ^ n1096 ;
  assign n51641 = n15502 ^ n12665 ^ 1'b0 ;
  assign n51642 = n20412 | n51641 ;
  assign n51643 = n51642 ^ n14146 ^ 1'b0 ;
  assign n51644 = ~n4670 & n21113 ;
  assign n51645 = n36145 ^ n23943 ^ 1'b0 ;
  assign n51646 = n43393 ^ n24268 ^ 1'b0 ;
  assign n51647 = ( n25118 & ~n38000 ) | ( n25118 & n51646 ) | ( ~n38000 & n51646 ) ;
  assign n51648 = n11400 & ~n43311 ;
  assign n51649 = ( n1520 & ~n4729 ) | ( n1520 & n9180 ) | ( ~n4729 & n9180 ) ;
  assign n51650 = n51649 ^ n13789 ^ 1'b0 ;
  assign n51651 = n32788 & ~n39050 ;
  assign n51652 = ( n36105 & n43053 ) | ( n36105 & n51651 ) | ( n43053 & n51651 ) ;
  assign n51653 = n23974 ^ n16894 ^ n12884 ;
  assign n51654 = n5625 & ~n22975 ;
  assign n51655 = n51654 ^ n36001 ^ n31579 ;
  assign n51656 = ( n46959 & n51653 ) | ( n46959 & n51655 ) | ( n51653 & n51655 ) ;
  assign n51657 = ( n5761 & n27511 ) | ( n5761 & n36380 ) | ( n27511 & n36380 ) ;
  assign n51658 = n43567 ^ n39728 ^ 1'b0 ;
  assign n51659 = n51657 | n51658 ;
  assign n51665 = n38201 ^ n10005 ^ 1'b0 ;
  assign n51660 = ~n5219 & n12950 ;
  assign n51661 = n51660 ^ n1246 ^ 1'b0 ;
  assign n51662 = ~n16701 & n41118 ;
  assign n51663 = ~n51661 & n51662 ;
  assign n51664 = n6318 & ~n51663 ;
  assign n51666 = n51665 ^ n51664 ^ 1'b0 ;
  assign n51667 = n5667 | n16969 ;
  assign n51668 = n48451 | n51667 ;
  assign n51670 = n3777 | n18919 ;
  assign n51669 = ~n2840 & n19984 ;
  assign n51671 = n51670 ^ n51669 ^ 1'b0 ;
  assign n51672 = n51671 ^ n22989 ^ 1'b0 ;
  assign n51673 = n2937 | n38558 ;
  assign n51674 = n51673 ^ n46781 ^ n35511 ;
  assign n51675 = ( n2767 & n24960 ) | ( n2767 & ~n42380 ) | ( n24960 & ~n42380 ) ;
  assign n51676 = n51027 ^ n37166 ^ n31864 ;
  assign n51677 = ( n466 & n22654 ) | ( n466 & ~n36608 ) | ( n22654 & ~n36608 ) ;
  assign n51678 = n46379 ^ n15028 ^ n11230 ;
  assign n51679 = n51678 ^ n13016 ^ n11619 ;
  assign n51680 = n8854 & n51679 ;
  assign n51681 = n50058 ^ n12910 ^ n12230 ;
  assign n51682 = n8675 & n51681 ;
  assign n51683 = n51682 ^ n47641 ^ n10443 ;
  assign n51684 = n25183 | n31647 ;
  assign n51685 = n28242 & ~n51684 ;
  assign n51686 = n51685 ^ n6624 ^ 1'b0 ;
  assign n51687 = ~n3826 & n51686 ;
  assign n51688 = n33713 & ~n51687 ;
  assign n51689 = n30893 ^ n24183 ^ 1'b0 ;
  assign n51690 = n42865 ^ n33467 ^ n19231 ;
  assign n51691 = ~n46555 & n51690 ;
  assign n51692 = n10448 & n43320 ;
  assign n51693 = n34203 & n51692 ;
  assign n51694 = ( n31073 & n37747 ) | ( n31073 & n51693 ) | ( n37747 & n51693 ) ;
  assign n51695 = n30172 ^ n28362 ^ 1'b0 ;
  assign n51696 = n17812 & ~n51695 ;
  assign n51697 = ( n2875 & ~n3181 ) | ( n2875 & n24463 ) | ( ~n3181 & n24463 ) ;
  assign n51698 = ( n4132 & n20738 ) | ( n4132 & ~n51697 ) | ( n20738 & ~n51697 ) ;
  assign n51699 = ~n51696 & n51698 ;
  assign n51700 = n51135 ^ n26080 ^ 1'b0 ;
  assign n51701 = n27788 & ~n51700 ;
  assign n51702 = ~n24124 & n51701 ;
  assign n51703 = n51702 ^ n15229 ^ 1'b0 ;
  assign n51704 = ( n2341 & ~n28791 ) | ( n2341 & n41867 ) | ( ~n28791 & n41867 ) ;
  assign n51705 = n50098 ^ n47977 ^ n46788 ;
  assign n51706 = n51705 ^ n10060 ^ 1'b0 ;
  assign n51707 = n51706 ^ n5847 ^ 1'b0 ;
  assign n51708 = ~n863 & n4804 ;
  assign n51709 = n40400 | n51708 ;
  assign n51710 = n27789 ^ n15972 ^ n5211 ;
  assign n51711 = n51710 ^ n45484 ^ n37785 ;
  assign n51712 = n24945 & ~n50871 ;
  assign n51713 = ( n15280 & n26566 ) | ( n15280 & ~n51712 ) | ( n26566 & ~n51712 ) ;
  assign n51714 = ( ~n7149 & n25014 ) | ( ~n7149 & n51713 ) | ( n25014 & n51713 ) ;
  assign n51715 = ~n29236 & n47419 ;
  assign n51716 = ( ~n18405 & n25891 ) | ( ~n18405 & n51715 ) | ( n25891 & n51715 ) ;
  assign n51717 = n5203 & ~n8595 ;
  assign n51718 = ( n17437 & ~n32661 ) | ( n17437 & n51717 ) | ( ~n32661 & n51717 ) ;
  assign n51719 = ( n28772 & n32900 ) | ( n28772 & n51215 ) | ( n32900 & n51215 ) ;
  assign n51720 = ~n4959 & n51719 ;
  assign n51721 = n48905 & n51720 ;
  assign n51722 = ~n4584 & n28677 ;
  assign n51723 = ~n16043 & n51722 ;
  assign n51724 = ( ~n3156 & n6102 ) | ( ~n3156 & n24857 ) | ( n6102 & n24857 ) ;
  assign n51725 = n22279 | n51724 ;
  assign n51726 = n25812 ^ n21590 ^ n6243 ;
  assign n51727 = n46393 ^ n38417 ^ n12132 ;
  assign n51728 = n24807 & n28051 ;
  assign n51729 = n40440 ^ n40381 ^ n12388 ;
  assign n51730 = ( n13954 & n51728 ) | ( n13954 & n51729 ) | ( n51728 & n51729 ) ;
  assign n51731 = n46542 ^ n17649 ^ n2357 ;
  assign n51732 = n51731 ^ n19970 ^ n653 ;
  assign n51733 = n31656 ^ n13699 ^ n12575 ;
  assign n51734 = ( n12863 & ~n15510 ) | ( n12863 & n25099 ) | ( ~n15510 & n25099 ) ;
  assign n51735 = n7763 | n14945 ;
  assign n51736 = n14654 ^ n9306 ^ 1'b0 ;
  assign n51737 = n51735 & ~n51736 ;
  assign n51738 = ( ~n29651 & n36069 ) | ( ~n29651 & n51737 ) | ( n36069 & n51737 ) ;
  assign n51739 = n13986 & ~n51738 ;
  assign n51740 = n51739 ^ n45959 ^ 1'b0 ;
  assign n51741 = n14838 & ~n20344 ;
  assign n51742 = ~n16336 & n27991 ;
  assign n51743 = n51741 & n51742 ;
  assign n51744 = ( n4911 & n48572 ) | ( n4911 & n51574 ) | ( n48572 & n51574 ) ;
  assign n51745 = ( n4010 & n29890 ) | ( n4010 & ~n51744 ) | ( n29890 & ~n51744 ) ;
  assign n51746 = n4768 | n51745 ;
  assign n51747 = n25466 & ~n42157 ;
  assign n51748 = n47439 ^ n20581 ^ n15178 ;
  assign n51749 = ( ~n19148 & n22812 ) | ( ~n19148 & n35153 ) | ( n22812 & n35153 ) ;
  assign n51750 = ( n7225 & n10834 ) | ( n7225 & ~n49531 ) | ( n10834 & ~n49531 ) ;
  assign n51751 = n9755 & ~n30019 ;
  assign n51752 = n51751 ^ n35353 ^ 1'b0 ;
  assign n51753 = ( n36501 & ~n51252 ) | ( n36501 & n51752 ) | ( ~n51252 & n51752 ) ;
  assign n51754 = n18024 ^ n9189 ^ n1819 ;
  assign n51755 = n51754 ^ n21812 ^ n12575 ;
  assign n51756 = ( n24208 & n36238 ) | ( n24208 & n51755 ) | ( n36238 & n51755 ) ;
  assign n51757 = n51756 ^ n20014 ^ 1'b0 ;
  assign n51758 = ( ~n32685 & n39093 ) | ( ~n32685 & n51000 ) | ( n39093 & n51000 ) ;
  assign n51759 = n2880 | n34487 ;
  assign n51760 = n24202 ^ n11079 ^ 1'b0 ;
  assign n51761 = n37432 & ~n51760 ;
  assign n51762 = n51761 ^ n44310 ^ n9067 ;
  assign n51763 = ( n25575 & n51759 ) | ( n25575 & ~n51762 ) | ( n51759 & ~n51762 ) ;
  assign n51764 = n51763 ^ n18871 ^ 1'b0 ;
  assign n51765 = n19259 | n51764 ;
  assign n51766 = ( ~n14700 & n19558 ) | ( ~n14700 & n30171 ) | ( n19558 & n30171 ) ;
  assign n51767 = n48948 ^ n41771 ^ n12938 ;
  assign n51768 = n6398 ^ n6223 ^ 1'b0 ;
  assign n51769 = ~n44236 & n48822 ;
  assign n51770 = ( n15457 & n19831 ) | ( n15457 & n51769 ) | ( n19831 & n51769 ) ;
  assign n51771 = ( n3250 & n10894 ) | ( n3250 & ~n49334 ) | ( n10894 & ~n49334 ) ;
  assign n51772 = n46164 ^ n28416 ^ n3987 ;
  assign n51773 = n34829 & ~n42959 ;
  assign n51774 = n43301 ^ n36736 ^ 1'b0 ;
  assign n51775 = n1610 | n51774 ;
  assign n51776 = n30978 & ~n51775 ;
  assign n51777 = n14698 | n50939 ;
  assign n51779 = ( ~n13062 & n45525 ) | ( ~n13062 & n49435 ) | ( n45525 & n49435 ) ;
  assign n51778 = n2157 | n29563 ;
  assign n51780 = n51779 ^ n51778 ^ 1'b0 ;
  assign n51781 = n18198 & ~n29584 ;
  assign n51787 = n11019 & ~n29924 ;
  assign n51783 = ( ~n10486 & n20506 ) | ( ~n10486 & n39772 ) | ( n20506 & n39772 ) ;
  assign n51784 = n51783 ^ n17917 ^ 1'b0 ;
  assign n51785 = ( n2380 & ~n23612 ) | ( n2380 & n51784 ) | ( ~n23612 & n51784 ) ;
  assign n51782 = ( n15683 & n44520 ) | ( n15683 & ~n46400 ) | ( n44520 & ~n46400 ) ;
  assign n51786 = n51785 ^ n51782 ^ n8019 ;
  assign n51788 = n51787 ^ n51786 ^ n17977 ;
  assign n51789 = n25609 ^ n24178 ^ n5002 ;
  assign n51790 = n27369 ^ n1394 ^ 1'b0 ;
  assign n51791 = n51790 ^ n16787 ^ n9324 ;
  assign n51792 = ( n15470 & ~n28918 ) | ( n15470 & n51791 ) | ( ~n28918 & n51791 ) ;
  assign n51793 = n8362 | n30431 ;
  assign n51794 = ( n4959 & ~n49874 ) | ( n4959 & n51793 ) | ( ~n49874 & n51793 ) ;
  assign n51795 = n1761 | n20458 ;
  assign n51796 = ( n35194 & ~n51794 ) | ( n35194 & n51795 ) | ( ~n51794 & n51795 ) ;
  assign n51797 = ( ~n16881 & n23332 ) | ( ~n16881 & n26085 ) | ( n23332 & n26085 ) ;
  assign n51798 = n4176 & ~n51797 ;
  assign n51799 = n51797 & n51798 ;
  assign n51800 = n51799 ^ n17786 ^ 1'b0 ;
  assign n51801 = n45072 & ~n51800 ;
  assign n51802 = ( n4649 & n8755 ) | ( n4649 & ~n17869 ) | ( n8755 & ~n17869 ) ;
  assign n51803 = ( n37901 & n51801 ) | ( n37901 & ~n51802 ) | ( n51801 & ~n51802 ) ;
  assign n51804 = n23826 ^ n21721 ^ n12295 ;
  assign n51805 = n27011 & n51804 ;
  assign n51806 = n51805 ^ n23671 ^ 1'b0 ;
  assign n51807 = ( ~n6097 & n34302 ) | ( ~n6097 & n41438 ) | ( n34302 & n41438 ) ;
  assign n51808 = n14310 ^ n7735 ^ n5415 ;
  assign n51809 = n45700 ^ n1575 ^ 1'b0 ;
  assign n51810 = ~n40530 & n51809 ;
  assign n51811 = n30886 ^ n25187 ^ n7560 ;
  assign n51812 = ( n1914 & n51810 ) | ( n1914 & ~n51811 ) | ( n51810 & ~n51811 ) ;
  assign n51813 = n49964 ^ n17940 ^ n16002 ;
  assign n51814 = ( n3680 & n13060 ) | ( n3680 & n21479 ) | ( n13060 & n21479 ) ;
  assign n51815 = ~n12430 & n17539 ;
  assign n51816 = n51815 ^ n22221 ^ n1104 ;
  assign n51817 = n51816 ^ n34983 ^ n10051 ;
  assign n51818 = n9300 ^ n8997 ^ 1'b0 ;
  assign n51819 = ( n19878 & ~n20282 ) | ( n19878 & n51818 ) | ( ~n20282 & n51818 ) ;
  assign n51820 = n44704 ^ n15869 ^ 1'b0 ;
  assign n51821 = n45348 & ~n51820 ;
  assign n51822 = n51819 & n51821 ;
  assign n51823 = n39124 & n43369 ;
  assign n51824 = n51823 ^ n36673 ^ 1'b0 ;
  assign n51825 = n6505 | n7757 ;
  assign n51826 = n25053 & ~n51825 ;
  assign n51827 = n1954 & ~n20595 ;
  assign n51828 = n18797 & n51827 ;
  assign n51829 = n12551 & n19166 ;
  assign n51830 = n27099 & n51829 ;
  assign n51831 = ( n51826 & ~n51828 ) | ( n51826 & n51830 ) | ( ~n51828 & n51830 ) ;
  assign n51832 = n14670 ^ n10618 ^ n10004 ;
  assign n51833 = n46194 ^ n30579 ^ n14127 ;
  assign n51834 = n24143 & ~n32459 ;
  assign n51835 = n51834 ^ n27415 ^ n10125 ;
  assign n51836 = ( n22468 & n29299 ) | ( n22468 & n32066 ) | ( n29299 & n32066 ) ;
  assign n51837 = ( n32124 & ~n34199 ) | ( n32124 & n44874 ) | ( ~n34199 & n44874 ) ;
  assign n51838 = n51837 ^ n49732 ^ n10758 ;
  assign n51839 = n10781 ^ n2125 ^ 1'b0 ;
  assign n51840 = n32350 & ~n51839 ;
  assign n51841 = ~n3751 & n48331 ;
  assign n51842 = n5216 & n51841 ;
  assign n51843 = n12590 | n35817 ;
  assign n51844 = n51843 ^ n4628 ^ 1'b0 ;
  assign n51845 = n12949 & n44773 ;
  assign n51846 = n51845 ^ n8422 ^ 1'b0 ;
  assign n51847 = ( ~n16432 & n23994 ) | ( ~n16432 & n35195 ) | ( n23994 & n35195 ) ;
  assign n51848 = ( n1121 & n45027 ) | ( n1121 & n51847 ) | ( n45027 & n51847 ) ;
  assign n51849 = n1982 & ~n22907 ;
  assign n51850 = n51849 ^ n15222 ^ 1'b0 ;
  assign n51851 = n30709 ^ n10897 ^ n5756 ;
  assign n51852 = n21608 & n48337 ;
  assign n51853 = ( n10349 & ~n36968 ) | ( n10349 & n40096 ) | ( ~n36968 & n40096 ) ;
  assign n51854 = n1033 | n35914 ;
  assign n51855 = n14577 & ~n28542 ;
  assign n51856 = n33749 ^ n6861 ^ 1'b0 ;
  assign n51857 = n38701 | n47072 ;
  assign n51858 = n51856 | n51857 ;
  assign n51859 = n51858 ^ n22423 ^ 1'b0 ;
  assign n51860 = n51855 & n51859 ;
  assign n51861 = n2243 | n5403 ;
  assign n51862 = n578 & n32920 ;
  assign n51863 = n51862 ^ n45265 ^ 1'b0 ;
  assign n51864 = ( n16242 & n42649 ) | ( n16242 & ~n51863 ) | ( n42649 & ~n51863 ) ;
  assign n51865 = n49141 ^ n19158 ^ n18243 ;
  assign n51866 = n3117 ^ n2553 ^ 1'b0 ;
  assign n51867 = n12025 & ~n51866 ;
  assign n51868 = n51867 ^ n26343 ^ n7430 ;
  assign n51869 = n51868 ^ n9394 ^ n6651 ;
  assign n51870 = ( ~n10449 & n16289 ) | ( ~n10449 & n19782 ) | ( n16289 & n19782 ) ;
  assign n51871 = n22811 ^ n6749 ^ 1'b0 ;
  assign n51872 = n2619 & ~n51871 ;
  assign n51873 = ( n23879 & ~n51870 ) | ( n23879 & n51872 ) | ( ~n51870 & n51872 ) ;
  assign n51874 = ( n12691 & n51296 ) | ( n12691 & n51873 ) | ( n51296 & n51873 ) ;
  assign n51875 = n46231 ^ n10897 ^ 1'b0 ;
  assign n51876 = ~n39603 & n51875 ;
  assign n51877 = ~n7815 & n17186 ;
  assign n51878 = n10223 & n51877 ;
  assign n51879 = n51878 ^ n43860 ^ 1'b0 ;
  assign n51880 = n51876 & ~n51879 ;
  assign n51881 = n11597 & ~n51880 ;
  assign n51882 = ( n2308 & n14815 ) | ( n2308 & n33601 ) | ( n14815 & n33601 ) ;
  assign n51883 = ~n19264 & n38272 ;
  assign n51884 = ~x132 & n51883 ;
  assign n51885 = n8065 | n28774 ;
  assign n51886 = n38503 & ~n51885 ;
  assign n51887 = n28007 & ~n51886 ;
  assign n51888 = n19964 & n51887 ;
  assign n51889 = ~n19493 & n37678 ;
  assign n51890 = ~n24699 & n51889 ;
  assign n51891 = n36237 ^ n10414 ^ 1'b0 ;
  assign n51892 = n17336 & ~n51891 ;
  assign n51893 = n38747 & n51892 ;
  assign n51894 = ( ~n25767 & n51890 ) | ( ~n25767 & n51893 ) | ( n51890 & n51893 ) ;
  assign n51895 = n49746 ^ n25769 ^ n20109 ;
  assign n51896 = n51895 ^ n13641 ^ 1'b0 ;
  assign n51897 = n6469 ^ n1775 ^ x125 ;
  assign n51898 = n31180 ^ n23237 ^ 1'b0 ;
  assign n51899 = ~n51897 & n51898 ;
  assign n51900 = ( n27917 & ~n49155 ) | ( n27917 & n51899 ) | ( ~n49155 & n51899 ) ;
  assign n51902 = n11428 | n49198 ;
  assign n51901 = ( n10676 & n10974 ) | ( n10676 & ~n27002 ) | ( n10974 & ~n27002 ) ;
  assign n51903 = n51902 ^ n51901 ^ n16191 ;
  assign n51904 = ~n11325 & n45173 ;
  assign n51905 = ~n4468 & n16319 ;
  assign n51906 = n51905 ^ n30022 ^ 1'b0 ;
  assign n51907 = n51906 ^ n8402 ^ 1'b0 ;
  assign n51908 = n51907 ^ n11895 ^ n3072 ;
  assign n51910 = n2024 & ~n13928 ;
  assign n51911 = n24155 & n51910 ;
  assign n51909 = n6980 | n22277 ;
  assign n51912 = n51911 ^ n51909 ^ 1'b0 ;
  assign n51916 = ( n24633 & n25085 ) | ( n24633 & n25157 ) | ( n25085 & n25157 ) ;
  assign n51917 = n51916 ^ n38242 ^ 1'b0 ;
  assign n51913 = n32591 ^ n5080 ^ 1'b0 ;
  assign n51914 = n5069 & ~n51913 ;
  assign n51915 = n37787 & n51914 ;
  assign n51918 = n51917 ^ n51915 ^ 1'b0 ;
  assign n51919 = n40209 ^ n9281 ^ n4682 ;
  assign n51920 = n51919 ^ n4649 ^ 1'b0 ;
  assign n51921 = n9914 & n51920 ;
  assign n51922 = n31536 ^ n1536 ^ 1'b0 ;
  assign n51923 = n30436 | n51922 ;
  assign n51924 = n12292 ^ n7249 ^ 1'b0 ;
  assign n51925 = n38382 & n51924 ;
  assign n51926 = n23205 | n51925 ;
  assign n51927 = n51923 | n51926 ;
  assign n51928 = ( n8814 & ~n19609 ) | ( n8814 & n36964 ) | ( ~n19609 & n36964 ) ;
  assign n51929 = n6810 ^ n635 ^ 1'b0 ;
  assign n51930 = ( n35926 & n48999 ) | ( n35926 & ~n51929 ) | ( n48999 & ~n51929 ) ;
  assign n51931 = ( n12300 & n51928 ) | ( n12300 & n51930 ) | ( n51928 & n51930 ) ;
  assign n51932 = n51931 ^ n14064 ^ n12929 ;
  assign n51933 = n39494 ^ n37932 ^ n34865 ;
  assign n51934 = n14593 & ~n22915 ;
  assign n51935 = n51934 ^ n8045 ^ 1'b0 ;
  assign n51936 = n51935 ^ n14440 ^ n6674 ;
  assign n51937 = ( n29387 & n51933 ) | ( n29387 & n51936 ) | ( n51933 & n51936 ) ;
  assign n51938 = n422 & n23193 ;
  assign n51939 = n44182 ^ n37044 ^ n3732 ;
  assign n51941 = ( n10410 & n38126 ) | ( n10410 & n41548 ) | ( n38126 & n41548 ) ;
  assign n51940 = n36593 ^ n33326 ^ n30401 ;
  assign n51942 = n51941 ^ n51940 ^ n9952 ;
  assign n51943 = ( n16985 & n51126 ) | ( n16985 & n51942 ) | ( n51126 & n51942 ) ;
  assign n51944 = ( ~n6054 & n31329 ) | ( ~n6054 & n51943 ) | ( n31329 & n51943 ) ;
  assign n51945 = n5197 & ~n14253 ;
  assign n51946 = n19144 & n51945 ;
  assign n51947 = n36421 ^ n10865 ^ 1'b0 ;
  assign n51948 = n34747 | n51947 ;
  assign n51949 = n36133 ^ n8529 ^ n6472 ;
  assign n51950 = ( n41633 & ~n41883 ) | ( n41633 & n51949 ) | ( ~n41883 & n51949 ) ;
  assign n51951 = n38843 ^ n11439 ^ n4601 ;
  assign n51952 = n51951 ^ n49240 ^ n41631 ;
  assign n51953 = ( n13730 & n44794 ) | ( n13730 & ~n50231 ) | ( n44794 & ~n50231 ) ;
  assign n51954 = n18069 & ~n47348 ;
  assign n51955 = n51954 ^ n4992 ^ 1'b0 ;
  assign n51956 = n51955 ^ n46600 ^ n31052 ;
  assign n51957 = n32362 ^ n9200 ^ n1090 ;
  assign n51958 = n51957 ^ n43411 ^ 1'b0 ;
  assign n51959 = ( n2079 & ~n15430 ) | ( n2079 & n17505 ) | ( ~n15430 & n17505 ) ;
  assign n51960 = n51959 ^ n34596 ^ 1'b0 ;
  assign n51961 = x111 & n51960 ;
  assign n51962 = n19061 ^ n5374 ^ n1173 ;
  assign n51963 = n51962 ^ n47237 ^ 1'b0 ;
  assign n51964 = n24194 ^ n3085 ^ 1'b0 ;
  assign n51965 = n51963 | n51964 ;
  assign n51966 = ( n32883 & n51961 ) | ( n32883 & n51965 ) | ( n51961 & n51965 ) ;
  assign n51967 = ( n2666 & n19224 ) | ( n2666 & ~n26509 ) | ( n19224 & ~n26509 ) ;
  assign n51968 = ( n5172 & ~n11117 ) | ( n5172 & n51967 ) | ( ~n11117 & n51967 ) ;
  assign n51969 = n51968 ^ n49658 ^ n7114 ;
  assign n51970 = n25148 ^ n24079 ^ 1'b0 ;
  assign n51971 = n41515 | n51970 ;
  assign n51972 = n10973 ^ n2820 ^ 1'b0 ;
  assign n51973 = n36783 | n51972 ;
  assign n51974 = n23614 & ~n51973 ;
  assign n51975 = n51974 ^ n4408 ^ 1'b0 ;
  assign n51976 = ( n32125 & n41701 ) | ( n32125 & ~n47705 ) | ( n41701 & ~n47705 ) ;
  assign n51977 = n32540 ^ n308 ^ 1'b0 ;
  assign n51978 = ~n36778 & n51977 ;
  assign n51979 = n51978 ^ n49087 ^ n41907 ;
  assign n51980 = n48757 ^ n4018 ^ 1'b0 ;
  assign n51981 = ~n7415 & n28580 ;
  assign n51982 = n51981 ^ n5831 ^ 1'b0 ;
  assign n51983 = ( ~n1406 & n32748 ) | ( ~n1406 & n43732 ) | ( n32748 & n43732 ) ;
  assign n51984 = n16687 ^ n1903 ^ 1'b0 ;
  assign n51985 = n51984 ^ n20119 ^ n14144 ;
  assign n51986 = n20212 & n37162 ;
  assign n51987 = n51986 ^ n27532 ^ 1'b0 ;
  assign n51988 = ( ~n23479 & n28373 ) | ( ~n23479 & n37800 ) | ( n28373 & n37800 ) ;
  assign n51989 = n42388 ^ n21238 ^ n6077 ;
  assign n51990 = ( n7650 & n18061 ) | ( n7650 & n23759 ) | ( n18061 & n23759 ) ;
  assign n51991 = n51990 ^ n50673 ^ n17118 ;
  assign n51992 = n17925 ^ n17048 ^ n8370 ;
  assign n51993 = n51992 ^ n51349 ^ n12362 ;
  assign n51994 = n1498 & ~n2697 ;
  assign n51995 = ~n36653 & n51994 ;
  assign n51996 = n15061 | n51995 ;
  assign n51998 = n43226 ^ n8944 ^ 1'b0 ;
  assign n51997 = n24794 ^ n21238 ^ n5600 ;
  assign n51999 = n51998 ^ n51997 ^ 1'b0 ;
  assign n52000 = n9766 | n51999 ;
  assign n52001 = n52000 ^ n46677 ^ 1'b0 ;
  assign n52002 = ~x211 & n48810 ;
  assign n52003 = n19563 | n38289 ;
  assign n52004 = n43419 ^ n28941 ^ n330 ;
  assign n52005 = n52004 ^ n18282 ^ n10517 ;
  assign n52006 = n51728 ^ n5981 ^ n4873 ;
  assign n52007 = n39223 ^ n28917 ^ n17889 ;
  assign n52008 = ( n40257 & ~n46882 ) | ( n40257 & n52007 ) | ( ~n46882 & n52007 ) ;
  assign n52009 = n22242 | n31374 ;
  assign n52010 = n2522 & ~n24876 ;
  assign n52012 = n7573 & ~n10741 ;
  assign n52011 = ( ~n5724 & n10958 ) | ( ~n5724 & n13322 ) | ( n10958 & n13322 ) ;
  assign n52013 = n52012 ^ n52011 ^ n17830 ;
  assign n52014 = n52013 ^ n17005 ^ n11914 ;
  assign n52015 = ( n35252 & n41583 ) | ( n35252 & ~n52014 ) | ( n41583 & ~n52014 ) ;
  assign n52016 = n19378 & n46560 ;
  assign n52017 = ( n26064 & n38391 ) | ( n26064 & ~n38433 ) | ( n38391 & ~n38433 ) ;
  assign n52018 = ( ~n6167 & n8791 ) | ( ~n6167 & n16926 ) | ( n8791 & n16926 ) ;
  assign n52019 = ( n11163 & ~n12212 ) | ( n11163 & n52018 ) | ( ~n12212 & n52018 ) ;
  assign n52020 = n52019 ^ n17067 ^ n16034 ;
  assign n52021 = n43723 ^ n9458 ^ 1'b0 ;
  assign n52022 = ( n15436 & ~n25950 ) | ( n15436 & n50228 ) | ( ~n25950 & n50228 ) ;
  assign n52023 = ( n40209 & n44632 ) | ( n40209 & ~n52022 ) | ( n44632 & ~n52022 ) ;
  assign n52027 = ( n8306 & n14964 ) | ( n8306 & ~n30792 ) | ( n14964 & ~n30792 ) ;
  assign n52026 = n14586 & n50002 ;
  assign n52024 = n32626 ^ n2963 ^ 1'b0 ;
  assign n52025 = n47088 | n52024 ;
  assign n52028 = n52027 ^ n52026 ^ n52025 ;
  assign n52029 = n18911 ^ n17849 ^ n15615 ;
  assign n52030 = ( n18002 & ~n24239 ) | ( n18002 & n31813 ) | ( ~n24239 & n31813 ) ;
  assign n52031 = n52030 ^ n30682 ^ n26008 ;
  assign n52032 = ( ~n46766 & n52029 ) | ( ~n46766 & n52031 ) | ( n52029 & n52031 ) ;
  assign n52033 = n46372 ^ n3163 ^ x32 ;
  assign n52035 = n35122 ^ n1588 ^ 1'b0 ;
  assign n52036 = n39456 & n52035 ;
  assign n52037 = n38043 ^ n22876 ^ 1'b0 ;
  assign n52038 = n29513 & n52037 ;
  assign n52039 = ( n4168 & ~n52036 ) | ( n4168 & n52038 ) | ( ~n52036 & n52038 ) ;
  assign n52034 = n1078 & n14053 ;
  assign n52040 = n52039 ^ n52034 ^ 1'b0 ;
  assign n52041 = n13973 | n45373 ;
  assign n52042 = n9629 & ~n52041 ;
  assign n52043 = ~n29261 & n43096 ;
  assign n52045 = ( n9736 & n10797 ) | ( n9736 & ~n20271 ) | ( n10797 & ~n20271 ) ;
  assign n52044 = ( n19274 & ~n23098 ) | ( n19274 & n23328 ) | ( ~n23098 & n23328 ) ;
  assign n52046 = n52045 ^ n52044 ^ n11915 ;
  assign n52047 = ~n12093 & n46428 ;
  assign n52048 = n47156 ^ n26476 ^ n26008 ;
  assign n52049 = n45067 ^ n3710 ^ 1'b0 ;
  assign n52050 = ( n46761 & n52048 ) | ( n46761 & n52049 ) | ( n52048 & n52049 ) ;
  assign n52051 = ( n1244 & ~n4019 ) | ( n1244 & n39530 ) | ( ~n4019 & n39530 ) ;
  assign n52052 = n31708 ^ n12217 ^ 1'b0 ;
  assign n52053 = n30915 ^ n24205 ^ 1'b0 ;
  assign n52054 = n15314 ^ n3278 ^ 1'b0 ;
  assign n52055 = ~n9818 & n52054 ;
  assign n52056 = n8085 ^ n1622 ^ 1'b0 ;
  assign n52057 = n36825 ^ n2875 ^ 1'b0 ;
  assign n52058 = n52056 & n52057 ;
  assign n52059 = n33294 ^ n22958 ^ 1'b0 ;
  assign n52060 = n44322 ^ n18356 ^ 1'b0 ;
  assign n52061 = n52060 ^ n24443 ^ n12957 ;
  assign n52062 = n37285 ^ n13031 ^ 1'b0 ;
  assign n52063 = ( n12930 & n13636 ) | ( n12930 & n36629 ) | ( n13636 & n36629 ) ;
  assign n52064 = n16779 & ~n52063 ;
  assign n52065 = ( n1819 & n5370 ) | ( n1819 & ~n13363 ) | ( n5370 & ~n13363 ) ;
  assign n52066 = n8826 & ~n52065 ;
  assign n52067 = ( n21226 & n33146 ) | ( n21226 & ~n52066 ) | ( n33146 & ~n52066 ) ;
  assign n52068 = ( n4614 & n34297 ) | ( n4614 & ~n38552 ) | ( n34297 & ~n38552 ) ;
  assign n52069 = n34852 ^ n7306 ^ 1'b0 ;
  assign n52070 = n3840 & ~n52069 ;
  assign n52071 = n4442 & n17762 ;
  assign n52072 = ~n330 & n52071 ;
  assign n52073 = ~n2971 & n11331 ;
  assign n52074 = n52073 ^ n21157 ^ 1'b0 ;
  assign n52075 = n1450 & n27531 ;
  assign n52076 = n21884 ^ n9458 ^ n9179 ;
  assign n52077 = n52076 ^ n34401 ^ 1'b0 ;
  assign n52078 = ~n31240 & n38843 ;
  assign n52079 = ( n1386 & n7385 ) | ( n1386 & ~n49997 ) | ( n7385 & ~n49997 ) ;
  assign n52080 = n52079 ^ n12860 ^ 1'b0 ;
  assign n52081 = n51152 ^ n46243 ^ 1'b0 ;
  assign n52082 = ( n30786 & n51267 ) | ( n30786 & ~n52081 ) | ( n51267 & ~n52081 ) ;
  assign n52083 = n52082 ^ n16481 ^ 1'b0 ;
  assign n52084 = n39303 ^ n22422 ^ 1'b0 ;
  assign n52085 = ~n29120 & n52084 ;
  assign n52086 = n52085 ^ n38973 ^ n19947 ;
  assign n52087 = ~n4571 & n16592 ;
  assign n52088 = n10645 & n52087 ;
  assign n52089 = n13675 ^ n8196 ^ 1'b0 ;
  assign n52090 = ~n8159 & n52089 ;
  assign n52091 = ( ~n529 & n11556 ) | ( ~n529 & n52090 ) | ( n11556 & n52090 ) ;
  assign n52092 = ~n12011 & n20627 ;
  assign n52093 = n29649 & n52092 ;
  assign n52094 = n52093 ^ n3897 ^ 1'b0 ;
  assign n52095 = n52091 | n52094 ;
  assign n52096 = n25614 ^ n19924 ^ 1'b0 ;
  assign n52097 = ( ~n3580 & n50418 ) | ( ~n3580 & n52096 ) | ( n50418 & n52096 ) ;
  assign n52098 = n28491 | n52097 ;
  assign n52099 = n17610 & ~n52098 ;
  assign n52103 = ( n1816 & n42786 ) | ( n1816 & n46569 ) | ( n42786 & n46569 ) ;
  assign n52104 = n52103 ^ n31773 ^ 1'b0 ;
  assign n52100 = n22617 ^ n495 ^ 1'b0 ;
  assign n52101 = n6518 | n52100 ;
  assign n52102 = ( n13723 & n32591 ) | ( n13723 & n52101 ) | ( n32591 & n52101 ) ;
  assign n52105 = n52104 ^ n52102 ^ n19850 ;
  assign n52106 = ( n31510 & n34930 ) | ( n31510 & ~n37514 ) | ( n34930 & ~n37514 ) ;
  assign n52107 = n51342 ^ n34976 ^ n19370 ;
  assign n52108 = n13706 ^ n13135 ^ n2453 ;
  assign n52109 = ( n10184 & ~n14222 ) | ( n10184 & n18031 ) | ( ~n14222 & n18031 ) ;
  assign n52110 = ( ~n43895 & n52108 ) | ( ~n43895 & n52109 ) | ( n52108 & n52109 ) ;
  assign n52111 = n52110 ^ n13869 ^ n1965 ;
  assign n52112 = n19193 ^ n12003 ^ n2897 ;
  assign n52113 = ( n8771 & ~n8845 ) | ( n8771 & n52112 ) | ( ~n8845 & n52112 ) ;
  assign n52114 = ~n15004 & n25503 ;
  assign n52115 = n4197 & ~n19184 ;
  assign n52116 = ~n52114 & n52115 ;
  assign n52117 = n6473 & ~n43635 ;
  assign n52118 = ~n45507 & n52117 ;
  assign n52119 = n35340 ^ n2358 ^ 1'b0 ;
  assign n52120 = n4658 | n25509 ;
  assign n52121 = n9472 | n12392 ;
  assign n52122 = ( n2809 & n10835 ) | ( n2809 & n28075 ) | ( n10835 & n28075 ) ;
  assign n52123 = n14199 ^ n8716 ^ 1'b0 ;
  assign n52124 = ~n52122 & n52123 ;
  assign n52125 = n52124 ^ n9886 ^ 1'b0 ;
  assign n52126 = n35753 ^ n33291 ^ n31098 ;
  assign n52127 = ~n20450 & n25938 ;
  assign n52128 = ~n10495 & n52127 ;
  assign n52129 = n52128 ^ n19469 ^ 1'b0 ;
  assign n52130 = ( n1001 & ~n16881 ) | ( n1001 & n45612 ) | ( ~n16881 & n45612 ) ;
  assign n52131 = ( n15804 & n29248 ) | ( n15804 & ~n35764 ) | ( n29248 & ~n35764 ) ;
  assign n52132 = n52131 ^ n20529 ^ 1'b0 ;
  assign n52133 = n52130 & n52132 ;
  assign n52134 = n5911 & n9847 ;
  assign n52135 = ~n50817 & n52134 ;
  assign n52136 = n25315 & ~n52135 ;
  assign n52137 = n7073 ^ n2021 ^ 1'b0 ;
  assign n52138 = ~n2827 & n52137 ;
  assign n52139 = ( ~n1339 & n3086 ) | ( ~n1339 & n20348 ) | ( n3086 & n20348 ) ;
  assign n52140 = n52139 ^ n28624 ^ n3427 ;
  assign n52141 = n36062 ^ n29754 ^ 1'b0 ;
  assign n52142 = ~n52140 & n52141 ;
  assign n52143 = n16756 ^ n10285 ^ n6757 ;
  assign n52144 = ~n1775 & n52143 ;
  assign n52145 = n52144 ^ n35196 ^ n5416 ;
  assign n52146 = n4272 | n52145 ;
  assign n52147 = n21268 & ~n49992 ;
  assign n52148 = n52147 ^ n24924 ^ 1'b0 ;
  assign n52149 = n52148 ^ n36961 ^ n16927 ;
  assign n52150 = n16894 ^ n3854 ^ 1'b0 ;
  assign n52151 = n52150 ^ n52122 ^ n25918 ;
  assign n52152 = n5210 ^ n3423 ^ n763 ;
  assign n52153 = n52152 ^ n24254 ^ n9552 ;
  assign n52154 = ~n16575 & n52153 ;
  assign n52155 = n52154 ^ n41200 ^ 1'b0 ;
  assign n52156 = ( ~n4537 & n29319 ) | ( ~n4537 & n52155 ) | ( n29319 & n52155 ) ;
  assign n52157 = n40076 ^ n15571 ^ n1449 ;
  assign n52158 = n20525 ^ n11066 ^ n3452 ;
  assign n52159 = n52158 ^ n20908 ^ n2615 ;
  assign n52160 = ~n22529 & n52159 ;
  assign n52161 = ( ~n8169 & n9444 ) | ( ~n8169 & n19995 ) | ( n9444 & n19995 ) ;
  assign n52162 = n41514 ^ n29633 ^ 1'b0 ;
  assign n52163 = ( n13513 & n52161 ) | ( n13513 & ~n52162 ) | ( n52161 & ~n52162 ) ;
  assign n52170 = n14586 ^ n14412 ^ n8577 ;
  assign n52171 = n52170 ^ n35039 ^ 1'b0 ;
  assign n52164 = ( n4106 & n7268 ) | ( n4106 & ~n7898 ) | ( n7268 & ~n7898 ) ;
  assign n52165 = n376 | n24592 ;
  assign n52166 = n37811 & ~n52165 ;
  assign n52167 = n52166 ^ n25950 ^ n6182 ;
  assign n52168 = ( n10067 & n52164 ) | ( n10067 & n52167 ) | ( n52164 & n52167 ) ;
  assign n52169 = n10204 & ~n52168 ;
  assign n52172 = n52171 ^ n52169 ^ 1'b0 ;
  assign n52173 = n4570 & n30907 ;
  assign n52174 = ( n14266 & ~n23755 ) | ( n14266 & n27742 ) | ( ~n23755 & n27742 ) ;
  assign n52175 = n9128 & ~n17891 ;
  assign n52176 = n52175 ^ n18209 ^ 1'b0 ;
  assign n52177 = n27242 ^ n18029 ^ n7868 ;
  assign n52178 = n51119 ^ n31810 ^ n31662 ;
  assign n52179 = ( n1459 & n48656 ) | ( n1459 & ~n52178 ) | ( n48656 & ~n52178 ) ;
  assign n52180 = n30158 ^ n12243 ^ n6089 ;
  assign n52181 = n15149 & ~n35021 ;
  assign n52182 = n52180 & n52181 ;
  assign n52183 = n52182 ^ n34233 ^ 1'b0 ;
  assign n52184 = ( n696 & n9591 ) | ( n696 & n40779 ) | ( n9591 & n40779 ) ;
  assign n52185 = ( n1635 & n30106 ) | ( n1635 & ~n50535 ) | ( n30106 & ~n50535 ) ;
  assign n52186 = n49958 ^ n20331 ^ n9441 ;
  assign n52187 = n52186 ^ n33540 ^ n15381 ;
  assign n52188 = ~n8253 & n52187 ;
  assign n52189 = ( ~n37218 & n49140 ) | ( ~n37218 & n52188 ) | ( n49140 & n52188 ) ;
  assign n52190 = n52189 ^ n8556 ^ n2914 ;
  assign n52191 = ( n51811 & ~n52185 ) | ( n51811 & n52190 ) | ( ~n52185 & n52190 ) ;
  assign n52192 = n8099 ^ n7200 ^ n2802 ;
  assign n52193 = ( n2531 & n5106 ) | ( n2531 & n45413 ) | ( n5106 & n45413 ) ;
  assign n52194 = ( n41945 & n52192 ) | ( n41945 & n52193 ) | ( n52192 & n52193 ) ;
  assign n52195 = n13258 | n45777 ;
  assign n52198 = n21945 ^ n20466 ^ n12876 ;
  assign n52196 = n11710 & n29934 ;
  assign n52197 = n52196 ^ n6439 ^ 1'b0 ;
  assign n52199 = n52198 ^ n52197 ^ n24832 ;
  assign n52200 = n36357 ^ n7938 ^ 1'b0 ;
  assign n52201 = n52199 & ~n52200 ;
  assign n52202 = n12276 ^ n621 ^ 1'b0 ;
  assign n52203 = n15114 & n52202 ;
  assign n52204 = ~n24967 & n26966 ;
  assign n52205 = ~n52203 & n52204 ;
  assign n52206 = n27506 & n32895 ;
  assign n52207 = n25206 ^ n16796 ^ 1'b0 ;
  assign n52208 = n1080 | n3261 ;
  assign n52209 = n8248 & ~n52208 ;
  assign n52210 = ( ~n3106 & n4570 ) | ( ~n3106 & n52209 ) | ( n4570 & n52209 ) ;
  assign n52211 = n52210 ^ n24569 ^ n1862 ;
  assign n52212 = n31020 & ~n32925 ;
  assign n52213 = n37892 & n52212 ;
  assign n52214 = n52213 ^ n46766 ^ n14471 ;
  assign n52215 = ( n1009 & n2952 ) | ( n1009 & ~n23082 ) | ( n2952 & ~n23082 ) ;
  assign n52216 = n52215 ^ n41757 ^ n37337 ;
  assign n52217 = n3497 & ~n8931 ;
  assign n52218 = n52217 ^ n10568 ^ 1'b0 ;
  assign n52219 = ( n287 & n4407 ) | ( n287 & n52218 ) | ( n4407 & n52218 ) ;
  assign n52220 = n52219 ^ n47142 ^ n2583 ;
  assign n52221 = n34226 ^ n32599 ^ n10986 ;
  assign n52222 = n38167 ^ n25663 ^ 1'b0 ;
  assign n52223 = n49993 & ~n52222 ;
  assign n52225 = ( n3955 & n10945 ) | ( n3955 & ~n12907 ) | ( n10945 & ~n12907 ) ;
  assign n52224 = n30882 & n30987 ;
  assign n52226 = n52225 ^ n52224 ^ 1'b0 ;
  assign n52227 = ~n39241 & n43859 ;
  assign n52228 = n39094 & n52227 ;
  assign n52229 = n43213 | n52228 ;
  assign n52230 = n52229 ^ n35556 ^ 1'b0 ;
  assign n52231 = n19193 ^ n5970 ^ n4281 ;
  assign n52232 = ( ~n8427 & n8555 ) | ( ~n8427 & n20872 ) | ( n8555 & n20872 ) ;
  assign n52233 = n21151 | n52232 ;
  assign n52234 = n24175 ^ n6346 ^ 1'b0 ;
  assign n52235 = n29550 & n52234 ;
  assign n52236 = ( ~n15556 & n52233 ) | ( ~n15556 & n52235 ) | ( n52233 & n52235 ) ;
  assign n52237 = n6660 ^ n6042 ^ n585 ;
  assign n52247 = n44939 ^ n26095 ^ n10999 ;
  assign n52244 = n18709 ^ n8340 ^ 1'b0 ;
  assign n52245 = n52244 ^ n44635 ^ n38683 ;
  assign n52246 = n52245 ^ n9890 ^ 1'b0 ;
  assign n52238 = n42026 ^ n19611 ^ n17707 ;
  assign n52239 = n31607 ^ n11498 ^ 1'b0 ;
  assign n52240 = n21426 | n52239 ;
  assign n52241 = n48439 & ~n52240 ;
  assign n52242 = ~n52238 & n52241 ;
  assign n52243 = ( ~n25967 & n50980 ) | ( ~n25967 & n52242 ) | ( n50980 & n52242 ) ;
  assign n52248 = n52247 ^ n52246 ^ n52243 ;
  assign n52249 = ~n3303 & n25949 ;
  assign n52250 = n18791 ^ n7367 ^ n2506 ;
  assign n52251 = n52250 ^ n28186 ^ n22987 ;
  assign n52252 = ( n787 & n29566 ) | ( n787 & ~n45848 ) | ( n29566 & ~n45848 ) ;
  assign n52253 = n16414 & n22048 ;
  assign n52254 = n32951 ^ n7424 ^ 1'b0 ;
  assign n52255 = n598 & n52254 ;
  assign n52256 = n43266 & n52255 ;
  assign n52257 = n52256 ^ n26590 ^ 1'b0 ;
  assign n52258 = n27144 & ~n46523 ;
  assign n52259 = n52258 ^ n20950 ^ 1'b0 ;
  assign n52260 = n18699 ^ n15227 ^ n3748 ;
  assign n52261 = n16104 ^ n2113 ^ 1'b0 ;
  assign n52262 = n24382 ^ n5716 ^ 1'b0 ;
  assign n52263 = n52262 ^ n37207 ^ 1'b0 ;
  assign n52264 = ( n5298 & n7132 ) | ( n5298 & ~n12463 ) | ( n7132 & ~n12463 ) ;
  assign n52265 = n27762 ^ n18865 ^ n4335 ;
  assign n52266 = ( n28458 & n52264 ) | ( n28458 & n52265 ) | ( n52264 & n52265 ) ;
  assign n52267 = n24631 & n52266 ;
  assign n52270 = ~n32147 & n47957 ;
  assign n52271 = n52270 ^ n11985 ^ 1'b0 ;
  assign n52268 = n43522 ^ n25533 ^ n9930 ;
  assign n52269 = n18127 & ~n52268 ;
  assign n52272 = n52271 ^ n52269 ^ n18119 ;
  assign n52273 = n11060 ^ n4986 ^ 1'b0 ;
  assign n52274 = ( ~n18760 & n24852 ) | ( ~n18760 & n52273 ) | ( n24852 & n52273 ) ;
  assign n52275 = n10740 & n42479 ;
  assign n52276 = ( n20845 & ~n30238 ) | ( n20845 & n52275 ) | ( ~n30238 & n52275 ) ;
  assign n52277 = n3562 | n24770 ;
  assign n52278 = n52277 ^ n26106 ^ 1'b0 ;
  assign n52279 = n52278 ^ n4497 ^ 1'b0 ;
  assign n52280 = n38776 ^ n14755 ^ 1'b0 ;
  assign n52281 = n12334 | n52280 ;
  assign n52282 = n31018 ^ n12562 ^ n4177 ;
  assign n52283 = ( n16707 & ~n25988 ) | ( n16707 & n52282 ) | ( ~n25988 & n52282 ) ;
  assign n52284 = n26085 ^ n16991 ^ n6499 ;
  assign n52285 = n52284 ^ n20873 ^ n11081 ;
  assign n52287 = n14198 ^ n5289 ^ 1'b0 ;
  assign n52288 = n1182 & n52287 ;
  assign n52286 = n423 & ~n40152 ;
  assign n52289 = n52288 ^ n52286 ^ 1'b0 ;
  assign n52290 = ( ~n43957 & n52285 ) | ( ~n43957 & n52289 ) | ( n52285 & n52289 ) ;
  assign n52291 = ~n20180 & n31790 ;
  assign n52292 = ( n12128 & ~n49203 ) | ( n12128 & n52291 ) | ( ~n49203 & n52291 ) ;
  assign n52293 = n45843 ^ n11044 ^ n817 ;
  assign n52294 = ( x46 & n2303 ) | ( x46 & n52293 ) | ( n2303 & n52293 ) ;
  assign n52295 = n23984 ^ n3234 ^ 1'b0 ;
  assign n52296 = n41220 ^ n1593 ^ 1'b0 ;
  assign n52297 = ~n14491 & n35392 ;
  assign n52298 = n52297 ^ n39168 ^ 1'b0 ;
  assign n52303 = n7467 ^ n5673 ^ 1'b0 ;
  assign n52304 = n10008 | n52303 ;
  assign n52305 = ( n5554 & ~n7886 ) | ( n5554 & n52304 ) | ( ~n7886 & n52304 ) ;
  assign n52301 = n8923 & ~n32189 ;
  assign n52302 = n31444 & ~n52301 ;
  assign n52306 = n52305 ^ n52302 ^ 1'b0 ;
  assign n52299 = ( n12743 & n20811 ) | ( n12743 & ~n23425 ) | ( n20811 & ~n23425 ) ;
  assign n52300 = n269 & ~n52299 ;
  assign n52307 = n52306 ^ n52300 ^ 1'b0 ;
  assign n52308 = n26665 ^ n5958 ^ 1'b0 ;
  assign n52309 = n51460 & n52308 ;
  assign n52310 = ~n5311 & n12360 ;
  assign n52311 = n28159 | n52310 ;
  assign n52312 = ( n16152 & ~n27297 ) | ( n16152 & n47356 ) | ( ~n27297 & n47356 ) ;
  assign n52313 = ( n41441 & ~n41586 ) | ( n41441 & n52312 ) | ( ~n41586 & n52312 ) ;
  assign n52314 = n39584 ^ n39358 ^ n11520 ;
  assign n52315 = n26159 ^ n25174 ^ n15377 ;
  assign n52316 = ( n50167 & ~n52314 ) | ( n50167 & n52315 ) | ( ~n52314 & n52315 ) ;
  assign n52319 = n50332 ^ n45946 ^ 1'b0 ;
  assign n52317 = n30293 ^ n8542 ^ 1'b0 ;
  assign n52318 = n23981 & ~n52317 ;
  assign n52320 = n52319 ^ n52318 ^ 1'b0 ;
  assign n52321 = n11027 & n52320 ;
  assign n52322 = n28492 ^ n26763 ^ n9670 ;
  assign n52324 = n3883 & ~n13061 ;
  assign n52323 = n51136 ^ n24125 ^ n20916 ;
  assign n52325 = n52324 ^ n52323 ^ 1'b0 ;
  assign n52326 = ( x240 & ~n39236 ) | ( x240 & n52325 ) | ( ~n39236 & n52325 ) ;
  assign n52327 = n2978 | n41330 ;
  assign n52328 = n52327 ^ n32402 ^ n9785 ;
  assign n52329 = ( n5235 & ~n10667 ) | ( n5235 & n24257 ) | ( ~n10667 & n24257 ) ;
  assign n52330 = n39952 ^ n546 ^ 1'b0 ;
  assign n52331 = n11997 & n52330 ;
  assign n52332 = ~n22115 & n30363 ;
  assign n52333 = n52332 ^ n46810 ^ 1'b0 ;
  assign n52334 = n970 & ~n3990 ;
  assign n52335 = n39811 & n52334 ;
  assign n52336 = ( n15194 & ~n29128 ) | ( n15194 & n31159 ) | ( ~n29128 & n31159 ) ;
  assign n52337 = n52336 ^ n47273 ^ n11406 ;
  assign n52340 = n15756 ^ n15372 ^ n3532 ;
  assign n52338 = n51543 ^ n14113 ^ 1'b0 ;
  assign n52339 = n30642 & ~n52338 ;
  assign n52341 = n52340 ^ n52339 ^ n28079 ;
  assign n52342 = n38566 ^ n22819 ^ 1'b0 ;
  assign n52343 = ~n12341 & n52342 ;
  assign n52344 = n42503 ^ n32807 ^ n9524 ;
  assign n52345 = n40634 ^ n5090 ^ n3562 ;
  assign n52346 = n52345 ^ n37326 ^ n2457 ;
  assign n52347 = n52346 ^ n47039 ^ n5556 ;
  assign n52348 = ( n5338 & n12873 ) | ( n5338 & n16666 ) | ( n12873 & n16666 ) ;
  assign n52349 = ~n3990 & n7036 ;
  assign n52350 = n52349 ^ n46517 ^ 1'b0 ;
  assign n52351 = n39947 & ~n41797 ;
  assign n52352 = ~n6849 & n26430 ;
  assign n52353 = n52352 ^ n1077 ^ 1'b0 ;
  assign n52354 = n2067 & ~n41821 ;
  assign n52357 = ~n10330 & n17425 ;
  assign n52358 = ~n7608 & n52357 ;
  assign n52359 = n22403 & ~n52358 ;
  assign n52355 = n46025 ^ n26354 ^ 1'b0 ;
  assign n52356 = n18996 & n52355 ;
  assign n52360 = n52359 ^ n52356 ^ n46440 ;
  assign n52362 = n3028 & ~n45820 ;
  assign n52361 = n32629 ^ n21976 ^ n21777 ;
  assign n52363 = n52362 ^ n52361 ^ n44555 ;
  assign n52364 = n22916 ^ n19462 ^ 1'b0 ;
  assign n52365 = ( n5399 & n36645 ) | ( n5399 & n52364 ) | ( n36645 & n52364 ) ;
  assign n52366 = ( ~n4441 & n6237 ) | ( ~n4441 & n28065 ) | ( n6237 & n28065 ) ;
  assign n52367 = n52366 ^ n2300 ^ 1'b0 ;
  assign n52368 = n52367 ^ n51366 ^ n10478 ;
  assign n52372 = ( n5525 & n18746 ) | ( n5525 & n20956 ) | ( n18746 & n20956 ) ;
  assign n52369 = n9679 & ~n27072 ;
  assign n52370 = ~n34341 & n52369 ;
  assign n52371 = n41848 & ~n52370 ;
  assign n52373 = n52372 ^ n52371 ^ 1'b0 ;
  assign n52374 = n52373 ^ n40094 ^ 1'b0 ;
  assign n52375 = n34458 & n52374 ;
  assign n52376 = n4025 | n36546 ;
  assign n52377 = n49966 | n52376 ;
  assign n52378 = n17150 ^ n16273 ^ 1'b0 ;
  assign n52379 = n23349 & ~n52378 ;
  assign n52380 = ( n2152 & n11859 ) | ( n2152 & n13800 ) | ( n11859 & n13800 ) ;
  assign n52381 = n52379 | n52380 ;
  assign n52382 = n6368 | n24014 ;
  assign n52383 = n52382 ^ n15449 ^ 1'b0 ;
  assign n52384 = n52383 ^ n41395 ^ n27014 ;
  assign n52385 = n23281 ^ n9396 ^ n731 ;
  assign n52386 = n30585 ^ n1946 ^ 1'b0 ;
  assign n52387 = ~n20041 & n48066 ;
  assign n52388 = ~n52386 & n52387 ;
  assign n52389 = ( n598 & n5310 ) | ( n598 & n44464 ) | ( n5310 & n44464 ) ;
  assign n52390 = ( n25481 & n52388 ) | ( n25481 & ~n52389 ) | ( n52388 & ~n52389 ) ;
  assign n52391 = ~n3379 & n13207 ;
  assign n52392 = n1892 & n52391 ;
  assign n52393 = ( ~n7357 & n27857 ) | ( ~n7357 & n52392 ) | ( n27857 & n52392 ) ;
  assign n52394 = n23761 ^ n13703 ^ n3852 ;
  assign n52395 = ( ~n3719 & n52393 ) | ( ~n3719 & n52394 ) | ( n52393 & n52394 ) ;
  assign n52396 = n52395 ^ n38949 ^ n12299 ;
  assign n52397 = ( n23292 & ~n33137 ) | ( n23292 & n43797 ) | ( ~n33137 & n43797 ) ;
  assign n52398 = n42904 ^ n36814 ^ n8907 ;
  assign n52399 = ( ~n2052 & n23290 ) | ( ~n2052 & n52398 ) | ( n23290 & n52398 ) ;
  assign n52400 = ( ~n24248 & n25941 ) | ( ~n24248 & n52399 ) | ( n25941 & n52399 ) ;
  assign n52402 = ( n3789 & ~n9146 ) | ( n3789 & n19337 ) | ( ~n9146 & n19337 ) ;
  assign n52403 = ( n9256 & n17294 ) | ( n9256 & ~n52402 ) | ( n17294 & ~n52402 ) ;
  assign n52401 = ( x0 & ~n10888 ) | ( x0 & n27879 ) | ( ~n10888 & n27879 ) ;
  assign n52404 = n52403 ^ n52401 ^ n27363 ;
  assign n52405 = n2979 & ~n8931 ;
  assign n52406 = n52405 ^ n36912 ^ 1'b0 ;
  assign n52407 = n1760 | n42147 ;
  assign n52408 = ~n37048 & n39909 ;
  assign n52409 = n52408 ^ n2449 ^ 1'b0 ;
  assign n52410 = n9924 ^ n3995 ^ n3945 ;
  assign n52411 = ( n2708 & ~n29293 ) | ( n2708 & n52410 ) | ( ~n29293 & n52410 ) ;
  assign n52412 = ( ~n10656 & n37809 ) | ( ~n10656 & n41420 ) | ( n37809 & n41420 ) ;
  assign n52413 = ( ~n32676 & n35466 ) | ( ~n32676 & n52412 ) | ( n35466 & n52412 ) ;
  assign n52414 = ( n33314 & ~n41934 ) | ( n33314 & n52413 ) | ( ~n41934 & n52413 ) ;
  assign n52415 = n52414 ^ n51374 ^ n13358 ;
  assign n52416 = n38468 ^ n22567 ^ n13532 ;
  assign n52417 = n14994 | n26668 ;
  assign n52418 = n2382 & ~n52417 ;
  assign n52419 = ( ~n38092 & n42351 ) | ( ~n38092 & n52418 ) | ( n42351 & n52418 ) ;
  assign n52420 = n23065 & n36888 ;
  assign n52421 = n20937 & ~n48021 ;
  assign n52422 = n52421 ^ n20119 ^ 1'b0 ;
  assign n52423 = n52422 ^ n6687 ^ 1'b0 ;
  assign n52424 = ( ~n30813 & n34807 ) | ( ~n30813 & n43433 ) | ( n34807 & n43433 ) ;
  assign n52425 = ( n44174 & n48649 ) | ( n44174 & ~n52424 ) | ( n48649 & ~n52424 ) ;
  assign n52426 = n10421 | n42549 ;
  assign n52427 = n52426 ^ n16417 ^ 1'b0 ;
  assign n52428 = n18612 ^ n13801 ^ 1'b0 ;
  assign n52429 = n6616 | n52428 ;
  assign n52430 = n17232 ^ n6495 ^ 1'b0 ;
  assign n52431 = n17548 & n52430 ;
  assign n52432 = ( n2208 & n47015 ) | ( n2208 & n52431 ) | ( n47015 & n52431 ) ;
  assign n52433 = n23289 ^ n15439 ^ n8512 ;
  assign n52434 = n8165 & n52433 ;
  assign n52435 = n52432 & n52434 ;
  assign n52436 = n11983 ^ n4883 ^ n2819 ;
  assign n52437 = ~n9610 & n52436 ;
  assign n52438 = n52437 ^ n50112 ^ n14528 ;
  assign n52439 = ( n2161 & n9499 ) | ( n2161 & ~n20033 ) | ( n9499 & ~n20033 ) ;
  assign n52440 = ( n7375 & n46778 ) | ( n7375 & ~n52439 ) | ( n46778 & ~n52439 ) ;
  assign n52441 = n19971 ^ n17917 ^ n8167 ;
  assign n52443 = n8208 & ~n43824 ;
  assign n52444 = n52443 ^ n1343 ^ 1'b0 ;
  assign n52442 = n7748 & ~n17655 ;
  assign n52445 = n52444 ^ n52442 ^ 1'b0 ;
  assign n52446 = n20693 | n52445 ;
  assign n52447 = ( n18729 & n35534 ) | ( n18729 & ~n40152 ) | ( n35534 & ~n40152 ) ;
  assign n52448 = n51616 ^ n26379 ^ n16978 ;
  assign n52449 = n8880 & n52448 ;
  assign n52450 = ~n26580 & n52449 ;
  assign n52451 = ~n1730 & n11792 ;
  assign n52452 = n52451 ^ n25752 ^ 1'b0 ;
  assign n52453 = n31410 & ~n52452 ;
  assign n52454 = n4177 ^ n1625 ^ 1'b0 ;
  assign n52455 = n13972 & ~n22783 ;
  assign n52456 = n18679 & n52455 ;
  assign n52457 = ( n40232 & n52454 ) | ( n40232 & ~n52456 ) | ( n52454 & ~n52456 ) ;
  assign n52458 = ( n15441 & ~n41504 ) | ( n15441 & n41843 ) | ( ~n41504 & n41843 ) ;
  assign n52459 = n52458 ^ n25535 ^ 1'b0 ;
  assign n52460 = n41623 ^ n15074 ^ 1'b0 ;
  assign n52461 = n6632 | n16511 ;
  assign n52462 = n6730 & n14044 ;
  assign n52464 = n30636 & n51815 ;
  assign n52463 = n39745 & n40354 ;
  assign n52465 = n52464 ^ n52463 ^ 1'b0 ;
  assign n52466 = ( n12050 & n20094 ) | ( n12050 & ~n38538 ) | ( n20094 & ~n38538 ) ;
  assign n52467 = ~n31760 & n52466 ;
  assign n52468 = n22682 & ~n43980 ;
  assign n52469 = n52468 ^ n37556 ^ 1'b0 ;
  assign n52470 = n21572 ^ n5721 ^ 1'b0 ;
  assign n52471 = n10784 ^ n7078 ^ 1'b0 ;
  assign n52472 = n52471 ^ n20699 ^ n7148 ;
  assign n52473 = ( n19288 & ~n52470 ) | ( n19288 & n52472 ) | ( ~n52470 & n52472 ) ;
  assign n52474 = n52473 ^ n39484 ^ 1'b0 ;
  assign n52475 = ( n19725 & ~n22940 ) | ( n19725 & n52474 ) | ( ~n22940 & n52474 ) ;
  assign n52476 = n37802 ^ n14581 ^ n9165 ;
  assign n52477 = n19337 | n52476 ;
  assign n52478 = n732 & ~n9769 ;
  assign n52479 = ( n6106 & n24083 ) | ( n6106 & n33769 ) | ( n24083 & n33769 ) ;
  assign n52480 = n24521 | n37038 ;
  assign n52481 = ( n8175 & n17312 ) | ( n8175 & n52480 ) | ( n17312 & n52480 ) ;
  assign n52482 = ( x181 & n32534 ) | ( x181 & n38201 ) | ( n32534 & n38201 ) ;
  assign n52483 = n52482 ^ n35956 ^ n29569 ;
  assign n52484 = n38171 | n40839 ;
  assign n52485 = ~n11588 & n52484 ;
  assign n52486 = n52485 ^ n5918 ^ 1'b0 ;
  assign n52488 = ~n32948 & n33648 ;
  assign n52489 = ~n43961 & n52488 ;
  assign n52487 = n28476 & ~n50182 ;
  assign n52490 = n52489 ^ n52487 ^ 1'b0 ;
  assign n52491 = ( n4502 & n14601 ) | ( n4502 & n45526 ) | ( n14601 & n45526 ) ;
  assign n52492 = n6604 | n52491 ;
  assign n52493 = n331 & ~n52492 ;
  assign n52494 = ( n5597 & n13514 ) | ( n5597 & ~n47161 ) | ( n13514 & ~n47161 ) ;
  assign n52495 = n27033 & ~n52494 ;
  assign n52496 = ( ~n21627 & n22174 ) | ( ~n21627 & n30961 ) | ( n22174 & n30961 ) ;
  assign n52497 = n34569 ^ n21629 ^ n13107 ;
  assign n52498 = ( n6117 & n40163 ) | ( n6117 & ~n52497 ) | ( n40163 & ~n52497 ) ;
  assign n52499 = n14635 & n25108 ;
  assign n52500 = ( n30334 & n42548 ) | ( n30334 & ~n52499 ) | ( n42548 & ~n52499 ) ;
  assign n52501 = n4428 & ~n8732 ;
  assign n52502 = ( n4867 & n34842 ) | ( n4867 & n52501 ) | ( n34842 & n52501 ) ;
  assign n52503 = n52502 ^ n13744 ^ n1267 ;
  assign n52504 = ( n14341 & ~n21040 ) | ( n14341 & n24227 ) | ( ~n21040 & n24227 ) ;
  assign n52505 = ~n5613 & n8325 ;
  assign n52506 = n52505 ^ n39095 ^ 1'b0 ;
  assign n52507 = n29937 | n34971 ;
  assign n52508 = n48753 ^ n36026 ^ n4271 ;
  assign n52509 = n19321 | n26605 ;
  assign n52510 = ~n23236 & n23587 ;
  assign n52511 = ~n26380 & n52510 ;
  assign n52512 = ( n18082 & ~n52509 ) | ( n18082 & n52511 ) | ( ~n52509 & n52511 ) ;
  assign n52513 = ( ~n828 & n34147 ) | ( ~n828 & n52512 ) | ( n34147 & n52512 ) ;
  assign n52514 = n10927 | n37067 ;
  assign n52515 = n52514 ^ n23442 ^ 1'b0 ;
  assign n52517 = ( n6049 & n29038 ) | ( n6049 & ~n42525 ) | ( n29038 & ~n42525 ) ;
  assign n52516 = n28821 | n40577 ;
  assign n52518 = n52517 ^ n52516 ^ n30585 ;
  assign n52519 = n36280 ^ n24424 ^ 1'b0 ;
  assign n52520 = n52519 ^ n47534 ^ 1'b0 ;
  assign n52521 = n52520 ^ n9859 ^ 1'b0 ;
  assign n52522 = n20631 ^ n5503 ^ 1'b0 ;
  assign n52523 = ~n23987 & n52522 ;
  assign n52524 = n52523 ^ n47482 ^ n7326 ;
  assign n52525 = ( ~n14648 & n22537 ) | ( ~n14648 & n48190 ) | ( n22537 & n48190 ) ;
  assign n52526 = n9454 & n34511 ;
  assign n52528 = ( n10040 & n19568 ) | ( n10040 & n21917 ) | ( n19568 & n21917 ) ;
  assign n52527 = n17800 & ~n19828 ;
  assign n52529 = n52528 ^ n52527 ^ 1'b0 ;
  assign n52530 = n52529 ^ n21949 ^ 1'b0 ;
  assign n52531 = n17999 ^ n12820 ^ n706 ;
  assign n52532 = n52531 ^ n32310 ^ n1897 ;
  assign n52533 = n19574 | n22310 ;
  assign n52534 = n25242 & ~n52533 ;
  assign n52535 = n7503 ^ n6436 ^ 1'b0 ;
  assign n52536 = n52534 | n52535 ;
  assign n52537 = n52536 ^ n41744 ^ 1'b0 ;
  assign n52538 = ( ~n2331 & n18625 ) | ( ~n2331 & n46810 ) | ( n18625 & n46810 ) ;
  assign n52539 = ~n5401 & n52538 ;
  assign n52540 = n51023 ^ n32266 ^ 1'b0 ;
  assign n52541 = ( n8614 & n11472 ) | ( n8614 & ~n52540 ) | ( n11472 & ~n52540 ) ;
  assign n52542 = n47036 ^ n31765 ^ n9810 ;
  assign n52543 = n25554 ^ n7799 ^ n6604 ;
  assign n52544 = n44513 | n52543 ;
  assign n52545 = n9362 | n52544 ;
  assign n52546 = n26661 & ~n52545 ;
  assign n52547 = ( n12207 & ~n18740 ) | ( n12207 & n52546 ) | ( ~n18740 & n52546 ) ;
  assign n52548 = ( n1467 & n5028 ) | ( n1467 & ~n9494 ) | ( n5028 & ~n9494 ) ;
  assign n52549 = n52548 ^ n29126 ^ 1'b0 ;
  assign n52551 = n13772 | n35639 ;
  assign n52550 = n7092 | n34143 ;
  assign n52552 = n52551 ^ n52550 ^ 1'b0 ;
  assign n52553 = n11712 & ~n51729 ;
  assign n52554 = n29205 & n52553 ;
  assign n52555 = ( ~n3467 & n10241 ) | ( ~n3467 & n23783 ) | ( n10241 & n23783 ) ;
  assign n52556 = ( ~n37513 & n38382 ) | ( ~n37513 & n52555 ) | ( n38382 & n52555 ) ;
  assign n52557 = n52556 ^ n34193 ^ n2510 ;
  assign n52559 = x228 & x253 ;
  assign n52560 = n20946 & n52559 ;
  assign n52558 = ( n6401 & n7395 ) | ( n6401 & ~n8660 ) | ( n7395 & ~n8660 ) ;
  assign n52561 = n52560 ^ n52558 ^ n20566 ;
  assign n52562 = ~n1871 & n16066 ;
  assign n52563 = n52562 ^ n30991 ^ 1'b0 ;
  assign n52564 = n52563 ^ n22568 ^ n8403 ;
  assign n52565 = n24590 ^ n15265 ^ n3342 ;
  assign n52566 = n5409 ^ n3334 ^ 1'b0 ;
  assign n52567 = n15449 & ~n52566 ;
  assign n52568 = ( n21774 & n28088 ) | ( n21774 & ~n52567 ) | ( n28088 & ~n52567 ) ;
  assign n52569 = ( n6365 & n23397 ) | ( n6365 & n52568 ) | ( n23397 & n52568 ) ;
  assign n52570 = n30706 ^ n11920 ^ n3290 ;
  assign n52571 = n52570 ^ n43098 ^ n7946 ;
  assign n52572 = ( n6161 & ~n40179 ) | ( n6161 & n52571 ) | ( ~n40179 & n52571 ) ;
  assign n52573 = n52569 & ~n52572 ;
  assign n52574 = n47245 | n48206 ;
  assign n52575 = n21140 | n52574 ;
  assign n52576 = ( n29955 & n35512 ) | ( n29955 & n52575 ) | ( n35512 & n52575 ) ;
  assign n52577 = ~n7789 & n29433 ;
  assign n52578 = n30533 & ~n52577 ;
  assign n52579 = n26338 ^ n11532 ^ n922 ;
  assign n52580 = n21750 ^ n1012 ^ 1'b0 ;
  assign n52581 = n52579 | n52580 ;
  assign n52582 = n43264 ^ n13917 ^ n9649 ;
  assign n52583 = n8722 & n52582 ;
  assign n52584 = n19240 & n19708 ;
  assign n52585 = ~n52583 & n52584 ;
  assign n52586 = n6024 | n23655 ;
  assign n52587 = n52586 ^ n49126 ^ 1'b0 ;
  assign n52588 = ( n8218 & n15703 ) | ( n8218 & n16105 ) | ( n15703 & n16105 ) ;
  assign n52589 = n52588 ^ n48130 ^ n32186 ;
  assign n52590 = ( n12531 & ~n33762 ) | ( n12531 & n51663 ) | ( ~n33762 & n51663 ) ;
  assign n52591 = n52590 ^ n35309 ^ 1'b0 ;
  assign n52592 = n2569 & n9191 ;
  assign n52594 = ( n4722 & n9413 ) | ( n4722 & n15903 ) | ( n9413 & n15903 ) ;
  assign n52595 = n398 & n52594 ;
  assign n52593 = n9666 & ~n43350 ;
  assign n52596 = n52595 ^ n52593 ^ 1'b0 ;
  assign n52597 = ( n24895 & n52592 ) | ( n24895 & n52596 ) | ( n52592 & n52596 ) ;
  assign n52598 = n27486 ^ n20113 ^ 1'b0 ;
  assign n52599 = ~n14558 & n26880 ;
  assign n52600 = ( n2438 & n52598 ) | ( n2438 & ~n52599 ) | ( n52598 & ~n52599 ) ;
  assign n52601 = ( n7365 & n27129 ) | ( n7365 & ~n52600 ) | ( n27129 & ~n52600 ) ;
  assign n52602 = n16230 & n25016 ;
  assign n52603 = n7069 & n52602 ;
  assign n52604 = n35362 ^ n13614 ^ 1'b0 ;
  assign n52605 = n25074 ^ n9694 ^ 1'b0 ;
  assign n52606 = ( n11631 & n17609 ) | ( n11631 & ~n52605 ) | ( n17609 & ~n52605 ) ;
  assign n52607 = n45096 ^ n18349 ^ 1'b0 ;
  assign n52608 = n21391 & ~n52413 ;
  assign n52609 = n7307 & n45619 ;
  assign n52610 = n52609 ^ n7326 ^ 1'b0 ;
  assign n52611 = n11081 & n52610 ;
  assign n52612 = n52611 ^ n35294 ^ 1'b0 ;
  assign n52613 = n21996 & n23271 ;
  assign n52614 = ( ~n15828 & n36035 ) | ( ~n15828 & n36878 ) | ( n36035 & n36878 ) ;
  assign n52615 = ( n6702 & ~n19092 ) | ( n6702 & n52614 ) | ( ~n19092 & n52614 ) ;
  assign n52616 = n46692 ^ n12551 ^ 1'b0 ;
  assign n52617 = n2437 & n52616 ;
  assign n52618 = n22030 & n52617 ;
  assign n52619 = n44259 & n46373 ;
  assign n52620 = n10381 & n52619 ;
  assign n52621 = n52620 ^ n38768 ^ 1'b0 ;
  assign n52622 = n28954 ^ n7753 ^ 1'b0 ;
  assign n52623 = n9554 & ~n52622 ;
  assign n52624 = n52623 ^ n44013 ^ n2010 ;
  assign n52625 = ( n15415 & n17369 ) | ( n15415 & ~n51574 ) | ( n17369 & ~n51574 ) ;
  assign n52626 = ~n304 & n29096 ;
  assign n52627 = n19817 & n52626 ;
  assign n52628 = n52627 ^ n3278 ^ 1'b0 ;
  assign n52629 = n1695 | n32634 ;
  assign n52630 = n8459 & ~n52629 ;
  assign n52631 = ( ~n4915 & n6927 ) | ( ~n4915 & n30260 ) | ( n6927 & n30260 ) ;
  assign n52632 = n793 & n14818 ;
  assign n52633 = n52631 & n52632 ;
  assign n52634 = n39531 ^ n27531 ^ n8403 ;
  assign n52635 = n52634 ^ n13338 ^ n2526 ;
  assign n52636 = n7288 | n12057 ;
  assign n52637 = n10202 | n52636 ;
  assign n52638 = n52637 ^ n5465 ^ 1'b0 ;
  assign n52639 = n18680 ^ n5032 ^ 1'b0 ;
  assign n52640 = n28052 & ~n31212 ;
  assign n52641 = n52640 ^ n44112 ^ 1'b0 ;
  assign n52642 = n52641 ^ n43802 ^ n2804 ;
  assign n52643 = ( ~n12415 & n12749 ) | ( ~n12415 & n15797 ) | ( n12749 & n15797 ) ;
  assign n52644 = n39065 & ~n52643 ;
  assign n52645 = ( n16481 & ~n30675 ) | ( n16481 & n52644 ) | ( ~n30675 & n52644 ) ;
  assign n52646 = ~n22559 & n36773 ;
  assign n52647 = ~n35170 & n52646 ;
  assign n52648 = n13815 & n17718 ;
  assign n52649 = n52648 ^ n36019 ^ 1'b0 ;
  assign n52650 = n36766 ^ n14136 ^ n8190 ;
  assign n52651 = ( n51176 & ~n51967 ) | ( n51176 & n52650 ) | ( ~n51967 & n52650 ) ;
  assign n52652 = ( n3031 & n23624 ) | ( n3031 & n41114 ) | ( n23624 & n41114 ) ;
  assign n52653 = ( n10487 & n20095 ) | ( n10487 & n48533 ) | ( n20095 & n48533 ) ;
  assign n52654 = n40079 ^ n4621 ^ 1'b0 ;
  assign n52655 = ( ~n12394 & n18733 ) | ( ~n12394 & n48801 ) | ( n18733 & n48801 ) ;
  assign n52656 = n19846 & ~n35464 ;
  assign n52657 = n52655 & n52656 ;
  assign n52658 = n52657 ^ n30749 ^ n12229 ;
  assign n52659 = n35081 ^ n28996 ^ 1'b0 ;
  assign n52660 = n17226 & ~n52659 ;
  assign n52661 = n52660 ^ n10200 ^ 1'b0 ;
  assign n52662 = n51596 & n52661 ;
  assign n52663 = n45148 ^ n38443 ^ 1'b0 ;
  assign n52664 = n15720 & n52663 ;
  assign n52665 = ~n550 & n991 ;
  assign n52666 = n52665 ^ n46909 ^ 1'b0 ;
  assign n52667 = n22200 & n25814 ;
  assign n52668 = n18153 ^ n16680 ^ 1'b0 ;
  assign n52669 = ~n10212 & n52668 ;
  assign n52670 = ( n10749 & ~n15274 ) | ( n10749 & n52669 ) | ( ~n15274 & n52669 ) ;
  assign n52672 = n14808 ^ n3781 ^ n1284 ;
  assign n52671 = n4211 | n9350 ;
  assign n52673 = n52672 ^ n52671 ^ n15189 ;
  assign n52674 = n32679 ^ n11526 ^ n4635 ;
  assign n52675 = n52674 ^ n37639 ^ n7764 ;
  assign n52676 = n13106 & n37652 ;
  assign n52677 = n798 & n52676 ;
  assign n52678 = n52677 ^ n49403 ^ 1'b0 ;
  assign n52681 = n26486 ^ n25887 ^ n21918 ;
  assign n52679 = n20939 ^ n14594 ^ x191 ;
  assign n52680 = n52679 ^ n45916 ^ n14772 ;
  assign n52682 = n52681 ^ n52680 ^ n32002 ;
  assign n52683 = n9425 & ~n35141 ;
  assign n52684 = ( n12796 & n13599 ) | ( n12796 & ~n52683 ) | ( n13599 & ~n52683 ) ;
  assign n52685 = ~n6821 & n52684 ;
  assign n52686 = n29155 ^ n12231 ^ 1'b0 ;
  assign n52687 = ~n20622 & n52686 ;
  assign n52688 = n52687 ^ n23234 ^ 1'b0 ;
  assign n52690 = ( ~n645 & n7127 ) | ( ~n645 & n33964 ) | ( n7127 & n33964 ) ;
  assign n52689 = n6107 | n10659 ;
  assign n52691 = n52690 ^ n52689 ^ 1'b0 ;
  assign n52692 = n11494 | n15172 ;
  assign n52693 = n26461 | n52692 ;
  assign n52694 = ( n17798 & n26490 ) | ( n17798 & ~n27664 ) | ( n26490 & ~n27664 ) ;
  assign n52695 = n15537 & n52694 ;
  assign n52696 = n52695 ^ n44902 ^ n24416 ;
  assign n52697 = ( ~n11148 & n18996 ) | ( ~n11148 & n23318 ) | ( n18996 & n23318 ) ;
  assign n52698 = ( n10074 & n29628 ) | ( n10074 & ~n52697 ) | ( n29628 & ~n52697 ) ;
  assign n52699 = n46724 ^ n42770 ^ 1'b0 ;
  assign n52700 = n41583 ^ n31065 ^ n823 ;
  assign n52701 = n42136 | n52700 ;
  assign n52702 = n51661 ^ n2715 ^ 1'b0 ;
  assign n52703 = n30002 ^ n22002 ^ n2606 ;
  assign n52704 = n52703 ^ n35353 ^ n20647 ;
  assign n52705 = n46975 ^ n39853 ^ 1'b0 ;
  assign n52706 = n8276 & ~n50621 ;
  assign n52713 = n40955 ^ n39605 ^ n3508 ;
  assign n52711 = n18188 | n48924 ;
  assign n52707 = n35759 & n38053 ;
  assign n52708 = n52707 ^ n20894 ^ 1'b0 ;
  assign n52709 = n52708 ^ n35061 ^ n8798 ;
  assign n52710 = n52709 ^ n12808 ^ 1'b0 ;
  assign n52712 = n52711 ^ n52710 ^ n5571 ;
  assign n52714 = n52713 ^ n52712 ^ 1'b0 ;
  assign n52715 = n52706 & n52714 ;
  assign n52716 = ~n13983 & n35819 ;
  assign n52717 = n52716 ^ n30366 ^ 1'b0 ;
  assign n52718 = n2179 & n19302 ;
  assign n52719 = n39043 ^ n20932 ^ n6320 ;
  assign n52720 = ( n664 & n6271 ) | ( n664 & ~n9195 ) | ( n6271 & ~n9195 ) ;
  assign n52723 = n12430 ^ n8197 ^ 1'b0 ;
  assign n52724 = ( ~n2132 & n8316 ) | ( ~n2132 & n52723 ) | ( n8316 & n52723 ) ;
  assign n52721 = n14203 & ~n24853 ;
  assign n52722 = n52721 ^ n20941 ^ 1'b0 ;
  assign n52725 = n52724 ^ n52722 ^ n19011 ;
  assign n52726 = ( n31192 & n40081 ) | ( n31192 & n45820 ) | ( n40081 & n45820 ) ;
  assign n52727 = n34542 ^ n27975 ^ 1'b0 ;
  assign n52728 = n40654 | n52727 ;
  assign n52729 = n9472 | n29071 ;
  assign n52730 = n31426 & ~n52729 ;
  assign n52731 = n34000 ^ n24007 ^ 1'b0 ;
  assign n52732 = ~n25846 & n52731 ;
  assign n52733 = n26174 & ~n48903 ;
  assign n52734 = ~n10609 & n52733 ;
  assign n52735 = n43558 ^ n29125 ^ n21628 ;
  assign n52736 = n5275 | n52735 ;
  assign n52737 = ( ~n13334 & n40245 ) | ( ~n13334 & n52736 ) | ( n40245 & n52736 ) ;
  assign n52738 = n46917 & n51500 ;
  assign n52739 = n3699 & n52738 ;
  assign n52740 = ( n5990 & n6158 ) | ( n5990 & n52739 ) | ( n6158 & n52739 ) ;
  assign n52741 = ( n5467 & n26023 ) | ( n5467 & n52740 ) | ( n26023 & n52740 ) ;
  assign n52742 = n15775 ^ n11317 ^ 1'b0 ;
  assign n52743 = n52742 ^ n23905 ^ n13180 ;
  assign n52744 = n6966 & n45036 ;
  assign n52745 = n45802 ^ n24980 ^ n8710 ;
  assign n52746 = ( n11526 & n38906 ) | ( n11526 & n52745 ) | ( n38906 & n52745 ) ;
  assign n52747 = ( n9830 & ~n9838 ) | ( n9830 & n40543 ) | ( ~n9838 & n40543 ) ;
  assign n52748 = ( ~n16774 & n29860 ) | ( ~n16774 & n52747 ) | ( n29860 & n52747 ) ;
  assign n52751 = n30058 ^ n15065 ^ n12406 ;
  assign n52749 = n38757 ^ n26976 ^ n22599 ;
  assign n52750 = n3310 & n52749 ;
  assign n52752 = n52751 ^ n52750 ^ n38853 ;
  assign n52753 = n33128 ^ n961 ^ 1'b0 ;
  assign n52754 = n4614 & n52753 ;
  assign n52755 = n24451 ^ n16931 ^ n3489 ;
  assign n52756 = n52755 ^ n33971 ^ 1'b0 ;
  assign n52757 = ( n21884 & n39901 ) | ( n21884 & n52756 ) | ( n39901 & n52756 ) ;
  assign n52758 = n13887 & ~n17999 ;
  assign n52759 = ~n52757 & n52758 ;
  assign n52760 = n19578 & n41498 ;
  assign n52761 = n31521 & n52760 ;
  assign n52762 = ( n1958 & n37755 ) | ( n1958 & ~n50535 ) | ( n37755 & ~n50535 ) ;
  assign n52763 = n52762 ^ n47333 ^ n18896 ;
  assign n52764 = x238 & n44131 ;
  assign n52765 = n22634 ^ n21025 ^ n11917 ;
  assign n52766 = n52765 ^ n49703 ^ n7946 ;
  assign n52767 = n22424 ^ n21731 ^ n18889 ;
  assign n52770 = n14626 ^ n12704 ^ 1'b0 ;
  assign n52771 = n9271 | n52770 ;
  assign n52768 = ( n10639 & n12975 ) | ( n10639 & n33244 ) | ( n12975 & n33244 ) ;
  assign n52769 = n52768 ^ n37182 ^ n31161 ;
  assign n52772 = n52771 ^ n52769 ^ n15889 ;
  assign n52773 = ( n22003 & n28295 ) | ( n22003 & ~n52772 ) | ( n28295 & ~n52772 ) ;
  assign n52774 = n14630 & n17454 ;
  assign n52775 = n52774 ^ n23047 ^ n7312 ;
  assign n52776 = ( n4169 & n4207 ) | ( n4169 & n52775 ) | ( n4207 & n52775 ) ;
  assign n52777 = n52776 ^ n20724 ^ n6445 ;
  assign n52778 = n17426 ^ n13712 ^ 1'b0 ;
  assign n52780 = n38115 ^ n21750 ^ 1'b0 ;
  assign n52779 = n5153 & n44502 ;
  assign n52781 = n52780 ^ n52779 ^ 1'b0 ;
  assign n52782 = n24680 & n43278 ;
  assign n52783 = n12445 ^ n4957 ^ 1'b0 ;
  assign n52785 = n19271 & n34353 ;
  assign n52786 = n52785 ^ n40819 ^ n4298 ;
  assign n52787 = n2527 | n52786 ;
  assign n52784 = n17944 | n37718 ;
  assign n52788 = n52787 ^ n52784 ^ n35264 ;
  assign n52789 = n5859 & ~n14523 ;
  assign n52790 = ~n31871 & n46261 ;
  assign n52791 = n44489 ^ n28723 ^ n1871 ;
  assign n52792 = ( n18484 & n22446 ) | ( n18484 & ~n47118 ) | ( n22446 & ~n47118 ) ;
  assign n52793 = ( n38874 & n52791 ) | ( n38874 & ~n52792 ) | ( n52791 & ~n52792 ) ;
  assign n52794 = n30956 & n50658 ;
  assign n52795 = n52794 ^ n51516 ^ n5639 ;
  assign n52796 = ( n49296 & n52793 ) | ( n49296 & n52795 ) | ( n52793 & n52795 ) ;
  assign n52797 = n44319 ^ n10805 ^ 1'b0 ;
  assign n52798 = n29250 | n52797 ;
  assign n52799 = ( n1209 & n40149 ) | ( n1209 & n52798 ) | ( n40149 & n52798 ) ;
  assign n52800 = ( n40972 & n45573 ) | ( n40972 & ~n52799 ) | ( n45573 & ~n52799 ) ;
  assign n52801 = ( ~n3526 & n12020 ) | ( ~n3526 & n20497 ) | ( n12020 & n20497 ) ;
  assign n52805 = n28817 ^ n28453 ^ n24517 ;
  assign n52802 = n3917 & n23374 ;
  assign n52803 = ~n7173 & n52802 ;
  assign n52804 = n29327 | n52803 ;
  assign n52806 = n52805 ^ n52804 ^ 1'b0 ;
  assign n52808 = n24641 ^ n9986 ^ n343 ;
  assign n52807 = n10233 & ~n43740 ;
  assign n52809 = n52808 ^ n52807 ^ 1'b0 ;
  assign n52810 = ( ~n6604 & n18760 ) | ( ~n6604 & n52809 ) | ( n18760 & n52809 ) ;
  assign n52811 = ( n4668 & n24150 ) | ( n4668 & ~n52810 ) | ( n24150 & ~n52810 ) ;
  assign n52812 = ~n4585 & n11175 ;
  assign n52813 = n52811 & n52812 ;
  assign n52815 = ~n3276 & n12268 ;
  assign n52816 = n52815 ^ n3472 ^ 1'b0 ;
  assign n52817 = n52816 ^ n19398 ^ n15114 ;
  assign n52814 = n18689 & n48505 ;
  assign n52818 = n52817 ^ n52814 ^ 1'b0 ;
  assign n52819 = ( n10625 & n18859 ) | ( n10625 & n28394 ) | ( n18859 & n28394 ) ;
  assign n52820 = ~n15598 & n52819 ;
  assign n52821 = ~n991 & n52820 ;
  assign n52822 = n7839 & n34916 ;
  assign n52823 = n52822 ^ n11722 ^ 1'b0 ;
  assign n52824 = ( ~n1700 & n3279 ) | ( ~n1700 & n52823 ) | ( n3279 & n52823 ) ;
  assign n52825 = ( n13416 & ~n33118 ) | ( n13416 & n52824 ) | ( ~n33118 & n52824 ) ;
  assign n52828 = n32521 ^ n9185 ^ n2508 ;
  assign n52826 = n36424 & n45113 ;
  assign n52827 = n52826 ^ n15194 ^ 1'b0 ;
  assign n52829 = n52828 ^ n52827 ^ n6465 ;
  assign n52830 = n16773 ^ n12082 ^ n2381 ;
  assign n52832 = n13267 ^ n4529 ^ n4164 ;
  assign n52833 = n52832 ^ n24092 ^ n2521 ;
  assign n52834 = n52833 ^ n18206 ^ n4700 ;
  assign n52831 = n38703 ^ n21679 ^ n4248 ;
  assign n52835 = n52834 ^ n52831 ^ 1'b0 ;
  assign n52837 = ~n3737 & n22886 ;
  assign n52838 = n52837 ^ n16197 ^ 1'b0 ;
  assign n52836 = n10903 | n15486 ;
  assign n52839 = n52838 ^ n52836 ^ 1'b0 ;
  assign n52840 = ~n30971 & n52839 ;
  assign n52842 = n9364 | n11536 ;
  assign n52843 = n3927 & ~n52842 ;
  assign n52841 = ( ~n12907 & n15624 ) | ( ~n12907 & n46560 ) | ( n15624 & n46560 ) ;
  assign n52844 = n52843 ^ n52841 ^ n38348 ;
  assign n52845 = n9153 & n18598 ;
  assign n52846 = n33127 & n52845 ;
  assign n52847 = n52846 ^ n32472 ^ 1'b0 ;
  assign n52848 = ( n15228 & ~n28643 ) | ( n15228 & n52847 ) | ( ~n28643 & n52847 ) ;
  assign n52849 = n51884 ^ n2824 ^ 1'b0 ;
  assign n52850 = n18242 & n52849 ;
  assign n52851 = x181 & ~n8588 ;
  assign n52852 = n27971 ^ n17151 ^ n3757 ;
  assign n52853 = n52852 ^ n35930 ^ 1'b0 ;
  assign n52854 = n13614 & n52853 ;
  assign n52855 = n52854 ^ n6593 ^ 1'b0 ;
  assign n52856 = n13145 & ~n52855 ;
  assign n52857 = n9691 | n28744 ;
  assign n52858 = n29797 ^ n645 ^ 1'b0 ;
  assign n52859 = ( n9560 & ~n50479 ) | ( n9560 & n52858 ) | ( ~n50479 & n52858 ) ;
  assign n52860 = ~n5878 & n50484 ;
  assign n52861 = ~n11373 & n21950 ;
  assign n52862 = ~n16267 & n52861 ;
  assign n52863 = ( ~n8134 & n19987 ) | ( ~n8134 & n52862 ) | ( n19987 & n52862 ) ;
  assign n52864 = n23753 ^ n1355 ^ 1'b0 ;
  assign n52865 = ( ~n6282 & n12429 ) | ( ~n6282 & n52864 ) | ( n12429 & n52864 ) ;
  assign n52866 = n21717 ^ n10471 ^ n10431 ;
  assign n52867 = ( n21354 & n27076 ) | ( n21354 & n28076 ) | ( n27076 & n28076 ) ;
  assign n52868 = n38027 ^ n33910 ^ n33738 ;
  assign n52869 = ( n52866 & n52867 ) | ( n52866 & n52868 ) | ( n52867 & n52868 ) ;
  assign n52870 = n52869 ^ n45849 ^ n29900 ;
  assign n52871 = n9048 & n44290 ;
  assign n52873 = n10573 | n23010 ;
  assign n52874 = n9370 & ~n52873 ;
  assign n52872 = n20049 ^ n6602 ^ 1'b0 ;
  assign n52875 = n52874 ^ n52872 ^ n17126 ;
  assign n52876 = n52875 ^ n7294 ^ n5332 ;
  assign n52877 = ( ~n19387 & n52871 ) | ( ~n19387 & n52876 ) | ( n52871 & n52876 ) ;
  assign n52878 = n29261 ^ n27844 ^ n5557 ;
  assign n52879 = ( n44671 & ~n45974 ) | ( n44671 & n52878 ) | ( ~n45974 & n52878 ) ;
  assign n52880 = n21964 ^ n1170 ^ 1'b0 ;
  assign n52881 = n1691 & ~n52880 ;
  assign n52882 = n25335 ^ n23267 ^ 1'b0 ;
  assign n52883 = ~n41337 & n52882 ;
  assign n52884 = n5635 & ~n50385 ;
  assign n52885 = n28592 & n52884 ;
  assign n52886 = n4032 & n42917 ;
  assign n52887 = n8387 ^ n6495 ^ n3120 ;
  assign n52888 = n52887 ^ n39367 ^ n18155 ;
  assign n52889 = n52888 ^ n36028 ^ n462 ;
  assign n52890 = ( n11448 & n13564 ) | ( n11448 & n33130 ) | ( n13564 & n33130 ) ;
  assign n52891 = ( n12335 & ~n25520 ) | ( n12335 & n45378 ) | ( ~n25520 & n45378 ) ;
  assign n52893 = ( ~n415 & n5386 ) | ( ~n415 & n9148 ) | ( n5386 & n9148 ) ;
  assign n52894 = ( n993 & ~n9930 ) | ( n993 & n52893 ) | ( ~n9930 & n52893 ) ;
  assign n52892 = ( n6684 & n22073 ) | ( n6684 & n30621 ) | ( n22073 & n30621 ) ;
  assign n52895 = n52894 ^ n52892 ^ n42390 ;
  assign n52896 = ( n1200 & n24086 ) | ( n1200 & ~n43343 ) | ( n24086 & ~n43343 ) ;
  assign n52897 = ( n15780 & ~n24675 ) | ( n15780 & n52896 ) | ( ~n24675 & n52896 ) ;
  assign n52898 = n36886 ^ n12103 ^ 1'b0 ;
  assign n52899 = n42483 ^ n8846 ^ n1230 ;
  assign n52900 = n50569 ^ n21326 ^ 1'b0 ;
  assign n52901 = n52899 | n52900 ;
  assign n52902 = n21510 ^ n8171 ^ n4257 ;
  assign n52903 = n52902 ^ n14026 ^ x43 ;
  assign n52904 = n41245 ^ n9629 ^ 1'b0 ;
  assign n52905 = n21683 ^ n17053 ^ 1'b0 ;
  assign n52906 = ~n52904 & n52905 ;
  assign n52907 = n52906 ^ n1096 ^ 1'b0 ;
  assign n52908 = n52907 ^ n15873 ^ 1'b0 ;
  assign n52909 = n52908 ^ n52712 ^ n16254 ;
  assign n52910 = n51080 ^ n42460 ^ 1'b0 ;
  assign n52911 = n18963 & ~n40122 ;
  assign n52912 = n52911 ^ n23293 ^ 1'b0 ;
  assign n52913 = n52912 ^ n6956 ^ 1'b0 ;
  assign n52914 = n52572 ^ n2447 ^ 1'b0 ;
  assign n52915 = n28419 ^ n2643 ^ 1'b0 ;
  assign n52916 = ( n7492 & n9018 ) | ( n7492 & n33619 ) | ( n9018 & n33619 ) ;
  assign n52917 = n52916 ^ n16245 ^ 1'b0 ;
  assign n52918 = ~n13335 & n52917 ;
  assign n52919 = n52916 ^ n43536 ^ 1'b0 ;
  assign n52920 = ( n13193 & ~n14755 ) | ( n13193 & n43422 ) | ( ~n14755 & n43422 ) ;
  assign n52923 = n46764 ^ n23683 ^ 1'b0 ;
  assign n52924 = n34367 | n52923 ;
  assign n52921 = n23331 ^ n11614 ^ n498 ;
  assign n52922 = n52921 ^ n22714 ^ n11378 ;
  assign n52925 = n52924 ^ n52922 ^ n9324 ;
  assign n52926 = n44896 ^ n23809 ^ n15456 ;
  assign n52927 = n7853 & ~n42574 ;
  assign n52928 = ~n2341 & n9802 ;
  assign n52929 = n37606 ^ n28560 ^ n7926 ;
  assign n52930 = ~n18702 & n52929 ;
  assign n52931 = n52930 ^ n36403 ^ 1'b0 ;
  assign n52932 = n42837 ^ n14544 ^ 1'b0 ;
  assign n52933 = n26518 ^ n19813 ^ 1'b0 ;
  assign n52934 = n52932 | n52933 ;
  assign n52935 = n4060 | n40598 ;
  assign n52936 = n52935 ^ n20826 ^ 1'b0 ;
  assign n52937 = n21298 ^ n15345 ^ n9490 ;
  assign n52938 = ( ~n10836 & n34168 ) | ( ~n10836 & n52937 ) | ( n34168 & n52937 ) ;
  assign n52939 = n52938 ^ n12245 ^ 1'b0 ;
  assign n52940 = n32035 & ~n52939 ;
  assign n52941 = n15983 & n52940 ;
  assign n52942 = n52941 ^ n27406 ^ 1'b0 ;
  assign n52944 = ( n16242 & n16433 ) | ( n16242 & ~n51058 ) | ( n16433 & ~n51058 ) ;
  assign n52945 = ( n7761 & n7999 ) | ( n7761 & ~n52944 ) | ( n7999 & ~n52944 ) ;
  assign n52943 = n23226 ^ n18791 ^ n16782 ;
  assign n52946 = n52945 ^ n52943 ^ n40921 ;
  assign n52947 = n5341 & ~n27669 ;
  assign n52948 = ~n16316 & n52947 ;
  assign n52949 = ( ~n21765 & n48094 ) | ( ~n21765 & n52948 ) | ( n48094 & n52948 ) ;
  assign n52950 = n52949 ^ n32720 ^ 1'b0 ;
  assign n52951 = n21529 ^ n10401 ^ 1'b0 ;
  assign n52952 = n52951 ^ n45646 ^ n13824 ;
  assign n52953 = n46940 ^ n20440 ^ 1'b0 ;
  assign n52954 = n52953 ^ n35811 ^ n12075 ;
  assign n52955 = ( n27104 & ~n43293 ) | ( n27104 & n52954 ) | ( ~n43293 & n52954 ) ;
  assign n52956 = n2125 & ~n6420 ;
  assign n52957 = ( n3819 & n9211 ) | ( n3819 & ~n52956 ) | ( n9211 & ~n52956 ) ;
  assign n52958 = ( n9749 & ~n48404 ) | ( n9749 & n52957 ) | ( ~n48404 & n52957 ) ;
  assign n52959 = n24657 ^ n18185 ^ 1'b0 ;
  assign n52960 = n4568 & n27108 ;
  assign n52961 = n52960 ^ n2360 ^ 1'b0 ;
  assign n52962 = n7387 & n18889 ;
  assign n52963 = n50010 & n52962 ;
  assign n52964 = n33143 ^ n15100 ^ x81 ;
  assign n52965 = n16325 ^ n1553 ^ 1'b0 ;
  assign n52966 = ( ~n3677 & n4501 ) | ( ~n3677 & n10024 ) | ( n4501 & n10024 ) ;
  assign n52967 = ( n14325 & n25349 ) | ( n14325 & n52966 ) | ( n25349 & n52966 ) ;
  assign n52968 = ( n52964 & n52965 ) | ( n52964 & n52967 ) | ( n52965 & n52967 ) ;
  assign n52969 = n32798 ^ n32223 ^ n6148 ;
  assign n52970 = ( ~n25558 & n43559 ) | ( ~n25558 & n47146 ) | ( n43559 & n47146 ) ;
  assign n52971 = n19806 & n44394 ;
  assign n52972 = n43738 ^ n12002 ^ n7313 ;
  assign n52973 = n52972 ^ n47368 ^ 1'b0 ;
  assign n52974 = n41531 ^ n31007 ^ n18257 ;
  assign n52975 = ( ~n45096 & n48965 ) | ( ~n45096 & n52974 ) | ( n48965 & n52974 ) ;
  assign n52976 = n6735 | n36068 ;
  assign n52977 = ( ~n14267 & n15628 ) | ( ~n14267 & n23933 ) | ( n15628 & n23933 ) ;
  assign n52978 = n52977 ^ n28794 ^ n20758 ;
  assign n52979 = ~n47325 & n52978 ;
  assign n52980 = n7553 | n9391 ;
  assign n52981 = n29228 & ~n41785 ;
  assign n52982 = n52981 ^ n22509 ^ 1'b0 ;
  assign n52983 = n46880 ^ n38089 ^ n3319 ;
  assign n52984 = ~n26825 & n29427 ;
  assign n52985 = n48683 ^ n22600 ^ n15354 ;
  assign n52986 = ( n15450 & n17229 ) | ( n15450 & ~n49155 ) | ( n17229 & ~n49155 ) ;
  assign n52987 = ~n2150 & n51419 ;
  assign n52988 = n26306 & n52987 ;
  assign n52989 = ( n23540 & ~n51933 ) | ( n23540 & n52988 ) | ( ~n51933 & n52988 ) ;
  assign n52990 = n52989 ^ n16069 ^ n2941 ;
  assign n52991 = n45995 ^ n21490 ^ n14976 ;
  assign n52992 = n47547 ^ n40718 ^ n32319 ;
  assign n52995 = n6810 & ~n12186 ;
  assign n52993 = ~n6927 & n26770 ;
  assign n52994 = ~n11355 & n52993 ;
  assign n52996 = n52995 ^ n52994 ^ 1'b0 ;
  assign n52997 = n19592 ^ n16402 ^ n1612 ;
  assign n52998 = n48404 ^ n42711 ^ 1'b0 ;
  assign n52999 = n52997 & ~n52998 ;
  assign n53000 = ~n24038 & n32610 ;
  assign n53001 = ( n7827 & ~n15954 ) | ( n7827 & n53000 ) | ( ~n15954 & n53000 ) ;
  assign n53002 = ( n6512 & n9202 ) | ( n6512 & ~n10305 ) | ( n9202 & ~n10305 ) ;
  assign n53003 = n47787 ^ n14960 ^ 1'b0 ;
  assign n53004 = n53003 ^ n10570 ^ n5432 ;
  assign n53005 = ( n6450 & n25350 ) | ( n6450 & ~n44972 ) | ( n25350 & ~n44972 ) ;
  assign n53006 = n17476 & ~n21748 ;
  assign n53007 = n53006 ^ n21303 ^ n2377 ;
  assign n53008 = n25207 ^ n23451 ^ 1'b0 ;
  assign n53009 = n43489 | n53008 ;
  assign n53010 = n42159 ^ n12259 ^ 1'b0 ;
  assign n53011 = ~n12742 & n53010 ;
  assign n53012 = n53011 ^ n28941 ^ 1'b0 ;
  assign n53013 = ( ~n45125 & n53009 ) | ( ~n45125 & n53012 ) | ( n53009 & n53012 ) ;
  assign n53014 = n25177 ^ n8034 ^ 1'b0 ;
  assign n53015 = n53014 ^ n33230 ^ n4855 ;
  assign n53016 = n53015 ^ n45507 ^ n29586 ;
  assign n53017 = ~n23943 & n50681 ;
  assign n53018 = n53017 ^ n38446 ^ 1'b0 ;
  assign n53019 = n11575 ^ n8830 ^ n5760 ;
  assign n53022 = n21768 ^ n10863 ^ n5579 ;
  assign n53020 = n30501 ^ n23940 ^ n1567 ;
  assign n53021 = n10423 & n53020 ;
  assign n53023 = n53022 ^ n53021 ^ 1'b0 ;
  assign n53024 = n53019 & n53023 ;
  assign n53025 = n48679 ^ n37645 ^ n16894 ;
  assign n53026 = n53025 ^ n17584 ^ n15503 ;
  assign n53027 = n7359 ^ n6083 ^ 1'b0 ;
  assign n53028 = n11520 | n53027 ;
  assign n53029 = n6375 ^ n1422 ^ 1'b0 ;
  assign n53030 = ~n53028 & n53029 ;
  assign n53031 = n53030 ^ n49995 ^ n38276 ;
  assign n53032 = ( ~n16839 & n26622 ) | ( ~n16839 & n45777 ) | ( n26622 & n45777 ) ;
  assign n53033 = ( n17446 & n22338 ) | ( n17446 & ~n51256 ) | ( n22338 & ~n51256 ) ;
  assign n53034 = n19953 ^ n8630 ^ n7178 ;
  assign n53035 = n53034 ^ n18619 ^ n2848 ;
  assign n53036 = ( ~n18322 & n39053 ) | ( ~n18322 & n53035 ) | ( n39053 & n53035 ) ;
  assign n53037 = n43398 ^ n39353 ^ n10144 ;
  assign n53038 = ( n6139 & n12889 ) | ( n6139 & ~n53037 ) | ( n12889 & ~n53037 ) ;
  assign n53039 = n13748 & n22708 ;
  assign n53040 = n20174 & n53039 ;
  assign n53041 = n33343 & n44220 ;
  assign n53042 = n10677 & n53041 ;
  assign n53044 = n3441 | n4537 ;
  assign n53045 = n27296 | n53044 ;
  assign n53043 = n30441 ^ n22036 ^ n5991 ;
  assign n53046 = n53045 ^ n53043 ^ n47083 ;
  assign n53047 = n24724 & ~n53046 ;
  assign n53052 = n19441 ^ n4774 ^ n3137 ;
  assign n53049 = ( n9640 & n12755 ) | ( n9640 & ~n33766 ) | ( n12755 & ~n33766 ) ;
  assign n53050 = n53049 ^ n30897 ^ n12044 ;
  assign n53048 = n11622 | n22200 ;
  assign n53051 = n53050 ^ n53048 ^ 1'b0 ;
  assign n53053 = n53052 ^ n53051 ^ n31750 ;
  assign n53054 = n16707 ^ n12819 ^ n9746 ;
  assign n53055 = ( n969 & n18487 ) | ( n969 & n33458 ) | ( n18487 & n33458 ) ;
  assign n53056 = x187 & ~n47229 ;
  assign n53057 = n53056 ^ n29037 ^ 1'b0 ;
  assign n53058 = ( n20272 & n53055 ) | ( n20272 & n53057 ) | ( n53055 & n53057 ) ;
  assign n53059 = ( n312 & n4079 ) | ( n312 & ~n10776 ) | ( n4079 & ~n10776 ) ;
  assign n53060 = ( n1985 & n6968 ) | ( n1985 & ~n20601 ) | ( n6968 & ~n20601 ) ;
  assign n53061 = ( ~n44017 & n53059 ) | ( ~n44017 & n53060 ) | ( n53059 & n53060 ) ;
  assign n53062 = n53061 ^ n17889 ^ n17378 ;
  assign n53063 = n27129 ^ n16130 ^ 1'b0 ;
  assign n53064 = n38783 ^ n34823 ^ n18825 ;
  assign n53065 = ( n15298 & n38924 ) | ( n15298 & n53064 ) | ( n38924 & n53064 ) ;
  assign n53066 = n53065 ^ n48744 ^ n10326 ;
  assign n53067 = n32843 ^ n22246 ^ 1'b0 ;
  assign n53068 = ~n18348 & n53067 ;
  assign n53069 = ~n5216 & n16429 ;
  assign n53070 = n53069 ^ n28614 ^ 1'b0 ;
  assign n53071 = n40839 ^ n29418 ^ 1'b0 ;
  assign n53072 = n44905 ^ n42800 ^ n30123 ;
  assign n53073 = n11553 ^ n4523 ^ 1'b0 ;
  assign n53074 = n53073 ^ n25637 ^ 1'b0 ;
  assign n53075 = n4951 | n22427 ;
  assign n53076 = n53075 ^ n21737 ^ n4362 ;
  assign n53077 = n52004 ^ n15868 ^ n6437 ;
  assign n53078 = n47380 ^ x184 ^ 1'b0 ;
  assign n53079 = n52531 & n53078 ;
  assign n53080 = ( ~n13094 & n19260 ) | ( ~n13094 & n20973 ) | ( n19260 & n20973 ) ;
  assign n53081 = ( ~n21473 & n35272 ) | ( ~n21473 & n53080 ) | ( n35272 & n53080 ) ;
  assign n53082 = ( n3857 & n13589 ) | ( n3857 & ~n21264 ) | ( n13589 & ~n21264 ) ;
  assign n53083 = n53082 ^ n18597 ^ 1'b0 ;
  assign n53084 = n33294 ^ n12044 ^ 1'b0 ;
  assign n53085 = n53084 ^ n47953 ^ n14270 ;
  assign n53086 = n53085 ^ n14741 ^ 1'b0 ;
  assign n53087 = n29663 & n53086 ;
  assign n53088 = n15885 | n21729 ;
  assign n53089 = n46736 | n53088 ;
  assign n53090 = n16829 | n26817 ;
  assign n53091 = n36108 ^ n4583 ^ 1'b0 ;
  assign n53092 = n53091 ^ n50839 ^ n8310 ;
  assign n53093 = ( n984 & n10635 ) | ( n984 & n29681 ) | ( n10635 & n29681 ) ;
  assign n53094 = n53093 ^ n27296 ^ n3397 ;
  assign n53095 = ( n32138 & n42704 ) | ( n32138 & n53094 ) | ( n42704 & n53094 ) ;
  assign n53096 = n1469 & n16810 ;
  assign n53097 = n3385 & ~n46287 ;
  assign n53098 = ( n28168 & n53096 ) | ( n28168 & n53097 ) | ( n53096 & n53097 ) ;
  assign n53099 = n53098 ^ n29135 ^ n11617 ;
  assign n53100 = n46677 ^ n45444 ^ n13263 ;
  assign n53101 = n15281 ^ n7265 ^ 1'b0 ;
  assign n53102 = ( n19246 & n41612 ) | ( n19246 & n53101 ) | ( n41612 & n53101 ) ;
  assign n53103 = n15017 ^ n7726 ^ 1'b0 ;
  assign n53104 = ~n482 & n2221 ;
  assign n53105 = n53104 ^ n11210 ^ 1'b0 ;
  assign n53106 = n53105 ^ n29838 ^ 1'b0 ;
  assign n53108 = ( n2527 & ~n4101 ) | ( n2527 & n21763 ) | ( ~n4101 & n21763 ) ;
  assign n53107 = n44752 & ~n47859 ;
  assign n53109 = n53108 ^ n53107 ^ 1'b0 ;
  assign n53110 = n42819 ^ n30884 ^ n28549 ;
  assign n53111 = n19712 ^ n2976 ^ 1'b0 ;
  assign n53112 = n35090 & n53111 ;
  assign n53113 = n43119 & n53112 ;
  assign n53115 = n12036 ^ n5719 ^ 1'b0 ;
  assign n53116 = n26070 & ~n53115 ;
  assign n53114 = ~n35174 & n45641 ;
  assign n53117 = n53116 ^ n53114 ^ n20233 ;
  assign n53118 = n11919 ^ n7240 ^ n3547 ;
  assign n53119 = n13581 ^ n2827 ^ 1'b0 ;
  assign n53120 = n19943 & ~n53119 ;
  assign n53121 = n53120 ^ n34907 ^ n33214 ;
  assign n53122 = n7143 | n19155 ;
  assign n53123 = n53122 ^ n3023 ^ 1'b0 ;
  assign n53124 = ( n4410 & n36411 ) | ( n4410 & ~n53123 ) | ( n36411 & ~n53123 ) ;
  assign n53125 = n53124 ^ n46066 ^ n2288 ;
  assign n53126 = ( n1542 & ~n15296 ) | ( n1542 & n51053 ) | ( ~n15296 & n51053 ) ;
  assign n53127 = n26000 ^ n24979 ^ 1'b0 ;
  assign n53128 = n2843 & n53127 ;
  assign n53129 = n8148 & n12911 ;
  assign n53130 = n5630 & n53129 ;
  assign n53131 = n41120 ^ n23159 ^ n19303 ;
  assign n53132 = n37043 & n37824 ;
  assign n53133 = ( n17569 & n34102 ) | ( n17569 & n43813 ) | ( n34102 & n43813 ) ;
  assign n53134 = n951 & n50354 ;
  assign n53135 = ~n17850 & n30382 ;
  assign n53136 = n42102 & n53135 ;
  assign n53137 = n4331 & n53136 ;
  assign n53138 = ~n41785 & n52856 ;
  assign n53139 = n53138 ^ n27284 ^ 1'b0 ;
  assign n53141 = ~n20541 & n23725 ;
  assign n53142 = n10276 & n53141 ;
  assign n53143 = n37821 & ~n53142 ;
  assign n53140 = n7187 & ~n44465 ;
  assign n53144 = n53143 ^ n53140 ^ 1'b0 ;
  assign n53145 = ( n4155 & ~n4619 ) | ( n4155 & n42826 ) | ( ~n4619 & n42826 ) ;
  assign n53146 = n45510 & n53145 ;
  assign n53147 = n53146 ^ n22316 ^ 1'b0 ;
  assign n53148 = n33305 & ~n36761 ;
  assign n53149 = n53148 ^ n34747 ^ 1'b0 ;
  assign n53150 = n9810 ^ n5917 ^ 1'b0 ;
  assign n53151 = n34546 | n53150 ;
  assign n53152 = ( n18691 & n22602 ) | ( n18691 & ~n51628 ) | ( n22602 & ~n51628 ) ;
  assign n53153 = n49153 ^ n21600 ^ 1'b0 ;
  assign n53154 = ( n4518 & n12795 ) | ( n4518 & n43256 ) | ( n12795 & n43256 ) ;
  assign n53156 = n3044 & n7402 ;
  assign n53157 = n53156 ^ n14474 ^ 1'b0 ;
  assign n53155 = n42102 ^ n798 ^ 1'b0 ;
  assign n53158 = n53157 ^ n53155 ^ n38660 ;
  assign n53159 = ( n6706 & n7500 ) | ( n6706 & ~n26896 ) | ( n7500 & ~n26896 ) ;
  assign n53160 = ( n9343 & n17049 ) | ( n9343 & ~n53159 ) | ( n17049 & ~n53159 ) ;
  assign n53161 = n41595 ^ n30539 ^ 1'b0 ;
  assign n53162 = n26918 & ~n53161 ;
  assign n53165 = n29498 ^ n17880 ^ n5837 ;
  assign n53163 = ( n12433 & n18423 ) | ( n12433 & n51291 ) | ( n18423 & n51291 ) ;
  assign n53164 = n53163 ^ n46194 ^ n1218 ;
  assign n53166 = n53165 ^ n53164 ^ n41218 ;
  assign n53167 = n53162 & n53166 ;
  assign n53168 = n53167 ^ n44911 ^ 1'b0 ;
  assign n53169 = n5828 & ~n47442 ;
  assign n53170 = n21081 & ~n53169 ;
  assign n53171 = ~n41370 & n53170 ;
  assign n53172 = n16212 ^ n14336 ^ 1'b0 ;
  assign n53173 = n33640 ^ n14359 ^ n11554 ;
  assign n53174 = n26003 | n46254 ;
  assign n53175 = ( ~n23300 & n30899 ) | ( ~n23300 & n53174 ) | ( n30899 & n53174 ) ;
  assign n53176 = n15452 | n28796 ;
  assign n53177 = n37377 | n53176 ;
  assign n53178 = ~n1597 & n23589 ;
  assign n53182 = ( n3438 & n13145 ) | ( n3438 & n29770 ) | ( n13145 & n29770 ) ;
  assign n53183 = n8297 | n53182 ;
  assign n53184 = n49575 | n53183 ;
  assign n53179 = n18932 & ~n35167 ;
  assign n53180 = n22653 ^ n5368 ^ 1'b0 ;
  assign n53181 = n53179 & n53180 ;
  assign n53185 = n53184 ^ n53181 ^ n16421 ;
  assign n53186 = ( n53177 & n53178 ) | ( n53177 & n53185 ) | ( n53178 & n53185 ) ;
  assign n53189 = n30288 & ~n31936 ;
  assign n53187 = n16654 ^ n559 ^ 1'b0 ;
  assign n53188 = n18437 | n53187 ;
  assign n53190 = n53189 ^ n53188 ^ n38118 ;
  assign n53191 = ( n6395 & n15593 ) | ( n6395 & n23591 ) | ( n15593 & n23591 ) ;
  assign n53192 = ( n14545 & n33549 ) | ( n14545 & n53191 ) | ( n33549 & n53191 ) ;
  assign n53193 = ( n6179 & n43060 ) | ( n6179 & n53192 ) | ( n43060 & n53192 ) ;
  assign n53194 = ( n1646 & n11505 ) | ( n1646 & ~n16022 ) | ( n11505 & ~n16022 ) ;
  assign n53195 = ( n22002 & n26560 ) | ( n22002 & n53194 ) | ( n26560 & n53194 ) ;
  assign n53196 = ~n12674 & n19164 ;
  assign n53197 = n21518 & n53196 ;
  assign n53198 = ( ~n15575 & n15689 ) | ( ~n15575 & n53197 ) | ( n15689 & n53197 ) ;
  assign n53199 = ( ~n7209 & n53195 ) | ( ~n7209 & n53198 ) | ( n53195 & n53198 ) ;
  assign n53200 = n26618 & n50451 ;
  assign n53201 = n21994 & n31291 ;
  assign n53202 = n53201 ^ n25120 ^ 1'b0 ;
  assign n53203 = n3450 & ~n15691 ;
  assign n53204 = ~n53202 & n53203 ;
  assign n53205 = n13990 | n53204 ;
  assign n53206 = n21351 & n28102 ;
  assign n53207 = n53206 ^ n23080 ^ n10395 ;
  assign n53208 = n31498 ^ n8822 ^ n3422 ;
  assign n53209 = ( n1655 & n5722 ) | ( n1655 & n17313 ) | ( n5722 & n17313 ) ;
  assign n53210 = ( ~x209 & n53208 ) | ( ~x209 & n53209 ) | ( n53208 & n53209 ) ;
  assign n53211 = n4213 ^ n2058 ^ 1'b0 ;
  assign n53212 = n6608 & ~n53211 ;
  assign n53213 = n53212 ^ n30710 ^ n2139 ;
  assign n53214 = n53213 ^ n10683 ^ n1683 ;
  assign n53215 = ( n36440 & n44881 ) | ( n36440 & ~n50681 ) | ( n44881 & ~n50681 ) ;
  assign n53216 = n50074 ^ n35693 ^ 1'b0 ;
  assign n53217 = n27419 & n53216 ;
  assign n53218 = n53217 ^ n35582 ^ 1'b0 ;
  assign n53219 = n4889 & ~n32241 ;
  assign n53220 = n53219 ^ n34837 ^ n1341 ;
  assign n53221 = n53220 ^ n41493 ^ n10088 ;
  assign n53222 = n3088 & ~n4291 ;
  assign n53223 = ( n4625 & ~n8145 ) | ( n4625 & n17542 ) | ( ~n8145 & n17542 ) ;
  assign n53224 = ( n21799 & n53222 ) | ( n21799 & ~n53223 ) | ( n53222 & ~n53223 ) ;
  assign n53225 = n8503 | n15596 ;
  assign n53226 = n53225 ^ n26316 ^ 1'b0 ;
  assign n53227 = ~n9553 & n23940 ;
  assign n53228 = n53227 ^ n49424 ^ 1'b0 ;
  assign n53229 = n10989 ^ n2588 ^ x34 ;
  assign n53230 = n53229 ^ n27215 ^ n13205 ;
  assign n53231 = n12066 ^ n9787 ^ 1'b0 ;
  assign n53232 = ( n24879 & n53230 ) | ( n24879 & n53231 ) | ( n53230 & n53231 ) ;
  assign n53233 = n6695 & n53232 ;
  assign n53235 = n29209 ^ n10618 ^ 1'b0 ;
  assign n53234 = n14251 & ~n24863 ;
  assign n53236 = n53235 ^ n53234 ^ n3218 ;
  assign n53237 = n4036 & ~n53236 ;
  assign n53238 = n5599 & ~n23664 ;
  assign n53242 = n32328 ^ n19315 ^ n6850 ;
  assign n53239 = n27068 & n30734 ;
  assign n53240 = ~n18050 & n53239 ;
  assign n53241 = n53240 ^ n21995 ^ n19512 ;
  assign n53243 = n53242 ^ n53241 ^ n31389 ;
  assign n53244 = n23233 & n51986 ;
  assign n53245 = ( n49093 & n53243 ) | ( n49093 & ~n53244 ) | ( n53243 & ~n53244 ) ;
  assign n53249 = n31965 ^ n18512 ^ 1'b0 ;
  assign n53250 = n1632 & ~n53249 ;
  assign n53246 = n19491 ^ n5490 ^ n5154 ;
  assign n53247 = ( n14260 & ~n20792 ) | ( n14260 & n53246 ) | ( ~n20792 & n53246 ) ;
  assign n53248 = n37607 & n53247 ;
  assign n53251 = n53250 ^ n53248 ^ 1'b0 ;
  assign n53252 = n53251 ^ n28976 ^ 1'b0 ;
  assign n53254 = n4011 | n4208 ;
  assign n53255 = n53254 ^ n12240 ^ 1'b0 ;
  assign n53256 = n40577 ^ n34546 ^ n21096 ;
  assign n53257 = ( n18602 & ~n53255 ) | ( n18602 & n53256 ) | ( ~n53255 & n53256 ) ;
  assign n53253 = n27973 ^ n21941 ^ n1175 ;
  assign n53258 = n53257 ^ n53253 ^ n53189 ;
  assign n53259 = ~n38952 & n49919 ;
  assign n53260 = ~n22184 & n53259 ;
  assign n53261 = ( n1946 & n43028 ) | ( n1946 & ~n53260 ) | ( n43028 & ~n53260 ) ;
  assign n53262 = n8908 | n13267 ;
  assign n53263 = n53262 ^ n25662 ^ 1'b0 ;
  assign n53264 = n26728 ^ n5913 ^ n4598 ;
  assign n53265 = n27494 ^ n9518 ^ 1'b0 ;
  assign n53266 = n53265 ^ n18580 ^ n13834 ;
  assign n53269 = n22933 ^ n4372 ^ 1'b0 ;
  assign n53270 = ~n20624 & n53269 ;
  assign n53267 = ~n2905 & n12964 ;
  assign n53268 = n53267 ^ n9575 ^ 1'b0 ;
  assign n53271 = n53270 ^ n53268 ^ n6437 ;
  assign n53272 = ( n30584 & n53266 ) | ( n30584 & n53271 ) | ( n53266 & n53271 ) ;
  assign n53273 = ~n4175 & n7924 ;
  assign n53274 = n53273 ^ n52712 ^ n27140 ;
  assign n53275 = n3548 & ~n52372 ;
  assign n53276 = n49042 ^ n35938 ^ n34548 ;
  assign n53277 = n37544 ^ n14661 ^ n4717 ;
  assign n53278 = ( n12733 & ~n21238 ) | ( n12733 & n26675 ) | ( ~n21238 & n26675 ) ;
  assign n53279 = n28791 ^ n13578 ^ 1'b0 ;
  assign n53280 = n53279 ^ n19000 ^ 1'b0 ;
  assign n53281 = ~n9719 & n53280 ;
  assign n53282 = n2044 | n9345 ;
  assign n53283 = n53282 ^ n23979 ^ 1'b0 ;
  assign n53284 = n23343 ^ n17342 ^ 1'b0 ;
  assign n53285 = n13080 & ~n15335 ;
  assign n53286 = n53285 ^ n11783 ^ 1'b0 ;
  assign n53287 = ( n39282 & n43425 ) | ( n39282 & n53286 ) | ( n43425 & n53286 ) ;
  assign n53288 = ~n40715 & n53287 ;
  assign n53289 = ( ~n934 & n3268 ) | ( ~n934 & n11081 ) | ( n3268 & n11081 ) ;
  assign n53290 = ~n17838 & n25508 ;
  assign n53291 = n53290 ^ n24248 ^ 1'b0 ;
  assign n53293 = n33806 ^ n15900 ^ n422 ;
  assign n53292 = n37657 ^ n24420 ^ n2125 ;
  assign n53294 = n53293 ^ n53292 ^ 1'b0 ;
  assign n53295 = ( n13214 & n27887 ) | ( n13214 & ~n28357 ) | ( n27887 & ~n28357 ) ;
  assign n53296 = ( n21538 & ~n38432 ) | ( n21538 & n41441 ) | ( ~n38432 & n41441 ) ;
  assign n53297 = n53295 & ~n53296 ;
  assign n53298 = n17344 ^ n7905 ^ x235 ;
  assign n53299 = n53298 ^ n51042 ^ n8571 ;
  assign n53300 = n35693 ^ n1737 ^ 1'b0 ;
  assign n53301 = n23106 | n53300 ;
  assign n53304 = ( n1251 & n2701 ) | ( n1251 & n11074 ) | ( n2701 & n11074 ) ;
  assign n53302 = n5089 | n22171 ;
  assign n53303 = n53302 ^ n16519 ^ 1'b0 ;
  assign n53305 = n53304 ^ n53303 ^ n768 ;
  assign n53306 = ( n39376 & ~n46810 ) | ( n39376 & n53305 ) | ( ~n46810 & n53305 ) ;
  assign n53307 = ( ~n740 & n4889 ) | ( ~n740 & n45995 ) | ( n4889 & n45995 ) ;
  assign n53308 = n19481 ^ n1061 ^ 1'b0 ;
  assign n53309 = n18059 & n53308 ;
  assign n53310 = n53309 ^ n37732 ^ 1'b0 ;
  assign n53315 = n48160 ^ n23026 ^ n8175 ;
  assign n53311 = ( n347 & n22872 ) | ( n347 & n39659 ) | ( n22872 & n39659 ) ;
  assign n53312 = n7112 ^ n6649 ^ 1'b0 ;
  assign n53313 = n53311 & ~n53312 ;
  assign n53314 = ~n15725 & n53313 ;
  assign n53316 = n53315 ^ n53314 ^ 1'b0 ;
  assign n53317 = ~n2472 & n46259 ;
  assign n53318 = n53317 ^ n15149 ^ 1'b0 ;
  assign n53319 = n53318 ^ n52424 ^ n22140 ;
  assign n53320 = n52473 ^ n29060 ^ n19875 ;
  assign n53321 = n7850 | n40075 ;
  assign n53322 = ( n1146 & n22235 ) | ( n1146 & n53321 ) | ( n22235 & n53321 ) ;
  assign n53323 = x219 & n11815 ;
  assign n53324 = ~n22138 & n53323 ;
  assign n53325 = n3106 | n13146 ;
  assign n53326 = n53325 ^ n18905 ^ 1'b0 ;
  assign n53327 = n16128 ^ n822 ^ 1'b0 ;
  assign n53328 = n9274 & ~n53327 ;
  assign n53329 = ~n1037 & n53328 ;
  assign n53330 = n33669 & n53329 ;
  assign n53331 = ( n31751 & ~n44278 ) | ( n31751 & n53330 ) | ( ~n44278 & n53330 ) ;
  assign n53332 = n10707 ^ n5834 ^ n5171 ;
  assign n53333 = ( n10881 & ~n32772 ) | ( n10881 & n53332 ) | ( ~n32772 & n53332 ) ;
  assign n53334 = n3452 & ~n14764 ;
  assign n53335 = n1961 | n53334 ;
  assign n53336 = ( n8369 & ~n36892 ) | ( n8369 & n46123 ) | ( ~n36892 & n46123 ) ;
  assign n53337 = ( n5461 & ~n5649 ) | ( n5461 & n16203 ) | ( ~n5649 & n16203 ) ;
  assign n53338 = n53337 ^ n35512 ^ 1'b0 ;
  assign n53339 = ( n5383 & ~n30086 ) | ( n5383 & n50149 ) | ( ~n30086 & n50149 ) ;
  assign n53340 = ( n4969 & n18672 ) | ( n4969 & n30830 ) | ( n18672 & n30830 ) ;
  assign n53342 = n19394 ^ n499 ^ x180 ;
  assign n53343 = n53342 ^ n23415 ^ n4397 ;
  assign n53344 = ( n8189 & n46512 ) | ( n8189 & n53343 ) | ( n46512 & n53343 ) ;
  assign n53345 = n13432 | n53344 ;
  assign n53341 = n856 & ~n29399 ;
  assign n53346 = n53345 ^ n53341 ^ n51554 ;
  assign n53347 = n51759 ^ n13080 ^ n1653 ;
  assign n53348 = n24469 | n53347 ;
  assign n53349 = n17743 | n53348 ;
  assign n53350 = n20835 | n43066 ;
  assign n53351 = n13485 | n53350 ;
  assign n53352 = n53351 ^ n15581 ^ 1'b0 ;
  assign n53353 = ( n27965 & ~n42449 ) | ( n27965 & n53352 ) | ( ~n42449 & n53352 ) ;
  assign n53355 = ( ~n12540 & n25590 ) | ( ~n12540 & n42044 ) | ( n25590 & n42044 ) ;
  assign n53354 = n455 & n6754 ;
  assign n53356 = n53355 ^ n53354 ^ n44356 ;
  assign n53357 = ( n4749 & n6960 ) | ( n4749 & ~n53356 ) | ( n6960 & ~n53356 ) ;
  assign n53358 = n53357 ^ n42788 ^ n7655 ;
  assign n53359 = n50900 ^ n36414 ^ n18246 ;
  assign n53360 = n18156 ^ n16534 ^ 1'b0 ;
  assign n53361 = ( n993 & n31727 ) | ( n993 & n53360 ) | ( n31727 & n53360 ) ;
  assign n53362 = n53361 ^ n23601 ^ n15145 ;
  assign n53363 = ( ~n6310 & n7995 ) | ( ~n6310 & n26064 ) | ( n7995 & n26064 ) ;
  assign n53364 = n19856 ^ n14084 ^ 1'b0 ;
  assign n53365 = ( n4000 & ~n7035 ) | ( n4000 & n43150 ) | ( ~n7035 & n43150 ) ;
  assign n53366 = ( n5453 & ~n24469 ) | ( n5453 & n53365 ) | ( ~n24469 & n53365 ) ;
  assign n53367 = n9557 ^ n4503 ^ 1'b0 ;
  assign n53368 = ~n20296 & n42945 ;
  assign n53369 = ( n53366 & n53367 ) | ( n53366 & n53368 ) | ( n53367 & n53368 ) ;
  assign n53370 = n2680 & n24294 ;
  assign n53371 = ~n31725 & n53370 ;
  assign n53372 = ~n16923 & n18742 ;
  assign n53373 = n53372 ^ n43604 ^ 1'b0 ;
  assign n53374 = n15061 & ~n45166 ;
  assign n53375 = n41804 & n53374 ;
  assign n53376 = n5511 | n53375 ;
  assign n53377 = n32376 & ~n53376 ;
  assign n53380 = n29363 ^ n24711 ^ 1'b0 ;
  assign n53381 = n3574 & n53380 ;
  assign n53378 = n4176 & n39974 ;
  assign n53379 = n53378 ^ n391 ^ 1'b0 ;
  assign n53382 = n53381 ^ n53379 ^ n1822 ;
  assign n53383 = ( n29504 & n35031 ) | ( n29504 & ~n48646 ) | ( n35031 & ~n48646 ) ;
  assign n53384 = ( ~n3950 & n14830 ) | ( ~n3950 & n33479 ) | ( n14830 & n33479 ) ;
  assign n53385 = n23641 | n53384 ;
  assign n53386 = ( n14250 & n18533 ) | ( n14250 & n33917 ) | ( n18533 & n33917 ) ;
  assign n53387 = n24412 ^ n12689 ^ 1'b0 ;
  assign n53388 = n16607 & n26831 ;
  assign n53389 = n53388 ^ n33362 ^ 1'b0 ;
  assign n53390 = n53389 ^ n7062 ^ n2438 ;
  assign n53391 = n53390 ^ n11660 ^ n8419 ;
  assign n53392 = n49654 ^ n13917 ^ 1'b0 ;
  assign n53393 = n5875 & ~n53392 ;
  assign n53394 = n14880 ^ n5609 ^ 1'b0 ;
  assign n53395 = n38691 ^ n12741 ^ 1'b0 ;
  assign n53396 = ~n44840 & n49134 ;
  assign n53397 = ~n53395 & n53396 ;
  assign n53398 = ( ~n2960 & n28387 ) | ( ~n2960 & n32819 ) | ( n28387 & n32819 ) ;
  assign n53399 = ( x232 & n1351 ) | ( x232 & n23461 ) | ( n1351 & n23461 ) ;
  assign n53400 = n45323 ^ n7237 ^ 1'b0 ;
  assign n53401 = n53400 ^ n52180 ^ n9796 ;
  assign n53402 = n8196 ^ n1694 ^ n973 ;
  assign n53403 = ( ~n19064 & n20048 ) | ( ~n19064 & n34575 ) | ( n20048 & n34575 ) ;
  assign n53404 = n37321 ^ n4147 ^ n1182 ;
  assign n53405 = n53404 ^ n30668 ^ n7469 ;
  assign n53406 = ( ~n31065 & n44558 ) | ( ~n31065 & n53405 ) | ( n44558 & n53405 ) ;
  assign n53407 = ( ~n3754 & n53403 ) | ( ~n3754 & n53406 ) | ( n53403 & n53406 ) ;
  assign n53408 = n19617 ^ n17304 ^ n13084 ;
  assign n53409 = n48599 ^ n40195 ^ n23786 ;
  assign n53410 = n52366 & ~n53409 ;
  assign n53411 = ~n9105 & n27891 ;
  assign n53412 = n53411 ^ n16138 ^ 1'b0 ;
  assign n53413 = n53412 ^ n19261 ^ 1'b0 ;
  assign n53414 = n11345 & ~n53413 ;
  assign n53415 = n36878 ^ n7145 ^ 1'b0 ;
  assign n53416 = ( n12986 & n25788 ) | ( n12986 & ~n28384 ) | ( n25788 & ~n28384 ) ;
  assign n53417 = n25827 ^ n22286 ^ n21644 ;
  assign n53418 = n53417 ^ n46809 ^ n20894 ;
  assign n53419 = ( n3094 & n27036 ) | ( n3094 & ~n44027 ) | ( n27036 & ~n44027 ) ;
  assign n53420 = n45339 ^ n33523 ^ n32900 ;
  assign n53421 = n53420 ^ n17653 ^ 1'b0 ;
  assign n53422 = n4322 & n17294 ;
  assign n53423 = n40616 & ~n53422 ;
  assign n53424 = n53423 ^ n16770 ^ 1'b0 ;
  assign n53425 = ( n3536 & ~n7393 ) | ( n3536 & n53424 ) | ( ~n7393 & n53424 ) ;
  assign n53426 = ( n38592 & n51761 ) | ( n38592 & ~n53425 ) | ( n51761 & ~n53425 ) ;
  assign n53427 = n53426 ^ n50354 ^ n8259 ;
  assign n53428 = n21970 ^ n2181 ^ 1'b0 ;
  assign n53429 = n1526 & ~n53428 ;
  assign n53430 = n17563 | n41977 ;
  assign n53431 = n53430 ^ n14449 ^ 1'b0 ;
  assign n53432 = ( ~n6095 & n53429 ) | ( ~n6095 & n53431 ) | ( n53429 & n53431 ) ;
  assign n53433 = ( n21447 & ~n53427 ) | ( n21447 & n53432 ) | ( ~n53427 & n53432 ) ;
  assign n53434 = ( n16043 & ~n28637 ) | ( n16043 & n32425 ) | ( ~n28637 & n32425 ) ;
  assign n53435 = n7134 ^ n3048 ^ 1'b0 ;
  assign n53436 = n5599 | n53435 ;
  assign n53437 = ( n24741 & n36624 ) | ( n24741 & n53436 ) | ( n36624 & n53436 ) ;
  assign n53438 = n34753 & ~n49345 ;
  assign n53439 = n2975 | n4547 ;
  assign n53440 = n38555 | n53439 ;
  assign n53441 = n811 | n10970 ;
  assign n53442 = n53441 ^ n25741 ^ 1'b0 ;
  assign n53443 = ~n16967 & n33907 ;
  assign n53444 = n15330 & ~n53443 ;
  assign n53445 = ~n36454 & n53444 ;
  assign n53446 = n21333 ^ n9176 ^ 1'b0 ;
  assign n53447 = n42545 & n53446 ;
  assign n53448 = n24019 & ~n53447 ;
  assign n53449 = n5574 ^ n5243 ^ 1'b0 ;
  assign n53452 = ~n9717 & n28691 ;
  assign n53453 = n13831 & n53452 ;
  assign n53450 = n16599 & n17387 ;
  assign n53451 = n53450 ^ n3839 ^ 1'b0 ;
  assign n53454 = n53453 ^ n53451 ^ 1'b0 ;
  assign n53455 = n12074 ^ n1003 ^ 1'b0 ;
  assign n53456 = n31928 ^ n31589 ^ n11455 ;
  assign n53457 = n53456 ^ n34107 ^ n31755 ;
  assign n53458 = ( n7219 & n8834 ) | ( n7219 & ~n45004 ) | ( n8834 & ~n45004 ) ;
  assign n53459 = n35252 ^ n2036 ^ 1'b0 ;
  assign n53460 = n12690 ^ n1205 ^ 1'b0 ;
  assign n53461 = n24395 & n53460 ;
  assign n53462 = n53461 ^ n12828 ^ 1'b0 ;
  assign n53463 = ~n1809 & n53462 ;
  assign n53464 = n37716 ^ n1632 ^ 1'b0 ;
  assign n53465 = n22418 ^ n735 ^ 1'b0 ;
  assign n53466 = n33011 | n53465 ;
  assign n53467 = n35515 ^ n26963 ^ 1'b0 ;
  assign n53468 = n51706 & n53467 ;
  assign n53469 = ( n4586 & n14822 ) | ( n4586 & ~n33763 ) | ( n14822 & ~n33763 ) ;
  assign n53470 = ( ~n19235 & n33163 ) | ( ~n19235 & n53469 ) | ( n33163 & n53469 ) ;
  assign n53472 = n17882 ^ n4752 ^ 1'b0 ;
  assign n53471 = n17856 ^ n17197 ^ n9771 ;
  assign n53473 = n53472 ^ n53471 ^ n5947 ;
  assign n53474 = ( n8427 & n28218 ) | ( n8427 & ~n53473 ) | ( n28218 & ~n53473 ) ;
  assign n53475 = n42590 ^ n19568 ^ 1'b0 ;
  assign n53476 = ( ~x44 & n30573 ) | ( ~x44 & n51936 ) | ( n30573 & n51936 ) ;
  assign n53477 = ( n2782 & ~n4748 ) | ( n2782 & n8229 ) | ( ~n4748 & n8229 ) ;
  assign n53478 = n53477 ^ n42553 ^ n25827 ;
  assign n53479 = n53478 ^ n12743 ^ n2911 ;
  assign n53480 = n1242 & ~n21329 ;
  assign n53481 = n53480 ^ n33203 ^ n14571 ;
  assign n53482 = n12513 & n13719 ;
  assign n53483 = ( n1457 & n8726 ) | ( n1457 & n26285 ) | ( n8726 & n26285 ) ;
  assign n53484 = n19564 ^ n19359 ^ n18568 ;
  assign n53485 = ~n53483 & n53484 ;
  assign n53486 = n38286 ^ n17273 ^ 1'b0 ;
  assign n53487 = n27553 ^ n9625 ^ 1'b0 ;
  assign n53488 = n53486 & n53487 ;
  assign n53489 = n9323 & n53488 ;
  assign n53490 = ~n53485 & n53489 ;
  assign n53492 = n8831 | n16010 ;
  assign n53493 = n10127 | n53492 ;
  assign n53494 = n53493 ^ n26680 ^ 1'b0 ;
  assign n53491 = n17647 | n30584 ;
  assign n53495 = n53494 ^ n53491 ^ 1'b0 ;
  assign n53496 = ( n8939 & n27632 ) | ( n8939 & n33430 ) | ( n27632 & n33430 ) ;
  assign n53497 = ( x108 & n7227 ) | ( x108 & ~n10628 ) | ( n7227 & ~n10628 ) ;
  assign n53498 = n53497 ^ n17064 ^ 1'b0 ;
  assign n53499 = ~n53496 & n53498 ;
  assign n53500 = n17913 & n19107 ;
  assign n53501 = ( ~n6828 & n7448 ) | ( ~n6828 & n37921 ) | ( n7448 & n37921 ) ;
  assign n53502 = n17583 ^ n14946 ^ n6898 ;
  assign n53503 = ( ~n5468 & n21456 ) | ( ~n5468 & n53502 ) | ( n21456 & n53502 ) ;
  assign n53504 = n44899 ^ n12219 ^ n11382 ;
  assign n53505 = n21806 ^ n15290 ^ n3000 ;
  assign n53506 = ( x121 & n32753 ) | ( x121 & n53505 ) | ( n32753 & n53505 ) ;
  assign n53507 = ( n29982 & ~n45284 ) | ( n29982 & n47012 ) | ( ~n45284 & n47012 ) ;
  assign n53508 = ( n1118 & ~n35866 ) | ( n1118 & n42649 ) | ( ~n35866 & n42649 ) ;
  assign n53509 = ~n1631 & n25465 ;
  assign n53510 = n53509 ^ n4736 ^ 1'b0 ;
  assign n53511 = n2042 & ~n4240 ;
  assign n53512 = n5339 & n53511 ;
  assign n53513 = ( n4426 & ~n30763 ) | ( n4426 & n53512 ) | ( ~n30763 & n53512 ) ;
  assign n53514 = n53513 ^ n5662 ^ 1'b0 ;
  assign n53515 = n37113 | n53514 ;
  assign n53516 = ~n298 & n3089 ;
  assign n53517 = ( n4710 & n5765 ) | ( n4710 & n53516 ) | ( n5765 & n53516 ) ;
  assign n53518 = ( n17649 & n38871 ) | ( n17649 & n53517 ) | ( n38871 & n53517 ) ;
  assign n53519 = ( ~n13988 & n21888 ) | ( ~n13988 & n28261 ) | ( n21888 & n28261 ) ;
  assign n53520 = ( n32883 & n43567 ) | ( n32883 & n53519 ) | ( n43567 & n53519 ) ;
  assign n53521 = ( n3584 & n15995 ) | ( n3584 & n50862 ) | ( n15995 & n50862 ) ;
  assign n53522 = n52081 ^ n33134 ^ 1'b0 ;
  assign n53523 = n11995 & ~n38392 ;
  assign n53524 = n53523 ^ n32436 ^ n31442 ;
  assign n53525 = n43035 ^ n13026 ^ n1504 ;
  assign n53526 = n14678 & ~n22592 ;
  assign n53527 = n53526 ^ n47079 ^ n34283 ;
  assign n53528 = n53527 ^ n35556 ^ n13427 ;
  assign n53529 = ( ~n10634 & n14927 ) | ( ~n10634 & n53528 ) | ( n14927 & n53528 ) ;
  assign n53533 = n12905 ^ n8172 ^ n4867 ;
  assign n53530 = n16721 & n27108 ;
  assign n53531 = n53530 ^ n31839 ^ 1'b0 ;
  assign n53532 = n39850 & n53531 ;
  assign n53534 = n53533 ^ n53532 ^ 1'b0 ;
  assign n53535 = n20666 ^ n11004 ^ x221 ;
  assign n53536 = n21535 ^ n9747 ^ n8644 ;
  assign n53537 = n53536 ^ n7461 ^ n6834 ;
  assign n53538 = n53537 ^ n46116 ^ 1'b0 ;
  assign n53539 = ~n53535 & n53538 ;
  assign n53540 = n27688 ^ n24818 ^ n10791 ;
  assign n53541 = n28953 ^ n27357 ^ 1'b0 ;
  assign n53542 = ~n53540 & n53541 ;
  assign n53543 = n43905 ^ n2615 ^ 1'b0 ;
  assign n53545 = ( n6911 & n14592 ) | ( n6911 & ~n52065 ) | ( n14592 & ~n52065 ) ;
  assign n53544 = ( n28331 & ~n29864 ) | ( n28331 & n48932 ) | ( ~n29864 & n48932 ) ;
  assign n53546 = n53545 ^ n53544 ^ n3872 ;
  assign n53547 = n1046 | n16267 ;
  assign n53548 = n53547 ^ n9228 ^ 1'b0 ;
  assign n53549 = n35280 ^ n18882 ^ n15896 ;
  assign n53552 = ( ~n11300 & n13270 ) | ( ~n11300 & n25431 ) | ( n13270 & n25431 ) ;
  assign n53550 = ( ~n947 & n5247 ) | ( ~n947 & n24647 ) | ( n5247 & n24647 ) ;
  assign n53551 = ( ~n35970 & n37495 ) | ( ~n35970 & n53550 ) | ( n37495 & n53550 ) ;
  assign n53553 = n53552 ^ n53551 ^ n38827 ;
  assign n53554 = ( n35309 & n53549 ) | ( n35309 & ~n53553 ) | ( n53549 & ~n53553 ) ;
  assign n53555 = n32755 ^ n5331 ^ n3049 ;
  assign n53556 = n11907 ^ n11536 ^ 1'b0 ;
  assign n53557 = n6770 & ~n20579 ;
  assign n53558 = n1315 & n53557 ;
  assign n53559 = n7149 & ~n31881 ;
  assign n53560 = ~n22461 & n53559 ;
  assign n53561 = ~n15368 & n43369 ;
  assign n53562 = n53561 ^ n29424 ^ 1'b0 ;
  assign n53563 = ( n8889 & n20609 ) | ( n8889 & n44093 ) | ( n20609 & n44093 ) ;
  assign n53564 = n53563 ^ n20855 ^ n5613 ;
  assign n53565 = n8115 | n31549 ;
  assign n53567 = x225 & n30317 ;
  assign n53566 = n43738 ^ n26693 ^ n2749 ;
  assign n53568 = n53567 ^ n53566 ^ n25846 ;
  assign n53569 = ( ~n4247 & n7421 ) | ( ~n4247 & n37584 ) | ( n7421 & n37584 ) ;
  assign n53570 = ( n24329 & ~n34167 ) | ( n24329 & n53569 ) | ( ~n34167 & n53569 ) ;
  assign n53571 = n53570 ^ n5318 ^ 1'b0 ;
  assign n53572 = ( ~n5111 & n13603 ) | ( ~n5111 & n19955 ) | ( n13603 & n19955 ) ;
  assign n53574 = ( n4074 & n15274 ) | ( n4074 & ~n17166 ) | ( n15274 & ~n17166 ) ;
  assign n53575 = n53574 ^ n21777 ^ 1'b0 ;
  assign n53576 = n11260 & n53575 ;
  assign n53573 = ~n38449 & n39758 ;
  assign n53577 = n53576 ^ n53573 ^ n3536 ;
  assign n53578 = n26087 ^ n25493 ^ n2663 ;
  assign n53579 = n34983 | n38239 ;
  assign n53580 = n5875 & n46572 ;
  assign n53581 = n22621 & n53580 ;
  assign n53582 = n7022 & ~n46140 ;
  assign n53583 = n28196 & ~n53582 ;
  assign n53584 = n38560 | n51828 ;
  assign n53585 = n34986 ^ n33252 ^ n6419 ;
  assign n53586 = n17595 & ~n30757 ;
  assign n53587 = n29645 & n48745 ;
  assign n53588 = ( n28249 & n39133 ) | ( n28249 & n51393 ) | ( n39133 & n51393 ) ;
  assign n53589 = n8941 ^ n8482 ^ n8472 ;
  assign n53590 = ( n5309 & ~n8970 ) | ( n5309 & n53589 ) | ( ~n8970 & n53589 ) ;
  assign n53591 = n53590 ^ n37904 ^ n19576 ;
  assign n53592 = n32159 ^ n14514 ^ 1'b0 ;
  assign n53593 = n18240 ^ n3635 ^ n1490 ;
  assign n53594 = ( n34097 & n53592 ) | ( n34097 & n53593 ) | ( n53592 & n53593 ) ;
  assign n53595 = n45116 ^ n5343 ^ 1'b0 ;
  assign n53596 = n36956 | n53595 ;
  assign n53597 = ~n1444 & n2111 ;
  assign n53598 = n53597 ^ n1564 ^ 1'b0 ;
  assign n53600 = n48371 ^ n25482 ^ n18018 ;
  assign n53599 = n10655 & ~n12150 ;
  assign n53601 = n53600 ^ n53599 ^ 1'b0 ;
  assign n53602 = ( n19479 & n37231 ) | ( n19479 & ~n43612 ) | ( n37231 & ~n43612 ) ;
  assign n53603 = n13193 & n39222 ;
  assign n53604 = n44846 ^ n38380 ^ n27375 ;
  assign n53605 = n36912 ^ n21547 ^ 1'b0 ;
  assign n53606 = n53604 & ~n53605 ;
  assign n53607 = n53606 ^ n33362 ^ n811 ;
  assign n53608 = n53607 ^ n36133 ^ n5250 ;
  assign n53609 = n11345 & n37201 ;
  assign n53610 = n16869 & ~n28008 ;
  assign n53611 = ~n21634 & n53610 ;
  assign n53612 = ( n8277 & n15855 ) | ( n8277 & ~n27732 ) | ( n15855 & ~n27732 ) ;
  assign n53613 = ( ~n28289 & n53611 ) | ( ~n28289 & n53612 ) | ( n53611 & n53612 ) ;
  assign n53614 = ( n18150 & n53609 ) | ( n18150 & n53613 ) | ( n53609 & n53613 ) ;
  assign n53615 = ( n35199 & n36305 ) | ( n35199 & n50034 ) | ( n36305 & n50034 ) ;
  assign n53616 = n4273 ^ n2681 ^ n1336 ;
  assign n53617 = n23259 ^ n10800 ^ 1'b0 ;
  assign n53618 = n26097 & n53617 ;
  assign n53619 = n53618 ^ n19228 ^ n17177 ;
  assign n53620 = n53619 ^ n14765 ^ n2086 ;
  assign n53621 = n53620 ^ n52234 ^ n34293 ;
  assign n53622 = n18869 ^ n10235 ^ 1'b0 ;
  assign n53623 = x240 & ~n53622 ;
  assign n53624 = n53623 ^ n25249 ^ 1'b0 ;
  assign n53625 = ~n1485 & n22342 ;
  assign n53626 = n11976 & ~n21721 ;
  assign n53627 = ~n14861 & n53626 ;
  assign n53628 = ( ~n5980 & n8806 ) | ( ~n5980 & n52579 ) | ( n8806 & n52579 ) ;
  assign n53629 = ( x162 & n3809 ) | ( x162 & n20679 ) | ( n3809 & n20679 ) ;
  assign n53630 = n53629 ^ n40589 ^ n25405 ;
  assign n53631 = n7304 | n33387 ;
  assign n53632 = n11186 | n53631 ;
  assign n53633 = n53632 ^ n23744 ^ n5494 ;
  assign n53637 = ( ~n8922 & n24562 ) | ( ~n8922 & n47272 ) | ( n24562 & n47272 ) ;
  assign n53634 = n11974 | n32677 ;
  assign n53635 = n5505 | n53634 ;
  assign n53636 = n53635 ^ n43261 ^ n20885 ;
  assign n53638 = n53637 ^ n53636 ^ n30880 ;
  assign n53639 = ( n3748 & n5083 ) | ( n3748 & n6271 ) | ( n5083 & n6271 ) ;
  assign n53640 = ( n34621 & n44616 ) | ( n34621 & ~n53639 ) | ( n44616 & ~n53639 ) ;
  assign n53641 = n40291 ^ n35389 ^ n7508 ;
  assign n53642 = n53641 ^ n42124 ^ 1'b0 ;
  assign n53643 = n12969 & ~n14190 ;
  assign n53644 = n53643 ^ n9869 ^ 1'b0 ;
  assign n53645 = n51950 & n53644 ;
  assign n53646 = n53645 ^ n16283 ^ 1'b0 ;
  assign n53647 = ~n15435 & n23120 ;
  assign n53648 = n15650 & n53647 ;
  assign n53649 = ~n19658 & n43536 ;
  assign n53650 = n53648 & n53649 ;
  assign n53651 = n27088 | n27261 ;
  assign n53652 = n53651 ^ n13196 ^ 1'b0 ;
  assign n53653 = n46270 ^ n1256 ^ 1'b0 ;
  assign n53654 = ~n52977 & n53653 ;
  assign n53655 = n25099 ^ n14866 ^ n9815 ;
  assign n53656 = ( n19625 & n26132 ) | ( n19625 & n43852 ) | ( n26132 & n43852 ) ;
  assign n53657 = n53656 ^ n22898 ^ 1'b0 ;
  assign n53658 = n29959 ^ n20337 ^ x45 ;
  assign n53659 = n23664 | n33723 ;
  assign n53660 = ~n2638 & n19685 ;
  assign n53661 = n6799 & ~n49265 ;
  assign n53662 = ( n29348 & ~n53660 ) | ( n29348 & n53661 ) | ( ~n53660 & n53661 ) ;
  assign n53663 = n44072 ^ n1755 ^ 1'b0 ;
  assign n53664 = ~n975 & n12360 ;
  assign n53665 = ~n1442 & n53664 ;
  assign n53666 = n53665 ^ n38982 ^ n2485 ;
  assign n53667 = n32045 & n38624 ;
  assign n53668 = n53667 ^ n13096 ^ 1'b0 ;
  assign n53669 = ~n6701 & n13838 ;
  assign n53670 = n53669 ^ n2692 ^ 1'b0 ;
  assign n53671 = n50586 ^ n40565 ^ n9320 ;
  assign n53672 = n7160 & ~n53671 ;
  assign n53673 = n53672 ^ n8172 ^ 1'b0 ;
  assign n53674 = n23424 | n45749 ;
  assign n53675 = n16400 | n50737 ;
  assign n53676 = ~n18865 & n31410 ;
  assign n53677 = ~n10353 & n33303 ;
  assign n53678 = n53677 ^ n46352 ^ 1'b0 ;
  assign n53679 = ( n11658 & n27366 ) | ( n11658 & ~n53678 ) | ( n27366 & ~n53678 ) ;
  assign n53680 = n22396 ^ n16443 ^ n5399 ;
  assign n53685 = ( ~n2097 & n17091 ) | ( ~n2097 & n19655 ) | ( n17091 & n19655 ) ;
  assign n53682 = n1464 | n3771 ;
  assign n53683 = n53682 ^ n28600 ^ 1'b0 ;
  assign n53681 = ( n9390 & ~n21595 ) | ( n9390 & n36883 ) | ( ~n21595 & n36883 ) ;
  assign n53684 = n53683 ^ n53681 ^ n28028 ;
  assign n53686 = n53685 ^ n53684 ^ n18735 ;
  assign n53687 = ( n12344 & n16893 ) | ( n12344 & ~n27644 ) | ( n16893 & ~n27644 ) ;
  assign n53688 = ( x249 & n10409 ) | ( x249 & ~n53687 ) | ( n10409 & ~n53687 ) ;
  assign n53689 = ( n12199 & n16338 ) | ( n12199 & ~n53688 ) | ( n16338 & ~n53688 ) ;
  assign n53690 = ~n29668 & n33854 ;
  assign n53691 = n53690 ^ n49408 ^ n39905 ;
  assign n53692 = n14021 & ~n23164 ;
  assign n53693 = n53692 ^ n39853 ^ 1'b0 ;
  assign n53694 = ( ~n2960 & n11855 ) | ( ~n2960 & n13460 ) | ( n11855 & n13460 ) ;
  assign n53695 = n24104 | n53694 ;
  assign n53696 = n53695 ^ n10550 ^ 1'b0 ;
  assign n53697 = ( n552 & ~n7709 ) | ( n552 & n35120 ) | ( ~n7709 & n35120 ) ;
  assign n53698 = n11868 & n16025 ;
  assign n53699 = ~n53697 & n53698 ;
  assign n53700 = n35643 ^ n13114 ^ 1'b0 ;
  assign n53701 = ~x4 & n53700 ;
  assign n53702 = ( n13033 & n18424 ) | ( n13033 & n53701 ) | ( n18424 & n53701 ) ;
  assign n53703 = n6890 | n14762 ;
  assign n53704 = ~n2273 & n53703 ;
  assign n53705 = n49333 ^ n39462 ^ n27555 ;
  assign n53706 = n47291 ^ n46239 ^ n3866 ;
  assign n53707 = ( n36525 & n38198 ) | ( n36525 & ~n50886 ) | ( n38198 & ~n50886 ) ;
  assign n53708 = n36363 ^ n3517 ^ n2426 ;
  assign n53709 = n3747 | n17457 ;
  assign n53710 = n33487 ^ n15125 ^ 1'b0 ;
  assign n53711 = n13586 & ~n53710 ;
  assign n53712 = ~n26128 & n26971 ;
  assign n53713 = ~n19532 & n53712 ;
  assign n53714 = ~n8593 & n51070 ;
  assign n53715 = n53714 ^ n17678 ^ 1'b0 ;
  assign n53716 = n10448 ^ n5795 ^ n2223 ;
  assign n53717 = ~n24545 & n53716 ;
  assign n53718 = n43041 & n53717 ;
  assign n53719 = n37276 ^ n28600 ^ 1'b0 ;
  assign n53720 = n33766 ^ n13779 ^ n9376 ;
  assign n53721 = n45892 ^ n25219 ^ n21840 ;
  assign n53722 = n35456 ^ n8798 ^ 1'b0 ;
  assign n53723 = ~n40631 & n53722 ;
  assign n53724 = ~n24428 & n53723 ;
  assign n53725 = n39941 ^ n19359 ^ n16004 ;
  assign n53729 = n22363 ^ n7613 ^ 1'b0 ;
  assign n53728 = n6520 & n10315 ;
  assign n53726 = n896 & ~n29310 ;
  assign n53727 = n53726 ^ n23488 ^ 1'b0 ;
  assign n53730 = n53729 ^ n53728 ^ n53727 ;
  assign n53731 = n20946 | n32661 ;
  assign n53732 = n53731 ^ n32930 ^ 1'b0 ;
  assign n53733 = n33018 ^ n3342 ^ n1719 ;
  assign n53734 = n742 | n16691 ;
  assign n53735 = n1708 | n53734 ;
  assign n53736 = n53735 ^ n19176 ^ n8269 ;
  assign n53737 = n53736 ^ n53043 ^ n37518 ;
  assign n53738 = ( n19065 & n53733 ) | ( n19065 & ~n53737 ) | ( n53733 & ~n53737 ) ;
  assign n53739 = ( n2625 & n18538 ) | ( n2625 & n40500 ) | ( n18538 & n40500 ) ;
  assign n53740 = n53739 ^ n21509 ^ 1'b0 ;
  assign n53741 = n53738 | n53740 ;
  assign n53742 = n2310 & ~n27023 ;
  assign n53743 = n40529 ^ n10492 ^ 1'b0 ;
  assign n53744 = n27726 | n29501 ;
  assign n53745 = n53744 ^ n595 ^ 1'b0 ;
  assign n53746 = ( n39060 & n41707 ) | ( n39060 & n53745 ) | ( n41707 & n53745 ) ;
  assign n53747 = n22617 ^ n9408 ^ n1905 ;
  assign n53748 = ( n5612 & n23854 ) | ( n5612 & ~n27423 ) | ( n23854 & ~n27423 ) ;
  assign n53749 = n37303 & n50425 ;
  assign n53756 = n46505 ^ n24976 ^ n6613 ;
  assign n53752 = n12738 & ~n14649 ;
  assign n53753 = n53752 ^ n13703 ^ 1'b0 ;
  assign n53754 = n2999 & ~n53753 ;
  assign n53755 = n53754 ^ n47042 ^ 1'b0 ;
  assign n53750 = n40594 ^ n22975 ^ 1'b0 ;
  assign n53751 = n53750 ^ n33905 ^ n6789 ;
  assign n53757 = n53756 ^ n53755 ^ n53751 ;
  assign n53758 = ( n9795 & ~n10950 ) | ( n9795 & n32809 ) | ( ~n10950 & n32809 ) ;
  assign n53759 = n16764 | n53758 ;
  assign n53760 = n16460 & n53759 ;
  assign n53761 = n53760 ^ n21780 ^ 1'b0 ;
  assign n53762 = n1330 ^ n1233 ^ 1'b0 ;
  assign n53763 = ( ~n32940 & n39137 ) | ( ~n32940 & n49517 ) | ( n39137 & n49517 ) ;
  assign n53764 = n53763 ^ n50190 ^ x190 ;
  assign n53765 = ( n368 & ~n39671 ) | ( n368 & n53764 ) | ( ~n39671 & n53764 ) ;
  assign n53766 = n35981 ^ n7932 ^ n7417 ;
  assign n53767 = n4946 | n7907 ;
  assign n53768 = n33901 | n53767 ;
  assign n53769 = ~n33801 & n41836 ;
  assign n53770 = ( ~n20570 & n53768 ) | ( ~n20570 & n53769 ) | ( n53768 & n53769 ) ;
  assign n53771 = n26933 ^ n23183 ^ 1'b0 ;
  assign n53772 = n47773 ^ n43748 ^ n3156 ;
  assign n53773 = n1226 & ~n20215 ;
  assign n53774 = n15628 ^ n9364 ^ n3487 ;
  assign n53775 = n53774 ^ n11947 ^ n6118 ;
  assign n53776 = ~n9458 & n51094 ;
  assign n53777 = ~n358 & n53776 ;
  assign n53778 = n19986 ^ n11998 ^ 1'b0 ;
  assign n53779 = ~n43957 & n53778 ;
  assign n53780 = n13594 ^ n9324 ^ 1'b0 ;
  assign n53783 = n4651 ^ n2887 ^ n2152 ;
  assign n53781 = n4594 & n19272 ;
  assign n53782 = n53781 ^ n11779 ^ 1'b0 ;
  assign n53784 = n53783 ^ n53782 ^ n46326 ;
  assign n53785 = n53784 ^ n31048 ^ n4072 ;
  assign n53786 = n8870 ^ n5593 ^ 1'b0 ;
  assign n53787 = n19248 | n53786 ;
  assign n53788 = ~n1240 & n20728 ;
  assign n53789 = ( ~n8216 & n53787 ) | ( ~n8216 & n53788 ) | ( n53787 & n53788 ) ;
  assign n53790 = ~n20178 & n22095 ;
  assign n53791 = ( n26488 & n31591 ) | ( n26488 & ~n53790 ) | ( n31591 & ~n53790 ) ;
  assign n53792 = ( n18115 & n32851 ) | ( n18115 & ~n53791 ) | ( n32851 & ~n53791 ) ;
  assign n53793 = n31711 ^ n16892 ^ n13493 ;
  assign n53794 = n33646 ^ n13563 ^ n11260 ;
  assign n53795 = ( ~n30334 & n49684 ) | ( ~n30334 & n53794 ) | ( n49684 & n53794 ) ;
  assign n53796 = n51926 ^ n34901 ^ 1'b0 ;
  assign n53797 = x77 & ~n53796 ;
  assign n53798 = n53797 ^ n18300 ^ n7398 ;
  assign n53799 = n15038 & ~n36860 ;
  assign n53800 = n25328 | n40255 ;
  assign n53801 = n53800 ^ n9897 ^ 1'b0 ;
  assign n53802 = n20889 & n32169 ;
  assign n53803 = n53802 ^ n9788 ^ 1'b0 ;
  assign n53804 = ( n3061 & n12961 ) | ( n3061 & n13457 ) | ( n12961 & n13457 ) ;
  assign n53805 = ( n3837 & n15672 ) | ( n3837 & ~n53804 ) | ( n15672 & ~n53804 ) ;
  assign n53806 = ( n14712 & ~n41248 ) | ( n14712 & n53805 ) | ( ~n41248 & n53805 ) ;
  assign n53807 = ~n19361 & n53806 ;
  assign n53808 = n52793 ^ n33367 ^ n32405 ;
  assign n53809 = n2429 & ~n7349 ;
  assign n53810 = n53809 ^ n3188 ^ 1'b0 ;
  assign n53811 = n4827 | n16175 ;
  assign n53812 = n53810 & ~n53811 ;
  assign n53813 = n53812 ^ n15321 ^ n9825 ;
  assign n53814 = ( n6167 & ~n18246 ) | ( n6167 & n47229 ) | ( ~n18246 & n47229 ) ;
  assign n53815 = ( n23333 & n28341 ) | ( n23333 & ~n53814 ) | ( n28341 & ~n53814 ) ;
  assign n53816 = n48306 ^ n27042 ^ n19144 ;
  assign n53817 = n53816 ^ n23803 ^ n18181 ;
  assign n53818 = ~n28188 & n38358 ;
  assign n53819 = n53818 ^ n25413 ^ 1'b0 ;
  assign n53820 = n4973 & n37616 ;
  assign n53821 = n53820 ^ n29112 ^ 1'b0 ;
  assign n53822 = ( ~n16991 & n53819 ) | ( ~n16991 & n53821 ) | ( n53819 & n53821 ) ;
  assign n53823 = n45961 ^ n12911 ^ n9807 ;
  assign n53824 = n3824 & n53823 ;
  assign n53826 = n41324 ^ n17754 ^ n3292 ;
  assign n53827 = n53826 ^ n21479 ^ 1'b0 ;
  assign n53828 = n7375 & n53827 ;
  assign n53829 = ( n7839 & n44275 ) | ( n7839 & ~n53828 ) | ( n44275 & ~n53828 ) ;
  assign n53830 = n45634 ^ n11087 ^ 1'b0 ;
  assign n53831 = n42461 | n53830 ;
  assign n53832 = n8830 | n53831 ;
  assign n53833 = n53829 | n53832 ;
  assign n53825 = n19626 & n40234 ;
  assign n53834 = n53833 ^ n53825 ^ 1'b0 ;
  assign n53835 = n47533 | n47905 ;
  assign n53836 = n17118 ^ n2833 ^ 1'b0 ;
  assign n53837 = n53835 & ~n53836 ;
  assign n53838 = n4024 & n50234 ;
  assign n53839 = n10443 & n53838 ;
  assign n53842 = n21062 ^ n8245 ^ 1'b0 ;
  assign n53843 = n26000 & ~n53842 ;
  assign n53840 = n10786 ^ n3642 ^ n3577 ;
  assign n53841 = ( n4705 & n23702 ) | ( n4705 & n53840 ) | ( n23702 & n53840 ) ;
  assign n53844 = n53843 ^ n53841 ^ n33880 ;
  assign n53846 = n52523 ^ n37514 ^ n31224 ;
  assign n53845 = n14037 ^ n13205 ^ n5533 ;
  assign n53847 = n53846 ^ n53845 ^ n44369 ;
  assign n53848 = ( n11756 & ~n29676 ) | ( n11756 & n44949 ) | ( ~n29676 & n44949 ) ;
  assign n53849 = n23417 ^ n5248 ^ 1'b0 ;
  assign n53850 = n5468 & ~n53849 ;
  assign n53851 = ( n532 & n49779 ) | ( n532 & ~n53850 ) | ( n49779 & ~n53850 ) ;
  assign n53852 = ( n21328 & n28777 ) | ( n21328 & n53851 ) | ( n28777 & n53851 ) ;
  assign n53853 = n16181 & n33360 ;
  assign n53854 = n33033 & n53853 ;
  assign n53855 = n37200 ^ n25787 ^ n15422 ;
  assign n53856 = ( n32156 & n36369 ) | ( n32156 & n53855 ) | ( n36369 & n53855 ) ;
  assign n53857 = n51509 ^ n43365 ^ n5533 ;
  assign n53858 = ~n8454 & n10699 ;
  assign n53859 = ( n5617 & n6693 ) | ( n5617 & n27559 ) | ( n6693 & n27559 ) ;
  assign n53860 = n21860 & n24474 ;
  assign n53861 = n53859 & n53860 ;
  assign n53862 = ( n15326 & n15415 ) | ( n15326 & ~n16687 ) | ( n15415 & ~n16687 ) ;
  assign n53863 = n53862 ^ n35598 ^ n23722 ;
  assign n53864 = n53863 ^ n12085 ^ n5427 ;
  assign n53866 = n5279 & n25261 ;
  assign n53865 = n28376 ^ n23595 ^ n11428 ;
  assign n53867 = n53866 ^ n53865 ^ n1714 ;
  assign n53868 = ( ~n1705 & n10187 ) | ( ~n1705 & n36881 ) | ( n10187 & n36881 ) ;
  assign n53876 = n2228 & ~n25623 ;
  assign n53877 = n42460 & n53876 ;
  assign n53870 = ( n5159 & n6015 ) | ( n5159 & ~n8067 ) | ( n6015 & ~n8067 ) ;
  assign n53871 = n53870 ^ n48059 ^ n19257 ;
  assign n53869 = ( n17345 & n18418 ) | ( n17345 & ~n33003 ) | ( n18418 & ~n33003 ) ;
  assign n53872 = n53871 ^ n53869 ^ n5710 ;
  assign n53873 = ( n15314 & n35755 ) | ( n15314 & n53872 ) | ( n35755 & n53872 ) ;
  assign n53874 = n11586 | n53873 ;
  assign n53875 = n20026 & ~n53874 ;
  assign n53878 = n53877 ^ n53875 ^ n34222 ;
  assign n53879 = n53868 & ~n53878 ;
  assign n53880 = n40784 ^ n16063 ^ 1'b0 ;
  assign n53881 = ( ~n20486 & n20904 ) | ( ~n20486 & n53880 ) | ( n20904 & n53880 ) ;
  assign n53884 = n41510 ^ n9406 ^ 1'b0 ;
  assign n53882 = n2474 & n11372 ;
  assign n53883 = n53882 ^ n24380 ^ n14944 ;
  assign n53885 = n53884 ^ n53883 ^ n32564 ;
  assign n53886 = ( n5588 & n12034 ) | ( n5588 & ~n53469 ) | ( n12034 & ~n53469 ) ;
  assign n53887 = ( ~n3938 & n14621 ) | ( ~n3938 & n15455 ) | ( n14621 & n15455 ) ;
  assign n53888 = ( n17226 & ~n23431 ) | ( n17226 & n47045 ) | ( ~n23431 & n47045 ) ;
  assign n53889 = n6689 & n53888 ;
  assign n53890 = ~n28297 & n53889 ;
  assign n53891 = n3540 | n33146 ;
  assign n53892 = n39812 & ~n53891 ;
  assign n53893 = n17946 ^ n4610 ^ 1'b0 ;
  assign n53894 = n22960 ^ n480 ^ 1'b0 ;
  assign n53895 = n19991 & ~n53894 ;
  assign n53896 = n53895 ^ n39975 ^ 1'b0 ;
  assign n53897 = n53896 ^ n21562 ^ n19826 ;
  assign n53900 = ~n929 & n18709 ;
  assign n53901 = ~n42417 & n53900 ;
  assign n53898 = ( n4589 & n9346 ) | ( n4589 & ~n16950 ) | ( n9346 & ~n16950 ) ;
  assign n53899 = n53898 ^ n37123 ^ n33461 ;
  assign n53902 = n53901 ^ n53899 ^ n20097 ;
  assign n53903 = ( n7939 & n8390 ) | ( n7939 & ~n36215 ) | ( n8390 & ~n36215 ) ;
  assign n53904 = n53903 ^ n9920 ^ 1'b0 ;
  assign n53905 = n51483 ^ n20435 ^ n1237 ;
  assign n53907 = n19252 ^ n15876 ^ 1'b0 ;
  assign n53908 = n46919 | n53907 ;
  assign n53906 = ( n6927 & ~n43496 ) | ( n6927 & n49140 ) | ( ~n43496 & n49140 ) ;
  assign n53909 = n53908 ^ n53906 ^ 1'b0 ;
  assign n53912 = ( n5922 & ~n15182 ) | ( n5922 & n16063 ) | ( ~n15182 & n16063 ) ;
  assign n53910 = n3856 & n11472 ;
  assign n53911 = n53910 ^ n3165 ^ n1344 ;
  assign n53913 = n53912 ^ n53911 ^ n32341 ;
  assign n53914 = n8395 & n47157 ;
  assign n53915 = ~n18044 & n53914 ;
  assign n53916 = n53304 & ~n53915 ;
  assign n53917 = n40575 ^ n20850 ^ 1'b0 ;
  assign n53918 = n32098 & ~n53917 ;
  assign n53919 = n356 & n16764 ;
  assign n53920 = n53919 ^ n3555 ^ 1'b0 ;
  assign n53921 = n2369 | n50332 ;
  assign n53922 = n23856 & ~n30792 ;
  assign n53923 = n25049 & n53922 ;
  assign n53924 = n53923 ^ n32747 ^ 1'b0 ;
  assign n53925 = n26861 & ~n53924 ;
  assign n53926 = n28987 ^ n25671 ^ n2565 ;
  assign n53927 = ( n33106 & n53925 ) | ( n33106 & ~n53926 ) | ( n53925 & ~n53926 ) ;
  assign n53928 = ( n5834 & n50633 ) | ( n5834 & ~n53927 ) | ( n50633 & ~n53927 ) ;
  assign n53929 = ( ~n45134 & n46094 ) | ( ~n45134 & n53928 ) | ( n46094 & n53928 ) ;
  assign n53930 = n24490 ^ n13015 ^ n9476 ;
  assign n53931 = ( n5761 & n18521 ) | ( n5761 & n24347 ) | ( n18521 & n24347 ) ;
  assign n53932 = n7930 ^ n3811 ^ 1'b0 ;
  assign n53933 = n53932 ^ n52289 ^ 1'b0 ;
  assign n53934 = n24870 & n35363 ;
  assign n53935 = ~n33877 & n53934 ;
  assign n53936 = ~n8627 & n16841 ;
  assign n53937 = n53935 & n53936 ;
  assign n53938 = n33276 ^ n5079 ^ 1'b0 ;
  assign n53939 = n15486 ^ n12456 ^ 1'b0 ;
  assign n53944 = n34095 ^ n18839 ^ n11651 ;
  assign n53942 = n25615 | n40849 ;
  assign n53943 = n53942 ^ n21391 ^ 1'b0 ;
  assign n53940 = n46874 ^ n32127 ^ 1'b0 ;
  assign n53941 = n53940 ^ n32362 ^ n11334 ;
  assign n53945 = n53944 ^ n53943 ^ n53941 ;
  assign n53946 = ( n7443 & n22113 ) | ( n7443 & ~n36786 ) | ( n22113 & ~n36786 ) ;
  assign n53947 = ( ~n12199 & n36912 ) | ( ~n12199 & n37220 ) | ( n36912 & n37220 ) ;
  assign n53948 = ( ~n1368 & n10075 ) | ( ~n1368 & n41981 ) | ( n10075 & n41981 ) ;
  assign n53949 = n34048 ^ n33763 ^ n11826 ;
  assign n53950 = ( n299 & n53948 ) | ( n299 & ~n53949 ) | ( n53948 & ~n53949 ) ;
  assign n53951 = ~n32953 & n51106 ;
  assign n53952 = ~n5796 & n53951 ;
  assign n53953 = n53952 ^ n9634 ^ 1'b0 ;
  assign n53954 = n39853 ^ n30033 ^ 1'b0 ;
  assign n53955 = n53954 ^ n45646 ^ 1'b0 ;
  assign n53956 = ( n13196 & ~n20590 ) | ( n13196 & n28141 ) | ( ~n20590 & n28141 ) ;
  assign n53957 = n53956 ^ n30626 ^ n8791 ;
  assign n53958 = n23156 ^ n2342 ^ 1'b0 ;
  assign n53959 = ~n47310 & n53958 ;
  assign n53960 = ( n30385 & n33622 ) | ( n30385 & n53959 ) | ( n33622 & n53959 ) ;
  assign n53961 = n43458 ^ n21880 ^ n21867 ;
  assign n53962 = n53961 ^ n34700 ^ n24297 ;
  assign n53963 = n10725 | n35539 ;
  assign n53964 = n15345 | n30417 ;
  assign n53965 = ~n34744 & n53964 ;
  assign n53966 = n53965 ^ n17388 ^ 1'b0 ;
  assign n53967 = ( ~n16448 & n36321 ) | ( ~n16448 & n53966 ) | ( n36321 & n53966 ) ;
  assign n53968 = n13551 & n13846 ;
  assign n53969 = n29142 & n53968 ;
  assign n53970 = n53969 ^ n23889 ^ n2771 ;
  assign n53971 = ( n1653 & ~n6576 ) | ( n1653 & n14678 ) | ( ~n6576 & n14678 ) ;
  assign n53972 = ( ~n9271 & n14629 ) | ( ~n9271 & n53971 ) | ( n14629 & n53971 ) ;
  assign n53973 = ~n5130 & n10176 ;
  assign n53974 = ~n40934 & n53973 ;
  assign n53975 = ( n1892 & ~n24977 ) | ( n1892 & n48873 ) | ( ~n24977 & n48873 ) ;
  assign n53976 = ~n22453 & n40336 ;
  assign n53977 = ~n53975 & n53976 ;
  assign n53978 = n53977 ^ n27872 ^ 1'b0 ;
  assign n53979 = n35019 ^ n16168 ^ n4878 ;
  assign n53980 = ( n34984 & n53978 ) | ( n34984 & n53979 ) | ( n53978 & n53979 ) ;
  assign n53981 = n3296 & ~n5703 ;
  assign n53982 = n45279 ^ n35346 ^ 1'b0 ;
  assign n53983 = ~n53981 & n53982 ;
  assign n53984 = n46099 ^ n34953 ^ n8161 ;
  assign n53985 = ( ~n29405 & n53983 ) | ( ~n29405 & n53984 ) | ( n53983 & n53984 ) ;
  assign n53986 = n46653 ^ n41145 ^ n7458 ;
  assign n53987 = n37007 ^ n32581 ^ n18041 ;
  assign n53988 = n34818 ^ n9888 ^ 1'b0 ;
  assign n53989 = n30565 & n53988 ;
  assign n53990 = ( n16007 & ~n53987 ) | ( n16007 & n53989 ) | ( ~n53987 & n53989 ) ;
  assign n53991 = ( ~n16748 & n23561 ) | ( ~n16748 & n51159 ) | ( n23561 & n51159 ) ;
  assign n53992 = n53991 ^ n32748 ^ n11695 ;
  assign n53993 = n39044 ^ n35797 ^ n27323 ;
  assign n53994 = ~n3723 & n9350 ;
  assign n53995 = n16766 | n53994 ;
  assign n53996 = n10363 & n11146 ;
  assign n53997 = ~n30486 & n53996 ;
  assign n53998 = n51975 ^ n9952 ^ 1'b0 ;
  assign n53999 = n43007 ^ n24275 ^ n3528 ;
  assign n54000 = ~n3099 & n53999 ;
  assign n54004 = n31383 ^ n27887 ^ n14204 ;
  assign n54003 = n28331 & ~n41350 ;
  assign n54001 = n3034 | n24103 ;
  assign n54002 = n54001 ^ n10415 ^ 1'b0 ;
  assign n54005 = n54004 ^ n54003 ^ n54002 ;
  assign n54006 = n18938 & n35579 ;
  assign n54007 = n33880 ^ n14898 ^ 1'b0 ;
  assign n54008 = n26026 & ~n54007 ;
  assign n54009 = n15243 & n19194 ;
  assign n54010 = ~n27864 & n54009 ;
  assign n54011 = ( ~n34233 & n54008 ) | ( ~n34233 & n54010 ) | ( n54008 & n54010 ) ;
  assign n54012 = n42836 ^ n18739 ^ n3659 ;
  assign n54013 = ( n18805 & ~n23681 ) | ( n18805 & n54012 ) | ( ~n23681 & n54012 ) ;
  assign n54014 = n26285 ^ n20999 ^ n4019 ;
  assign n54015 = n28029 & n38345 ;
  assign n54016 = ~n22844 & n54015 ;
  assign n54017 = n441 | n54016 ;
  assign n54018 = n54014 & ~n54017 ;
  assign n54019 = n54018 ^ n31399 ^ 1'b0 ;
  assign n54020 = n54019 ^ n42596 ^ n25338 ;
  assign n54021 = n2132 | n11832 ;
  assign n54022 = n1219 & n54021 ;
  assign n54023 = n54022 ^ n34731 ^ 1'b0 ;
  assign n54024 = n25431 ^ n4247 ^ 1'b0 ;
  assign n54025 = n6925 | n54024 ;
  assign n54026 = n32497 ^ n1419 ^ 1'b0 ;
  assign n54027 = n19650 & n54026 ;
  assign n54028 = n54027 ^ n36947 ^ 1'b0 ;
  assign n54029 = n48219 ^ n44029 ^ n39105 ;
  assign n54030 = n43543 ^ n17335 ^ 1'b0 ;
  assign n54031 = n25002 | n31277 ;
  assign n54032 = n31502 | n54031 ;
  assign n54033 = ( ~n17194 & n37446 ) | ( ~n17194 & n54032 ) | ( n37446 & n54032 ) ;
  assign n54034 = n10755 & ~n16156 ;
  assign n54035 = ( n6735 & n46120 ) | ( n6735 & ~n54034 ) | ( n46120 & ~n54034 ) ;
  assign n54036 = ( n13838 & n18643 ) | ( n13838 & n22380 ) | ( n18643 & n22380 ) ;
  assign n54037 = n24575 | n46899 ;
  assign n54038 = n54037 ^ n17343 ^ 1'b0 ;
  assign n54039 = ( n27793 & n54036 ) | ( n27793 & ~n54038 ) | ( n54036 & ~n54038 ) ;
  assign n54040 = ~n23763 & n46715 ;
  assign n54041 = n5912 | n9255 ;
  assign n54042 = n45168 ^ n9195 ^ 1'b0 ;
  assign n54043 = ( n7478 & n54041 ) | ( n7478 & n54042 ) | ( n54041 & n54042 ) ;
  assign n54044 = ( n20910 & n21847 ) | ( n20910 & n54043 ) | ( n21847 & n54043 ) ;
  assign n54045 = ( n53379 & ~n54040 ) | ( n53379 & n54044 ) | ( ~n54040 & n54044 ) ;
  assign n54046 = n16343 & n44769 ;
  assign n54047 = n21411 & n54046 ;
  assign n54048 = n24957 ^ n9278 ^ x179 ;
  assign n54049 = n21430 ^ n7439 ^ 1'b0 ;
  assign n54050 = ( n8609 & n43137 ) | ( n8609 & ~n54049 ) | ( n43137 & ~n54049 ) ;
  assign n54051 = ~n16930 & n52954 ;
  assign n54052 = n31543 | n47565 ;
  assign n54053 = n5939 & ~n54052 ;
  assign n54054 = n2170 & ~n25554 ;
  assign n54055 = ~n2104 & n54054 ;
  assign n54056 = n22915 | n54055 ;
  assign n54057 = n54056 ^ n9919 ^ 1'b0 ;
  assign n54058 = ( ~n8073 & n13972 ) | ( ~n8073 & n31945 ) | ( n13972 & n31945 ) ;
  assign n54059 = ( n45995 & ~n54057 ) | ( n45995 & n54058 ) | ( ~n54057 & n54058 ) ;
  assign n54060 = n16918 & n54059 ;
  assign n54061 = n54053 | n54060 ;
  assign n54062 = n47082 ^ n33931 ^ n418 ;
  assign n54063 = n511 & ~n36159 ;
  assign n54064 = ( n32926 & n41832 ) | ( n32926 & n54063 ) | ( n41832 & n54063 ) ;
  assign n54065 = ( n4177 & n26179 ) | ( n4177 & ~n43343 ) | ( n26179 & ~n43343 ) ;
  assign n54066 = n24060 ^ n4057 ^ 1'b0 ;
  assign n54067 = n43154 & ~n54066 ;
  assign n54068 = n14029 ^ n12599 ^ n5477 ;
  assign n54069 = n54068 ^ n36334 ^ n8547 ;
  assign n54070 = ( n24466 & n29539 ) | ( n24466 & ~n54069 ) | ( n29539 & ~n54069 ) ;
  assign n54071 = n54070 ^ n28727 ^ n15032 ;
  assign n54072 = n9659 ^ n1354 ^ 1'b0 ;
  assign n54073 = ~n54071 & n54072 ;
  assign n54074 = ~n5193 & n52091 ;
  assign n54075 = n10969 | n21343 ;
  assign n54076 = n4554 & ~n54075 ;
  assign n54077 = n25542 ^ n21543 ^ n16483 ;
  assign n54078 = ( n10308 & n32361 ) | ( n10308 & ~n54077 ) | ( n32361 & ~n54077 ) ;
  assign n54079 = n30931 ^ n9429 ^ 1'b0 ;
  assign n54080 = n49733 ^ n18402 ^ n14572 ;
  assign n54081 = ( n6299 & ~n35834 ) | ( n6299 & n54080 ) | ( ~n35834 & n54080 ) ;
  assign n54082 = n28073 ^ n11182 ^ 1'b0 ;
  assign n54083 = ( ~n6926 & n26684 ) | ( ~n6926 & n54082 ) | ( n26684 & n54082 ) ;
  assign n54084 = n29967 ^ n24444 ^ n9250 ;
  assign n54085 = n16687 ^ n2143 ^ 1'b0 ;
  assign n54086 = n54085 ^ n28547 ^ 1'b0 ;
  assign n54087 = ( n25754 & ~n48893 ) | ( n25754 & n54086 ) | ( ~n48893 & n54086 ) ;
  assign n54088 = n31421 ^ n23264 ^ n9128 ;
  assign n54089 = n1955 & n54088 ;
  assign n54090 = n44380 ^ n27572 ^ 1'b0 ;
  assign n54091 = n25205 | n54090 ;
  assign n54092 = n41648 ^ n26865 ^ n11649 ;
  assign n54093 = n5471 ^ n4335 ^ 1'b0 ;
  assign n54094 = ~n54092 & n54093 ;
  assign n54097 = ( n1408 & ~n15407 ) | ( n1408 & n34412 ) | ( ~n15407 & n34412 ) ;
  assign n54098 = ~n40361 & n54097 ;
  assign n54099 = ~n13493 & n54098 ;
  assign n54095 = n6915 & ~n46493 ;
  assign n54096 = n54095 ^ n22529 ^ 1'b0 ;
  assign n54100 = n54099 ^ n54096 ^ n3309 ;
  assign n54101 = n10711 ^ n7278 ^ 1'b0 ;
  assign n54102 = n10684 & ~n26525 ;
  assign n54103 = n54102 ^ n22535 ^ n19368 ;
  assign n54104 = ( n14146 & ~n24606 ) | ( n14146 & n43226 ) | ( ~n24606 & n43226 ) ;
  assign n54105 = n54104 ^ n19252 ^ n14040 ;
  assign n54109 = n5557 & n27715 ;
  assign n54110 = n54109 ^ n18188 ^ 1'b0 ;
  assign n54106 = n41066 ^ n31591 ^ 1'b0 ;
  assign n54107 = ~n1653 & n32347 ;
  assign n54108 = ~n54106 & n54107 ;
  assign n54111 = n54110 ^ n54108 ^ n2313 ;
  assign n54112 = n40810 ^ n22358 ^ n3230 ;
  assign n54113 = ( n1121 & ~n39641 ) | ( n1121 & n54112 ) | ( ~n39641 & n54112 ) ;
  assign n54114 = n13808 ^ n2379 ^ 1'b0 ;
  assign n54115 = n34471 | n54114 ;
  assign n54118 = n28910 ^ n22563 ^ n365 ;
  assign n54116 = n2091 | n41287 ;
  assign n54117 = n20838 & ~n54116 ;
  assign n54119 = n54118 ^ n54117 ^ 1'b0 ;
  assign n54120 = ( n21630 & n43021 ) | ( n21630 & n54119 ) | ( n43021 & n54119 ) ;
  assign n54121 = n54120 ^ n51714 ^ 1'b0 ;
  assign n54122 = n36840 & n54121 ;
  assign n54126 = n26286 ^ n14789 ^ n2200 ;
  assign n54123 = n52143 ^ n22989 ^ 1'b0 ;
  assign n54124 = ~x4 & n54123 ;
  assign n54125 = n15129 & n54124 ;
  assign n54127 = n54126 ^ n54125 ^ 1'b0 ;
  assign n54128 = n22130 ^ n18252 ^ 1'b0 ;
  assign n54129 = n36995 & ~n54128 ;
  assign n54130 = ~n18583 & n22190 ;
  assign n54131 = n18739 ^ n9618 ^ 1'b0 ;
  assign n54132 = ~n54130 & n54131 ;
  assign n54133 = n54132 ^ n40863 ^ n25123 ;
  assign n54134 = n54133 ^ n14595 ^ 1'b0 ;
  assign n54135 = ( ~n3583 & n10447 ) | ( ~n3583 & n54134 ) | ( n10447 & n54134 ) ;
  assign n54136 = n5773 | n50260 ;
  assign n54137 = n7442 & ~n54136 ;
  assign n54138 = n54137 ^ n30106 ^ n15429 ;
  assign n54139 = n54138 ^ n44929 ^ n4856 ;
  assign n54140 = n53142 ^ n30344 ^ 1'b0 ;
  assign n54141 = n9966 | n40733 ;
  assign n54142 = n54141 ^ n31594 ^ 1'b0 ;
  assign n54143 = ( n22325 & n48167 ) | ( n22325 & ~n54142 ) | ( n48167 & ~n54142 ) ;
  assign n54144 = n54143 ^ n30970 ^ n4771 ;
  assign n54145 = n42250 ^ n4588 ^ 1'b0 ;
  assign n54146 = n21104 ^ n19217 ^ 1'b0 ;
  assign n54147 = n393 & n54146 ;
  assign n54148 = ( n9589 & ~n40035 ) | ( n9589 & n41752 ) | ( ~n40035 & n41752 ) ;
  assign n54149 = ~n23628 & n54148 ;
  assign n54150 = ( n7035 & ~n29311 ) | ( n7035 & n54149 ) | ( ~n29311 & n54149 ) ;
  assign n54151 = n54150 ^ n32345 ^ n3631 ;
  assign n54152 = ~n24119 & n39711 ;
  assign n54153 = n6427 & n48804 ;
  assign n54154 = n47149 ^ n5909 ^ 1'b0 ;
  assign n54155 = n40893 & n54154 ;
  assign n54156 = n44705 ^ n22682 ^ 1'b0 ;
  assign n54157 = ( n43535 & ~n54155 ) | ( n43535 & n54156 ) | ( ~n54155 & n54156 ) ;
  assign n54158 = n48630 ^ n32902 ^ n22507 ;
  assign n54159 = ~n40725 & n54158 ;
  assign n54160 = n49388 ^ n33178 ^ n7802 ;
  assign n54161 = ( ~n8369 & n21545 ) | ( ~n8369 & n23247 ) | ( n21545 & n23247 ) ;
  assign n54162 = ( n34311 & n38558 ) | ( n34311 & n54161 ) | ( n38558 & n54161 ) ;
  assign n54163 = n36539 ^ n7409 ^ 1'b0 ;
  assign n54164 = x254 & ~n54163 ;
  assign n54165 = n54164 ^ n17977 ^ 1'b0 ;
  assign n54166 = n54165 ^ n823 ^ n410 ;
  assign n54167 = n18186 & ~n54166 ;
  assign n54171 = ( ~n626 & n18753 ) | ( ~n626 & n20630 ) | ( n18753 & n20630 ) ;
  assign n54172 = ( n20729 & n27508 ) | ( n20729 & n54171 ) | ( n27508 & n54171 ) ;
  assign n54173 = n54172 ^ n2842 ^ 1'b0 ;
  assign n54168 = n19882 ^ n11798 ^ 1'b0 ;
  assign n54169 = n8573 & n54168 ;
  assign n54170 = n54169 ^ n11156 ^ n6640 ;
  assign n54174 = n54173 ^ n54170 ^ n10778 ;
  assign n54175 = n54174 ^ n25117 ^ n21263 ;
  assign n54176 = ( n21549 & n41633 ) | ( n21549 & ~n54175 ) | ( n41633 & ~n54175 ) ;
  assign n54177 = n5180 | n50223 ;
  assign n54178 = n18348 & ~n54177 ;
  assign n54179 = n54178 ^ n14097 ^ n9212 ;
  assign n54181 = ~n20288 & n35295 ;
  assign n54180 = n2725 & n26075 ;
  assign n54182 = n54181 ^ n54180 ^ 1'b0 ;
  assign n54183 = n2880 ^ n2479 ^ 1'b0 ;
  assign n54184 = n32605 & n54183 ;
  assign n54185 = n15964 & n54184 ;
  assign n54186 = n54185 ^ n23939 ^ 1'b0 ;
  assign n54187 = n24590 & n50397 ;
  assign n54188 = n18986 & n54187 ;
  assign n54189 = n21491 & n27369 ;
  assign n54190 = n42508 ^ n23745 ^ n7345 ;
  assign n54191 = ( n891 & n50586 ) | ( n891 & ~n54190 ) | ( n50586 & ~n54190 ) ;
  assign n54192 = ( n6873 & n18664 ) | ( n6873 & ~n46489 ) | ( n18664 & ~n46489 ) ;
  assign n54193 = n47324 ^ n42765 ^ n36250 ;
  assign n54194 = n27353 ^ n13724 ^ n5145 ;
  assign n54195 = n54194 ^ n29518 ^ n3362 ;
  assign n54196 = n53182 ^ n30560 ^ 1'b0 ;
  assign n54197 = ~n45790 & n54196 ;
  assign n54198 = ( n10634 & n54195 ) | ( n10634 & ~n54197 ) | ( n54195 & ~n54197 ) ;
  assign n54199 = ( n28042 & n31465 ) | ( n28042 & n33917 ) | ( n31465 & n33917 ) ;
  assign n54200 = ( n23375 & n42990 ) | ( n23375 & ~n54199 ) | ( n42990 & ~n54199 ) ;
  assign n54202 = n17199 & n25566 ;
  assign n54203 = n54202 ^ n49791 ^ 1'b0 ;
  assign n54201 = ( n18774 & ~n23579 ) | ( n18774 & n45670 ) | ( ~n23579 & n45670 ) ;
  assign n54204 = n54203 ^ n54201 ^ n19821 ;
  assign n54205 = ( n15594 & ~n19886 ) | ( n15594 & n23587 ) | ( ~n19886 & n23587 ) ;
  assign n54206 = n54205 ^ n50899 ^ n33593 ;
  assign n54207 = n32240 | n49145 ;
  assign n54208 = n54207 ^ n50340 ^ 1'b0 ;
  assign n54209 = ( n25650 & ~n31539 ) | ( n25650 & n39797 ) | ( ~n31539 & n39797 ) ;
  assign n54210 = x190 & n1801 ;
  assign n54211 = n54209 & n54210 ;
  assign n54212 = n45622 ^ n7444 ^ 1'b0 ;
  assign n54213 = ~n54211 & n54212 ;
  assign n54214 = n11076 ^ n3044 ^ n2536 ;
  assign n54215 = ( n8080 & n20535 ) | ( n8080 & ~n20980 ) | ( n20535 & ~n20980 ) ;
  assign n54216 = n14772 | n15757 ;
  assign n54217 = n54216 ^ n36542 ^ 1'b0 ;
  assign n54218 = n54215 & n54217 ;
  assign n54219 = n43756 ^ n22644 ^ n17600 ;
  assign n54220 = n53484 ^ n45017 ^ n15585 ;
  assign n54221 = n42217 ^ n39367 ^ n7236 ;
  assign n54222 = ( n4980 & n44293 ) | ( n4980 & n54221 ) | ( n44293 & n54221 ) ;
  assign n54223 = ( n15518 & ~n29572 ) | ( n15518 & n41099 ) | ( ~n29572 & n41099 ) ;
  assign n54224 = n33770 & ~n54223 ;
  assign n54225 = n21990 & n43508 ;
  assign n54226 = n54225 ^ n14862 ^ 1'b0 ;
  assign n54227 = n54226 ^ n43574 ^ n12701 ;
  assign n54228 = ~n2800 & n17621 ;
  assign n54229 = n54228 ^ n31649 ^ 1'b0 ;
  assign n54230 = ~n1586 & n8798 ;
  assign n54231 = n54230 ^ n13092 ^ 1'b0 ;
  assign n54232 = n22423 & n37635 ;
  assign n54233 = ~n38467 & n54232 ;
  assign n54234 = n7617 | n34122 ;
  assign n54235 = ( ~n2752 & n27553 ) | ( ~n2752 & n41598 ) | ( n27553 & n41598 ) ;
  assign n54236 = ~n4332 & n6302 ;
  assign n54237 = ~x217 & n54236 ;
  assign n54238 = n41800 ^ n12036 ^ n7625 ;
  assign n54239 = n54238 ^ n47397 ^ 1'b0 ;
  assign n54240 = n47472 ^ n40692 ^ n5813 ;
  assign n54241 = ( ~n29736 & n44663 ) | ( ~n29736 & n54240 ) | ( n44663 & n54240 ) ;
  assign n54242 = ( n54237 & ~n54239 ) | ( n54237 & n54241 ) | ( ~n54239 & n54241 ) ;
  assign n54243 = n20376 & n45245 ;
  assign n54244 = ( n5206 & n8593 ) | ( n5206 & n22382 ) | ( n8593 & n22382 ) ;
  assign n54245 = ~n35347 & n45468 ;
  assign n54246 = n54245 ^ n39310 ^ 1'b0 ;
  assign n54247 = ( n29192 & ~n54244 ) | ( n29192 & n54246 ) | ( ~n54244 & n54246 ) ;
  assign n54248 = n54247 ^ n28988 ^ n24264 ;
  assign n54249 = n14445 & ~n42098 ;
  assign n54250 = n42098 ^ n10090 ^ n6797 ;
  assign n54251 = ( n5676 & n22396 ) | ( n5676 & n54250 ) | ( n22396 & n54250 ) ;
  assign n54252 = n54251 ^ n8991 ^ 1'b0 ;
  assign n54253 = ( ~n5118 & n54249 ) | ( ~n5118 & n54252 ) | ( n54249 & n54252 ) ;
  assign n54254 = ( n1614 & n35402 ) | ( n1614 & ~n36242 ) | ( n35402 & ~n36242 ) ;
  assign n54255 = n54254 ^ n15140 ^ 1'b0 ;
  assign n54256 = n14524 ^ n4440 ^ 1'b0 ;
  assign n54257 = ~n54255 & n54256 ;
  assign n54258 = n48640 & n54257 ;
  assign n54259 = n30139 ^ n24862 ^ 1'b0 ;
  assign n54260 = n2025 & n29316 ;
  assign n54261 = n7282 & n54260 ;
  assign n54262 = n44769 ^ n29564 ^ n13364 ;
  assign n54263 = n54262 ^ n46627 ^ 1'b0 ;
  assign n54264 = n32024 | n54263 ;
  assign n54265 = n760 & n18002 ;
  assign n54266 = ~n13578 & n54265 ;
  assign n54267 = ( n30387 & n34599 ) | ( n30387 & n50815 ) | ( n34599 & n50815 ) ;
  assign n54268 = n52291 ^ n41324 ^ n41046 ;
  assign n54269 = n27378 | n37785 ;
  assign n54270 = n49646 ^ n47567 ^ n38089 ;
  assign n54275 = ( n3991 & n9170 ) | ( n3991 & n9180 ) | ( n9170 & n9180 ) ;
  assign n54274 = n16921 ^ n11789 ^ n11447 ;
  assign n54271 = ( n10045 & n17900 ) | ( n10045 & ~n20916 ) | ( n17900 & ~n20916 ) ;
  assign n54272 = n23724 | n54271 ;
  assign n54273 = n54272 ^ n38471 ^ n24925 ;
  assign n54276 = n54275 ^ n54274 ^ n54273 ;
  assign n54277 = n52824 ^ n19321 ^ n6441 ;
  assign n54278 = n54277 ^ n14485 ^ n4182 ;
  assign n54279 = n26056 ^ n9180 ^ n3605 ;
  assign n54280 = n54279 ^ n52724 ^ n49646 ;
  assign n54281 = n54280 ^ n29335 ^ n4676 ;
  assign n54282 = n9760 ^ n8228 ^ 1'b0 ;
  assign n54283 = n6175 | n54282 ;
  assign n54284 = ( n15995 & n20637 ) | ( n15995 & ~n37080 ) | ( n20637 & ~n37080 ) ;
  assign n54285 = n54284 ^ n27460 ^ n24352 ;
  assign n54286 = ~n22056 & n26117 ;
  assign n54287 = n54285 & n54286 ;
  assign n54289 = n14053 & n14418 ;
  assign n54288 = n15448 ^ n5346 ^ n2929 ;
  assign n54290 = n54289 ^ n54288 ^ 1'b0 ;
  assign n54291 = n54290 ^ n6571 ^ 1'b0 ;
  assign n54292 = n26937 ^ n12557 ^ 1'b0 ;
  assign n54293 = ~n15281 & n54292 ;
  assign n54294 = n54293 ^ n20789 ^ n12497 ;
  assign n54295 = ( n20885 & n27607 ) | ( n20885 & n32926 ) | ( n27607 & n32926 ) ;
  assign n54296 = n8307 | n54295 ;
  assign n54297 = n54294 & ~n54296 ;
  assign n54298 = n41663 ^ n17304 ^ n16914 ;
  assign n54299 = n14038 ^ n12173 ^ n10164 ;
  assign n54300 = n23421 ^ n15849 ^ n10570 ;
  assign n54301 = n53639 ^ n38241 ^ 1'b0 ;
  assign n54302 = n54301 ^ n46117 ^ n29401 ;
  assign n54303 = n42520 ^ n34218 ^ n9233 ;
  assign n54304 = n54303 ^ n30010 ^ n12049 ;
  assign n54305 = n25870 & ~n41656 ;
  assign n54306 = n54305 ^ n17408 ^ 1'b0 ;
  assign n54307 = x222 | n54306 ;
  assign n54308 = ~n7355 & n9785 ;
  assign n54309 = n54308 ^ n7115 ^ 1'b0 ;
  assign n54310 = ( ~n23291 & n54307 ) | ( ~n23291 & n54309 ) | ( n54307 & n54309 ) ;
  assign n54311 = ( n31792 & n44345 ) | ( n31792 & n54310 ) | ( n44345 & n54310 ) ;
  assign n54312 = n44095 ^ n8395 ^ 1'b0 ;
  assign n54313 = ( n27742 & ~n37907 ) | ( n27742 & n54312 ) | ( ~n37907 & n54312 ) ;
  assign n54314 = n7362 ^ n4651 ^ 1'b0 ;
  assign n54315 = ~n36583 & n54314 ;
  assign n54316 = n14425 | n31363 ;
  assign n54317 = n42509 & ~n54316 ;
  assign n54318 = n26518 & ~n34438 ;
  assign n54319 = ~n36105 & n54318 ;
  assign n54320 = n26286 | n49045 ;
  assign n54321 = n54320 ^ n35469 ^ n2406 ;
  assign n54322 = n54321 ^ n2142 ^ 1'b0 ;
  assign n54323 = n54322 ^ n32305 ^ n11800 ;
  assign n54324 = ~n4915 & n31590 ;
  assign n54325 = n54324 ^ n49500 ^ 1'b0 ;
  assign n54326 = ( n16402 & ~n16768 ) | ( n16402 & n54325 ) | ( ~n16768 & n54325 ) ;
  assign n54327 = n33003 ^ n23908 ^ 1'b0 ;
  assign n54328 = ( n26614 & n35732 ) | ( n26614 & ~n44570 ) | ( n35732 & ~n44570 ) ;
  assign n54329 = ( n10235 & n54327 ) | ( n10235 & ~n54328 ) | ( n54327 & ~n54328 ) ;
  assign n54330 = n54329 ^ n51629 ^ n27593 ;
  assign n54331 = ( ~n11536 & n15470 ) | ( ~n11536 & n26139 ) | ( n15470 & n26139 ) ;
  assign n54332 = n35416 ^ n24208 ^ n2980 ;
  assign n54333 = ( ~n13045 & n37614 ) | ( ~n13045 & n49819 ) | ( n37614 & n49819 ) ;
  assign n54334 = ( ~n23818 & n37779 ) | ( ~n23818 & n54333 ) | ( n37779 & n54333 ) ;
  assign n54335 = n54334 ^ n30181 ^ 1'b0 ;
  assign n54336 = n54332 & n54335 ;
  assign n54337 = n54336 ^ n6887 ^ n5818 ;
  assign n54338 = n7643 & n20247 ;
  assign n54339 = ( ~n2051 & n46436 ) | ( ~n2051 & n54338 ) | ( n46436 & n54338 ) ;
  assign n54340 = n51558 ^ n6928 ^ n6820 ;
  assign n54341 = n9496 & ~n25794 ;
  assign n54342 = n38411 ^ n32178 ^ 1'b0 ;
  assign n54343 = ~n19588 & n54342 ;
  assign n54344 = ( n2101 & n42091 ) | ( n2101 & n49871 ) | ( n42091 & n49871 ) ;
  assign n54345 = ( n6648 & n18308 ) | ( n6648 & n24514 ) | ( n18308 & n24514 ) ;
  assign n54346 = n54345 ^ n30955 ^ n6352 ;
  assign n54347 = n54346 ^ n28696 ^ n16250 ;
  assign n54348 = ( n8145 & n15352 ) | ( n8145 & n25355 ) | ( n15352 & n25355 ) ;
  assign n54349 = ( n10043 & ~n12055 ) | ( n10043 & n16373 ) | ( ~n12055 & n16373 ) ;
  assign n54353 = n20119 ^ n5729 ^ n585 ;
  assign n54350 = n8031 ^ n1485 ^ 1'b0 ;
  assign n54351 = n54350 ^ n24167 ^ 1'b0 ;
  assign n54352 = n20478 & ~n54351 ;
  assign n54354 = n54353 ^ n54352 ^ n34163 ;
  assign n54355 = n54354 ^ n35903 ^ n8762 ;
  assign n54356 = ( n14402 & ~n21467 ) | ( n14402 & n28082 ) | ( ~n21467 & n28082 ) ;
  assign n54359 = n17557 ^ n10204 ^ n4446 ;
  assign n54360 = ( x109 & n37359 ) | ( x109 & ~n54359 ) | ( n37359 & ~n54359 ) ;
  assign n54357 = ( n672 & n4862 ) | ( n672 & n37129 ) | ( n4862 & n37129 ) ;
  assign n54358 = ( ~n20458 & n21506 ) | ( ~n20458 & n54357 ) | ( n21506 & n54357 ) ;
  assign n54361 = n54360 ^ n54358 ^ n16312 ;
  assign n54362 = ~n273 & n15405 ;
  assign n54363 = n54362 ^ n10471 ^ 1'b0 ;
  assign n54364 = n1760 & ~n13146 ;
  assign n54365 = n54364 ^ n24980 ^ 1'b0 ;
  assign n54366 = n7346 ^ n6821 ^ 1'b0 ;
  assign n54367 = ~n54365 & n54366 ;
  assign n54368 = ~n16214 & n39135 ;
  assign n54369 = ~x233 & n54368 ;
  assign n54370 = ( n3902 & n8707 ) | ( n3902 & ~n21880 ) | ( n8707 & ~n21880 ) ;
  assign n54371 = ( n2352 & ~n14391 ) | ( n2352 & n54370 ) | ( ~n14391 & n54370 ) ;
  assign n54372 = ~n21007 & n54371 ;
  assign n54373 = n43610 & n54372 ;
  assign n54374 = n54133 ^ n20711 ^ n17749 ;
  assign n54375 = n54374 ^ n6544 ^ n5759 ;
  assign n54376 = ( ~n4571 & n26097 ) | ( ~n4571 & n33063 ) | ( n26097 & n33063 ) ;
  assign n54377 = n54376 ^ n10439 ^ x219 ;
  assign n54378 = n54377 ^ n36806 ^ n31455 ;
  assign n54379 = ( ~n5782 & n10831 ) | ( ~n5782 & n30071 ) | ( n10831 & n30071 ) ;
  assign n54380 = ( n13265 & n30309 ) | ( n13265 & ~n54379 ) | ( n30309 & ~n54379 ) ;
  assign n54383 = n8854 ^ x235 ^ 1'b0 ;
  assign n54381 = ~n1582 & n37729 ;
  assign n54382 = n54381 ^ n28813 ^ 1'b0 ;
  assign n54384 = n54383 ^ n54382 ^ 1'b0 ;
  assign n54385 = n54384 ^ n24588 ^ 1'b0 ;
  assign n54386 = n23984 ^ n14644 ^ n7050 ;
  assign n54387 = ( n8342 & ~n21199 ) | ( n8342 & n23754 ) | ( ~n21199 & n23754 ) ;
  assign n54388 = n6715 & ~n23237 ;
  assign n54389 = ~n3969 & n54388 ;
  assign n54390 = n54389 ^ n913 ^ 1'b0 ;
  assign n54391 = n16147 & ~n54390 ;
  assign n54392 = n19736 ^ n19354 ^ 1'b0 ;
  assign n54393 = n24275 | n54392 ;
  assign n54394 = n1112 | n54393 ;
  assign n54395 = n2894 | n17284 ;
  assign n54396 = n30174 | n54395 ;
  assign n54397 = ~n3108 & n15997 ;
  assign n54398 = ( n16690 & n30157 ) | ( n16690 & n32439 ) | ( n30157 & n32439 ) ;
  assign n54399 = n54398 ^ n43947 ^ n14943 ;
  assign n54400 = ( n29380 & ~n32834 ) | ( n29380 & n34692 ) | ( ~n32834 & n34692 ) ;
  assign n54401 = n12242 & n26681 ;
  assign n54402 = n10144 ^ n1951 ^ 1'b0 ;
  assign n54403 = ~n7072 & n54402 ;
  assign n54404 = n2301 & ~n19684 ;
  assign n54405 = ~n54403 & n54404 ;
  assign n54406 = ( n14998 & n36284 ) | ( n14998 & n54405 ) | ( n36284 & n54405 ) ;
  assign n54408 = n36587 ^ n19003 ^ n10352 ;
  assign n54407 = n18037 ^ n1104 ^ 1'b0 ;
  assign n54409 = n54408 ^ n54407 ^ n28723 ;
  assign n54410 = n53209 ^ n42072 ^ 1'b0 ;
  assign n54411 = n18167 & ~n54410 ;
  assign n54412 = n54411 ^ n28647 ^ n25451 ;
  assign n54413 = n24037 ^ n3838 ^ 1'b0 ;
  assign n54414 = n42237 & n54413 ;
  assign n54415 = n24571 ^ n9075 ^ 1'b0 ;
  assign n54416 = n14544 & ~n54415 ;
  assign n54417 = ( n9842 & ~n11221 ) | ( n9842 & n46682 ) | ( ~n11221 & n46682 ) ;
  assign n54418 = n16942 & n24620 ;
  assign n54419 = ( n13245 & ~n44120 ) | ( n13245 & n54418 ) | ( ~n44120 & n54418 ) ;
  assign n54420 = ~n13339 & n21789 ;
  assign n54421 = n54420 ^ n33219 ^ n29375 ;
  assign n54422 = n54421 ^ n31477 ^ n16959 ;
  assign n54423 = n54178 ^ n36265 ^ n6768 ;
  assign n54424 = ( n1697 & ~n16426 ) | ( n1697 & n34645 ) | ( ~n16426 & n34645 ) ;
  assign n54425 = ( n14892 & n27612 ) | ( n14892 & n40307 ) | ( n27612 & n40307 ) ;
  assign n54426 = n19366 ^ n6709 ^ 1'b0 ;
  assign n54427 = ~n10735 & n54426 ;
  assign n54428 = n54427 ^ n26051 ^ n1031 ;
  assign n54429 = n54428 ^ n28473 ^ n20309 ;
  assign n54430 = n16548 ^ n6188 ^ n5309 ;
  assign n54431 = n54430 ^ n49051 ^ n14282 ;
  assign n54432 = n10011 & ~n54431 ;
  assign n54433 = n54432 ^ n36412 ^ 1'b0 ;
  assign n54434 = n46448 ^ n28462 ^ n27706 ;
  assign n54435 = n21217 ^ n308 ^ 1'b0 ;
  assign n54436 = n17170 & n54435 ;
  assign n54437 = ( ~n7262 & n49489 ) | ( ~n7262 & n54436 ) | ( n49489 & n54436 ) ;
  assign n54438 = n28698 ^ n18778 ^ 1'b0 ;
  assign n54439 = ( n3326 & n35288 ) | ( n3326 & ~n54438 ) | ( n35288 & ~n54438 ) ;
  assign n54442 = n5062 | n27520 ;
  assign n54443 = n14490 | n54442 ;
  assign n54444 = n54443 ^ n6736 ^ n3726 ;
  assign n54445 = ( n735 & n7164 ) | ( n735 & ~n10700 ) | ( n7164 & ~n10700 ) ;
  assign n54446 = n54445 ^ n42251 ^ 1'b0 ;
  assign n54447 = n54444 | n54446 ;
  assign n54440 = n27286 ^ n23640 ^ n19486 ;
  assign n54441 = n54440 ^ n38639 ^ n23168 ;
  assign n54448 = n54447 ^ n54441 ^ n2356 ;
  assign n54449 = n43643 ^ n37911 ^ n17906 ;
  assign n54450 = ( n12112 & ~n13247 ) | ( n12112 & n22489 ) | ( ~n13247 & n22489 ) ;
  assign n54451 = n31155 & n39324 ;
  assign n54452 = n54451 ^ n20256 ^ 1'b0 ;
  assign n54453 = n17619 & ~n35174 ;
  assign n54454 = ( n2928 & n30294 ) | ( n2928 & ~n32544 ) | ( n30294 & ~n32544 ) ;
  assign n54455 = n54454 ^ n31829 ^ n13567 ;
  assign n54456 = ( ~n7349 & n19233 ) | ( ~n7349 & n54124 ) | ( n19233 & n54124 ) ;
  assign n54457 = ( n14835 & ~n22553 ) | ( n14835 & n42557 ) | ( ~n22553 & n42557 ) ;
  assign n54460 = ( n1823 & n14286 ) | ( n1823 & ~n29846 ) | ( n14286 & ~n29846 ) ;
  assign n54461 = ( n4728 & ~n9793 ) | ( n4728 & n14879 ) | ( ~n9793 & n14879 ) ;
  assign n54462 = n54461 ^ n4872 ^ 1'b0 ;
  assign n54463 = n54460 & n54462 ;
  assign n54458 = ( ~n1001 & n10103 ) | ( ~n1001 & n30263 ) | ( n10103 & n30263 ) ;
  assign n54459 = ~n13084 & n54458 ;
  assign n54464 = n54463 ^ n54459 ^ n13139 ;
  assign n54465 = ( n17142 & ~n28097 ) | ( n17142 & n32698 ) | ( ~n28097 & n32698 ) ;
  assign n54466 = n23466 ^ n5418 ^ n1309 ;
  assign n54468 = n20123 | n48663 ;
  assign n54467 = n16538 & n22246 ;
  assign n54469 = n54468 ^ n54467 ^ n17710 ;
  assign n54470 = n43518 ^ n38775 ^ 1'b0 ;
  assign n54471 = n9686 | n54470 ;
  assign n54473 = n13105 ^ n4042 ^ 1'b0 ;
  assign n54474 = n6772 | n54473 ;
  assign n54472 = n33572 & ~n34639 ;
  assign n54475 = n54474 ^ n54472 ^ 1'b0 ;
  assign n54476 = ( n1907 & n28340 ) | ( n1907 & n37606 ) | ( n28340 & n37606 ) ;
  assign n54477 = n44911 ^ n30032 ^ n21579 ;
  assign n54478 = ~n16421 & n31589 ;
  assign n54479 = n1719 & n54478 ;
  assign n54480 = ( ~n28983 & n39516 ) | ( ~n28983 & n54479 ) | ( n39516 & n54479 ) ;
  assign n54481 = n44485 ^ n42647 ^ 1'b0 ;
  assign n54486 = n27662 ^ n20311 ^ n4190 ;
  assign n54485 = n18414 ^ n16193 ^ 1'b0 ;
  assign n54483 = n27955 ^ n7139 ^ n5603 ;
  assign n54482 = n41981 & ~n49800 ;
  assign n54484 = n54483 ^ n54482 ^ 1'b0 ;
  assign n54487 = n54486 ^ n54485 ^ n54484 ;
  assign n54488 = n36088 ^ n26750 ^ 1'b0 ;
  assign n54489 = n28597 ^ n19296 ^ n10298 ;
  assign n54490 = n30781 & ~n54489 ;
  assign n54491 = n54490 ^ n40430 ^ 1'b0 ;
  assign n54492 = n54491 ^ n40217 ^ n6026 ;
  assign n54493 = n38055 ^ n31063 ^ 1'b0 ;
  assign n54494 = ~n11520 & n54493 ;
  assign n54495 = ( n1690 & n21372 ) | ( n1690 & ~n22280 ) | ( n21372 & ~n22280 ) ;
  assign n54496 = ~n6664 & n54495 ;
  assign n54497 = n10634 & n54496 ;
  assign n54498 = n52775 ^ n34797 ^ n28878 ;
  assign n54499 = n54498 ^ n49652 ^ n32086 ;
  assign n54500 = n7448 ^ n4579 ^ 1'b0 ;
  assign n54501 = ( ~n4432 & n8635 ) | ( ~n4432 & n36278 ) | ( n8635 & n36278 ) ;
  assign n54502 = n21771 | n42556 ;
  assign n54503 = n5208 | n54502 ;
  assign n54504 = n54503 ^ n31028 ^ n29836 ;
  assign n54505 = n6474 & ~n43601 ;
  assign n54506 = n15494 & ~n17672 ;
  assign n54507 = ~n5500 & n54506 ;
  assign n54508 = ( n35381 & n41493 ) | ( n35381 & ~n54507 ) | ( n41493 & ~n54507 ) ;
  assign n54510 = n26880 ^ n970 ^ 1'b0 ;
  assign n54509 = n17646 & n22844 ;
  assign n54511 = n54510 ^ n54509 ^ 1'b0 ;
  assign n54512 = n36357 & n47455 ;
  assign n54513 = ~n25631 & n54512 ;
  assign n54514 = n54513 ^ n40805 ^ 1'b0 ;
  assign n54515 = n41350 & ~n54514 ;
  assign n54516 = n11144 | n12703 ;
  assign n54517 = n32935 ^ n12836 ^ n1493 ;
  assign n54518 = n25629 ^ n1804 ^ n894 ;
  assign n54519 = n54517 & ~n54518 ;
  assign n54520 = ( n2268 & n6042 ) | ( n2268 & n54519 ) | ( n6042 & n54519 ) ;
  assign n54521 = n42404 ^ n19300 ^ n18896 ;
  assign n54522 = n6716 & ~n20835 ;
  assign n54523 = ( ~n15656 & n34703 ) | ( ~n15656 & n54522 ) | ( n34703 & n54522 ) ;
  assign n54527 = n39001 & n42599 ;
  assign n54524 = n17962 & n22680 ;
  assign n54525 = ~n16634 & n54524 ;
  assign n54526 = n54525 ^ n9903 ^ n489 ;
  assign n54528 = n54527 ^ n54526 ^ n14729 ;
  assign n54529 = ( ~n3701 & n23662 ) | ( ~n3701 & n38514 ) | ( n23662 & n38514 ) ;
  assign n54530 = n1627 | n45211 ;
  assign n54531 = n54530 ^ n33073 ^ 1'b0 ;
  assign n54532 = n54531 ^ n39166 ^ n4175 ;
  assign n54533 = ( ~n32871 & n33089 ) | ( ~n32871 & n46832 ) | ( n33089 & n46832 ) ;
  assign n54534 = n22106 & ~n42786 ;
  assign n54535 = n54534 ^ n29159 ^ 1'b0 ;
  assign n54536 = n4554 & ~n4837 ;
  assign n54537 = ~n30788 & n54536 ;
  assign n54538 = n22513 & n26849 ;
  assign n54539 = ~n19059 & n53471 ;
  assign n54540 = ( n656 & n16125 ) | ( n656 & ~n53923 ) | ( n16125 & ~n53923 ) ;
  assign n54541 = n24310 ^ n19073 ^ n997 ;
  assign n54542 = n41051 ^ n21757 ^ n10364 ;
  assign n54543 = n54542 ^ n36954 ^ n29430 ;
  assign n54544 = ( n24770 & n54541 ) | ( n24770 & n54543 ) | ( n54541 & n54543 ) ;
  assign n54545 = n26954 ^ n16729 ^ n3600 ;
  assign n54546 = n54545 ^ n26296 ^ n20150 ;
  assign n54547 = n54546 ^ n16717 ^ n14909 ;
  assign n54548 = ( n27859 & n44110 ) | ( n27859 & n54547 ) | ( n44110 & n54547 ) ;
  assign n54549 = ( n21600 & ~n35733 ) | ( n21600 & n39225 ) | ( ~n35733 & n39225 ) ;
  assign n54550 = n32527 ^ n11045 ^ x203 ;
  assign n54551 = n5344 & ~n27353 ;
  assign n54552 = n54551 ^ n27858 ^ 1'b0 ;
  assign n54553 = n54550 & ~n54552 ;
  assign n54554 = ( n7039 & n8150 ) | ( n7039 & ~n21365 ) | ( n8150 & ~n21365 ) ;
  assign n54555 = n13233 ^ n7377 ^ 1'b0 ;
  assign n54556 = n45936 | n54555 ;
  assign n54557 = ( n27728 & n54554 ) | ( n27728 & n54556 ) | ( n54554 & n54556 ) ;
  assign n54558 = n54557 ^ n17160 ^ 1'b0 ;
  assign n54559 = n15540 | n49874 ;
  assign n54560 = n54559 ^ n25299 ^ 1'b0 ;
  assign n54561 = n54560 ^ n36968 ^ n15912 ;
  assign n54562 = ~n6762 & n49490 ;
  assign n54563 = ~n20234 & n54562 ;
  assign n54564 = ~n4824 & n51855 ;
  assign n54565 = n54564 ^ n29872 ^ 1'b0 ;
  assign n54566 = ( n19342 & n30919 ) | ( n19342 & ~n39412 ) | ( n30919 & ~n39412 ) ;
  assign n54567 = n27261 ^ n23505 ^ n14057 ;
  assign n54568 = n30383 ^ n22866 ^ 1'b0 ;
  assign n54569 = n21293 & ~n54568 ;
  assign n54570 = n54569 ^ n47612 ^ n26332 ;
  assign n54571 = n38908 ^ n20850 ^ n8979 ;
  assign n54572 = ( n7199 & n8504 ) | ( n7199 & n54571 ) | ( n8504 & n54571 ) ;
  assign n54573 = n54572 ^ n42115 ^ n9228 ;
  assign n54574 = n30803 ^ n21532 ^ n20273 ;
  assign n54575 = n53184 ^ n45966 ^ n37285 ;
  assign n54576 = ( x24 & n16758 ) | ( x24 & ~n46243 ) | ( n16758 & ~n46243 ) ;
  assign n54577 = n35560 ^ n1511 ^ 1'b0 ;
  assign n54578 = n18068 & ~n54577 ;
  assign n54579 = ~n1322 & n3352 ;
  assign n54580 = n54579 ^ n32131 ^ 1'b0 ;
  assign n54581 = n13349 ^ n11912 ^ 1'b0 ;
  assign n54582 = n26650 & n54581 ;
  assign n54585 = ( n542 & ~n5970 ) | ( n542 & n23815 ) | ( ~n5970 & n23815 ) ;
  assign n54583 = n36967 ^ n6503 ^ n346 ;
  assign n54584 = n53279 & n54583 ;
  assign n54586 = n54585 ^ n54584 ^ n44857 ;
  assign n54587 = n44079 ^ n6544 ^ n5574 ;
  assign n54588 = ~n5336 & n7363 ;
  assign n54589 = ~n33650 & n54588 ;
  assign n54590 = ( ~n41574 & n54587 ) | ( ~n41574 & n54589 ) | ( n54587 & n54589 ) ;
  assign n54591 = ~n10464 & n31338 ;
  assign n54592 = ( n14402 & n47993 ) | ( n14402 & n54591 ) | ( n47993 & n54591 ) ;
  assign n54593 = n7954 | n26950 ;
  assign n54594 = n19091 | n54593 ;
  assign n54595 = n38939 ^ n21406 ^ n17982 ;
  assign n54596 = ( n32411 & ~n54594 ) | ( n32411 & n54595 ) | ( ~n54594 & n54595 ) ;
  assign n54597 = n25484 ^ n10550 ^ n7900 ;
  assign n54598 = n14577 | n40076 ;
  assign n54599 = ( ~n17917 & n50453 ) | ( ~n17917 & n54598 ) | ( n50453 & n54598 ) ;
  assign n54600 = n37430 ^ n18671 ^ n10886 ;
  assign n54601 = n54600 ^ n40373 ^ 1'b0 ;
  assign n54603 = n7593 | n44586 ;
  assign n54602 = n1682 & n42315 ;
  assign n54604 = n54603 ^ n54602 ^ 1'b0 ;
  assign n54605 = n27655 ^ n13993 ^ 1'b0 ;
  assign n54606 = n46265 | n54605 ;
  assign n54607 = n24476 ^ n11308 ^ n9855 ;
  assign n54608 = n54607 ^ n50896 ^ 1'b0 ;
  assign n54609 = n15541 & ~n54608 ;
  assign n54610 = ( n7035 & ~n31223 ) | ( n7035 & n51543 ) | ( ~n31223 & n51543 ) ;
  assign n54611 = n17962 ^ n5275 ^ 1'b0 ;
  assign n54612 = n54611 ^ n23374 ^ n2395 ;
  assign n54613 = n54612 ^ n21456 ^ n17421 ;
  assign n54614 = ( n3023 & n54610 ) | ( n3023 & ~n54613 ) | ( n54610 & ~n54613 ) ;
  assign n54615 = n31330 & ~n49019 ;
  assign n54616 = n28972 ^ n20824 ^ n6767 ;
  assign n54617 = n7617 ^ n7243 ^ n1407 ;
  assign n54618 = n54617 ^ n41793 ^ n10747 ;
  assign n54619 = ~n14518 & n17372 ;
  assign n54620 = n54542 ^ n5119 ^ 1'b0 ;
  assign n54622 = n35563 ^ n1893 ^ 1'b0 ;
  assign n54621 = n1588 & n43412 ;
  assign n54623 = n54622 ^ n54621 ^ 1'b0 ;
  assign n54624 = n11577 ^ n8936 ^ 1'b0 ;
  assign n54625 = ~n23669 & n54624 ;
  assign n54626 = n13245 | n48056 ;
  assign n54627 = n54626 ^ n10144 ^ 1'b0 ;
  assign n54628 = n4397 | n15899 ;
  assign n54629 = ( n25602 & n31933 ) | ( n25602 & n37931 ) | ( n31933 & n37931 ) ;
  assign n54630 = n39535 ^ n21259 ^ 1'b0 ;
  assign n54631 = n28422 ^ n3728 ^ n2801 ;
  assign n54632 = n24920 ^ n24559 ^ 1'b0 ;
  assign n54633 = n39911 & ~n54632 ;
  assign n54634 = ( n7171 & ~n8924 ) | ( n7171 & n54633 ) | ( ~n8924 & n54633 ) ;
  assign n54635 = ( n3881 & n22413 ) | ( n3881 & n42058 ) | ( n22413 & n42058 ) ;
  assign n54636 = ( ~n28235 & n29548 ) | ( ~n28235 & n54008 ) | ( n29548 & n54008 ) ;
  assign n54637 = n39997 ^ n37253 ^ n6281 ;
  assign n54638 = ( n15746 & n16348 ) | ( n15746 & n54637 ) | ( n16348 & n54637 ) ;
  assign n54639 = n22481 | n25996 ;
  assign n54640 = n38297 | n54639 ;
  assign n54641 = ( n12784 & ~n20342 ) | ( n12784 & n29539 ) | ( ~n20342 & n29539 ) ;
  assign n54642 = n48651 ^ n44324 ^ n24594 ;
  assign n54643 = ( n12663 & n39831 ) | ( n12663 & n54642 ) | ( n39831 & n54642 ) ;
  assign n54644 = n4017 ^ x226 ^ 1'b0 ;
  assign n54645 = ( n10112 & ~n17974 ) | ( n10112 & n54644 ) | ( ~n17974 & n54644 ) ;
  assign n54647 = ( n11591 & ~n17342 ) | ( n11591 & n36784 ) | ( ~n17342 & n36784 ) ;
  assign n54646 = ( ~n1710 & n4397 ) | ( ~n1710 & n51585 ) | ( n4397 & n51585 ) ;
  assign n54648 = n54647 ^ n54646 ^ n42038 ;
  assign n54649 = n48831 ^ n15782 ^ 1'b0 ;
  assign n54650 = n54165 ^ n41631 ^ n2846 ;
  assign n54651 = n46671 ^ n41545 ^ n39758 ;
  assign n54652 = n17778 | n17884 ;
  assign n54653 = n54652 ^ n44273 ^ 1'b0 ;
  assign n54657 = ~n7917 & n23640 ;
  assign n54658 = ~n27965 & n54657 ;
  assign n54654 = n25175 & n52366 ;
  assign n54655 = n54654 ^ n46346 ^ 1'b0 ;
  assign n54656 = n4903 | n54655 ;
  assign n54659 = n54658 ^ n54656 ^ 1'b0 ;
  assign n54660 = n12912 ^ n1035 ^ 1'b0 ;
  assign n54661 = n23646 & ~n54660 ;
  assign n54662 = n54661 ^ n32188 ^ n4545 ;
  assign n54663 = n6691 & n54662 ;
  assign n54664 = ( n4933 & n21172 ) | ( n4933 & n40625 ) | ( n21172 & n40625 ) ;
  assign n54665 = n47212 ^ n10565 ^ n10011 ;
  assign n54666 = n54665 ^ n16187 ^ n2247 ;
  assign n54667 = n24543 ^ n21503 ^ n8703 ;
  assign n54668 = n14428 & ~n26574 ;
  assign n54669 = n54668 ^ n4284 ^ 1'b0 ;
  assign n54670 = n54669 ^ n42587 ^ n36445 ;
  assign n54671 = n5524 & n42250 ;
  assign n54672 = n54671 ^ n18359 ^ 1'b0 ;
  assign n54673 = n40815 ^ n17145 ^ n7180 ;
  assign n54674 = ( n4654 & n32240 ) | ( n4654 & n54673 ) | ( n32240 & n54673 ) ;
  assign n54675 = ( n18209 & ~n54672 ) | ( n18209 & n54674 ) | ( ~n54672 & n54674 ) ;
  assign n54676 = ( ~n5873 & n11843 ) | ( ~n5873 & n29079 ) | ( n11843 & n29079 ) ;
  assign n54678 = n12289 & ~n12818 ;
  assign n54679 = n54678 ^ n6743 ^ 1'b0 ;
  assign n54677 = n3407 & ~n4352 ;
  assign n54680 = n54679 ^ n54677 ^ 1'b0 ;
  assign n54681 = n49995 ^ n22912 ^ 1'b0 ;
  assign n54682 = n38225 | n54681 ;
  assign n54683 = n6951 ^ n5657 ^ n5426 ;
  assign n54684 = ( ~n12270 & n33128 ) | ( ~n12270 & n54683 ) | ( n33128 & n54683 ) ;
  assign n54685 = n45908 ^ n19646 ^ n10488 ;
  assign n54686 = n33845 ^ n24244 ^ n6287 ;
  assign n54687 = n54686 ^ n21610 ^ n20148 ;
  assign n54688 = ( ~n513 & n8682 ) | ( ~n513 & n26613 ) | ( n8682 & n26613 ) ;
  assign n54689 = n23943 ^ n18544 ^ n857 ;
  assign n54690 = n54689 ^ n20286 ^ 1'b0 ;
  assign n54691 = n42043 ^ n3158 ^ n2824 ;
  assign n54692 = n10215 & n51058 ;
  assign n54693 = n16446 ^ n6722 ^ n6239 ;
  assign n54694 = n54693 ^ n24687 ^ n5531 ;
  assign n54695 = n25494 & n54694 ;
  assign n54696 = ~n11024 & n54695 ;
  assign n54697 = ~n1970 & n20341 ;
  assign n54698 = n27676 ^ n16379 ^ n15805 ;
  assign n54699 = n53217 & ~n54698 ;
  assign n54700 = ( ~n4771 & n15914 ) | ( ~n4771 & n37806 ) | ( n15914 & n37806 ) ;
  assign n54702 = n36912 ^ n14625 ^ 1'b0 ;
  assign n54703 = ( n8886 & n9692 ) | ( n8886 & ~n54702 ) | ( n9692 & ~n54702 ) ;
  assign n54701 = ( ~n2800 & n15485 ) | ( ~n2800 & n27691 ) | ( n15485 & n27691 ) ;
  assign n54704 = n54703 ^ n54701 ^ n15504 ;
  assign n54705 = n39487 ^ n9099 ^ 1'b0 ;
  assign n54708 = n37308 ^ n20260 ^ 1'b0 ;
  assign n54709 = n14853 & ~n54708 ;
  assign n54710 = n54709 ^ n9202 ^ 1'b0 ;
  assign n54706 = n41704 ^ n11554 ^ 1'b0 ;
  assign n54707 = n19829 & ~n54706 ;
  assign n54711 = n54710 ^ n54707 ^ n3829 ;
  assign n54712 = ( n11983 & n34200 ) | ( n11983 & n46769 ) | ( n34200 & n46769 ) ;
  assign n54713 = ( n17445 & ~n32953 ) | ( n17445 & n48609 ) | ( ~n32953 & n48609 ) ;
  assign n54714 = n54713 ^ n22797 ^ 1'b0 ;
  assign n54715 = n1142 & ~n17362 ;
  assign n54716 = n54715 ^ n20903 ^ n19869 ;
  assign n54717 = ( n40081 & n40508 ) | ( n40081 & ~n54716 ) | ( n40508 & ~n54716 ) ;
  assign n54718 = n35604 ^ n13495 ^ 1'b0 ;
  assign n54719 = n4376 | n54718 ;
  assign n54720 = ( n22756 & n27146 ) | ( n22756 & ~n54719 ) | ( n27146 & ~n54719 ) ;
  assign n54721 = n15010 & n49736 ;
  assign n54722 = ~n54720 & n54721 ;
  assign n54723 = n15477 ^ n14740 ^ 1'b0 ;
  assign n54724 = x38 & n54723 ;
  assign n54725 = n531 & ~n32271 ;
  assign n54726 = ~n54724 & n54725 ;
  assign n54727 = n5526 | n18384 ;
  assign n54728 = n54727 ^ n21743 ^ 1'b0 ;
  assign n54729 = n51180 & n54728 ;
  assign n54730 = n4880 & n9002 ;
  assign n54731 = n46029 & n54730 ;
  assign n54732 = n54731 ^ n52198 ^ n4876 ;
  assign n54733 = n8720 ^ n6448 ^ n2572 ;
  assign n54734 = n24203 & ~n54733 ;
  assign n54735 = ~n51911 & n54557 ;
  assign n54736 = ( ~n1376 & n18966 ) | ( ~n1376 & n42591 ) | ( n18966 & n42591 ) ;
  assign n54737 = n54736 ^ n42451 ^ n25149 ;
  assign n54738 = ( n7713 & n8793 ) | ( n7713 & ~n37855 ) | ( n8793 & ~n37855 ) ;
  assign n54739 = n54738 ^ n21540 ^ 1'b0 ;
  assign n54740 = n32240 ^ n16637 ^ n10088 ;
  assign n54741 = n54740 ^ n35104 ^ n2490 ;
  assign n54742 = ( n4333 & n21070 ) | ( n4333 & n28587 ) | ( n21070 & n28587 ) ;
  assign n54743 = n15563 ^ n2216 ^ 1'b0 ;
  assign n54744 = n46772 | n54743 ;
  assign n54745 = n12036 ^ n7529 ^ 1'b0 ;
  assign n54746 = n26803 & ~n54745 ;
  assign n54747 = ~n4858 & n9136 ;
  assign n54748 = n54747 ^ n14345 ^ 1'b0 ;
  assign n54749 = n19007 & ~n35815 ;
  assign n54752 = n17074 ^ n8145 ^ 1'b0 ;
  assign n54753 = n1172 & ~n54752 ;
  assign n54750 = n34345 ^ n18660 ^ 1'b0 ;
  assign n54751 = n54750 ^ n15071 ^ n9209 ;
  assign n54754 = n54753 ^ n54751 ^ n24854 ;
  assign n54755 = n21217 ^ n8039 ^ n7368 ;
  assign n54756 = n54755 ^ n18260 ^ 1'b0 ;
  assign n54757 = ( n4984 & n8503 ) | ( n4984 & ~n9237 ) | ( n8503 & ~n9237 ) ;
  assign n54758 = ( n578 & n42955 ) | ( n578 & n54757 ) | ( n42955 & n54757 ) ;
  assign n54759 = n42025 ^ n15110 ^ n12241 ;
  assign n54760 = ( n5679 & n9871 ) | ( n5679 & ~n14468 ) | ( n9871 & ~n14468 ) ;
  assign n54761 = ( n11821 & n14628 ) | ( n11821 & n54760 ) | ( n14628 & n54760 ) ;
  assign n54762 = n54761 ^ n16106 ^ n7314 ;
  assign n54763 = n54762 ^ n30174 ^ n25848 ;
  assign n54767 = ( n1372 & n5841 ) | ( n1372 & n27136 ) | ( n5841 & n27136 ) ;
  assign n54768 = n54767 ^ n41057 ^ 1'b0 ;
  assign n54766 = n17960 & n42131 ;
  assign n54769 = n54768 ^ n54766 ^ 1'b0 ;
  assign n54764 = n26109 & n37322 ;
  assign n54765 = n54764 ^ n5686 ^ 1'b0 ;
  assign n54770 = n54769 ^ n54765 ^ n32066 ;
  assign n54771 = n8450 & ~n27673 ;
  assign n54772 = ~n51546 & n54771 ;
  assign n54773 = n10109 | n28105 ;
  assign n54774 = n28105 & ~n54773 ;
  assign n54775 = n6189 | n54774 ;
  assign n54776 = ( n1274 & ~n13960 ) | ( n1274 & n32434 ) | ( ~n13960 & n32434 ) ;
  assign n54777 = ( n10560 & ~n54775 ) | ( n10560 & n54776 ) | ( ~n54775 & n54776 ) ;
  assign n54778 = n9018 & ~n54777 ;
  assign n54779 = ~n2366 & n54778 ;
  assign n54780 = n30728 ^ n8677 ^ n794 ;
  assign n54781 = n9749 & n54780 ;
  assign n54782 = ~n31688 & n54781 ;
  assign n54783 = n3673 ^ n912 ^ 1'b0 ;
  assign n54784 = n1142 & ~n54783 ;
  assign n54785 = n54784 ^ n21264 ^ n8679 ;
  assign n54786 = n27854 & ~n54785 ;
  assign n54787 = ( n497 & n36713 ) | ( n497 & n38298 ) | ( n36713 & n38298 ) ;
  assign n54788 = ( n833 & ~n9670 ) | ( n833 & n14907 ) | ( ~n9670 & n14907 ) ;
  assign n54789 = ~n6364 & n54788 ;
  assign n54793 = n10002 | n43436 ;
  assign n54794 = n10638 & ~n54793 ;
  assign n54795 = x172 & ~n44087 ;
  assign n54796 = n54794 & n54795 ;
  assign n54790 = n16251 ^ n15994 ^ n622 ;
  assign n54791 = n33703 ^ n11453 ^ 1'b0 ;
  assign n54792 = n54790 & ~n54791 ;
  assign n54797 = n54796 ^ n54792 ^ n45413 ;
  assign n54798 = ( n3212 & n9320 ) | ( n3212 & n31782 ) | ( n9320 & n31782 ) ;
  assign n54799 = n54798 ^ n24351 ^ n9982 ;
  assign n54800 = n54799 ^ n22735 ^ n8828 ;
  assign n54801 = n39716 ^ n18103 ^ n17346 ;
  assign n54803 = n24699 ^ n24607 ^ n20477 ;
  assign n54802 = n34413 ^ n29803 ^ 1'b0 ;
  assign n54804 = n54803 ^ n54802 ^ n16585 ;
  assign n54805 = n30254 ^ n30019 ^ 1'b0 ;
  assign n54806 = n54805 ^ n53052 ^ n36040 ;
  assign n54807 = n42523 | n49816 ;
  assign n54808 = n21767 | n26699 ;
  assign n54809 = n2699 & ~n5430 ;
  assign n54810 = n54809 ^ n19493 ^ 1'b0 ;
  assign n54811 = n46079 ^ n39092 ^ n16791 ;
  assign n54812 = ( n6182 & n10219 ) | ( n6182 & n12400 ) | ( n10219 & n12400 ) ;
  assign n54813 = n34122 ^ n11607 ^ n10719 ;
  assign n54814 = ( n14384 & n54812 ) | ( n14384 & n54813 ) | ( n54812 & n54813 ) ;
  assign n54815 = n4176 & n36583 ;
  assign n54816 = n54815 ^ n46033 ^ n11967 ;
  assign n54817 = n38827 ^ n10267 ^ n7290 ;
  assign n54818 = n38990 ^ n3274 ^ 1'b0 ;
  assign n54819 = n29494 & ~n54818 ;
  assign n54820 = n54819 ^ n24898 ^ n4101 ;
  assign n54821 = n20127 ^ n1546 ^ 1'b0 ;
  assign n54822 = ( n11423 & ~n21329 ) | ( n11423 & n26680 ) | ( ~n21329 & n26680 ) ;
  assign n54823 = n1830 | n2559 ;
  assign n54824 = n4102 & ~n54823 ;
  assign n54825 = n30059 ^ n20133 ^ 1'b0 ;
  assign n54826 = n12777 & n50943 ;
  assign n54827 = ( n1423 & n3787 ) | ( n1423 & ~n52301 ) | ( n3787 & ~n52301 ) ;
  assign n54828 = n54827 ^ n31415 ^ n24310 ;
  assign n54829 = n12831 & ~n27669 ;
  assign n54830 = n54829 ^ n34916 ^ 1'b0 ;
  assign n54831 = ( ~n2978 & n31903 ) | ( ~n2978 & n54830 ) | ( n31903 & n54830 ) ;
  assign n54832 = n54831 ^ n4865 ^ 1'b0 ;
  assign n54833 = n21262 ^ n18095 ^ n14097 ;
  assign n54834 = n54833 ^ n15213 ^ n7429 ;
  assign n54835 = n33259 ^ n10562 ^ n8907 ;
  assign n54836 = n43509 ^ n6788 ^ 1'b0 ;
  assign n54837 = ( n11894 & ~n40856 ) | ( n11894 & n54836 ) | ( ~n40856 & n54836 ) ;
  assign n54838 = n18234 ^ n12040 ^ 1'b0 ;
  assign n54839 = n54838 ^ n32570 ^ 1'b0 ;
  assign n54840 = n34358 ^ n28151 ^ n27496 ;
  assign n54841 = ( n372 & ~n21656 ) | ( n372 & n54840 ) | ( ~n21656 & n54840 ) ;
  assign n54842 = ( n2804 & n16413 ) | ( n2804 & ~n54841 ) | ( n16413 & ~n54841 ) ;
  assign n54843 = ( n10276 & n38773 ) | ( n10276 & ~n54842 ) | ( n38773 & ~n54842 ) ;
  assign n54847 = ( n6039 & n11210 ) | ( n6039 & n36936 ) | ( n11210 & n36936 ) ;
  assign n54848 = n54847 ^ n6533 ^ 1'b0 ;
  assign n54844 = n7689 ^ n1152 ^ 1'b0 ;
  assign n54845 = ~n19233 & n54844 ;
  assign n54846 = ~n4012 & n54845 ;
  assign n54849 = n54848 ^ n54846 ^ 1'b0 ;
  assign n54850 = ( ~n333 & n3853 ) | ( ~n333 & n42743 ) | ( n3853 & n42743 ) ;
  assign n54851 = ( n2162 & ~n37486 ) | ( n2162 & n54850 ) | ( ~n37486 & n54850 ) ;
  assign n54852 = n54851 ^ n41390 ^ n23630 ;
  assign n54853 = n7654 & n54032 ;
  assign n54854 = ~n54852 & n54853 ;
  assign n54855 = ~n12983 & n18765 ;
  assign n54856 = n6724 & n54855 ;
  assign n54857 = n17211 | n54856 ;
  assign n54858 = n9392 | n54857 ;
  assign n54859 = n11151 & ~n26535 ;
  assign n54860 = n2428 | n28558 ;
  assign n54861 = n54860 ^ n53097 ^ 1'b0 ;
  assign n54862 = ( ~n28505 & n54859 ) | ( ~n28505 & n54861 ) | ( n54859 & n54861 ) ;
  assign n54863 = n9890 ^ n1714 ^ 1'b0 ;
  assign n54864 = n13789 & ~n33263 ;
  assign n54866 = n17218 & ~n26307 ;
  assign n54867 = ~n18752 & n54866 ;
  assign n54865 = ( ~n8004 & n29993 ) | ( ~n8004 & n34884 ) | ( n29993 & n34884 ) ;
  assign n54868 = n54867 ^ n54865 ^ n24763 ;
  assign n54869 = ( n334 & n1656 ) | ( n334 & ~n47621 ) | ( n1656 & ~n47621 ) ;
  assign n54870 = ( n5918 & n22708 ) | ( n5918 & n28521 ) | ( n22708 & n28521 ) ;
  assign n54871 = ( ~n11612 & n36182 ) | ( ~n11612 & n54870 ) | ( n36182 & n54870 ) ;
  assign n54872 = n48897 ^ n45409 ^ 1'b0 ;
  assign n54873 = ~n17845 & n54872 ;
  assign n54874 = n52520 ^ n17463 ^ 1'b0 ;
  assign n54875 = ( n37406 & ~n54873 ) | ( n37406 & n54874 ) | ( ~n54873 & n54874 ) ;
  assign n54876 = n33983 | n49491 ;
  assign n54877 = n54876 ^ n5759 ^ 1'b0 ;
  assign n54878 = n10554 | n18681 ;
  assign n54879 = n54878 ^ n32659 ^ 1'b0 ;
  assign n54880 = ( ~n1200 & n26059 ) | ( ~n1200 & n37861 ) | ( n26059 & n37861 ) ;
  assign n54881 = n2868 & n54880 ;
  assign n54882 = ~n1426 & n4100 ;
  assign n54884 = n19853 ^ n14203 ^ 1'b0 ;
  assign n54883 = n13567 ^ n11653 ^ n8798 ;
  assign n54885 = n54884 ^ n54883 ^ n3110 ;
  assign n54886 = ( ~n15203 & n45769 ) | ( ~n15203 & n46691 ) | ( n45769 & n46691 ) ;
  assign n54887 = ( ~n9200 & n13186 ) | ( ~n9200 & n23607 ) | ( n13186 & n23607 ) ;
  assign n54888 = ( n33590 & n33708 ) | ( n33590 & n53763 ) | ( n33708 & n53763 ) ;
  assign n54889 = n5742 | n16268 ;
  assign n54890 = ( n3566 & n21741 ) | ( n3566 & n54889 ) | ( n21741 & n54889 ) ;
  assign n54891 = n11340 & n49913 ;
  assign n54892 = n54891 ^ n6119 ^ 1'b0 ;
  assign n54893 = n44159 ^ x93 ^ 1'b0 ;
  assign n54894 = n40708 & n54893 ;
  assign n54895 = n42812 ^ n42520 ^ n33236 ;
  assign n54896 = n31948 ^ n14644 ^ n7939 ;
  assign n54897 = n54896 ^ n39153 ^ 1'b0 ;
  assign n54898 = n46789 ^ n9650 ^ n8711 ;
  assign n54899 = n44437 ^ n43469 ^ n32676 ;
  assign n54900 = n27940 ^ n18664 ^ 1'b0 ;
  assign n54901 = ~n25085 & n40611 ;
  assign n54902 = n35717 & n54901 ;
  assign n54903 = ( ~n10950 & n35183 ) | ( ~n10950 & n54902 ) | ( n35183 & n54902 ) ;
  assign n54904 = ( n6376 & ~n20515 ) | ( n6376 & n54903 ) | ( ~n20515 & n54903 ) ;
  assign n54905 = n8869 & ~n24258 ;
  assign n54906 = n54905 ^ n46930 ^ 1'b0 ;
  assign n54907 = n3160 | n15241 ;
  assign n54908 = n54906 & ~n54907 ;
  assign n54909 = ( n7367 & ~n22745 ) | ( n7367 & n54908 ) | ( ~n22745 & n54908 ) ;
  assign n54910 = n5782 & ~n30984 ;
  assign n54911 = n54910 ^ n21338 ^ n10763 ;
  assign n54912 = n51791 ^ n41736 ^ n8269 ;
  assign n54913 = n54912 ^ n16250 ^ 1'b0 ;
  assign n54914 = n54913 ^ n48989 ^ n26669 ;
  assign n54915 = ~n54911 & n54914 ;
  assign n54916 = ~n9686 & n41247 ;
  assign n54917 = n39938 & n54916 ;
  assign n54918 = n544 | n30364 ;
  assign n54919 = n54918 ^ n22767 ^ 1'b0 ;
  assign n54920 = n18287 | n34621 ;
  assign n54921 = ( n3580 & n10917 ) | ( n3580 & ~n54920 ) | ( n10917 & ~n54920 ) ;
  assign n54922 = ~n18681 & n54921 ;
  assign n54923 = ( ~n2890 & n3300 ) | ( ~n2890 & n54922 ) | ( n3300 & n54922 ) ;
  assign n54924 = n20444 | n28917 ;
  assign n54925 = n54924 ^ n10109 ^ 1'b0 ;
  assign n54926 = n24947 & ~n54925 ;
  assign n54927 = n54926 ^ n25432 ^ 1'b0 ;
  assign n54928 = ( ~n25222 & n41378 ) | ( ~n25222 & n54927 ) | ( n41378 & n54927 ) ;
  assign n54929 = n54928 ^ n30445 ^ 1'b0 ;
  assign n54930 = n43607 ^ n43210 ^ n3919 ;
  assign n54932 = ~n8907 & n28505 ;
  assign n54933 = n2315 & n54932 ;
  assign n54931 = n45295 ^ n41020 ^ n6797 ;
  assign n54934 = n54933 ^ n54931 ^ n47717 ;
  assign n54935 = n9612 & n44334 ;
  assign n54936 = n54935 ^ n32193 ^ 1'b0 ;
  assign n54937 = n54936 ^ n49600 ^ n10475 ;
  assign n54938 = n26228 ^ n8094 ^ n7666 ;
  assign n54939 = n54938 ^ n15425 ^ 1'b0 ;
  assign n54940 = n48391 ^ n25954 ^ n7398 ;
  assign n54941 = n32445 ^ n7440 ^ 1'b0 ;
  assign n54942 = ( ~n4910 & n25485 ) | ( ~n4910 & n54941 ) | ( n25485 & n54941 ) ;
  assign n54943 = n54942 ^ n35185 ^ n2379 ;
  assign n54944 = ( ~n23472 & n46584 ) | ( ~n23472 & n54943 ) | ( n46584 & n54943 ) ;
  assign n54945 = ( n32085 & ~n54940 ) | ( n32085 & n54944 ) | ( ~n54940 & n54944 ) ;
  assign n54946 = n38124 ^ n13436 ^ 1'b0 ;
  assign n54947 = n39585 ^ n21592 ^ n3860 ;
  assign n54948 = n22472 ^ n5202 ^ 1'b0 ;
  assign n54949 = ~n54947 & n54948 ;
  assign n54950 = n3407 & n20341 ;
  assign n54951 = n54950 ^ n14001 ^ 1'b0 ;
  assign n54952 = n42365 ^ n8352 ^ 1'b0 ;
  assign n54953 = n36041 ^ n15950 ^ 1'b0 ;
  assign n54954 = n34256 ^ n22388 ^ 1'b0 ;
  assign n54955 = n12216 & ~n54954 ;
  assign n54956 = ( n32099 & n45374 ) | ( n32099 & n54955 ) | ( n45374 & n54955 ) ;
  assign n54957 = ( n1844 & ~n3483 ) | ( n1844 & n41583 ) | ( ~n3483 & n41583 ) ;
  assign n54958 = n30424 | n46512 ;
  assign n54959 = n54957 | n54958 ;
  assign n54960 = n4805 & n54959 ;
  assign n54961 = ( ~n10150 & n46910 ) | ( ~n10150 & n54960 ) | ( n46910 & n54960 ) ;
  assign n54964 = n1867 & n6883 ;
  assign n54965 = n54964 ^ n21367 ^ 1'b0 ;
  assign n54966 = n54965 ^ n24984 ^ n14344 ;
  assign n54963 = n10312 ^ n9701 ^ n341 ;
  assign n54967 = n54966 ^ n54963 ^ n49874 ;
  assign n54962 = ( ~n12280 & n15407 ) | ( ~n12280 & n25970 ) | ( n15407 & n25970 ) ;
  assign n54968 = n54967 ^ n54962 ^ 1'b0 ;
  assign n54970 = n16762 & n36081 ;
  assign n54971 = n54970 ^ n10755 ^ n8688 ;
  assign n54969 = ( n1524 & n39366 ) | ( n1524 & n50871 ) | ( n39366 & n50871 ) ;
  assign n54972 = n54971 ^ n54969 ^ n23881 ;
  assign n54973 = n42351 ^ n6965 ^ 1'b0 ;
  assign n54974 = n23952 | n54973 ;
  assign n54975 = n4015 ^ n3761 ^ n2402 ;
  assign n54976 = n8039 & n54975 ;
  assign n54977 = n54974 & n54976 ;
  assign n54978 = n23595 ^ n20378 ^ 1'b0 ;
  assign n54979 = n367 & n54978 ;
  assign n54980 = n16551 ^ n11792 ^ n8962 ;
  assign n54981 = ~n24607 & n54980 ;
  assign n54982 = n54981 ^ n12227 ^ 1'b0 ;
  assign n54983 = n54982 ^ n36981 ^ n21610 ;
  assign n54984 = n33849 ^ n19781 ^ n13914 ;
  assign n54985 = ( n20189 & n54983 ) | ( n20189 & ~n54984 ) | ( n54983 & ~n54984 ) ;
  assign n54986 = ( n16717 & n34382 ) | ( n16717 & n50889 ) | ( n34382 & n50889 ) ;
  assign n54987 = n54986 ^ n40878 ^ n8668 ;
  assign n54988 = ( n9911 & n16421 ) | ( n9911 & ~n24895 ) | ( n16421 & ~n24895 ) ;
  assign n54989 = ( ~n14051 & n16989 ) | ( ~n14051 & n24608 ) | ( n16989 & n24608 ) ;
  assign n54990 = n54989 ^ n45247 ^ 1'b0 ;
  assign n54991 = n36325 ^ n11317 ^ 1'b0 ;
  assign n54992 = ( n24076 & n25402 ) | ( n24076 & ~n54991 ) | ( n25402 & ~n54991 ) ;
  assign n54993 = n6255 ^ n2893 ^ 1'b0 ;
  assign n54994 = n3730 & ~n54993 ;
  assign n54995 = ( n38773 & n39513 ) | ( n38773 & n54994 ) | ( n39513 & n54994 ) ;
  assign n54996 = n6465 & ~n8955 ;
  assign n54997 = ( n6187 & n29204 ) | ( n6187 & n54996 ) | ( n29204 & n54996 ) ;
  assign n54998 = n39928 & n54997 ;
  assign n54999 = n54998 ^ n18155 ^ 1'b0 ;
  assign n55000 = ( n2427 & n6463 ) | ( n2427 & n41969 ) | ( n6463 & n41969 ) ;
  assign n55001 = ( n2248 & n20595 ) | ( n2248 & ~n55000 ) | ( n20595 & ~n55000 ) ;
  assign n55002 = n3469 | n55001 ;
  assign n55003 = n6871 | n55002 ;
  assign n55004 = n41301 ^ n29140 ^ n27117 ;
  assign n55005 = n55004 ^ n44737 ^ n30049 ;
  assign n55006 = n55005 ^ n47772 ^ 1'b0 ;
  assign n55007 = n30092 | n35464 ;
  assign n55008 = n22870 & ~n55007 ;
  assign n55009 = n17521 | n27830 ;
  assign n55010 = n14643 & ~n55009 ;
  assign n55011 = ( n15773 & ~n16557 ) | ( n15773 & n55010 ) | ( ~n16557 & n55010 ) ;
  assign n55012 = ( ~n21700 & n24484 ) | ( ~n21700 & n28666 ) | ( n24484 & n28666 ) ;
  assign n55013 = n5872 & ~n55012 ;
  assign n55014 = n48713 ^ n26497 ^ n9725 ;
  assign n55015 = ( n35197 & ~n43098 ) | ( n35197 & n55014 ) | ( ~n43098 & n55014 ) ;
  assign n55016 = n36132 ^ n27771 ^ n6896 ;
  assign n55017 = ~n4599 & n12577 ;
  assign n55018 = ( n2070 & n36140 ) | ( n2070 & n46827 ) | ( n36140 & n46827 ) ;
  assign n55019 = n15494 ^ n10306 ^ 1'b0 ;
  assign n55020 = n6246 & ~n31247 ;
  assign n55021 = n43023 & n55020 ;
  assign n55022 = ~n25860 & n50648 ;
  assign n55023 = ~n47957 & n55022 ;
  assign n55027 = ( n6545 & n39439 ) | ( n6545 & ~n46438 ) | ( n39439 & ~n46438 ) ;
  assign n55024 = n42223 ^ n29850 ^ 1'b0 ;
  assign n55025 = n29911 & ~n55024 ;
  assign n55026 = ~n29986 & n55025 ;
  assign n55028 = n55027 ^ n55026 ^ 1'b0 ;
  assign n55029 = ~n14527 & n17793 ;
  assign n55030 = n52366 ^ n29481 ^ n20399 ;
  assign n55031 = n835 | n5450 ;
  assign n55032 = n55031 ^ n20798 ^ n10254 ;
  assign n55033 = ( ~n5175 & n8099 ) | ( ~n5175 & n48818 ) | ( n8099 & n48818 ) ;
  assign n55034 = ( n13876 & ~n20690 ) | ( n13876 & n41952 ) | ( ~n20690 & n41952 ) ;
  assign n55035 = ( ~n7227 & n32641 ) | ( ~n7227 & n55034 ) | ( n32641 & n55034 ) ;
  assign n55036 = n49037 ^ n497 ^ 1'b0 ;
  assign n55037 = n34512 ^ n33553 ^ n2859 ;
  assign n55038 = n54790 & ~n55037 ;
  assign n55039 = n28496 ^ n27356 ^ n27226 ;
  assign n55040 = ~n14782 & n17486 ;
  assign n55041 = n55040 ^ n51289 ^ 1'b0 ;
  assign y0 = x37 ;
  assign y1 = x41 ;
  assign y2 = x64 ;
  assign y3 = x71 ;
  assign y4 = x86 ;
  assign y5 = x87 ;
  assign y6 = x89 ;
  assign y7 = x93 ;
  assign y8 = x96 ;
  assign y9 = x116 ;
  assign y10 = x120 ;
  assign y11 = x127 ;
  assign y12 = x128 ;
  assign y13 = x133 ;
  assign y14 = x141 ;
  assign y15 = x142 ;
  assign y16 = x144 ;
  assign y17 = x158 ;
  assign y18 = x172 ;
  assign y19 = x174 ;
  assign y20 = x177 ;
  assign y21 = x182 ;
  assign y22 = x184 ;
  assign y23 = x186 ;
  assign y24 = x189 ;
  assign y25 = x200 ;
  assign y26 = x208 ;
  assign y27 = x213 ;
  assign y28 = x214 ;
  assign y29 = x230 ;
  assign y30 = x236 ;
  assign y31 = x239 ;
  assign y32 = x240 ;
  assign y33 = x241 ;
  assign y34 = n257 ;
  assign y35 = ~n259 ;
  assign y36 = ~n261 ;
  assign y37 = n263 ;
  assign y38 = ~n266 ;
  assign y39 = ~n268 ;
  assign y40 = ~1'b0 ;
  assign y41 = n269 ;
  assign y42 = ~1'b0 ;
  assign y43 = ~n270 ;
  assign y44 = ~n273 ;
  assign y45 = ~1'b0 ;
  assign y46 = n279 ;
  assign y47 = n284 ;
  assign y48 = n286 ;
  assign y49 = n287 ;
  assign y50 = ~1'b0 ;
  assign y51 = ~n290 ;
  assign y52 = ~n293 ;
  assign y53 = ~n295 ;
  assign y54 = n301 ;
  assign y55 = ~n304 ;
  assign y56 = ~n308 ;
  assign y57 = n315 ;
  assign y58 = n320 ;
  assign y59 = ~n323 ;
  assign y60 = ~1'b0 ;
  assign y61 = n324 ;
  assign y62 = n328 ;
  assign y63 = ~1'b0 ;
  assign y64 = ~n329 ;
  assign y65 = n331 ;
  assign y66 = n332 ;
  assign y67 = ~n342 ;
  assign y68 = ~n343 ;
  assign y69 = n350 ;
  assign y70 = ~n352 ;
  assign y71 = n356 ;
  assign y72 = n357 ;
  assign y73 = n360 ;
  assign y74 = ~n363 ;
  assign y75 = ~n365 ;
  assign y76 = ~n369 ;
  assign y77 = n373 ;
  assign y78 = ~n376 ;
  assign y79 = n378 ;
  assign y80 = n381 ;
  assign y81 = ~n391 ;
  assign y82 = n396 ;
  assign y83 = ~n397 ;
  assign y84 = n398 ;
  assign y85 = ~n400 ;
  assign y86 = n404 ;
  assign y87 = ~n409 ;
  assign y88 = ~n415 ;
  assign y89 = ~n419 ;
  assign y90 = n424 ;
  assign y91 = ~n430 ;
  assign y92 = ~n431 ;
  assign y93 = ~n434 ;
  assign y94 = n440 ;
  assign y95 = ~1'b0 ;
  assign y96 = ~n441 ;
  assign y97 = ~n452 ;
  assign y98 = ~n453 ;
  assign y99 = ~n455 ;
  assign y100 = n458 ;
  assign y101 = n460 ;
  assign y102 = n461 ;
  assign y103 = ~n463 ;
  assign y104 = ~1'b0 ;
  assign y105 = 1'b0 ;
  assign y106 = ~n474 ;
  assign y107 = ~1'b0 ;
  assign y108 = n480 ;
  assign y109 = n482 ;
  assign y110 = ~n486 ;
  assign y111 = n490 ;
  assign y112 = n492 ;
  assign y113 = ~n495 ;
  assign y114 = n511 ;
  assign y115 = ~n527 ;
  assign y116 = n531 ;
  assign y117 = ~n535 ;
  assign y118 = ~n538 ;
  assign y119 = n540 ;
  assign y120 = n541 ;
  assign y121 = n546 ;
  assign y122 = n547 ;
  assign y123 = ~n549 ;
  assign y124 = ~n550 ;
  assign y125 = n555 ;
  assign y126 = n559 ;
  assign y127 = n560 ;
  assign y128 = ~n561 ;
  assign y129 = n563 ;
  assign y130 = ~1'b0 ;
  assign y131 = ~n570 ;
  assign y132 = n574 ;
  assign y133 = n585 ;
  assign y134 = n597 ;
  assign y135 = ~n604 ;
  assign y136 = n605 ;
  assign y137 = ~n612 ;
  assign y138 = ~1'b0 ;
  assign y139 = ~1'b0 ;
  assign y140 = ~n620 ;
  assign y141 = ~n621 ;
  assign y142 = ~n633 ;
  assign y143 = n634 ;
  assign y144 = ~x67 ;
  assign y145 = n643 ;
  assign y146 = ~n648 ;
  assign y147 = n653 ;
  assign y148 = ~n658 ;
  assign y149 = n661 ;
  assign y150 = ~n662 ;
  assign y151 = n669 ;
  assign y152 = ~n670 ;
  assign y153 = ~n672 ;
  assign y154 = n677 ;
  assign y155 = n681 ;
  assign y156 = n690 ;
  assign y157 = n692 ;
  assign y158 = n694 ;
  assign y159 = n704 ;
  assign y160 = n708 ;
  assign y161 = n735 ;
  assign y162 = ~1'b0 ;
  assign y163 = n745 ;
  assign y164 = ~n748 ;
  assign y165 = n751 ;
  assign y166 = ~n757 ;
  assign y167 = ~n764 ;
  assign y168 = ~n770 ;
  assign y169 = ~n773 ;
  assign y170 = ~n777 ;
  assign y171 = n783 ;
  assign y172 = n784 ;
  assign y173 = ~n786 ;
  assign y174 = ~n790 ;
  assign y175 = ~n791 ;
  assign y176 = n798 ;
  assign y177 = ~n802 ;
  assign y178 = ~1'b0 ;
  assign y179 = n803 ;
  assign y180 = ~1'b0 ;
  assign y181 = ~1'b0 ;
  assign y182 = n807 ;
  assign y183 = ~n811 ;
  assign y184 = n818 ;
  assign y185 = n820 ;
  assign y186 = ~n821 ;
  assign y187 = ~n822 ;
  assign y188 = ~n829 ;
  assign y189 = ~1'b0 ;
  assign y190 = n838 ;
  assign y191 = ~n850 ;
  assign y192 = n865 ;
  assign y193 = ~n869 ;
  assign y194 = ~1'b0 ;
  assign y195 = n870 ;
  assign y196 = ~n876 ;
  assign y197 = n886 ;
  assign y198 = ~n887 ;
  assign y199 = n890 ;
  assign y200 = ~n892 ;
  assign y201 = ~1'b0 ;
  assign y202 = n896 ;
  assign y203 = n897 ;
  assign y204 = ~n905 ;
  assign y205 = x212 ;
  assign y206 = ~n909 ;
  assign y207 = n913 ;
  assign y208 = ~n916 ;
  assign y209 = ~n920 ;
  assign y210 = n921 ;
  assign y211 = n925 ;
  assign y212 = ~n929 ;
  assign y213 = ~n930 ;
  assign y214 = ~n932 ;
  assign y215 = ~1'b0 ;
  assign y216 = n936 ;
  assign y217 = ~n939 ;
  assign y218 = ~n942 ;
  assign y219 = ~n945 ;
  assign y220 = n959 ;
  assign y221 = ~n963 ;
  assign y222 = ~n968 ;
  assign y223 = n970 ;
  assign y224 = n974 ;
  assign y225 = ~n979 ;
  assign y226 = n1007 ;
  assign y227 = ~n1009 ;
  assign y228 = ~1'b0 ;
  assign y229 = n1014 ;
  assign y230 = ~1'b0 ;
  assign y231 = n1018 ;
  assign y232 = ~n1022 ;
  assign y233 = ~n1026 ;
  assign y234 = n1029 ;
  assign y235 = ~n1032 ;
  assign y236 = ~n1033 ;
  assign y237 = n1034 ;
  assign y238 = ~n1039 ;
  assign y239 = n1047 ;
  assign y240 = ~n1057 ;
  assign y241 = n1067 ;
  assign y242 = n1071 ;
  assign y243 = ~n1076 ;
  assign y244 = n1078 ;
  assign y245 = ~n1080 ;
  assign y246 = ~n1088 ;
  assign y247 = ~n1095 ;
  assign y248 = n1102 ;
  assign y249 = ~n1106 ;
  assign y250 = ~n1109 ;
  assign y251 = ~n1114 ;
  assign y252 = ~n1126 ;
  assign y253 = ~n1127 ;
  assign y254 = ~n1134 ;
  assign y255 = n1135 ;
  assign y256 = ~n1136 ;
  assign y257 = ~n1143 ;
  assign y258 = ~n1149 ;
  assign y259 = ~n1152 ;
  assign y260 = n1159 ;
  assign y261 = ~1'b0 ;
  assign y262 = n1164 ;
  assign y263 = n1179 ;
  assign y264 = ~n1180 ;
  assign y265 = n1182 ;
  assign y266 = ~n1194 ;
  assign y267 = ~1'b0 ;
  assign y268 = n1198 ;
  assign y269 = ~n1201 ;
  assign y270 = ~n1204 ;
  assign y271 = n1206 ;
  assign y272 = n1208 ;
  assign y273 = ~n1214 ;
  assign y274 = n1219 ;
  assign y275 = ~1'b0 ;
  assign y276 = ~n1227 ;
  assign y277 = ~1'b0 ;
  assign y278 = n1230 ;
  assign y279 = n1233 ;
  assign y280 = n1241 ;
  assign y281 = n1245 ;
  assign y282 = n1247 ;
  assign y283 = n1256 ;
  assign y284 = ~n1264 ;
  assign y285 = n1265 ;
  assign y286 = ~1'b0 ;
  assign y287 = ~n1268 ;
  assign y288 = ~n1272 ;
  assign y289 = n1279 ;
  assign y290 = ~1'b0 ;
  assign y291 = ~n1290 ;
  assign y292 = n1291 ;
  assign y293 = n1297 ;
  assign y294 = n1316 ;
  assign y295 = n1321 ;
  assign y296 = ~n1322 ;
  assign y297 = n1323 ;
  assign y298 = ~n1339 ;
  assign y299 = n1352 ;
  assign y300 = n1357 ;
  assign y301 = ~1'b0 ;
  assign y302 = n1359 ;
  assign y303 = ~n1362 ;
  assign y304 = n1367 ;
  assign y305 = ~n1369 ;
  assign y306 = n1376 ;
  assign y307 = ~n1379 ;
  assign y308 = ~n1389 ;
  assign y309 = ~n1390 ;
  assign y310 = ~n501 ;
  assign y311 = n1401 ;
  assign y312 = ~n1404 ;
  assign y313 = ~n1409 ;
  assign y314 = n1418 ;
  assign y315 = ~n1424 ;
  assign y316 = n1425 ;
  assign y317 = n1428 ;
  assign y318 = ~n1433 ;
  assign y319 = n1434 ;
  assign y320 = ~n1440 ;
  assign y321 = n1442 ;
  assign y322 = n1455 ;
  assign y323 = ~1'b0 ;
  assign y324 = n1463 ;
  assign y325 = n1465 ;
  assign y326 = ~n1472 ;
  assign y327 = ~n1474 ;
  assign y328 = n1476 ;
  assign y329 = n1480 ;
  assign y330 = ~n1482 ;
  assign y331 = ~n1487 ;
  assign y332 = ~n1492 ;
  assign y333 = n1498 ;
  assign y334 = ~1'b0 ;
  assign y335 = ~1'b0 ;
  assign y336 = n1511 ;
  assign y337 = ~1'b0 ;
  assign y338 = n1514 ;
  assign y339 = ~n1517 ;
  assign y340 = n1519 ;
  assign y341 = n1529 ;
  assign y342 = ~n1550 ;
  assign y343 = ~n1556 ;
  assign y344 = n1560 ;
  assign y345 = ~n1571 ;
  assign y346 = n1572 ;
  assign y347 = ~n1575 ;
  assign y348 = n1577 ;
  assign y349 = n1581 ;
  assign y350 = n1588 ;
  assign y351 = ~1'b0 ;
  assign y352 = n1594 ;
  assign y353 = ~n1595 ;
  assign y354 = ~n1598 ;
  assign y355 = n1602 ;
  assign y356 = n1605 ;
  assign y357 = ~n1610 ;
  assign y358 = n1611 ;
  assign y359 = ~n1625 ;
  assign y360 = ~n1631 ;
  assign y361 = ~n1638 ;
  assign y362 = ~n1651 ;
  assign y363 = n1659 ;
  assign y364 = ~n1664 ;
  assign y365 = n1672 ;
  assign y366 = n1673 ;
  assign y367 = ~1'b0 ;
  assign y368 = n1680 ;
  assign y369 = ~n1681 ;
  assign y370 = ~n1695 ;
  assign y371 = ~n1700 ;
  assign y372 = ~n1706 ;
  assign y373 = n1708 ;
  assign y374 = n1711 ;
  assign y375 = n1713 ;
  assign y376 = ~n1716 ;
  assign y377 = n1717 ;
  assign y378 = n1737 ;
  assign y379 = n1741 ;
  assign y380 = ~n1743 ;
  assign y381 = ~1'b0 ;
  assign y382 = ~n1746 ;
  assign y383 = ~n1748 ;
  assign y384 = ~1'b0 ;
  assign y385 = n1752 ;
  assign y386 = n1753 ;
  assign y387 = ~n1764 ;
  assign y388 = n1773 ;
  assign y389 = n1776 ;
  assign y390 = ~n1777 ;
  assign y391 = n1780 ;
  assign y392 = ~n1789 ;
  assign y393 = n1790 ;
  assign y394 = ~n1803 ;
  assign y395 = n1804 ;
  assign y396 = ~n1807 ;
  assign y397 = ~n1811 ;
  assign y398 = n1820 ;
  assign y399 = n1823 ;
  assign y400 = n1827 ;
  assign y401 = ~n1830 ;
  assign y402 = ~n1833 ;
  assign y403 = n1835 ;
  assign y404 = n1840 ;
  assign y405 = ~1'b0 ;
  assign y406 = ~n1844 ;
  assign y407 = n1846 ;
  assign y408 = n1863 ;
  assign y409 = n1882 ;
  assign y410 = ~n1892 ;
  assign y411 = ~n1905 ;
  assign y412 = ~1'b0 ;
  assign y413 = ~n1910 ;
  assign y414 = n1934 ;
  assign y415 = ~n1935 ;
  assign y416 = n1938 ;
  assign y417 = ~n1950 ;
  assign y418 = n1954 ;
  assign y419 = ~n1956 ;
  assign y420 = n1977 ;
  assign y421 = ~n1996 ;
  assign y422 = n1998 ;
  assign y423 = ~n1999 ;
  assign y424 = ~n2005 ;
  assign y425 = ~n2008 ;
  assign y426 = ~n2009 ;
  assign y427 = ~n2015 ;
  assign y428 = ~n2019 ;
  assign y429 = ~1'b0 ;
  assign y430 = n2020 ;
  assign y431 = n2024 ;
  assign y432 = n2025 ;
  assign y433 = ~n2027 ;
  assign y434 = n2028 ;
  assign y435 = n2031 ;
  assign y436 = n2042 ;
  assign y437 = ~n2044 ;
  assign y438 = n2046 ;
  assign y439 = n2047 ;
  assign y440 = ~n2069 ;
  assign y441 = n2070 ;
  assign y442 = n2074 ;
  assign y443 = n2078 ;
  assign y444 = ~n2082 ;
  assign y445 = ~n2083 ;
  assign y446 = ~n2088 ;
  assign y447 = ~n2091 ;
  assign y448 = ~n2099 ;
  assign y449 = n2100 ;
  assign y450 = ~n2107 ;
  assign y451 = n2111 ;
  assign y452 = ~n2116 ;
  assign y453 = n2118 ;
  assign y454 = n2142 ;
  assign y455 = ~n2157 ;
  assign y456 = n2158 ;
  assign y457 = n2176 ;
  assign y458 = ~n2187 ;
  assign y459 = n2188 ;
  assign y460 = ~1'b0 ;
  assign y461 = ~n2194 ;
  assign y462 = ~n2206 ;
  assign y463 = ~n2208 ;
  assign y464 = ~1'b0 ;
  assign y465 = n2221 ;
  assign y466 = ~1'b0 ;
  assign y467 = ~n2222 ;
  assign y468 = ~1'b0 ;
  assign y469 = n2226 ;
  assign y470 = n2230 ;
  assign y471 = n2231 ;
  assign y472 = n2233 ;
  assign y473 = ~n2234 ;
  assign y474 = ~n2241 ;
  assign y475 = ~n2244 ;
  assign y476 = n2251 ;
  assign y477 = ~n2252 ;
  assign y478 = n2258 ;
  assign y479 = n2266 ;
  assign y480 = ~n2271 ;
  assign y481 = n2280 ;
  assign y482 = ~n2290 ;
  assign y483 = ~n2295 ;
  assign y484 = ~1'b0 ;
  assign y485 = n2301 ;
  assign y486 = n2302 ;
  assign y487 = n2306 ;
  assign y488 = ~n2311 ;
  assign y489 = n2328 ;
  assign y490 = ~n2333 ;
  assign y491 = n2343 ;
  assign y492 = ~n2353 ;
  assign y493 = n2364 ;
  assign y494 = ~n2370 ;
  assign y495 = n2371 ;
  assign y496 = ~n2379 ;
  assign y497 = n2385 ;
  assign y498 = ~n2397 ;
  assign y499 = ~1'b0 ;
  assign y500 = ~n2424 ;
  assign y501 = ~n2427 ;
  assign y502 = ~n2428 ;
  assign y503 = n2429 ;
  assign y504 = n2430 ;
  assign y505 = n2435 ;
  assign y506 = n2444 ;
  assign y507 = n2449 ;
  assign y508 = ~1'b0 ;
  assign y509 = ~n2451 ;
  assign y510 = ~n2472 ;
  assign y511 = ~n2479 ;
  assign y512 = ~n2480 ;
  assign y513 = ~n2486 ;
  assign y514 = ~n2491 ;
  assign y515 = ~n2496 ;
  assign y516 = ~n2515 ;
  assign y517 = ~n2516 ;
  assign y518 = ~1'b0 ;
  assign y519 = ~n2523 ;
  assign y520 = ~1'b0 ;
  assign y521 = n2525 ;
  assign y522 = ~n2530 ;
  assign y523 = n2531 ;
  assign y524 = n2546 ;
  assign y525 = n2550 ;
  assign y526 = n2556 ;
  assign y527 = n2558 ;
  assign y528 = ~n2560 ;
  assign y529 = ~n2569 ;
  assign y530 = n2570 ;
  assign y531 = ~n2579 ;
  assign y532 = n2586 ;
  assign y533 = ~n2599 ;
  assign y534 = ~n2608 ;
  assign y535 = ~n2610 ;
  assign y536 = n2618 ;
  assign y537 = n2620 ;
  assign y538 = ~1'b0 ;
  assign y539 = ~1'b0 ;
  assign y540 = n2622 ;
  assign y541 = ~1'b0 ;
  assign y542 = n2624 ;
  assign y543 = n2627 ;
  assign y544 = ~n2634 ;
  assign y545 = n2648 ;
  assign y546 = ~n2649 ;
  assign y547 = n2650 ;
  assign y548 = ~n2651 ;
  assign y549 = n2657 ;
  assign y550 = n2662 ;
  assign y551 = n2664 ;
  assign y552 = n2680 ;
  assign y553 = ~n2693 ;
  assign y554 = ~1'b0 ;
  assign y555 = n2699 ;
  assign y556 = ~n2706 ;
  assign y557 = ~n2710 ;
  assign y558 = n2712 ;
  assign y559 = n2730 ;
  assign y560 = n2738 ;
  assign y561 = ~n2739 ;
  assign y562 = n2742 ;
  assign y563 = ~n2746 ;
  assign y564 = ~n2756 ;
  assign y565 = ~n2758 ;
  assign y566 = ~n2759 ;
  assign y567 = n2765 ;
  assign y568 = n2773 ;
  assign y569 = ~n2779 ;
  assign y570 = ~n2782 ;
  assign y571 = ~n2789 ;
  assign y572 = n2791 ;
  assign y573 = ~n2797 ;
  assign y574 = ~n2800 ;
  assign y575 = ~1'b0 ;
  assign y576 = n2802 ;
  assign y577 = ~1'b0 ;
  assign y578 = ~n2807 ;
  assign y579 = ~n2820 ;
  assign y580 = ~n2823 ;
  assign y581 = ~n2825 ;
  assign y582 = ~n2828 ;
  assign y583 = ~n2830 ;
  assign y584 = ~n2840 ;
  assign y585 = n2491 ;
  assign y586 = n2844 ;
  assign y587 = ~n2847 ;
  assign y588 = ~n2848 ;
  assign y589 = n2856 ;
  assign y590 = ~n2859 ;
  assign y591 = ~n2861 ;
  assign y592 = n2862 ;
  assign y593 = n2863 ;
  assign y594 = n2864 ;
  assign y595 = ~n2866 ;
  assign y596 = ~n2869 ;
  assign y597 = n2885 ;
  assign y598 = ~n2897 ;
  assign y599 = ~1'b0 ;
  assign y600 = ~n2905 ;
  assign y601 = n2924 ;
  assign y602 = ~n903 ;
  assign y603 = ~n2926 ;
  assign y604 = ~n2929 ;
  assign y605 = ~n2933 ;
  assign y606 = ~n2937 ;
  assign y607 = n2939 ;
  assign y608 = n2947 ;
  assign y609 = ~n2949 ;
  assign y610 = n2951 ;
  assign y611 = n2956 ;
  assign y612 = n2963 ;
  assign y613 = ~n2965 ;
  assign y614 = ~n2971 ;
  assign y615 = ~n2973 ;
  assign y616 = n2976 ;
  assign y617 = ~1'b0 ;
  assign y618 = ~n2977 ;
  assign y619 = ~n2978 ;
  assign y620 = ~1'b0 ;
  assign y621 = ~n2985 ;
  assign y622 = n2987 ;
  assign y623 = n2999 ;
  assign y624 = ~n3004 ;
  assign y625 = ~n1588 ;
  assign y626 = n3007 ;
  assign y627 = n3009 ;
  assign y628 = ~n3014 ;
  assign y629 = ~n3016 ;
  assign y630 = ~n3019 ;
  assign y631 = n3028 ;
  assign y632 = n3035 ;
  assign y633 = ~n3036 ;
  assign y634 = n3042 ;
  assign y635 = ~n3046 ;
  assign y636 = ~n3051 ;
  assign y637 = n3056 ;
  assign y638 = ~n3060 ;
  assign y639 = n3063 ;
  assign y640 = ~n3073 ;
  assign y641 = n3076 ;
  assign y642 = n3077 ;
  assign y643 = n3085 ;
  assign y644 = ~1'b0 ;
  assign y645 = n3089 ;
  assign y646 = n3092 ;
  assign y647 = n3098 ;
  assign y648 = n3102 ;
  assign y649 = ~1'b0 ;
  assign y650 = ~n3106 ;
  assign y651 = n3108 ;
  assign y652 = ~n3109 ;
  assign y653 = ~n3119 ;
  assign y654 = ~n3124 ;
  assign y655 = ~n3129 ;
  assign y656 = n3137 ;
  assign y657 = n3141 ;
  assign y658 = n3142 ;
  assign y659 = n3146 ;
  assign y660 = n3149 ;
  assign y661 = n3157 ;
  assign y662 = ~1'b0 ;
  assign y663 = ~n3161 ;
  assign y664 = n3162 ;
  assign y665 = n3175 ;
  assign y666 = n3176 ;
  assign y667 = ~1'b0 ;
  assign y668 = n3182 ;
  assign y669 = n3189 ;
  assign y670 = n3190 ;
  assign y671 = ~n3195 ;
  assign y672 = ~n3208 ;
  assign y673 = ~n3218 ;
  assign y674 = ~1'b0 ;
  assign y675 = n3219 ;
  assign y676 = ~n3220 ;
  assign y677 = ~n3223 ;
  assign y678 = ~n3231 ;
  assign y679 = ~n3241 ;
  assign y680 = n3242 ;
  assign y681 = n3255 ;
  assign y682 = n3259 ;
  assign y683 = n3264 ;
  assign y684 = n3274 ;
  assign y685 = n3275 ;
  assign y686 = ~n3278 ;
  assign y687 = ~n3279 ;
  assign y688 = n3281 ;
  assign y689 = n3286 ;
  assign y690 = ~n3291 ;
  assign y691 = ~n3294 ;
  assign y692 = ~1'b0 ;
  assign y693 = ~n3307 ;
  assign y694 = n3310 ;
  assign y695 = ~n3311 ;
  assign y696 = ~1'b0 ;
  assign y697 = ~n3315 ;
  assign y698 = ~n3316 ;
  assign y699 = ~n3327 ;
  assign y700 = ~n3335 ;
  assign y701 = ~n3336 ;
  assign y702 = ~n3349 ;
  assign y703 = n3353 ;
  assign y704 = 1'b0 ;
  assign y705 = ~n3356 ;
  assign y706 = n3358 ;
  assign y707 = ~n3359 ;
  assign y708 = n3367 ;
  assign y709 = ~n3379 ;
  assign y710 = n3386 ;
  assign y711 = n3389 ;
  assign y712 = n3391 ;
  assign y713 = n3405 ;
  assign y714 = n3407 ;
  assign y715 = ~1'b0 ;
  assign y716 = n3416 ;
  assign y717 = n3420 ;
  assign y718 = n3423 ;
  assign y719 = n3430 ;
  assign y720 = ~n3435 ;
  assign y721 = n3446 ;
  assign y722 = ~n3447 ;
  assign y723 = ~1'b0 ;
  assign y724 = ~1'b0 ;
  assign y725 = ~n3448 ;
  assign y726 = ~1'b0 ;
  assign y727 = ~n3453 ;
  assign y728 = ~n3454 ;
  assign y729 = ~n3455 ;
  assign y730 = ~n3458 ;
  assign y731 = ~n3465 ;
  assign y732 = ~n3468 ;
  assign y733 = ~n3469 ;
  assign y734 = n3471 ;
  assign y735 = ~n3473 ;
  assign y736 = ~n3478 ;
  assign y737 = ~n3479 ;
  assign y738 = ~n3483 ;
  assign y739 = ~1'b0 ;
  assign y740 = n3511 ;
  assign y741 = ~n3512 ;
  assign y742 = ~n3518 ;
  assign y743 = n3522 ;
  assign y744 = ~n3535 ;
  assign y745 = ~n3537 ;
  assign y746 = ~n3540 ;
  assign y747 = n3545 ;
  assign y748 = ~n3551 ;
  assign y749 = n3553 ;
  assign y750 = n3574 ;
  assign y751 = ~n3578 ;
  assign y752 = ~n3581 ;
  assign y753 = ~n3588 ;
  assign y754 = ~n3593 ;
  assign y755 = ~n3594 ;
  assign y756 = n3595 ;
  assign y757 = n3603 ;
  assign y758 = ~n3607 ;
  assign y759 = n3609 ;
  assign y760 = ~n3611 ;
  assign y761 = ~n3613 ;
  assign y762 = ~n3615 ;
  assign y763 = ~n3622 ;
  assign y764 = ~n3630 ;
  assign y765 = n3632 ;
  assign y766 = ~n3643 ;
  assign y767 = ~n3646 ;
  assign y768 = ~n3648 ;
  assign y769 = ~n3656 ;
  assign y770 = n3658 ;
  assign y771 = ~n3675 ;
  assign y772 = n3679 ;
  assign y773 = n3690 ;
  assign y774 = ~n3706 ;
  assign y775 = ~1'b0 ;
  assign y776 = ~1'b0 ;
  assign y777 = ~n3707 ;
  assign y778 = ~n3708 ;
  assign y779 = ~n3711 ;
  assign y780 = n3717 ;
  assign y781 = ~n3720 ;
  assign y782 = ~n3721 ;
  assign y783 = ~n3734 ;
  assign y784 = ~1'b0 ;
  assign y785 = ~n3735 ;
  assign y786 = ~n3738 ;
  assign y787 = n3740 ;
  assign y788 = ~1'b0 ;
  assign y789 = ~n3741 ;
  assign y790 = n3742 ;
  assign y791 = n3745 ;
  assign y792 = n2266 ;
  assign y793 = ~1'b0 ;
  assign y794 = ~n3746 ;
  assign y795 = n3750 ;
  assign y796 = ~n3751 ;
  assign y797 = n3763 ;
  assign y798 = ~1'b0 ;
  assign y799 = ~1'b0 ;
  assign y800 = n3764 ;
  assign y801 = ~n3768 ;
  assign y802 = n3774 ;
  assign y803 = ~n3779 ;
  assign y804 = ~n3782 ;
  assign y805 = n3785 ;
  assign y806 = ~n3786 ;
  assign y807 = n3791 ;
  assign y808 = n3792 ;
  assign y809 = n3793 ;
  assign y810 = n3798 ;
  assign y811 = ~n3810 ;
  assign y812 = n3814 ;
  assign y813 = n3816 ;
  assign y814 = n3819 ;
  assign y815 = ~n3822 ;
  assign y816 = ~n3830 ;
  assign y817 = n3836 ;
  assign y818 = n3837 ;
  assign y819 = ~n3845 ;
  assign y820 = n3847 ;
  assign y821 = ~1'b0 ;
  assign y822 = ~n3848 ;
  assign y823 = ~n3865 ;
  assign y824 = ~1'b0 ;
  assign y825 = n3878 ;
  assign y826 = n3885 ;
  assign y827 = ~n3892 ;
  assign y828 = n3897 ;
  assign y829 = n3901 ;
  assign y830 = ~1'b0 ;
  assign y831 = ~1'b0 ;
  assign y832 = n3908 ;
  assign y833 = n3912 ;
  assign y834 = ~n3916 ;
  assign y835 = ~n3921 ;
  assign y836 = ~n3923 ;
  assign y837 = ~n3929 ;
  assign y838 = ~n3940 ;
  assign y839 = ~n3943 ;
  assign y840 = ~n3944 ;
  assign y841 = n3954 ;
  assign y842 = n3961 ;
  assign y843 = n3964 ;
  assign y844 = n3975 ;
  assign y845 = n3985 ;
  assign y846 = n3988 ;
  assign y847 = ~n3990 ;
  assign y848 = n3996 ;
  assign y849 = ~n3997 ;
  assign y850 = n3999 ;
  assign y851 = n4009 ;
  assign y852 = ~n4012 ;
  assign y853 = ~1'b0 ;
  assign y854 = n4014 ;
  assign y855 = ~n4016 ;
  assign y856 = ~1'b0 ;
  assign y857 = n4024 ;
  assign y858 = ~n4025 ;
  assign y859 = n4027 ;
  assign y860 = n4038 ;
  assign y861 = ~n4042 ;
  assign y862 = ~n4043 ;
  assign y863 = n4045 ;
  assign y864 = ~n4046 ;
  assign y865 = ~n4051 ;
  assign y866 = n4056 ;
  assign y867 = ~1'b0 ;
  assign y868 = ~n4057 ;
  assign y869 = ~n4060 ;
  assign y870 = n4064 ;
  assign y871 = n4066 ;
  assign y872 = ~n4067 ;
  assign y873 = ~n4075 ;
  assign y874 = ~n4079 ;
  assign y875 = n4091 ;
  assign y876 = n4093 ;
  assign y877 = n4097 ;
  assign y878 = ~n4104 ;
  assign y879 = ~1'b0 ;
  assign y880 = ~n4109 ;
  assign y881 = n4113 ;
  assign y882 = ~n4116 ;
  assign y883 = ~n4118 ;
  assign y884 = n4119 ;
  assign y885 = ~n4124 ;
  assign y886 = ~n4136 ;
  assign y887 = n4138 ;
  assign y888 = n3917 ;
  assign y889 = ~n4142 ;
  assign y890 = n4145 ;
  assign y891 = ~n4155 ;
  assign y892 = ~1'b0 ;
  assign y893 = n4161 ;
  assign y894 = ~1'b0 ;
  assign y895 = n4172 ;
  assign y896 = ~n4174 ;
  assign y897 = ~n4178 ;
  assign y898 = ~n4184 ;
  assign y899 = ~n4192 ;
  assign y900 = n4200 ;
  assign y901 = n4202 ;
  assign y902 = n4204 ;
  assign y903 = ~n4208 ;
  assign y904 = n4212 ;
  assign y905 = n4213 ;
  assign y906 = ~n4215 ;
  assign y907 = ~n4232 ;
  assign y908 = ~n4236 ;
  assign y909 = n4237 ;
  assign y910 = ~n4238 ;
  assign y911 = n4239 ;
  assign y912 = n4247 ;
  assign y913 = ~n4254 ;
  assign y914 = n4261 ;
  assign y915 = ~n4262 ;
  assign y916 = n4264 ;
  assign y917 = n4268 ;
  assign y918 = ~1'b0 ;
  assign y919 = ~n4269 ;
  assign y920 = n4278 ;
  assign y921 = n4285 ;
  assign y922 = n4289 ;
  assign y923 = ~n4292 ;
  assign y924 = ~n4298 ;
  assign y925 = ~n4307 ;
  assign y926 = n4316 ;
  assign y927 = ~n4319 ;
  assign y928 = n4324 ;
  assign y929 = ~n4327 ;
  assign y930 = ~n4329 ;
  assign y931 = ~n4335 ;
  assign y932 = ~n4337 ;
  assign y933 = ~n4338 ;
  assign y934 = n4339 ;
  assign y935 = ~n4350 ;
  assign y936 = ~n4351 ;
  assign y937 = ~n4352 ;
  assign y938 = ~n4358 ;
  assign y939 = ~n4361 ;
  assign y940 = ~n4369 ;
  assign y941 = ~n4372 ;
  assign y942 = n4373 ;
  assign y943 = n4380 ;
  assign y944 = n4400 ;
  assign y945 = ~n4401 ;
  assign y946 = n4405 ;
  assign y947 = ~n4406 ;
  assign y948 = ~n4413 ;
  assign y949 = ~n4414 ;
  assign y950 = ~n4415 ;
  assign y951 = ~n4423 ;
  assign y952 = n4424 ;
  assign y953 = ~1'b0 ;
  assign y954 = ~n4425 ;
  assign y955 = n4428 ;
  assign y956 = ~n4434 ;
  assign y957 = ~n4439 ;
  assign y958 = ~n4440 ;
  assign y959 = n4448 ;
  assign y960 = n4450 ;
  assign y961 = n4453 ;
  assign y962 = n4454 ;
  assign y963 = n4456 ;
  assign y964 = n4463 ;
  assign y965 = ~n4464 ;
  assign y966 = n4467 ;
  assign y967 = ~n4469 ;
  assign y968 = n4476 ;
  assign y969 = ~n4484 ;
  assign y970 = ~n4497 ;
  assign y971 = n4501 ;
  assign y972 = n4509 ;
  assign y973 = n4511 ;
  assign y974 = ~1'b0 ;
  assign y975 = ~n4519 ;
  assign y976 = ~n4521 ;
  assign y977 = n4525 ;
  assign y978 = ~n4530 ;
  assign y979 = ~n4535 ;
  assign y980 = n4536 ;
  assign y981 = ~n4540 ;
  assign y982 = ~1'b0 ;
  assign y983 = ~n4547 ;
  assign y984 = n4553 ;
  assign y985 = ~n4559 ;
  assign y986 = ~1'b0 ;
  assign y987 = n4566 ;
  assign y988 = n4568 ;
  assign y989 = ~1'b0 ;
  assign y990 = ~n4575 ;
  assign y991 = ~n4584 ;
  assign y992 = ~1'b0 ;
  assign y993 = ~n4585 ;
  assign y994 = ~n4595 ;
  assign y995 = ~n4607 ;
  assign y996 = n4611 ;
  assign y997 = ~n4612 ;
  assign y998 = ~n4620 ;
  assign y999 = ~1'b0 ;
  assign y1000 = ~n4629 ;
  assign y1001 = n4639 ;
  assign y1002 = ~n4647 ;
  assign y1003 = ~n4649 ;
  assign y1004 = n4650 ;
  assign y1005 = ~n4653 ;
  assign y1006 = ~n4659 ;
  assign y1007 = ~n4667 ;
  assign y1008 = ~n4669 ;
  assign y1009 = n4672 ;
  assign y1010 = ~1'b0 ;
  assign y1011 = n4678 ;
  assign y1012 = n4679 ;
  assign y1013 = ~n4681 ;
  assign y1014 = n4713 ;
  assign y1015 = ~n4718 ;
  assign y1016 = n4725 ;
  assign y1017 = ~n4730 ;
  assign y1018 = n4738 ;
  assign y1019 = ~1'b0 ;
  assign y1020 = ~n4751 ;
  assign y1021 = ~1'b0 ;
  assign y1022 = n4755 ;
  assign y1023 = ~n4762 ;
  assign y1024 = n4765 ;
  assign y1025 = ~n4767 ;
  assign y1026 = n4768 ;
  assign y1027 = ~n4769 ;
  assign y1028 = ~n4779 ;
  assign y1029 = ~n4784 ;
  assign y1030 = ~n4785 ;
  assign y1031 = ~n4786 ;
  assign y1032 = n4790 ;
  assign y1033 = n4793 ;
  assign y1034 = ~1'b0 ;
  assign y1035 = n4801 ;
  assign y1036 = n4804 ;
  assign y1037 = n4805 ;
  assign y1038 = n4811 ;
  assign y1039 = ~n4819 ;
  assign y1040 = ~n4824 ;
  assign y1041 = ~n4827 ;
  assign y1042 = ~n4837 ;
  assign y1043 = n4851 ;
  assign y1044 = n4860 ;
  assign y1045 = ~1'b0 ;
  assign y1046 = n4863 ;
  assign y1047 = ~n4869 ;
  assign y1048 = n4872 ;
  assign y1049 = ~n4879 ;
  assign y1050 = n4884 ;
  assign y1051 = n4888 ;
  assign y1052 = ~n4893 ;
  assign y1053 = n4897 ;
  assign y1054 = ~n4903 ;
  assign y1055 = ~n4908 ;
  assign y1056 = ~n4915 ;
  assign y1057 = ~n4917 ;
  assign y1058 = n4923 ;
  assign y1059 = ~n4930 ;
  assign y1060 = ~n4935 ;
  assign y1061 = ~n4939 ;
  assign y1062 = ~1'b0 ;
  assign y1063 = ~n4942 ;
  assign y1064 = ~n4959 ;
  assign y1065 = n4967 ;
  assign y1066 = n4973 ;
  assign y1067 = n4982 ;
  assign y1068 = n4986 ;
  assign y1069 = ~n4990 ;
  assign y1070 = n4991 ;
  assign y1071 = n4995 ;
  assign y1072 = ~n4997 ;
  assign y1073 = ~n4998 ;
  assign y1074 = ~n4999 ;
  assign y1075 = n5003 ;
  assign y1076 = ~n5004 ;
  assign y1077 = ~n5010 ;
  assign y1078 = ~n5013 ;
  assign y1079 = n5020 ;
  assign y1080 = ~1'b0 ;
  assign y1081 = n5024 ;
  assign y1082 = ~1'b0 ;
  assign y1083 = ~1'b0 ;
  assign y1084 = n5027 ;
  assign y1085 = n5030 ;
  assign y1086 = n5034 ;
  assign y1087 = n5037 ;
  assign y1088 = ~n5039 ;
  assign y1089 = n5043 ;
  assign y1090 = ~n5044 ;
  assign y1091 = ~n5048 ;
  assign y1092 = n5049 ;
  assign y1093 = ~n5050 ;
  assign y1094 = ~1'b0 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = n5053 ;
  assign y1097 = n5064 ;
  assign y1098 = ~n5066 ;
  assign y1099 = n5071 ;
  assign y1100 = ~1'b0 ;
  assign y1101 = n5075 ;
  assign y1102 = ~n5078 ;
  assign y1103 = n5088 ;
  assign y1104 = ~n5092 ;
  assign y1105 = ~n5098 ;
  assign y1106 = ~n5100 ;
  assign y1107 = n5104 ;
  assign y1108 = ~n5107 ;
  assign y1109 = ~n5109 ;
  assign y1110 = ~n5112 ;
  assign y1111 = n5123 ;
  assign y1112 = ~1'b0 ;
  assign y1113 = ~n5126 ;
  assign y1114 = n5134 ;
  assign y1115 = ~1'b0 ;
  assign y1116 = n5137 ;
  assign y1117 = n5153 ;
  assign y1118 = ~1'b0 ;
  assign y1119 = n5155 ;
  assign y1120 = ~n5157 ;
  assign y1121 = ~1'b0 ;
  assign y1122 = ~n5177 ;
  assign y1123 = ~n5180 ;
  assign y1124 = ~n5181 ;
  assign y1125 = n5186 ;
  assign y1126 = n5187 ;
  assign y1127 = n5190 ;
  assign y1128 = n5202 ;
  assign y1129 = n5203 ;
  assign y1130 = n5209 ;
  assign y1131 = ~n5213 ;
  assign y1132 = ~n5218 ;
  assign y1133 = n5225 ;
  assign y1134 = n5231 ;
  assign y1135 = 1'b0 ;
  assign y1136 = n5232 ;
  assign y1137 = n5238 ;
  assign y1138 = ~n5241 ;
  assign y1139 = ~n5245 ;
  assign y1140 = ~n5247 ;
  assign y1141 = ~n5258 ;
  assign y1142 = n5260 ;
  assign y1143 = ~1'b0 ;
  assign y1144 = ~n5273 ;
  assign y1145 = ~n5274 ;
  assign y1146 = ~n5276 ;
  assign y1147 = ~n5277 ;
  assign y1148 = n5286 ;
  assign y1149 = ~n5287 ;
  assign y1150 = ~n5309 ;
  assign y1151 = ~1'b0 ;
  assign y1152 = n5315 ;
  assign y1153 = n5319 ;
  assign y1154 = n5320 ;
  assign y1155 = n5323 ;
  assign y1156 = n5326 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = ~n5327 ;
  assign y1159 = n5330 ;
  assign y1160 = ~n5334 ;
  assign y1161 = ~n5349 ;
  assign y1162 = n5350 ;
  assign y1163 = ~n5357 ;
  assign y1164 = ~n5362 ;
  assign y1165 = n5366 ;
  assign y1166 = n5371 ;
  assign y1167 = ~n5374 ;
  assign y1168 = ~n5389 ;
  assign y1169 = n5393 ;
  assign y1170 = n5403 ;
  assign y1171 = n5407 ;
  assign y1172 = n5412 ;
  assign y1173 = ~n5414 ;
  assign y1174 = ~n5415 ;
  assign y1175 = n5419 ;
  assign y1176 = ~n5423 ;
  assign y1177 = ~1'b0 ;
  assign y1178 = ~1'b0 ;
  assign y1179 = n5433 ;
  assign y1180 = ~n5442 ;
  assign y1181 = ~n5459 ;
  assign y1182 = n5470 ;
  assign y1183 = ~n5477 ;
  assign y1184 = ~n5478 ;
  assign y1185 = n5504 ;
  assign y1186 = ~n5506 ;
  assign y1187 = ~n5511 ;
  assign y1188 = n5517 ;
  assign y1189 = ~n5522 ;
  assign y1190 = ~n5527 ;
  assign y1191 = ~n5536 ;
  assign y1192 = n5540 ;
  assign y1193 = n5543 ;
  assign y1194 = ~n5546 ;
  assign y1195 = n5547 ;
  assign y1196 = ~n5553 ;
  assign y1197 = n5561 ;
  assign y1198 = ~n5563 ;
  assign y1199 = ~n5567 ;
  assign y1200 = ~n5569 ;
  assign y1201 = ~n5570 ;
  assign y1202 = n5579 ;
  assign y1203 = ~1'b0 ;
  assign y1204 = ~n5580 ;
  assign y1205 = n5582 ;
  assign y1206 = ~1'b0 ;
  assign y1207 = n5597 ;
  assign y1208 = ~n5620 ;
  assign y1209 = ~n5626 ;
  assign y1210 = ~1'b0 ;
  assign y1211 = ~n5627 ;
  assign y1212 = ~n5632 ;
  assign y1213 = ~n5633 ;
  assign y1214 = n5634 ;
  assign y1215 = n5643 ;
  assign y1216 = n5645 ;
  assign y1217 = n5649 ;
  assign y1218 = ~n5657 ;
  assign y1219 = n5662 ;
  assign y1220 = ~n5663 ;
  assign y1221 = n5664 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = ~n5665 ;
  assign y1224 = n5669 ;
  assign y1225 = ~1'b0 ;
  assign y1226 = ~n5670 ;
  assign y1227 = n5671 ;
  assign y1228 = ~n5672 ;
  assign y1229 = ~1'b0 ;
  assign y1230 = n5673 ;
  assign y1231 = ~n5691 ;
  assign y1232 = ~n5694 ;
  assign y1233 = ~n5695 ;
  assign y1234 = n5701 ;
  assign y1235 = ~n5707 ;
  assign y1236 = ~n5718 ;
  assign y1237 = ~n5721 ;
  assign y1238 = ~n5730 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = n5736 ;
  assign y1241 = n5742 ;
  assign y1242 = ~n5748 ;
  assign y1243 = ~n5757 ;
  assign y1244 = ~1'b0 ;
  assign y1245 = n5766 ;
  assign y1246 = ~n5769 ;
  assign y1247 = ~n5773 ;
  assign y1248 = ~n5774 ;
  assign y1249 = ~n5775 ;
  assign y1250 = n5776 ;
  assign y1251 = n5778 ;
  assign y1252 = ~n530 ;
  assign y1253 = n5784 ;
  assign y1254 = ~n5792 ;
  assign y1255 = n5795 ;
  assign y1256 = ~n5796 ;
  assign y1257 = ~1'b0 ;
  assign y1258 = ~n5801 ;
  assign y1259 = ~n5802 ;
  assign y1260 = ~n5810 ;
  assign y1261 = n5817 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = n5824 ;
  assign y1264 = n5839 ;
  assign y1265 = ~n5840 ;
  assign y1266 = n5850 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~1'b0 ;
  assign y1269 = n5860 ;
  assign y1270 = n5861 ;
  assign y1271 = n5867 ;
  assign y1272 = ~n5881 ;
  assign y1273 = ~n5882 ;
  assign y1274 = ~1'b0 ;
  assign y1275 = ~n5887 ;
  assign y1276 = ~n5888 ;
  assign y1277 = n5898 ;
  assign y1278 = n5899 ;
  assign y1279 = n5909 ;
  assign y1280 = n5911 ;
  assign y1281 = ~n5917 ;
  assign y1282 = ~n5921 ;
  assign y1283 = ~1'b0 ;
  assign y1284 = n5930 ;
  assign y1285 = n5934 ;
  assign y1286 = ~n5944 ;
  assign y1287 = ~n5955 ;
  assign y1288 = ~n5957 ;
  assign y1289 = ~n5958 ;
  assign y1290 = n5963 ;
  assign y1291 = n5966 ;
  assign y1292 = ~n5969 ;
  assign y1293 = n5972 ;
  assign y1294 = ~n5985 ;
  assign y1295 = ~1'b0 ;
  assign y1296 = ~n5987 ;
  assign y1297 = n5988 ;
  assign y1298 = ~n6002 ;
  assign y1299 = ~n6003 ;
  assign y1300 = ~1'b0 ;
  assign y1301 = ~n6009 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = n6010 ;
  assign y1304 = n6021 ;
  assign y1305 = n6029 ;
  assign y1306 = ~n6034 ;
  assign y1307 = ~n6036 ;
  assign y1308 = n6046 ;
  assign y1309 = n6050 ;
  assign y1310 = n6071 ;
  assign y1311 = n6081 ;
  assign y1312 = n6090 ;
  assign y1313 = ~1'b0 ;
  assign y1314 = ~n6091 ;
  assign y1315 = n6102 ;
  assign y1316 = ~n6107 ;
  assign y1317 = ~1'b0 ;
  assign y1318 = ~n6112 ;
  assign y1319 = n6122 ;
  assign y1320 = ~n6123 ;
  assign y1321 = ~n6129 ;
  assign y1322 = ~1'b0 ;
  assign y1323 = ~1'b0 ;
  assign y1324 = n6130 ;
  assign y1325 = ~n6131 ;
  assign y1326 = n6136 ;
  assign y1327 = ~1'b0 ;
  assign y1328 = n6138 ;
  assign y1329 = n6141 ;
  assign y1330 = ~n6150 ;
  assign y1331 = n6153 ;
  assign y1332 = ~n6160 ;
  assign y1333 = ~n6166 ;
  assign y1334 = ~n6168 ;
  assign y1335 = n6173 ;
  assign y1336 = n6178 ;
  assign y1337 = ~n6181 ;
  assign y1338 = ~n6185 ;
  assign y1339 = n6189 ;
  assign y1340 = ~n6196 ;
  assign y1341 = n6209 ;
  assign y1342 = ~n6210 ;
  assign y1343 = ~1'b0 ;
  assign y1344 = ~n6216 ;
  assign y1345 = ~1'b0 ;
  assign y1346 = ~n6220 ;
  assign y1347 = ~n6227 ;
  assign y1348 = n6230 ;
  assign y1349 = n6236 ;
  assign y1350 = ~1'b0 ;
  assign y1351 = n6237 ;
  assign y1352 = ~1'b0 ;
  assign y1353 = n6239 ;
  assign y1354 = n6244 ;
  assign y1355 = n6250 ;
  assign y1356 = n6255 ;
  assign y1357 = ~n6262 ;
  assign y1358 = n6277 ;
  assign y1359 = n6283 ;
  assign y1360 = n6298 ;
  assign y1361 = ~n6301 ;
  assign y1362 = n6302 ;
  assign y1363 = n6304 ;
  assign y1364 = ~n6312 ;
  assign y1365 = n6321 ;
  assign y1366 = n6326 ;
  assign y1367 = n6327 ;
  assign y1368 = ~n6337 ;
  assign y1369 = ~n6339 ;
  assign y1370 = ~n6343 ;
  assign y1371 = ~n6345 ;
  assign y1372 = n6347 ;
  assign y1373 = n6351 ;
  assign y1374 = n6357 ;
  assign y1375 = n6366 ;
  assign y1376 = n6375 ;
  assign y1377 = n6379 ;
  assign y1378 = n6380 ;
  assign y1379 = ~n6388 ;
  assign y1380 = ~1'b0 ;
  assign y1381 = ~1'b0 ;
  assign y1382 = n6391 ;
  assign y1383 = n6396 ;
  assign y1384 = ~n6400 ;
  assign y1385 = n6407 ;
  assign y1386 = n6411 ;
  assign y1387 = n6415 ;
  assign y1388 = n6425 ;
  assign y1389 = n6427 ;
  assign y1390 = ~n6428 ;
  assign y1391 = ~n6431 ;
  assign y1392 = ~1'b0 ;
  assign y1393 = ~n6441 ;
  assign y1394 = ~n6451 ;
  assign y1395 = n6452 ;
  assign y1396 = ~n6456 ;
  assign y1397 = n6457 ;
  assign y1398 = ~n6459 ;
  assign y1399 = ~n6467 ;
  assign y1400 = n6468 ;
  assign y1401 = n6473 ;
  assign y1402 = n6476 ;
  assign y1403 = ~n6478 ;
  assign y1404 = n6479 ;
  assign y1405 = ~n6484 ;
  assign y1406 = ~n6496 ;
  assign y1407 = ~n6499 ;
  assign y1408 = ~n4339 ;
  assign y1409 = ~n6513 ;
  assign y1410 = ~n6523 ;
  assign y1411 = ~n6525 ;
  assign y1412 = n6537 ;
  assign y1413 = ~1'b0 ;
  assign y1414 = ~n6538 ;
  assign y1415 = n6566 ;
  assign y1416 = ~n6571 ;
  assign y1417 = n6572 ;
  assign y1418 = ~n6573 ;
  assign y1419 = n6576 ;
  assign y1420 = n6586 ;
  assign y1421 = ~n6587 ;
  assign y1422 = ~n6589 ;
  assign y1423 = n6592 ;
  assign y1424 = ~n6595 ;
  assign y1425 = ~n6598 ;
  assign y1426 = n6600 ;
  assign y1427 = ~1'b0 ;
  assign y1428 = ~n6604 ;
  assign y1429 = ~n6615 ;
  assign y1430 = ~1'b0 ;
  assign y1431 = ~n6624 ;
  assign y1432 = n6633 ;
  assign y1433 = n6643 ;
  assign y1434 = n6652 ;
  assign y1435 = ~n6664 ;
  assign y1436 = ~n6673 ;
  assign y1437 = n6675 ;
  assign y1438 = ~1'b0 ;
  assign y1439 = n6677 ;
  assign y1440 = ~n6682 ;
  assign y1441 = n6683 ;
  assign y1442 = n6689 ;
  assign y1443 = ~n6693 ;
  assign y1444 = ~n6701 ;
  assign y1445 = ~n6706 ;
  assign y1446 = n6708 ;
  assign y1447 = n6714 ;
  assign y1448 = n6715 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = n6718 ;
  assign y1451 = ~n6726 ;
  assign y1452 = n6731 ;
  assign y1453 = n6740 ;
  assign y1454 = ~1'b0 ;
  assign y1455 = n6754 ;
  assign y1456 = ~n6760 ;
  assign y1457 = ~n6761 ;
  assign y1458 = ~n6772 ;
  assign y1459 = ~n6775 ;
  assign y1460 = n6788 ;
  assign y1461 = ~n6792 ;
  assign y1462 = n6797 ;
  assign y1463 = ~n6801 ;
  assign y1464 = ~n6802 ;
  assign y1465 = ~n6815 ;
  assign y1466 = n6816 ;
  assign y1467 = n6819 ;
  assign y1468 = n6825 ;
  assign y1469 = ~n6833 ;
  assign y1470 = ~n6844 ;
  assign y1471 = ~1'b0 ;
  assign y1472 = n6845 ;
  assign y1473 = ~n6846 ;
  assign y1474 = n6852 ;
  assign y1475 = ~n6854 ;
  assign y1476 = n6858 ;
  assign y1477 = n6860 ;
  assign y1478 = ~n6863 ;
  assign y1479 = n6866 ;
  assign y1480 = ~n6870 ;
  assign y1481 = ~n6878 ;
  assign y1482 = n6883 ;
  assign y1483 = n6885 ;
  assign y1484 = ~n6889 ;
  assign y1485 = ~n6895 ;
  assign y1486 = ~n6900 ;
  assign y1487 = ~n6913 ;
  assign y1488 = ~n6920 ;
  assign y1489 = n6924 ;
  assign y1490 = n6940 ;
  assign y1491 = n6957 ;
  assign y1492 = ~n6961 ;
  assign y1493 = ~1'b0 ;
  assign y1494 = ~n6964 ;
  assign y1495 = ~n6965 ;
  assign y1496 = n6974 ;
  assign y1497 = n6975 ;
  assign y1498 = ~n6976 ;
  assign y1499 = ~n6978 ;
  assign y1500 = n6984 ;
  assign y1501 = n6993 ;
  assign y1502 = ~n6995 ;
  assign y1503 = ~n6996 ;
  assign y1504 = n7001 ;
  assign y1505 = ~n7024 ;
  assign y1506 = n7026 ;
  assign y1507 = n7038 ;
  assign y1508 = ~1'b0 ;
  assign y1509 = ~1'b0 ;
  assign y1510 = n7041 ;
  assign y1511 = ~n7060 ;
  assign y1512 = ~n7061 ;
  assign y1513 = ~n7072 ;
  assign y1514 = ~n7080 ;
  assign y1515 = ~n7083 ;
  assign y1516 = n7084 ;
  assign y1517 = ~n7090 ;
  assign y1518 = ~n7095 ;
  assign y1519 = n7098 ;
  assign y1520 = ~n7108 ;
  assign y1521 = n7109 ;
  assign y1522 = ~n7111 ;
  assign y1523 = n7113 ;
  assign y1524 = n7121 ;
  assign y1525 = ~n7122 ;
  assign y1526 = n7129 ;
  assign y1527 = n7137 ;
  assign y1528 = ~1'b0 ;
  assign y1529 = n7141 ;
  assign y1530 = ~n7143 ;
  assign y1531 = ~n7145 ;
  assign y1532 = n7149 ;
  assign y1533 = ~n7154 ;
  assign y1534 = n7160 ;
  assign y1535 = n7187 ;
  assign y1536 = ~1'b0 ;
  assign y1537 = n7190 ;
  assign y1538 = ~n7207 ;
  assign y1539 = x96 ;
  assign y1540 = ~1'b0 ;
  assign y1541 = ~n7208 ;
  assign y1542 = ~n7211 ;
  assign y1543 = n7214 ;
  assign y1544 = n7217 ;
  assign y1545 = n7221 ;
  assign y1546 = n7229 ;
  assign y1547 = ~n7235 ;
  assign y1548 = n7237 ;
  assign y1549 = n7245 ;
  assign y1550 = n7255 ;
  assign y1551 = n7256 ;
  assign y1552 = n7260 ;
  assign y1553 = ~n7261 ;
  assign y1554 = ~n7263 ;
  assign y1555 = ~n7272 ;
  assign y1556 = n7275 ;
  assign y1557 = ~n7276 ;
  assign y1558 = n7281 ;
  assign y1559 = ~n7289 ;
  assign y1560 = n7291 ;
  assign y1561 = n7295 ;
  assign y1562 = ~n7300 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~n7305 ;
  assign y1565 = n7308 ;
  assign y1566 = ~n7315 ;
  assign y1567 = ~n7319 ;
  assign y1568 = n7325 ;
  assign y1569 = n7330 ;
  assign y1570 = ~n7332 ;
  assign y1571 = ~n7344 ;
  assign y1572 = ~1'b0 ;
  assign y1573 = ~n7346 ;
  assign y1574 = ~n7352 ;
  assign y1575 = n7358 ;
  assign y1576 = ~n4417 ;
  assign y1577 = ~n7372 ;
  assign y1578 = ~n7373 ;
  assign y1579 = ~1'b0 ;
  assign y1580 = n7374 ;
  assign y1581 = ~n7377 ;
  assign y1582 = n7385 ;
  assign y1583 = n7387 ;
  assign y1584 = ~n7389 ;
  assign y1585 = ~n7409 ;
  assign y1586 = ~n7413 ;
  assign y1587 = ~n7415 ;
  assign y1588 = n7424 ;
  assign y1589 = ~n7436 ;
  assign y1590 = ~n7438 ;
  assign y1591 = n7455 ;
  assign y1592 = n7466 ;
  assign y1593 = n7471 ;
  assign y1594 = ~n7479 ;
  assign y1595 = ~n7482 ;
  assign y1596 = n7488 ;
  assign y1597 = ~n4633 ;
  assign y1598 = ~n7491 ;
  assign y1599 = ~1'b0 ;
  assign y1600 = n7505 ;
  assign y1601 = ~n7519 ;
  assign y1602 = ~n7522 ;
  assign y1603 = ~n7529 ;
  assign y1604 = ~1'b0 ;
  assign y1605 = ~n7530 ;
  assign y1606 = n7532 ;
  assign y1607 = n7547 ;
  assign y1608 = ~n7550 ;
  assign y1609 = n7554 ;
  assign y1610 = n7568 ;
  assign y1611 = n7573 ;
  assign y1612 = ~n7579 ;
  assign y1613 = ~n7584 ;
  assign y1614 = ~n7590 ;
  assign y1615 = ~n7598 ;
  assign y1616 = n7599 ;
  assign y1617 = n7607 ;
  assign y1618 = ~n7620 ;
  assign y1619 = ~n7622 ;
  assign y1620 = ~n7624 ;
  assign y1621 = n7628 ;
  assign y1622 = ~n7632 ;
  assign y1623 = n7634 ;
  assign y1624 = n7636 ;
  assign y1625 = n7637 ;
  assign y1626 = ~n7639 ;
  assign y1627 = n7640 ;
  assign y1628 = n7650 ;
  assign y1629 = n7654 ;
  assign y1630 = ~n7659 ;
  assign y1631 = n7672 ;
  assign y1632 = n7674 ;
  assign y1633 = ~n7685 ;
  assign y1634 = ~n7689 ;
  assign y1635 = n7692 ;
  assign y1636 = n7694 ;
  assign y1637 = n7697 ;
  assign y1638 = n7705 ;
  assign y1639 = n7707 ;
  assign y1640 = n7712 ;
  assign y1641 = n7717 ;
  assign y1642 = ~n7722 ;
  assign y1643 = ~1'b0 ;
  assign y1644 = ~n7727 ;
  assign y1645 = ~n284 ;
  assign y1646 = ~n7745 ;
  assign y1647 = n7748 ;
  assign y1648 = n7753 ;
  assign y1649 = ~n7755 ;
  assign y1650 = n7756 ;
  assign y1651 = ~n7757 ;
  assign y1652 = n7760 ;
  assign y1653 = ~n7765 ;
  assign y1654 = n7772 ;
  assign y1655 = n7783 ;
  assign y1656 = n7788 ;
  assign y1657 = ~n7789 ;
  assign y1658 = n7790 ;
  assign y1659 = n7791 ;
  assign y1660 = ~n7792 ;
  assign y1661 = ~n7797 ;
  assign y1662 = ~1'b0 ;
  assign y1663 = n7800 ;
  assign y1664 = n7803 ;
  assign y1665 = ~n7805 ;
  assign y1666 = ~1'b0 ;
  assign y1667 = ~n7812 ;
  assign y1668 = n7820 ;
  assign y1669 = n7829 ;
  assign y1670 = ~n7842 ;
  assign y1671 = ~1'b0 ;
  assign y1672 = n7843 ;
  assign y1673 = ~n7845 ;
  assign y1674 = ~n7847 ;
  assign y1675 = ~n7849 ;
  assign y1676 = ~n7859 ;
  assign y1677 = ~n7860 ;
  assign y1678 = n7862 ;
  assign y1679 = ~1'b0 ;
  assign y1680 = ~n7867 ;
  assign y1681 = n7870 ;
  assign y1682 = n7875 ;
  assign y1683 = ~1'b0 ;
  assign y1684 = n7876 ;
  assign y1685 = ~n7879 ;
  assign y1686 = n7880 ;
  assign y1687 = ~n7882 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = ~1'b0 ;
  assign y1690 = ~n7886 ;
  assign y1691 = ~n7892 ;
  assign y1692 = n7894 ;
  assign y1693 = n7896 ;
  assign y1694 = n7904 ;
  assign y1695 = ~n7908 ;
  assign y1696 = ~1'b0 ;
  assign y1697 = n7912 ;
  assign y1698 = n7913 ;
  assign y1699 = n7915 ;
  assign y1700 = ~n7917 ;
  assign y1701 = ~1'b0 ;
  assign y1702 = n7927 ;
  assign y1703 = ~1'b0 ;
  assign y1704 = ~n7938 ;
  assign y1705 = n7941 ;
  assign y1706 = n7949 ;
  assign y1707 = ~n7956 ;
  assign y1708 = n7957 ;
  assign y1709 = ~n7961 ;
  assign y1710 = n7962 ;
  assign y1711 = n7963 ;
  assign y1712 = ~n7968 ;
  assign y1713 = ~n7974 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = n7980 ;
  assign y1716 = n7983 ;
  assign y1717 = n7986 ;
  assign y1718 = ~n7988 ;
  assign y1719 = ~n7989 ;
  assign y1720 = n7991 ;
  assign y1721 = n7997 ;
  assign y1722 = n8000 ;
  assign y1723 = ~n8006 ;
  assign y1724 = n8013 ;
  assign y1725 = ~n8018 ;
  assign y1726 = ~n8027 ;
  assign y1727 = n8028 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = ~n8031 ;
  assign y1730 = ~n8036 ;
  assign y1731 = n8039 ;
  assign y1732 = n8042 ;
  assign y1733 = n8046 ;
  assign y1734 = n8051 ;
  assign y1735 = ~n8052 ;
  assign y1736 = ~n8053 ;
  assign y1737 = ~n8065 ;
  assign y1738 = n8066 ;
  assign y1739 = ~n8072 ;
  assign y1740 = n8074 ;
  assign y1741 = ~1'b0 ;
  assign y1742 = n8076 ;
  assign y1743 = ~1'b0 ;
  assign y1744 = ~n8079 ;
  assign y1745 = n8080 ;
  assign y1746 = ~n8082 ;
  assign y1747 = ~1'b0 ;
  assign y1748 = n8093 ;
  assign y1749 = n8098 ;
  assign y1750 = ~n8106 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = ~n8110 ;
  assign y1753 = ~n8121 ;
  assign y1754 = ~n8125 ;
  assign y1755 = ~n8132 ;
  assign y1756 = ~n8137 ;
  assign y1757 = n8143 ;
  assign y1758 = ~n8144 ;
  assign y1759 = n8146 ;
  assign y1760 = n8154 ;
  assign y1761 = ~1'b0 ;
  assign y1762 = n8165 ;
  assign y1763 = ~n8171 ;
  assign y1764 = n8174 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = n8195 ;
  assign y1767 = ~n8198 ;
  assign y1768 = ~n8199 ;
  assign y1769 = n8210 ;
  assign y1770 = n8219 ;
  assign y1771 = ~n8224 ;
  assign y1772 = ~n8225 ;
  assign y1773 = n8235 ;
  assign y1774 = ~n8236 ;
  assign y1775 = n8240 ;
  assign y1776 = n8258 ;
  assign y1777 = ~n8263 ;
  assign y1778 = ~n8272 ;
  assign y1779 = n8276 ;
  assign y1780 = ~n8289 ;
  assign y1781 = ~n8292 ;
  assign y1782 = ~n8297 ;
  assign y1783 = ~n8302 ;
  assign y1784 = ~n8305 ;
  assign y1785 = ~n8315 ;
  assign y1786 = ~n8319 ;
  assign y1787 = n8325 ;
  assign y1788 = n8329 ;
  assign y1789 = n8330 ;
  assign y1790 = n8339 ;
  assign y1791 = n8340 ;
  assign y1792 = ~1'b0 ;
  assign y1793 = ~n8347 ;
  assign y1794 = n8354 ;
  assign y1795 = n8355 ;
  assign y1796 = ~n8359 ;
  assign y1797 = ~n8362 ;
  assign y1798 = ~n8364 ;
  assign y1799 = ~1'b0 ;
  assign y1800 = ~n8376 ;
  assign y1801 = ~n7362 ;
  assign y1802 = n8381 ;
  assign y1803 = n8386 ;
  assign y1804 = n8387 ;
  assign y1805 = n8388 ;
  assign y1806 = n8392 ;
  assign y1807 = n8409 ;
  assign y1808 = ~1'b0 ;
  assign y1809 = n8413 ;
  assign y1810 = ~1'b0 ;
  assign y1811 = n8419 ;
  assign y1812 = ~n8420 ;
  assign y1813 = n8422 ;
  assign y1814 = ~1'b0 ;
  assign y1815 = ~n8425 ;
  assign y1816 = n8430 ;
  assign y1817 = n8439 ;
  assign y1818 = ~n8444 ;
  assign y1819 = n8450 ;
  assign y1820 = ~1'b0 ;
  assign y1821 = n8453 ;
  assign y1822 = ~n8461 ;
  assign y1823 = n8465 ;
  assign y1824 = ~n8477 ;
  assign y1825 = ~n8486 ;
  assign y1826 = ~n8491 ;
  assign y1827 = n8493 ;
  assign y1828 = n8495 ;
  assign y1829 = ~1'b0 ;
  assign y1830 = ~1'b0 ;
  assign y1831 = ~n8496 ;
  assign y1832 = n8498 ;
  assign y1833 = ~n8503 ;
  assign y1834 = n8508 ;
  assign y1835 = n8509 ;
  assign y1836 = n8514 ;
  assign y1837 = ~n8517 ;
  assign y1838 = n8524 ;
  assign y1839 = ~n8532 ;
  assign y1840 = n8536 ;
  assign y1841 = ~1'b0 ;
  assign y1842 = ~n8538 ;
  assign y1843 = n8540 ;
  assign y1844 = ~n8544 ;
  assign y1845 = ~n8545 ;
  assign y1846 = n8554 ;
  assign y1847 = ~n8566 ;
  assign y1848 = ~n8578 ;
  assign y1849 = ~n8583 ;
  assign y1850 = ~1'b0 ;
  assign y1851 = ~n8591 ;
  assign y1852 = ~n8593 ;
  assign y1853 = n8601 ;
  assign y1854 = n8607 ;
  assign y1855 = n8613 ;
  assign y1856 = ~1'b0 ;
  assign y1857 = n8616 ;
  assign y1858 = ~n8627 ;
  assign y1859 = n8637 ;
  assign y1860 = ~n8643 ;
  assign y1861 = n8648 ;
  assign y1862 = ~n8657 ;
  assign y1863 = ~n8661 ;
  assign y1864 = ~n8663 ;
  assign y1865 = ~n8664 ;
  assign y1866 = ~n8666 ;
  assign y1867 = ~n8671 ;
  assign y1868 = ~n8672 ;
  assign y1869 = n8675 ;
  assign y1870 = ~n8683 ;
  assign y1871 = ~1'b0 ;
  assign y1872 = n8702 ;
  assign y1873 = n8709 ;
  assign y1874 = n8712 ;
  assign y1875 = ~1'b0 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = ~n8716 ;
  assign y1878 = n8717 ;
  assign y1879 = n8730 ;
  assign y1880 = n8734 ;
  assign y1881 = ~n8745 ;
  assign y1882 = ~1'b0 ;
  assign y1883 = n8757 ;
  assign y1884 = ~n8758 ;
  assign y1885 = n8765 ;
  assign y1886 = ~n8768 ;
  assign y1887 = ~n8772 ;
  assign y1888 = ~1'b0 ;
  assign y1889 = ~n8776 ;
  assign y1890 = n8786 ;
  assign y1891 = ~n8794 ;
  assign y1892 = n8798 ;
  assign y1893 = n8805 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = ~n8806 ;
  assign y1896 = n8808 ;
  assign y1897 = ~n8809 ;
  assign y1898 = n8811 ;
  assign y1899 = n8817 ;
  assign y1900 = ~n8830 ;
  assign y1901 = ~1'b0 ;
  assign y1902 = ~n8831 ;
  assign y1903 = n8838 ;
  assign y1904 = ~n8843 ;
  assign y1905 = n8847 ;
  assign y1906 = ~n8848 ;
  assign y1907 = n8851 ;
  assign y1908 = ~n8852 ;
  assign y1909 = n8856 ;
  assign y1910 = n8868 ;
  assign y1911 = n8880 ;
  assign y1912 = n8892 ;
  assign y1913 = ~1'b0 ;
  assign y1914 = ~n8896 ;
  assign y1915 = ~n8897 ;
  assign y1916 = ~n8898 ;
  assign y1917 = ~n8905 ;
  assign y1918 = ~n8908 ;
  assign y1919 = n8910 ;
  assign y1920 = ~1'b0 ;
  assign y1921 = ~n8913 ;
  assign y1922 = ~n8921 ;
  assign y1923 = ~n8923 ;
  assign y1924 = ~n8931 ;
  assign y1925 = ~n8936 ;
  assign y1926 = ~n8307 ;
  assign y1927 = ~n8943 ;
  assign y1928 = n8946 ;
  assign y1929 = ~n8953 ;
  assign y1930 = ~n8958 ;
  assign y1931 = ~n8963 ;
  assign y1932 = ~n8969 ;
  assign y1933 = ~n8976 ;
  assign y1934 = ~n8980 ;
  assign y1935 = n8981 ;
  assign y1936 = ~n8988 ;
  assign y1937 = ~n8993 ;
  assign y1938 = ~n8999 ;
  assign y1939 = ~n9001 ;
  assign y1940 = n9002 ;
  assign y1941 = ~1'b0 ;
  assign y1942 = ~n9005 ;
  assign y1943 = n9008 ;
  assign y1944 = n9014 ;
  assign y1945 = n9018 ;
  assign y1946 = n9020 ;
  assign y1947 = n9025 ;
  assign y1948 = ~n9029 ;
  assign y1949 = ~1'b0 ;
  assign y1950 = ~n9032 ;
  assign y1951 = n9033 ;
  assign y1952 = n9034 ;
  assign y1953 = ~n9035 ;
  assign y1954 = ~n9037 ;
  assign y1955 = ~n9041 ;
  assign y1956 = ~n9045 ;
  assign y1957 = n9046 ;
  assign y1958 = ~n9049 ;
  assign y1959 = n9052 ;
  assign y1960 = n9057 ;
  assign y1961 = n9058 ;
  assign y1962 = n9068 ;
  assign y1963 = n9074 ;
  assign y1964 = ~n9075 ;
  assign y1965 = ~n9082 ;
  assign y1966 = ~n9084 ;
  assign y1967 = n9087 ;
  assign y1968 = ~n9089 ;
  assign y1969 = n9090 ;
  assign y1970 = ~1'b0 ;
  assign y1971 = ~n9094 ;
  assign y1972 = ~n9097 ;
  assign y1973 = n9098 ;
  assign y1974 = ~n9101 ;
  assign y1975 = n9125 ;
  assign y1976 = ~n9132 ;
  assign y1977 = n9136 ;
  assign y1978 = n9137 ;
  assign y1979 = ~n9139 ;
  assign y1980 = ~n9143 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = ~n9149 ;
  assign y1983 = n9153 ;
  assign y1984 = n9156 ;
  assign y1985 = n9157 ;
  assign y1986 = n9161 ;
  assign y1987 = n9163 ;
  assign y1988 = n9173 ;
  assign y1989 = ~n9175 ;
  assign y1990 = ~n9176 ;
  assign y1991 = ~n9178 ;
  assign y1992 = ~n9183 ;
  assign y1993 = n9189 ;
  assign y1994 = n9194 ;
  assign y1995 = n9210 ;
  assign y1996 = n9218 ;
  assign y1997 = n9220 ;
  assign y1998 = n9235 ;
  assign y1999 = ~1'b0 ;
  assign y2000 = n9240 ;
  assign y2001 = ~n9257 ;
  assign y2002 = n9262 ;
  assign y2003 = n9268 ;
  assign y2004 = ~n9275 ;
  assign y2005 = n9282 ;
  assign y2006 = ~n9289 ;
  assign y2007 = ~n9291 ;
  assign y2008 = ~1'b0 ;
  assign y2009 = ~n9296 ;
  assign y2010 = ~1'b0 ;
  assign y2011 = ~n9298 ;
  assign y2012 = ~n9300 ;
  assign y2013 = n9302 ;
  assign y2014 = n9304 ;
  assign y2015 = ~n9309 ;
  assign y2016 = n9323 ;
  assign y2017 = n9324 ;
  assign y2018 = ~n9326 ;
  assign y2019 = ~n9328 ;
  assign y2020 = n9332 ;
  assign y2021 = n2741 ;
  assign y2022 = n9338 ;
  assign y2023 = ~n9342 ;
  assign y2024 = n9348 ;
  assign y2025 = n9356 ;
  assign y2026 = n9360 ;
  assign y2027 = ~n9363 ;
  assign y2028 = n9368 ;
  assign y2029 = ~n9370 ;
  assign y2030 = ~n9373 ;
  assign y2031 = ~n9374 ;
  assign y2032 = n9378 ;
  assign y2033 = n9399 ;
  assign y2034 = n9412 ;
  assign y2035 = n9415 ;
  assign y2036 = n9435 ;
  assign y2037 = ~n9436 ;
  assign y2038 = ~n9437 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = n9442 ;
  assign y2041 = n9445 ;
  assign y2042 = ~n9458 ;
  assign y2043 = n9464 ;
  assign y2044 = n9469 ;
  assign y2045 = ~n9471 ;
  assign y2046 = ~n9475 ;
  assign y2047 = ~n9478 ;
  assign y2048 = ~n6676 ;
  assign y2049 = n9481 ;
  assign y2050 = ~n9488 ;
  assign y2051 = ~n9491 ;
  assign y2052 = ~n9492 ;
  assign y2053 = ~n9493 ;
  assign y2054 = ~n9506 ;
  assign y2055 = ~n9509 ;
  assign y2056 = n9519 ;
  assign y2057 = ~1'b0 ;
  assign y2058 = n9523 ;
  assign y2059 = ~n9526 ;
  assign y2060 = n9544 ;
  assign y2061 = n9547 ;
  assign y2062 = ~n9556 ;
  assign y2063 = ~1'b0 ;
  assign y2064 = ~n9562 ;
  assign y2065 = ~n9566 ;
  assign y2066 = n9569 ;
  assign y2067 = n9574 ;
  assign y2068 = ~n9584 ;
  assign y2069 = n9587 ;
  assign y2070 = n9606 ;
  assign y2071 = n9612 ;
  assign y2072 = ~n9618 ;
  assign y2073 = n9619 ;
  assign y2074 = ~n9627 ;
  assign y2075 = n9642 ;
  assign y2076 = n9649 ;
  assign y2077 = n9656 ;
  assign y2078 = n9657 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = n9658 ;
  assign y2081 = ~n9659 ;
  assign y2082 = n9661 ;
  assign y2083 = ~n9664 ;
  assign y2084 = ~n9668 ;
  assign y2085 = ~n9676 ;
  assign y2086 = n9678 ;
  assign y2087 = n9681 ;
  assign y2088 = n9689 ;
  assign y2089 = ~1'b0 ;
  assign y2090 = n9690 ;
  assign y2091 = ~n9691 ;
  assign y2092 = ~n9692 ;
  assign y2093 = ~1'b0 ;
  assign y2094 = ~n9700 ;
  assign y2095 = ~n9703 ;
  assign y2096 = ~n3505 ;
  assign y2097 = n9705 ;
  assign y2098 = n9723 ;
  assign y2099 = ~n9729 ;
  assign y2100 = ~1'b0 ;
  assign y2101 = ~n9731 ;
  assign y2102 = n9740 ;
  assign y2103 = n9741 ;
  assign y2104 = ~n9751 ;
  assign y2105 = ~n9757 ;
  assign y2106 = ~n9760 ;
  assign y2107 = n9762 ;
  assign y2108 = ~n9766 ;
  assign y2109 = n9773 ;
  assign y2110 = n9776 ;
  assign y2111 = ~n9784 ;
  assign y2112 = n9791 ;
  assign y2113 = n9792 ;
  assign y2114 = n9808 ;
  assign y2115 = ~n9814 ;
  assign y2116 = n9816 ;
  assign y2117 = ~n9820 ;
  assign y2118 = n9823 ;
  assign y2119 = n9827 ;
  assign y2120 = ~n9833 ;
  assign y2121 = n9836 ;
  assign y2122 = n9844 ;
  assign y2123 = n9846 ;
  assign y2124 = ~n9850 ;
  assign y2125 = n9852 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = n9854 ;
  assign y2128 = n9855 ;
  assign y2129 = ~n9868 ;
  assign y2130 = n9873 ;
  assign y2131 = ~1'b0 ;
  assign y2132 = ~n9885 ;
  assign y2133 = n9894 ;
  assign y2134 = n9897 ;
  assign y2135 = n9899 ;
  assign y2136 = n9906 ;
  assign y2137 = n9912 ;
  assign y2138 = n9915 ;
  assign y2139 = ~n9936 ;
  assign y2140 = ~n9937 ;
  assign y2141 = ~n9938 ;
  assign y2142 = n9945 ;
  assign y2143 = ~n9954 ;
  assign y2144 = n9958 ;
  assign y2145 = n9960 ;
  assign y2146 = ~n9961 ;
  assign y2147 = n9962 ;
  assign y2148 = n9964 ;
  assign y2149 = ~n9966 ;
  assign y2150 = ~n9967 ;
  assign y2151 = n9977 ;
  assign y2152 = ~n9990 ;
  assign y2153 = n9994 ;
  assign y2154 = n9996 ;
  assign y2155 = ~n10006 ;
  assign y2156 = ~n10008 ;
  assign y2157 = n10013 ;
  assign y2158 = ~1'b0 ;
  assign y2159 = ~n10017 ;
  assign y2160 = ~n10023 ;
  assign y2161 = ~1'b0 ;
  assign y2162 = ~n10024 ;
  assign y2163 = n10025 ;
  assign y2164 = n10027 ;
  assign y2165 = n10032 ;
  assign y2166 = n10038 ;
  assign y2167 = ~1'b0 ;
  assign y2168 = ~n10041 ;
  assign y2169 = n10047 ;
  assign y2170 = ~n10052 ;
  assign y2171 = ~n10053 ;
  assign y2172 = ~n10054 ;
  assign y2173 = n10057 ;
  assign y2174 = ~1'b0 ;
  assign y2175 = ~n10062 ;
  assign y2176 = ~n10064 ;
  assign y2177 = n10070 ;
  assign y2178 = ~n10080 ;
  assign y2179 = n10085 ;
  assign y2180 = ~n10089 ;
  assign y2181 = n10096 ;
  assign y2182 = ~n10107 ;
  assign y2183 = n10119 ;
  assign y2184 = n10128 ;
  assign y2185 = n10146 ;
  assign y2186 = ~n10151 ;
  assign y2187 = ~n10159 ;
  assign y2188 = n10162 ;
  assign y2189 = ~n10165 ;
  assign y2190 = n10171 ;
  assign y2191 = ~n10172 ;
  assign y2192 = ~n10173 ;
  assign y2193 = ~n10175 ;
  assign y2194 = n10176 ;
  assign y2195 = ~n10182 ;
  assign y2196 = n10188 ;
  assign y2197 = ~n10189 ;
  assign y2198 = n10191 ;
  assign y2199 = ~n10192 ;
  assign y2200 = n10200 ;
  assign y2201 = n10204 ;
  assign y2202 = ~1'b0 ;
  assign y2203 = ~n10225 ;
  assign y2204 = ~n10231 ;
  assign y2205 = n10233 ;
  assign y2206 = n10234 ;
  assign y2207 = n10246 ;
  assign y2208 = ~n10251 ;
  assign y2209 = ~n10256 ;
  assign y2210 = ~n10262 ;
  assign y2211 = ~n7120 ;
  assign y2212 = ~n10266 ;
  assign y2213 = ~1'b0 ;
  assign y2214 = n10270 ;
  assign y2215 = ~n10271 ;
  assign y2216 = n10272 ;
  assign y2217 = n10277 ;
  assign y2218 = n10283 ;
  assign y2219 = ~n10285 ;
  assign y2220 = ~1'b0 ;
  assign y2221 = ~n10302 ;
  assign y2222 = n10311 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = ~1'b0 ;
  assign y2225 = ~1'b0 ;
  assign y2226 = ~n10315 ;
  assign y2227 = ~n10330 ;
  assign y2228 = ~n10332 ;
  assign y2229 = n10342 ;
  assign y2230 = ~n10347 ;
  assign y2231 = ~n10353 ;
  assign y2232 = ~n10359 ;
  assign y2233 = ~n10360 ;
  assign y2234 = n10363 ;
  assign y2235 = n10366 ;
  assign y2236 = ~n10368 ;
  assign y2237 = ~n10375 ;
  assign y2238 = ~n10379 ;
  assign y2239 = n10386 ;
  assign y2240 = ~n10388 ;
  assign y2241 = ~n10393 ;
  assign y2242 = n10400 ;
  assign y2243 = ~n10402 ;
  assign y2244 = n10416 ;
  assign y2245 = n10423 ;
  assign y2246 = ~n10424 ;
  assign y2247 = n10425 ;
  assign y2248 = n10428 ;
  assign y2249 = ~n10435 ;
  assign y2250 = ~1'b0 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = n10436 ;
  assign y2253 = ~n10438 ;
  assign y2254 = n10453 ;
  assign y2255 = n10455 ;
  assign y2256 = ~n10456 ;
  assign y2257 = n10464 ;
  assign y2258 = n10468 ;
  assign y2259 = ~n10469 ;
  assign y2260 = ~n10474 ;
  assign y2261 = n10479 ;
  assign y2262 = n10483 ;
  assign y2263 = ~n10485 ;
  assign y2264 = ~n10499 ;
  assign y2265 = ~n10502 ;
  assign y2266 = ~n10508 ;
  assign y2267 = ~n10519 ;
  assign y2268 = n10520 ;
  assign y2269 = ~n10527 ;
  assign y2270 = n10528 ;
  assign y2271 = n10529 ;
  assign y2272 = ~n10532 ;
  assign y2273 = ~n10536 ;
  assign y2274 = n10542 ;
  assign y2275 = ~n10543 ;
  assign y2276 = ~n10546 ;
  assign y2277 = n10548 ;
  assign y2278 = ~n10554 ;
  assign y2279 = n10555 ;
  assign y2280 = n4277 ;
  assign y2281 = n10556 ;
  assign y2282 = ~n10566 ;
  assign y2283 = ~n10575 ;
  assign y2284 = n10580 ;
  assign y2285 = n10581 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n10585 ;
  assign y2288 = ~n10586 ;
  assign y2289 = ~1'b0 ;
  assign y2290 = n10591 ;
  assign y2291 = ~1'b0 ;
  assign y2292 = ~1'b0 ;
  assign y2293 = ~n10592 ;
  assign y2294 = n10595 ;
  assign y2295 = ~n10599 ;
  assign y2296 = n10603 ;
  assign y2297 = n10607 ;
  assign y2298 = n10613 ;
  assign y2299 = ~1'b0 ;
  assign y2300 = n10620 ;
  assign y2301 = ~n10636 ;
  assign y2302 = n10640 ;
  assign y2303 = n10655 ;
  assign y2304 = n10662 ;
  assign y2305 = ~n10669 ;
  assign y2306 = 1'b0 ;
  assign y2307 = ~n10673 ;
  assign y2308 = n10677 ;
  assign y2309 = n10679 ;
  assign y2310 = ~1'b0 ;
  assign y2311 = n10681 ;
  assign y2312 = ~n10693 ;
  assign y2313 = n10698 ;
  assign y2314 = ~n10708 ;
  assign y2315 = n10709 ;
  assign y2316 = n10710 ;
  assign y2317 = ~n10713 ;
  assign y2318 = ~n10714 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = ~n10715 ;
  assign y2321 = ~n10719 ;
  assign y2322 = ~n10728 ;
  assign y2323 = n10729 ;
  assign y2324 = ~n10730 ;
  assign y2325 = n10745 ;
  assign y2326 = n10757 ;
  assign y2327 = ~n10759 ;
  assign y2328 = ~n10761 ;
  assign y2329 = ~1'b0 ;
  assign y2330 = ~n10769 ;
  assign y2331 = ~n10772 ;
  assign y2332 = ~n10781 ;
  assign y2333 = ~n10785 ;
  assign y2334 = n10795 ;
  assign y2335 = ~n10802 ;
  assign y2336 = ~n10805 ;
  assign y2337 = n10809 ;
  assign y2338 = n7859 ;
  assign y2339 = n10811 ;
  assign y2340 = ~n10816 ;
  assign y2341 = ~1'b0 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = ~n10822 ;
  assign y2344 = n10824 ;
  assign y2345 = ~n10830 ;
  assign y2346 = n10832 ;
  assign y2347 = ~n10843 ;
  assign y2348 = n10851 ;
  assign y2349 = n10862 ;
  assign y2350 = ~n10866 ;
  assign y2351 = ~1'b0 ;
  assign y2352 = ~n10868 ;
  assign y2353 = ~n10869 ;
  assign y2354 = n10870 ;
  assign y2355 = ~n10872 ;
  assign y2356 = n10876 ;
  assign y2357 = ~n10877 ;
  assign y2358 = ~n10889 ;
  assign y2359 = n10900 ;
  assign y2360 = ~n10902 ;
  assign y2361 = ~n10905 ;
  assign y2362 = n10906 ;
  assign y2363 = n10908 ;
  assign y2364 = n10919 ;
  assign y2365 = n10920 ;
  assign y2366 = n10926 ;
  assign y2367 = n10931 ;
  assign y2368 = n10937 ;
  assign y2369 = n10961 ;
  assign y2370 = n10968 ;
  assign y2371 = ~n10971 ;
  assign y2372 = ~n10978 ;
  assign y2373 = ~n10988 ;
  assign y2374 = ~n10989 ;
  assign y2375 = n10995 ;
  assign y2376 = n11002 ;
  assign y2377 = ~1'b0 ;
  assign y2378 = ~n11005 ;
  assign y2379 = ~n11010 ;
  assign y2380 = ~n11014 ;
  assign y2381 = ~n11025 ;
  assign y2382 = ~n11026 ;
  assign y2383 = ~1'b0 ;
  assign y2384 = ~n11032 ;
  assign y2385 = n11036 ;
  assign y2386 = ~n11038 ;
  assign y2387 = ~n11042 ;
  assign y2388 = n11046 ;
  assign y2389 = ~1'b0 ;
  assign y2390 = ~n11056 ;
  assign y2391 = ~n11058 ;
  assign y2392 = ~n11061 ;
  assign y2393 = n11069 ;
  assign y2394 = n11079 ;
  assign y2395 = ~n11082 ;
  assign y2396 = n11087 ;
  assign y2397 = n11090 ;
  assign y2398 = n11095 ;
  assign y2399 = ~n11098 ;
  assign y2400 = ~n11100 ;
  assign y2401 = ~1'b0 ;
  assign y2402 = n11101 ;
  assign y2403 = n11111 ;
  assign y2404 = ~n11113 ;
  assign y2405 = n11115 ;
  assign y2406 = n11116 ;
  assign y2407 = ~n11118 ;
  assign y2408 = ~n11122 ;
  assign y2409 = n11135 ;
  assign y2410 = ~n11146 ;
  assign y2411 = n11159 ;
  assign y2412 = n11161 ;
  assign y2413 = ~n11168 ;
  assign y2414 = n11190 ;
  assign y2415 = n11194 ;
  assign y2416 = ~n11197 ;
  assign y2417 = ~1'b0 ;
  assign y2418 = ~n11200 ;
  assign y2419 = ~n11203 ;
  assign y2420 = ~1'b0 ;
  assign y2421 = ~n11204 ;
  assign y2422 = ~1'b0 ;
  assign y2423 = n11207 ;
  assign y2424 = ~1'b0 ;
  assign y2425 = ~n11211 ;
  assign y2426 = n11223 ;
  assign y2427 = n11225 ;
  assign y2428 = n11228 ;
  assign y2429 = ~n11234 ;
  assign y2430 = ~n11235 ;
  assign y2431 = ~n11239 ;
  assign y2432 = n11248 ;
  assign y2433 = ~n11254 ;
  assign y2434 = n11257 ;
  assign y2435 = ~n11260 ;
  assign y2436 = ~n11263 ;
  assign y2437 = ~n11265 ;
  assign y2438 = n11266 ;
  assign y2439 = ~n11273 ;
  assign y2440 = n11280 ;
  assign y2441 = n11288 ;
  assign y2442 = n11295 ;
  assign y2443 = n11297 ;
  assign y2444 = n11298 ;
  assign y2445 = n11308 ;
  assign y2446 = n11309 ;
  assign y2447 = n11321 ;
  assign y2448 = n11327 ;
  assign y2449 = n11329 ;
  assign y2450 = ~n11332 ;
  assign y2451 = n11333 ;
  assign y2452 = n11340 ;
  assign y2453 = n11344 ;
  assign y2454 = ~n11351 ;
  assign y2455 = n11352 ;
  assign y2456 = ~n11355 ;
  assign y2457 = ~n11360 ;
  assign y2458 = n11361 ;
  assign y2459 = ~n11365 ;
  assign y2460 = ~1'b0 ;
  assign y2461 = n11371 ;
  assign y2462 = ~n11381 ;
  assign y2463 = n11386 ;
  assign y2464 = ~n11387 ;
  assign y2465 = ~n11395 ;
  assign y2466 = n11398 ;
  assign y2467 = ~n11403 ;
  assign y2468 = n11405 ;
  assign y2469 = ~n11410 ;
  assign y2470 = ~n11425 ;
  assign y2471 = ~n11427 ;
  assign y2472 = ~n11435 ;
  assign y2473 = ~n11439 ;
  assign y2474 = n11444 ;
  assign y2475 = n11445 ;
  assign y2476 = ~n11446 ;
  assign y2477 = ~n11453 ;
  assign y2478 = ~n11463 ;
  assign y2479 = n11464 ;
  assign y2480 = n11473 ;
  assign y2481 = ~n11480 ;
  assign y2482 = n11484 ;
  assign y2483 = ~n11485 ;
  assign y2484 = ~n11489 ;
  assign y2485 = n11498 ;
  assign y2486 = ~1'b0 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = n11515 ;
  assign y2489 = n11519 ;
  assign y2490 = ~n11522 ;
  assign y2491 = n11528 ;
  assign y2492 = n11531 ;
  assign y2493 = ~n11532 ;
  assign y2494 = ~n11538 ;
  assign y2495 = ~n11539 ;
  assign y2496 = n11542 ;
  assign y2497 = ~1'b0 ;
  assign y2498 = ~n11546 ;
  assign y2499 = ~n11550 ;
  assign y2500 = ~n11552 ;
  assign y2501 = ~n11559 ;
  assign y2502 = n11561 ;
  assign y2503 = ~n11566 ;
  assign y2504 = n11579 ;
  assign y2505 = ~n11582 ;
  assign y2506 = ~1'b0 ;
  assign y2507 = ~n11584 ;
  assign y2508 = ~n11586 ;
  assign y2509 = ~1'b0 ;
  assign y2510 = ~n11588 ;
  assign y2511 = ~n11594 ;
  assign y2512 = n11600 ;
  assign y2513 = ~n11601 ;
  assign y2514 = ~n11602 ;
  assign y2515 = ~1'b0 ;
  assign y2516 = n11613 ;
  assign y2517 = ~n11616 ;
  assign y2518 = ~n11622 ;
  assign y2519 = ~1'b0 ;
  assign y2520 = ~n11624 ;
  assign y2521 = n11632 ;
  assign y2522 = n11635 ;
  assign y2523 = ~n11641 ;
  assign y2524 = n11649 ;
  assign y2525 = n11662 ;
  assign y2526 = ~n11663 ;
  assign y2527 = n11668 ;
  assign y2528 = n11677 ;
  assign y2529 = ~n11687 ;
  assign y2530 = n11691 ;
  assign y2531 = n11698 ;
  assign y2532 = ~n11700 ;
  assign y2533 = ~n11705 ;
  assign y2534 = ~1'b0 ;
  assign y2535 = n11707 ;
  assign y2536 = ~1'b0 ;
  assign y2537 = n11710 ;
  assign y2538 = n11712 ;
  assign y2539 = n11716 ;
  assign y2540 = n11720 ;
  assign y2541 = n11731 ;
  assign y2542 = ~n11733 ;
  assign y2543 = ~n11744 ;
  assign y2544 = n11759 ;
  assign y2545 = n11764 ;
  assign y2546 = n11765 ;
  assign y2547 = n11770 ;
  assign y2548 = ~1'b0 ;
  assign y2549 = ~1'b0 ;
  assign y2550 = ~1'b0 ;
  assign y2551 = n11771 ;
  assign y2552 = n11776 ;
  assign y2553 = n11778 ;
  assign y2554 = ~n11783 ;
  assign y2555 = n11791 ;
  assign y2556 = ~1'b0 ;
  assign y2557 = n11793 ;
  assign y2558 = ~n11796 ;
  assign y2559 = ~n11801 ;
  assign y2560 = ~n11806 ;
  assign y2561 = ~n11808 ;
  assign y2562 = n11815 ;
  assign y2563 = ~1'b0 ;
  assign y2564 = n11819 ;
  assign y2565 = n11823 ;
  assign y2566 = n11830 ;
  assign y2567 = ~n11836 ;
  assign y2568 = ~n11844 ;
  assign y2569 = ~n11847 ;
  assign y2570 = ~n11848 ;
  assign y2571 = ~n11849 ;
  assign y2572 = ~1'b0 ;
  assign y2573 = n11857 ;
  assign y2574 = ~n11859 ;
  assign y2575 = n11865 ;
  assign y2576 = ~1'b0 ;
  assign y2577 = ~n11869 ;
  assign y2578 = n3044 ;
  assign y2579 = ~1'b0 ;
  assign y2580 = n11874 ;
  assign y2581 = n11877 ;
  assign y2582 = n11898 ;
  assign y2583 = ~n11900 ;
  assign y2584 = n11903 ;
  assign y2585 = n11906 ;
  assign y2586 = n11910 ;
  assign y2587 = ~n11922 ;
  assign y2588 = ~n11925 ;
  assign y2589 = ~n11930 ;
  assign y2590 = ~n11937 ;
  assign y2591 = ~n11953 ;
  assign y2592 = n11957 ;
  assign y2593 = ~n11958 ;
  assign y2594 = n11966 ;
  assign y2595 = ~1'b0 ;
  assign y2596 = ~n11968 ;
  assign y2597 = n11973 ;
  assign y2598 = n11986 ;
  assign y2599 = ~n11993 ;
  assign y2600 = ~n11994 ;
  assign y2601 = n11995 ;
  assign y2602 = n11996 ;
  assign y2603 = ~1'b0 ;
  assign y2604 = ~n11998 ;
  assign y2605 = ~n12006 ;
  assign y2606 = ~n12018 ;
  assign y2607 = ~1'b0 ;
  assign y2608 = n12021 ;
  assign y2609 = n12023 ;
  assign y2610 = n12027 ;
  assign y2611 = ~n12031 ;
  assign y2612 = ~1'b0 ;
  assign y2613 = ~1'b0 ;
  assign y2614 = ~n12038 ;
  assign y2615 = n12039 ;
  assign y2616 = n12043 ;
  assign y2617 = ~n12048 ;
  assign y2618 = ~n12057 ;
  assign y2619 = n12058 ;
  assign y2620 = n12071 ;
  assign y2621 = ~n12080 ;
  assign y2622 = ~n12089 ;
  assign y2623 = ~n12099 ;
  assign y2624 = ~n12104 ;
  assign y2625 = ~1'b0 ;
  assign y2626 = n12110 ;
  assign y2627 = n12111 ;
  assign y2628 = ~n12115 ;
  assign y2629 = ~n12130 ;
  assign y2630 = ~n12140 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = ~n12144 ;
  assign y2633 = ~n12147 ;
  assign y2634 = ~n12148 ;
  assign y2635 = n12149 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = ~n12155 ;
  assign y2638 = n12174 ;
  assign y2639 = ~n12175 ;
  assign y2640 = ~1'b0 ;
  assign y2641 = ~n12179 ;
  assign y2642 = ~1'b0 ;
  assign y2643 = n12180 ;
  assign y2644 = n12181 ;
  assign y2645 = n12183 ;
  assign y2646 = ~n12186 ;
  assign y2647 = n12194 ;
  assign y2648 = n12198 ;
  assign y2649 = n12199 ;
  assign y2650 = ~n12203 ;
  assign y2651 = ~n12208 ;
  assign y2652 = n12210 ;
  assign y2653 = ~n12214 ;
  assign y2654 = ~1'b0 ;
  assign y2655 = ~n12224 ;
  assign y2656 = n12233 ;
  assign y2657 = n12245 ;
  assign y2658 = n12254 ;
  assign y2659 = ~n12255 ;
  assign y2660 = n12264 ;
  assign y2661 = ~n12266 ;
  assign y2662 = n12268 ;
  assign y2663 = n12271 ;
  assign y2664 = n12273 ;
  assign y2665 = n12288 ;
  assign y2666 = ~n12291 ;
  assign y2667 = ~1'b0 ;
  assign y2668 = ~n12292 ;
  assign y2669 = ~1'b0 ;
  assign y2670 = ~n12298 ;
  assign y2671 = n12305 ;
  assign y2672 = ~n12315 ;
  assign y2673 = ~n12322 ;
  assign y2674 = ~n12324 ;
  assign y2675 = ~n12325 ;
  assign y2676 = ~n12326 ;
  assign y2677 = ~1'b0 ;
  assign y2678 = ~n12329 ;
  assign y2679 = n12331 ;
  assign y2680 = ~n12332 ;
  assign y2681 = ~n12373 ;
  assign y2682 = ~n12377 ;
  assign y2683 = ~n12389 ;
  assign y2684 = ~n12404 ;
  assign y2685 = ~n12407 ;
  assign y2686 = n12411 ;
  assign y2687 = 1'b0 ;
  assign y2688 = ~n12414 ;
  assign y2689 = ~1'b0 ;
  assign y2690 = n12416 ;
  assign y2691 = ~n12418 ;
  assign y2692 = ~n12422 ;
  assign y2693 = ~1'b0 ;
  assign y2694 = ~n12425 ;
  assign y2695 = n12428 ;
  assign y2696 = ~1'b0 ;
  assign y2697 = n12434 ;
  assign y2698 = n12440 ;
  assign y2699 = ~n12445 ;
  assign y2700 = ~1'b0 ;
  assign y2701 = ~n12447 ;
  assign y2702 = ~n12453 ;
  assign y2703 = ~n12458 ;
  assign y2704 = ~n12461 ;
  assign y2705 = ~n12466 ;
  assign y2706 = ~n12470 ;
  assign y2707 = ~n12471 ;
  assign y2708 = n12477 ;
  assign y2709 = ~n12486 ;
  assign y2710 = n12490 ;
  assign y2711 = ~n12491 ;
  assign y2712 = n12495 ;
  assign y2713 = ~n12500 ;
  assign y2714 = ~n12503 ;
  assign y2715 = ~1'b0 ;
  assign y2716 = n12505 ;
  assign y2717 = ~n12508 ;
  assign y2718 = n12513 ;
  assign y2719 = ~1'b0 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = n12520 ;
  assign y2722 = n12529 ;
  assign y2723 = ~n12530 ;
  assign y2724 = n12531 ;
  assign y2725 = n12536 ;
  assign y2726 = n12540 ;
  assign y2727 = ~n12542 ;
  assign y2728 = ~n12546 ;
  assign y2729 = n12548 ;
  assign y2730 = ~n12555 ;
  assign y2731 = n12569 ;
  assign y2732 = n12573 ;
  assign y2733 = ~n12580 ;
  assign y2734 = ~n12585 ;
  assign y2735 = ~n12590 ;
  assign y2736 = n12591 ;
  assign y2737 = ~n12601 ;
  assign y2738 = ~1'b0 ;
  assign y2739 = ~n12605 ;
  assign y2740 = n12608 ;
  assign y2741 = ~n12610 ;
  assign y2742 = n12616 ;
  assign y2743 = ~n12619 ;
  assign y2744 = ~1'b0 ;
  assign y2745 = ~1'b0 ;
  assign y2746 = n12631 ;
  assign y2747 = n12638 ;
  assign y2748 = ~n12639 ;
  assign y2749 = n12648 ;
  assign y2750 = n12651 ;
  assign y2751 = ~n12654 ;
  assign y2752 = n12664 ;
  assign y2753 = n12667 ;
  assign y2754 = n12668 ;
  assign y2755 = ~n12671 ;
  assign y2756 = ~n12672 ;
  assign y2757 = ~1'b0 ;
  assign y2758 = ~n12674 ;
  assign y2759 = ~n12682 ;
  assign y2760 = ~n12694 ;
  assign y2761 = n12695 ;
  assign y2762 = ~n12706 ;
  assign y2763 = ~n12714 ;
  assign y2764 = ~1'b0 ;
  assign y2765 = ~n12715 ;
  assign y2766 = n12721 ;
  assign y2767 = n12735 ;
  assign y2768 = ~n12737 ;
  assign y2769 = ~n12744 ;
  assign y2770 = ~n12761 ;
  assign y2771 = n12766 ;
  assign y2772 = n12771 ;
  assign y2773 = n12775 ;
  assign y2774 = n12778 ;
  assign y2775 = ~1'b0 ;
  assign y2776 = n12779 ;
  assign y2777 = n12783 ;
  assign y2778 = n12785 ;
  assign y2779 = n12794 ;
  assign y2780 = n12798 ;
  assign y2781 = n12809 ;
  assign y2782 = ~n12813 ;
  assign y2783 = ~n12817 ;
  assign y2784 = n12821 ;
  assign y2785 = ~n12822 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = ~n12826 ;
  assign y2788 = n12828 ;
  assign y2789 = n12832 ;
  assign y2790 = n12834 ;
  assign y2791 = n12837 ;
  assign y2792 = ~n12839 ;
  assign y2793 = ~n12859 ;
  assign y2794 = n12866 ;
  assign y2795 = ~n12868 ;
  assign y2796 = ~n12871 ;
  assign y2797 = ~n12885 ;
  assign y2798 = n12891 ;
  assign y2799 = ~n12895 ;
  assign y2800 = ~1'b0 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = ~n12897 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = n12911 ;
  assign y2805 = n12912 ;
  assign y2806 = ~1'b0 ;
  assign y2807 = ~n12915 ;
  assign y2808 = ~n12916 ;
  assign y2809 = n12921 ;
  assign y2810 = n12930 ;
  assign y2811 = ~n12933 ;
  assign y2812 = ~1'b0 ;
  assign y2813 = ~1'b0 ;
  assign y2814 = ~n12935 ;
  assign y2815 = n12937 ;
  assign y2816 = n12941 ;
  assign y2817 = ~n12943 ;
  assign y2818 = n12964 ;
  assign y2819 = ~n12967 ;
  assign y2820 = n12973 ;
  assign y2821 = ~n12982 ;
  assign y2822 = ~n12983 ;
  assign y2823 = n12989 ;
  assign y2824 = ~n12991 ;
  assign y2825 = n12999 ;
  assign y2826 = n13005 ;
  assign y2827 = n13006 ;
  assign y2828 = ~n13011 ;
  assign y2829 = n13013 ;
  assign y2830 = ~n13018 ;
  assign y2831 = ~1'b0 ;
  assign y2832 = ~1'b0 ;
  assign y2833 = n13024 ;
  assign y2834 = ~1'b0 ;
  assign y2835 = n13025 ;
  assign y2836 = n13034 ;
  assign y2837 = ~n13035 ;
  assign y2838 = ~n13040 ;
  assign y2839 = n13048 ;
  assign y2840 = n13049 ;
  assign y2841 = n13051 ;
  assign y2842 = n13059 ;
  assign y2843 = n13064 ;
  assign y2844 = n13068 ;
  assign y2845 = n13075 ;
  assign y2846 = ~n13081 ;
  assign y2847 = ~n13083 ;
  assign y2848 = n13085 ;
  assign y2849 = ~n13088 ;
  assign y2850 = n13097 ;
  assign y2851 = n13099 ;
  assign y2852 = n13101 ;
  assign y2853 = ~n13107 ;
  assign y2854 = ~1'b0 ;
  assign y2855 = ~n13113 ;
  assign y2856 = n13118 ;
  assign y2857 = n13119 ;
  assign y2858 = n13120 ;
  assign y2859 = ~1'b0 ;
  assign y2860 = n13122 ;
  assign y2861 = n13124 ;
  assign y2862 = n13128 ;
  assign y2863 = ~n13129 ;
  assign y2864 = n13137 ;
  assign y2865 = n13141 ;
  assign y2866 = n13143 ;
  assign y2867 = n13153 ;
  assign y2868 = ~n13155 ;
  assign y2869 = ~n13157 ;
  assign y2870 = ~n13165 ;
  assign y2871 = n13167 ;
  assign y2872 = ~1'b0 ;
  assign y2873 = ~1'b0 ;
  assign y2874 = ~n13169 ;
  assign y2875 = ~1'b0 ;
  assign y2876 = n13174 ;
  assign y2877 = n13185 ;
  assign y2878 = n13188 ;
  assign y2879 = ~n13198 ;
  assign y2880 = ~n13199 ;
  assign y2881 = n13204 ;
  assign y2882 = n13214 ;
  assign y2883 = n13215 ;
  assign y2884 = n13222 ;
  assign y2885 = n13226 ;
  assign y2886 = ~n13229 ;
  assign y2887 = ~1'b0 ;
  assign y2888 = n13233 ;
  assign y2889 = n13236 ;
  assign y2890 = ~n13237 ;
  assign y2891 = ~n13253 ;
  assign y2892 = ~1'b0 ;
  assign y2893 = ~n13260 ;
  assign y2894 = n13261 ;
  assign y2895 = ~n13262 ;
  assign y2896 = n13287 ;
  assign y2897 = n13288 ;
  assign y2898 = ~n13289 ;
  assign y2899 = n13301 ;
  assign y2900 = ~n13305 ;
  assign y2901 = n13311 ;
  assign y2902 = ~n13312 ;
  assign y2903 = ~n13317 ;
  assign y2904 = ~n13323 ;
  assign y2905 = ~n13326 ;
  assign y2906 = n13327 ;
  assign y2907 = n13328 ;
  assign y2908 = ~n13330 ;
  assign y2909 = ~n13344 ;
  assign y2910 = n13350 ;
  assign y2911 = n13352 ;
  assign y2912 = ~n13360 ;
  assign y2913 = n13365 ;
  assign y2914 = ~n13377 ;
  assign y2915 = ~1'b0 ;
  assign y2916 = n13383 ;
  assign y2917 = ~1'b0 ;
  assign y2918 = n13389 ;
  assign y2919 = n13401 ;
  assign y2920 = n13402 ;
  assign y2921 = ~1'b0 ;
  assign y2922 = ~n13420 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = n13423 ;
  assign y2925 = ~n13431 ;
  assign y2926 = ~n13432 ;
  assign y2927 = n13440 ;
  assign y2928 = ~n13444 ;
  assign y2929 = ~n13445 ;
  assign y2930 = n13446 ;
  assign y2931 = ~n13452 ;
  assign y2932 = ~n13454 ;
  assign y2933 = n13456 ;
  assign y2934 = n13457 ;
  assign y2935 = ~n13462 ;
  assign y2936 = ~n13479 ;
  assign y2937 = ~n13485 ;
  assign y2938 = n13491 ;
  assign y2939 = ~n13495 ;
  assign y2940 = ~n13507 ;
  assign y2941 = n13509 ;
  assign y2942 = ~1'b0 ;
  assign y2943 = ~n13515 ;
  assign y2944 = ~1'b0 ;
  assign y2945 = ~n13517 ;
  assign y2946 = ~n13519 ;
  assign y2947 = ~n13520 ;
  assign y2948 = n13526 ;
  assign y2949 = ~n13528 ;
  assign y2950 = ~n13534 ;
  assign y2951 = ~n13535 ;
  assign y2952 = n13541 ;
  assign y2953 = ~n13544 ;
  assign y2954 = ~n13549 ;
  assign y2955 = n13557 ;
  assign y2956 = n13560 ;
  assign y2957 = ~n13561 ;
  assign y2958 = ~n13570 ;
  assign y2959 = n13571 ;
  assign y2960 = ~1'b0 ;
  assign y2961 = n13591 ;
  assign y2962 = ~n13598 ;
  assign y2963 = ~n13599 ;
  assign y2964 = ~n13604 ;
  assign y2965 = n13607 ;
  assign y2966 = ~n13612 ;
  assign y2967 = n13620 ;
  assign y2968 = ~n13623 ;
  assign y2969 = ~n13629 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = ~n13633 ;
  assign y2972 = ~n13638 ;
  assign y2973 = ~n13643 ;
  assign y2974 = ~n13649 ;
  assign y2975 = ~n13653 ;
  assign y2976 = ~1'b0 ;
  assign y2977 = ~n13656 ;
  assign y2978 = ~n13659 ;
  assign y2979 = ~n13662 ;
  assign y2980 = ~n13663 ;
  assign y2981 = ~1'b0 ;
  assign y2982 = n13669 ;
  assign y2983 = n13680 ;
  assign y2984 = n13685 ;
  assign y2985 = ~n13698 ;
  assign y2986 = ~n13702 ;
  assign y2987 = ~n13708 ;
  assign y2988 = ~1'b0 ;
  assign y2989 = n13714 ;
  assign y2990 = ~n13717 ;
  assign y2991 = ~n13728 ;
  assign y2992 = n13729 ;
  assign y2993 = n13738 ;
  assign y2994 = ~n13743 ;
  assign y2995 = n13748 ;
  assign y2996 = n13750 ;
  assign y2997 = n13753 ;
  assign y2998 = ~1'b0 ;
  assign y2999 = n13754 ;
  assign y3000 = n13755 ;
  assign y3001 = n13760 ;
  assign y3002 = ~1'b0 ;
  assign y3003 = n13770 ;
  assign y3004 = ~n13771 ;
  assign y3005 = ~n13772 ;
  assign y3006 = n13775 ;
  assign y3007 = ~n13778 ;
  assign y3008 = ~n13790 ;
  assign y3009 = ~n13797 ;
  assign y3010 = n13802 ;
  assign y3011 = n13807 ;
  assign y3012 = ~n13809 ;
  assign y3013 = n13816 ;
  assign y3014 = n13819 ;
  assign y3015 = ~n13820 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = n13830 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = ~n13835 ;
  assign y3020 = n13841 ;
  assign y3021 = n13846 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = n13848 ;
  assign y3024 = ~n13853 ;
  assign y3025 = n13857 ;
  assign y3026 = ~n13866 ;
  assign y3027 = n13868 ;
  assign y3028 = n13872 ;
  assign y3029 = n13881 ;
  assign y3030 = ~n13886 ;
  assign y3031 = n13887 ;
  assign y3032 = n13891 ;
  assign y3033 = ~n13897 ;
  assign y3034 = ~n2021 ;
  assign y3035 = n13898 ;
  assign y3036 = ~n13900 ;
  assign y3037 = ~1'b0 ;
  assign y3038 = ~n13901 ;
  assign y3039 = n13903 ;
  assign y3040 = n13905 ;
  assign y3041 = n13907 ;
  assign y3042 = n13915 ;
  assign y3043 = n13927 ;
  assign y3044 = n13937 ;
  assign y3045 = ~n13943 ;
  assign y3046 = n13946 ;
  assign y3047 = ~n13947 ;
  assign y3048 = n13952 ;
  assign y3049 = ~n13959 ;
  assign y3050 = n13965 ;
  assign y3051 = n13972 ;
  assign y3052 = ~n13973 ;
  assign y3053 = ~n13983 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = n13986 ;
  assign y3056 = ~n13990 ;
  assign y3057 = ~n13993 ;
  assign y3058 = n13997 ;
  assign y3059 = ~n14000 ;
  assign y3060 = n14003 ;
  assign y3061 = n14004 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = n14013 ;
  assign y3064 = n14018 ;
  assign y3065 = ~n14022 ;
  assign y3066 = ~n14028 ;
  assign y3067 = ~n14041 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = n14043 ;
  assign y3070 = ~n5684 ;
  assign y3071 = ~n14052 ;
  assign y3072 = n14055 ;
  assign y3073 = n14056 ;
  assign y3074 = n14068 ;
  assign y3075 = n14076 ;
  assign y3076 = ~n14077 ;
  assign y3077 = ~n14083 ;
  assign y3078 = n14091 ;
  assign y3079 = ~n14100 ;
  assign y3080 = n14101 ;
  assign y3081 = ~n14103 ;
  assign y3082 = n14107 ;
  assign y3083 = ~n14113 ;
  assign y3084 = ~n14125 ;
  assign y3085 = ~n14128 ;
  assign y3086 = n14147 ;
  assign y3087 = ~n12118 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = n14148 ;
  assign y3090 = ~n14163 ;
  assign y3091 = n14183 ;
  assign y3092 = ~n14190 ;
  assign y3093 = ~n14193 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = ~n14198 ;
  assign y3096 = n14207 ;
  assign y3097 = ~n14210 ;
  assign y3098 = ~1'b0 ;
  assign y3099 = ~n14211 ;
  assign y3100 = ~n14213 ;
  assign y3101 = ~n14219 ;
  assign y3102 = ~n14228 ;
  assign y3103 = ~n14229 ;
  assign y3104 = n14231 ;
  assign y3105 = n14239 ;
  assign y3106 = ~n14241 ;
  assign y3107 = ~1'b0 ;
  assign y3108 = ~n14247 ;
  assign y3109 = n14248 ;
  assign y3110 = ~n14253 ;
  assign y3111 = ~n14259 ;
  assign y3112 = ~n14265 ;
  assign y3113 = n14272 ;
  assign y3114 = ~n14274 ;
  assign y3115 = ~n14277 ;
  assign y3116 = n14289 ;
  assign y3117 = ~n14291 ;
  assign y3118 = ~n14293 ;
  assign y3119 = ~n14294 ;
  assign y3120 = n14298 ;
  assign y3121 = ~n14299 ;
  assign y3122 = ~n14315 ;
  assign y3123 = ~n14319 ;
  assign y3124 = n14322 ;
  assign y3125 = n14327 ;
  assign y3126 = ~1'b0 ;
  assign y3127 = n14330 ;
  assign y3128 = n14332 ;
  assign y3129 = n14333 ;
  assign y3130 = n14342 ;
  assign y3131 = ~n14347 ;
  assign y3132 = n14351 ;
  assign y3133 = n14354 ;
  assign y3134 = n14356 ;
  assign y3135 = ~n14358 ;
  assign y3136 = ~n14363 ;
  assign y3137 = n14365 ;
  assign y3138 = n14368 ;
  assign y3139 = ~n14370 ;
  assign y3140 = ~n1808 ;
  assign y3141 = n14373 ;
  assign y3142 = ~n14385 ;
  assign y3143 = ~n14386 ;
  assign y3144 = ~n14393 ;
  assign y3145 = ~n14394 ;
  assign y3146 = ~n14396 ;
  assign y3147 = n14403 ;
  assign y3148 = ~n14407 ;
  assign y3149 = n14412 ;
  assign y3150 = n14415 ;
  assign y3151 = ~n14417 ;
  assign y3152 = ~n14418 ;
  assign y3153 = ~n14425 ;
  assign y3154 = n14427 ;
  assign y3155 = ~n14431 ;
  assign y3156 = ~n14433 ;
  assign y3157 = n14439 ;
  assign y3158 = n14442 ;
  assign y3159 = ~n14450 ;
  assign y3160 = ~n14452 ;
  assign y3161 = n14457 ;
  assign y3162 = n14463 ;
  assign y3163 = ~n14464 ;
  assign y3164 = ~n14465 ;
  assign y3165 = ~n14478 ;
  assign y3166 = n14488 ;
  assign y3167 = ~n14494 ;
  assign y3168 = ~n14496 ;
  assign y3169 = ~n14499 ;
  assign y3170 = ~n14501 ;
  assign y3171 = n14503 ;
  assign y3172 = ~n14506 ;
  assign y3173 = ~n14511 ;
  assign y3174 = ~n14514 ;
  assign y3175 = ~n14524 ;
  assign y3176 = n14530 ;
  assign y3177 = n14538 ;
  assign y3178 = n14541 ;
  assign y3179 = n14542 ;
  assign y3180 = ~1'b0 ;
  assign y3181 = ~1'b0 ;
  assign y3182 = n14547 ;
  assign y3183 = 1'b0 ;
  assign y3184 = ~n14553 ;
  assign y3185 = n14559 ;
  assign y3186 = n14562 ;
  assign y3187 = n14565 ;
  assign y3188 = n14568 ;
  assign y3189 = n14574 ;
  assign y3190 = ~n14582 ;
  assign y3191 = ~1'b0 ;
  assign y3192 = ~n14591 ;
  assign y3193 = ~n12124 ;
  assign y3194 = n14597 ;
  assign y3195 = n14598 ;
  assign y3196 = n14607 ;
  assign y3197 = ~n14609 ;
  assign y3198 = n14614 ;
  assign y3199 = ~n14617 ;
  assign y3200 = ~n14627 ;
  assign y3201 = ~n14636 ;
  assign y3202 = ~n14638 ;
  assign y3203 = ~n14640 ;
  assign y3204 = ~n14642 ;
  assign y3205 = n14646 ;
  assign y3206 = n14647 ;
  assign y3207 = n14651 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = ~n14652 ;
  assign y3210 = n14654 ;
  assign y3211 = ~n14656 ;
  assign y3212 = ~n14659 ;
  assign y3213 = n14663 ;
  assign y3214 = n14671 ;
  assign y3215 = ~n14672 ;
  assign y3216 = ~n14677 ;
  assign y3217 = n14686 ;
  assign y3218 = ~n14689 ;
  assign y3219 = n14693 ;
  assign y3220 = ~n14694 ;
  assign y3221 = ~n14698 ;
  assign y3222 = ~n14706 ;
  assign y3223 = ~n14718 ;
  assign y3224 = ~n14724 ;
  assign y3225 = ~n14734 ;
  assign y3226 = n14741 ;
  assign y3227 = ~1'b0 ;
  assign y3228 = ~n14748 ;
  assign y3229 = ~n14758 ;
  assign y3230 = ~n14764 ;
  assign y3231 = ~1'b0 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = ~n14765 ;
  assign y3234 = n14771 ;
  assign y3235 = ~n14774 ;
  assign y3236 = ~n14778 ;
  assign y3237 = ~n14780 ;
  assign y3238 = n14791 ;
  assign y3239 = n14797 ;
  assign y3240 = n14800 ;
  assign y3241 = ~1'b0 ;
  assign y3242 = n14801 ;
  assign y3243 = ~n14802 ;
  assign y3244 = ~n14804 ;
  assign y3245 = ~n14806 ;
  assign y3246 = ~n14811 ;
  assign y3247 = n14812 ;
  assign y3248 = n14816 ;
  assign y3249 = n14818 ;
  assign y3250 = n14819 ;
  assign y3251 = ~n14826 ;
  assign y3252 = n14832 ;
  assign y3253 = ~1'b0 ;
  assign y3254 = n14833 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = n14840 ;
  assign y3257 = n14850 ;
  assign y3258 = n14853 ;
  assign y3259 = ~n14854 ;
  assign y3260 = n14855 ;
  assign y3261 = ~n14860 ;
  assign y3262 = n14867 ;
  assign y3263 = n14868 ;
  assign y3264 = ~1'b0 ;
  assign y3265 = ~n14869 ;
  assign y3266 = ~n14875 ;
  assign y3267 = ~n14876 ;
  assign y3268 = ~n14880 ;
  assign y3269 = n14882 ;
  assign y3270 = ~1'b0 ;
  assign y3271 = n14884 ;
  assign y3272 = ~n14885 ;
  assign y3273 = n14891 ;
  assign y3274 = n14895 ;
  assign y3275 = n14905 ;
  assign y3276 = ~n14910 ;
  assign y3277 = n14914 ;
  assign y3278 = ~1'b0 ;
  assign y3279 = ~n14919 ;
  assign y3280 = n14921 ;
  assign y3281 = n14922 ;
  assign y3282 = ~n14924 ;
  assign y3283 = n14939 ;
  assign y3284 = n14940 ;
  assign y3285 = ~n14947 ;
  assign y3286 = ~1'b0 ;
  assign y3287 = n14948 ;
  assign y3288 = ~n14951 ;
  assign y3289 = n14954 ;
  assign y3290 = n14961 ;
  assign y3291 = n14962 ;
  assign y3292 = ~n14963 ;
  assign y3293 = n14969 ;
  assign y3294 = ~n14971 ;
  assign y3295 = n14975 ;
  assign y3296 = n14978 ;
  assign y3297 = ~n14983 ;
  assign y3298 = ~n14985 ;
  assign y3299 = ~n14994 ;
  assign y3300 = ~n14997 ;
  assign y3301 = ~n15000 ;
  assign y3302 = n15001 ;
  assign y3303 = ~n15005 ;
  assign y3304 = ~n15011 ;
  assign y3305 = ~n10370 ;
  assign y3306 = ~n15018 ;
  assign y3307 = ~n15022 ;
  assign y3308 = ~n15029 ;
  assign y3309 = ~n15040 ;
  assign y3310 = ~1'b0 ;
  assign y3311 = ~1'b0 ;
  assign y3312 = n15046 ;
  assign y3313 = ~n15047 ;
  assign y3314 = n15052 ;
  assign y3315 = ~n15058 ;
  assign y3316 = ~n15060 ;
  assign y3317 = n15064 ;
  assign y3318 = ~1'b0 ;
  assign y3319 = ~n15066 ;
  assign y3320 = ~n15073 ;
  assign y3321 = n15076 ;
  assign y3322 = n15079 ;
  assign y3323 = n15081 ;
  assign y3324 = ~n15083 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~n15085 ;
  assign y3327 = ~n15087 ;
  assign y3328 = n15088 ;
  assign y3329 = n15091 ;
  assign y3330 = n15094 ;
  assign y3331 = ~1'b0 ;
  assign y3332 = n15100 ;
  assign y3333 = ~n15106 ;
  assign y3334 = ~n15127 ;
  assign y3335 = ~n15130 ;
  assign y3336 = ~1'b0 ;
  assign y3337 = ~n15137 ;
  assign y3338 = n15138 ;
  assign y3339 = ~n15139 ;
  assign y3340 = ~n15142 ;
  assign y3341 = ~n15152 ;
  assign y3342 = n15154 ;
  assign y3343 = ~n15160 ;
  assign y3344 = ~n15163 ;
  assign y3345 = ~1'b0 ;
  assign y3346 = n15168 ;
  assign y3347 = n15170 ;
  assign y3348 = ~n15172 ;
  assign y3349 = n15176 ;
  assign y3350 = n15179 ;
  assign y3351 = ~n15180 ;
  assign y3352 = ~n15183 ;
  assign y3353 = n15184 ;
  assign y3354 = ~n15188 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = n15194 ;
  assign y3357 = n15197 ;
  assign y3358 = ~n15201 ;
  assign y3359 = n15205 ;
  assign y3360 = n15206 ;
  assign y3361 = ~n15210 ;
  assign y3362 = ~n15215 ;
  assign y3363 = n15220 ;
  assign y3364 = ~n15234 ;
  assign y3365 = ~n15235 ;
  assign y3366 = n15242 ;
  assign y3367 = n15243 ;
  assign y3368 = ~n15246 ;
  assign y3369 = n15250 ;
  assign y3370 = n15253 ;
  assign y3371 = ~n15257 ;
  assign y3372 = n15259 ;
  assign y3373 = n15272 ;
  assign y3374 = ~n15277 ;
  assign y3375 = ~n15285 ;
  assign y3376 = n15289 ;
  assign y3377 = ~n15305 ;
  assign y3378 = ~n15306 ;
  assign y3379 = n15308 ;
  assign y3380 = ~n15314 ;
  assign y3381 = ~n15328 ;
  assign y3382 = n15330 ;
  assign y3383 = ~1'b0 ;
  assign y3384 = n15339 ;
  assign y3385 = ~n15341 ;
  assign y3386 = ~n15346 ;
  assign y3387 = n15350 ;
  assign y3388 = ~n15356 ;
  assign y3389 = ~1'b0 ;
  assign y3390 = ~n15367 ;
  assign y3391 = ~1'b0 ;
  assign y3392 = n15373 ;
  assign y3393 = ~n15382 ;
  assign y3394 = ~1'b0 ;
  assign y3395 = n15386 ;
  assign y3396 = ~n15391 ;
  assign y3397 = n15400 ;
  assign y3398 = n15401 ;
  assign y3399 = ~n15403 ;
  assign y3400 = n15409 ;
  assign y3401 = n15417 ;
  assign y3402 = n15423 ;
  assign y3403 = ~n15427 ;
  assign y3404 = ~n15432 ;
  assign y3405 = ~n15440 ;
  assign y3406 = ~n15443 ;
  assign y3407 = ~n15447 ;
  assign y3408 = n15451 ;
  assign y3409 = n15453 ;
  assign y3410 = ~n15454 ;
  assign y3411 = ~n15463 ;
  assign y3412 = n15468 ;
  assign y3413 = ~n15477 ;
  assign y3414 = ~n15479 ;
  assign y3415 = ~n15480 ;
  assign y3416 = n15482 ;
  assign y3417 = ~n15484 ;
  assign y3418 = n15487 ;
  assign y3419 = n15490 ;
  assign y3420 = ~n15492 ;
  assign y3421 = n15497 ;
  assign y3422 = ~n15501 ;
  assign y3423 = ~1'b0 ;
  assign y3424 = ~n15511 ;
  assign y3425 = ~n15512 ;
  assign y3426 = ~n15520 ;
  assign y3427 = n15521 ;
  assign y3428 = n15525 ;
  assign y3429 = n15528 ;
  assign y3430 = ~n15538 ;
  assign y3431 = ~n15539 ;
  assign y3432 = ~n15545 ;
  assign y3433 = n15554 ;
  assign y3434 = n15563 ;
  assign y3435 = ~n15565 ;
  assign y3436 = n716 ;
  assign y3437 = n15570 ;
  assign y3438 = ~1'b0 ;
  assign y3439 = ~n15572 ;
  assign y3440 = n15579 ;
  assign y3441 = 1'b0 ;
  assign y3442 = ~n15587 ;
  assign y3443 = n15590 ;
  assign y3444 = ~n15598 ;
  assign y3445 = ~n15603 ;
  assign y3446 = ~1'b0 ;
  assign y3447 = ~n15606 ;
  assign y3448 = n15609 ;
  assign y3449 = n15613 ;
  assign y3450 = ~n15620 ;
  assign y3451 = n15627 ;
  assign y3452 = ~n15631 ;
  assign y3453 = ~n15639 ;
  assign y3454 = ~n15645 ;
  assign y3455 = n15649 ;
  assign y3456 = n15653 ;
  assign y3457 = n15663 ;
  assign y3458 = n15665 ;
  assign y3459 = n15671 ;
  assign y3460 = ~n15673 ;
  assign y3461 = n15675 ;
  assign y3462 = n15676 ;
  assign y3463 = ~n15677 ;
  assign y3464 = ~n15679 ;
  assign y3465 = ~n15686 ;
  assign y3466 = ~n15692 ;
  assign y3467 = ~n15698 ;
  assign y3468 = n15705 ;
  assign y3469 = n15707 ;
  assign y3470 = n15714 ;
  assign y3471 = ~n15718 ;
  assign y3472 = ~n15722 ;
  assign y3473 = ~n15723 ;
  assign y3474 = n15740 ;
  assign y3475 = n15745 ;
  assign y3476 = ~n15757 ;
  assign y3477 = ~n15759 ;
  assign y3478 = ~n15763 ;
  assign y3479 = ~1'b0 ;
  assign y3480 = ~n15766 ;
  assign y3481 = n15775 ;
  assign y3482 = ~n15787 ;
  assign y3483 = ~n15793 ;
  assign y3484 = ~n15801 ;
  assign y3485 = n15802 ;
  assign y3486 = n15803 ;
  assign y3487 = ~n15805 ;
  assign y3488 = ~n15810 ;
  assign y3489 = n15815 ;
  assign y3490 = ~n15820 ;
  assign y3491 = ~n15826 ;
  assign y3492 = ~1'b0 ;
  assign y3493 = ~n15832 ;
  assign y3494 = n15839 ;
  assign y3495 = ~n15844 ;
  assign y3496 = ~n15848 ;
  assign y3497 = ~n15861 ;
  assign y3498 = ~n15863 ;
  assign y3499 = ~n15865 ;
  assign y3500 = ~1'b0 ;
  assign y3501 = ~n15871 ;
  assign y3502 = n15879 ;
  assign y3503 = ~n15885 ;
  assign y3504 = n15887 ;
  assign y3505 = ~n15888 ;
  assign y3506 = n15902 ;
  assign y3507 = ~n15906 ;
  assign y3508 = ~1'b0 ;
  assign y3509 = n15907 ;
  assign y3510 = n15909 ;
  assign y3511 = ~n15918 ;
  assign y3512 = n15924 ;
  assign y3513 = n15925 ;
  assign y3514 = ~n15927 ;
  assign y3515 = ~n15934 ;
  assign y3516 = n15939 ;
  assign y3517 = n15942 ;
  assign y3518 = ~n15946 ;
  assign y3519 = ~n15948 ;
  assign y3520 = ~n15951 ;
  assign y3521 = ~n15956 ;
  assign y3522 = ~n15958 ;
  assign y3523 = ~n15960 ;
  assign y3524 = n15961 ;
  assign y3525 = n15964 ;
  assign y3526 = n15969 ;
  assign y3527 = n15978 ;
  assign y3528 = n15982 ;
  assign y3529 = n15983 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = n15984 ;
  assign y3532 = n15989 ;
  assign y3533 = n16000 ;
  assign y3534 = ~n16008 ;
  assign y3535 = n16012 ;
  assign y3536 = n16015 ;
  assign y3537 = n16025 ;
  assign y3538 = ~n16026 ;
  assign y3539 = ~n16031 ;
  assign y3540 = ~n16040 ;
  assign y3541 = n16045 ;
  assign y3542 = ~n16052 ;
  assign y3543 = ~n16058 ;
  assign y3544 = n16060 ;
  assign y3545 = n16061 ;
  assign y3546 = ~1'b0 ;
  assign y3547 = n16072 ;
  assign y3548 = ~1'b0 ;
  assign y3549 = ~n16074 ;
  assign y3550 = n16075 ;
  assign y3551 = ~1'b0 ;
  assign y3552 = ~1'b0 ;
  assign y3553 = ~1'b0 ;
  assign y3554 = ~n16076 ;
  assign y3555 = ~n16085 ;
  assign y3556 = n16086 ;
  assign y3557 = n16088 ;
  assign y3558 = ~n16092 ;
  assign y3559 = ~1'b0 ;
  assign y3560 = n16096 ;
  assign y3561 = ~n16107 ;
  assign y3562 = ~n16108 ;
  assign y3563 = n16112 ;
  assign y3564 = ~n16116 ;
  assign y3565 = ~n16126 ;
  assign y3566 = ~n16131 ;
  assign y3567 = ~n16133 ;
  assign y3568 = ~n16140 ;
  assign y3569 = n16141 ;
  assign y3570 = ~n16142 ;
  assign y3571 = n16144 ;
  assign y3572 = ~n16165 ;
  assign y3573 = ~n16178 ;
  assign y3574 = n16183 ;
  assign y3575 = ~n16190 ;
  assign y3576 = ~n16191 ;
  assign y3577 = ~n16196 ;
  assign y3578 = ~n16202 ;
  assign y3579 = ~n16204 ;
  assign y3580 = ~n16214 ;
  assign y3581 = n16215 ;
  assign y3582 = ~n16217 ;
  assign y3583 = ~n16222 ;
  assign y3584 = ~n16223 ;
  assign y3585 = n16226 ;
  assign y3586 = ~n16229 ;
  assign y3587 = n16231 ;
  assign y3588 = n16232 ;
  assign y3589 = n16234 ;
  assign y3590 = n16235 ;
  assign y3591 = ~n16236 ;
  assign y3592 = n16239 ;
  assign y3593 = ~1'b0 ;
  assign y3594 = ~n16243 ;
  assign y3595 = n16245 ;
  assign y3596 = n16246 ;
  assign y3597 = n16247 ;
  assign y3598 = ~n16249 ;
  assign y3599 = n16259 ;
  assign y3600 = n16270 ;
  assign y3601 = n16277 ;
  assign y3602 = n16282 ;
  assign y3603 = ~n16286 ;
  assign y3604 = n16290 ;
  assign y3605 = ~1'b0 ;
  assign y3606 = ~n16291 ;
  assign y3607 = n16292 ;
  assign y3608 = n16298 ;
  assign y3609 = n16301 ;
  assign y3610 = ~n16302 ;
  assign y3611 = n16303 ;
  assign y3612 = ~n16304 ;
  assign y3613 = n16306 ;
  assign y3614 = n16307 ;
  assign y3615 = ~1'b0 ;
  assign y3616 = n16319 ;
  assign y3617 = ~1'b0 ;
  assign y3618 = ~n16323 ;
  assign y3619 = ~n16327 ;
  assign y3620 = ~n16329 ;
  assign y3621 = n16340 ;
  assign y3622 = n16342 ;
  assign y3623 = ~1'b0 ;
  assign y3624 = n16343 ;
  assign y3625 = ~n16347 ;
  assign y3626 = ~n16350 ;
  assign y3627 = ~n16353 ;
  assign y3628 = n16357 ;
  assign y3629 = n16366 ;
  assign y3630 = n16375 ;
  assign y3631 = ~1'b0 ;
  assign y3632 = ~n16384 ;
  assign y3633 = n16403 ;
  assign y3634 = n16406 ;
  assign y3635 = n16409 ;
  assign y3636 = ~n16410 ;
  assign y3637 = ~1'b0 ;
  assign y3638 = n16412 ;
  assign y3639 = n16423 ;
  assign y3640 = n16429 ;
  assign y3641 = ~1'b0 ;
  assign y3642 = n16430 ;
  assign y3643 = n16438 ;
  assign y3644 = n16440 ;
  assign y3645 = ~n16449 ;
  assign y3646 = ~n16450 ;
  assign y3647 = n16452 ;
  assign y3648 = n16460 ;
  assign y3649 = n16463 ;
  assign y3650 = ~n16466 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = ~n16468 ;
  assign y3653 = n16472 ;
  assign y3654 = ~1'b0 ;
  assign y3655 = n16477 ;
  assign y3656 = ~n16491 ;
  assign y3657 = ~n16502 ;
  assign y3658 = n16510 ;
  assign y3659 = n16512 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = ~1'b0 ;
  assign y3662 = ~n16525 ;
  assign y3663 = n16529 ;
  assign y3664 = ~n16541 ;
  assign y3665 = ~1'b0 ;
  assign y3666 = ~n16543 ;
  assign y3667 = ~1'b0 ;
  assign y3668 = ~n16555 ;
  assign y3669 = n16562 ;
  assign y3670 = n16563 ;
  assign y3671 = ~n16575 ;
  assign y3672 = ~n16580 ;
  assign y3673 = n16587 ;
  assign y3674 = n16589 ;
  assign y3675 = n16591 ;
  assign y3676 = n16592 ;
  assign y3677 = n16599 ;
  assign y3678 = ~n16605 ;
  assign y3679 = ~n16609 ;
  assign y3680 = n16614 ;
  assign y3681 = ~n16616 ;
  assign y3682 = n16617 ;
  assign y3683 = ~n16620 ;
  assign y3684 = n16626 ;
  assign y3685 = n16635 ;
  assign y3686 = n16637 ;
  assign y3687 = ~n16649 ;
  assign y3688 = ~n16653 ;
  assign y3689 = n16656 ;
  assign y3690 = ~n16657 ;
  assign y3691 = ~n16663 ;
  assign y3692 = n16664 ;
  assign y3693 = ~n16672 ;
  assign y3694 = n16673 ;
  assign y3695 = ~n16676 ;
  assign y3696 = ~n16677 ;
  assign y3697 = n16684 ;
  assign y3698 = ~n16686 ;
  assign y3699 = ~n16691 ;
  assign y3700 = ~n16699 ;
  assign y3701 = ~n16702 ;
  assign y3702 = ~n16705 ;
  assign y3703 = n16709 ;
  assign y3704 = ~n16715 ;
  assign y3705 = ~n16716 ;
  assign y3706 = n16721 ;
  assign y3707 = n16723 ;
  assign y3708 = n16727 ;
  assign y3709 = ~n16733 ;
  assign y3710 = n13740 ;
  assign y3711 = ~n16738 ;
  assign y3712 = ~n16747 ;
  assign y3713 = n16755 ;
  assign y3714 = ~n16763 ;
  assign y3715 = ~n16767 ;
  assign y3716 = n16781 ;
  assign y3717 = ~n16790 ;
  assign y3718 = ~n16797 ;
  assign y3719 = ~n16799 ;
  assign y3720 = ~n16805 ;
  assign y3721 = n16809 ;
  assign y3722 = n16813 ;
  assign y3723 = ~n16814 ;
  assign y3724 = n16820 ;
  assign y3725 = ~n16821 ;
  assign y3726 = n16822 ;
  assign y3727 = n16824 ;
  assign y3728 = ~n16828 ;
  assign y3729 = ~n16829 ;
  assign y3730 = n16836 ;
  assign y3731 = ~n16843 ;
  assign y3732 = n16848 ;
  assign y3733 = ~n16851 ;
  assign y3734 = n16857 ;
  assign y3735 = ~n16858 ;
  assign y3736 = ~n16865 ;
  assign y3737 = ~n16868 ;
  assign y3738 = n16869 ;
  assign y3739 = n16871 ;
  assign y3740 = n16873 ;
  assign y3741 = ~n16875 ;
  assign y3742 = n16878 ;
  assign y3743 = ~n16882 ;
  assign y3744 = ~n16885 ;
  assign y3745 = n16887 ;
  assign y3746 = ~n16897 ;
  assign y3747 = n16899 ;
  assign y3748 = n16901 ;
  assign y3749 = ~n16902 ;
  assign y3750 = n16906 ;
  assign y3751 = ~n16908 ;
  assign y3752 = n16912 ;
  assign y3753 = ~n16915 ;
  assign y3754 = ~n16922 ;
  assign y3755 = n16932 ;
  assign y3756 = ~n16935 ;
  assign y3757 = ~n16944 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = ~n16947 ;
  assign y3760 = ~n16948 ;
  assign y3761 = ~n16950 ;
  assign y3762 = ~1'b0 ;
  assign y3763 = ~n16952 ;
  assign y3764 = n16739 ;
  assign y3765 = ~1'b0 ;
  assign y3766 = n16957 ;
  assign y3767 = ~n16958 ;
  assign y3768 = ~n16961 ;
  assign y3769 = ~n16969 ;
  assign y3770 = ~1'b0 ;
  assign y3771 = n16974 ;
  assign y3772 = ~n16977 ;
  assign y3773 = ~n16980 ;
  assign y3774 = n16984 ;
  assign y3775 = n16986 ;
  assign y3776 = ~n16991 ;
  assign y3777 = ~1'b0 ;
  assign y3778 = ~n17004 ;
  assign y3779 = n17009 ;
  assign y3780 = ~n17016 ;
  assign y3781 = ~1'b0 ;
  assign y3782 = n17020 ;
  assign y3783 = ~n17021 ;
  assign y3784 = n17030 ;
  assign y3785 = ~1'b0 ;
  assign y3786 = ~n17036 ;
  assign y3787 = ~n17044 ;
  assign y3788 = ~n17053 ;
  assign y3789 = n17059 ;
  assign y3790 = n17063 ;
  assign y3791 = n17064 ;
  assign y3792 = n17069 ;
  assign y3793 = n17072 ;
  assign y3794 = n17086 ;
  assign y3795 = n17087 ;
  assign y3796 = n17089 ;
  assign y3797 = ~n17094 ;
  assign y3798 = n17095 ;
  assign y3799 = ~1'b0 ;
  assign y3800 = ~n17096 ;
  assign y3801 = ~1'b0 ;
  assign y3802 = ~n17105 ;
  assign y3803 = ~1'b0 ;
  assign y3804 = ~n17113 ;
  assign y3805 = ~n17118 ;
  assign y3806 = ~n17120 ;
  assign y3807 = n17129 ;
  assign y3808 = ~n17133 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~n17134 ;
  assign y3811 = n17145 ;
  assign y3812 = ~n17149 ;
  assign y3813 = n17150 ;
  assign y3814 = ~n17158 ;
  assign y3815 = n17159 ;
  assign y3816 = n17165 ;
  assign y3817 = ~n17168 ;
  assign y3818 = ~n17171 ;
  assign y3819 = ~n17178 ;
  assign y3820 = n17184 ;
  assign y3821 = ~n17195 ;
  assign y3822 = n17204 ;
  assign y3823 = ~n17207 ;
  assign y3824 = n17208 ;
  assign y3825 = ~n17211 ;
  assign y3826 = n17213 ;
  assign y3827 = n17216 ;
  assign y3828 = n17220 ;
  assign y3829 = ~n17221 ;
  assign y3830 = ~1'b0 ;
  assign y3831 = n17223 ;
  assign y3832 = n17231 ;
  assign y3833 = ~n17235 ;
  assign y3834 = ~n17236 ;
  assign y3835 = n17238 ;
  assign y3836 = ~n17242 ;
  assign y3837 = n17247 ;
  assign y3838 = n17252 ;
  assign y3839 = n17257 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~n17268 ;
  assign y3842 = ~n17269 ;
  assign y3843 = ~1'b0 ;
  assign y3844 = ~1'b0 ;
  assign y3845 = ~1'b0 ;
  assign y3846 = n17271 ;
  assign y3847 = n17272 ;
  assign y3848 = ~n17273 ;
  assign y3849 = n17275 ;
  assign y3850 = ~n17283 ;
  assign y3851 = ~n17284 ;
  assign y3852 = n17285 ;
  assign y3853 = n17296 ;
  assign y3854 = n17297 ;
  assign y3855 = ~n17303 ;
  assign y3856 = ~n17305 ;
  assign y3857 = n17307 ;
  assign y3858 = n17309 ;
  assign y3859 = ~n17310 ;
  assign y3860 = ~n17315 ;
  assign y3861 = n17317 ;
  assign y3862 = n17320 ;
  assign y3863 = ~n17326 ;
  assign y3864 = n17327 ;
  assign y3865 = n17337 ;
  assign y3866 = ~n17341 ;
  assign y3867 = ~n17348 ;
  assign y3868 = n17355 ;
  assign y3869 = ~n17361 ;
  assign y3870 = ~n17365 ;
  assign y3871 = ~n17367 ;
  assign y3872 = ~n17374 ;
  assign y3873 = n17375 ;
  assign y3874 = ~n17377 ;
  assign y3875 = ~n4945 ;
  assign y3876 = ~n17382 ;
  assign y3877 = n17384 ;
  assign y3878 = ~n17385 ;
  assign y3879 = n17392 ;
  assign y3880 = ~n17400 ;
  assign y3881 = ~n17402 ;
  assign y3882 = n17403 ;
  assign y3883 = n17409 ;
  assign y3884 = n17411 ;
  assign y3885 = n17412 ;
  assign y3886 = ~1'b0 ;
  assign y3887 = n17415 ;
  assign y3888 = ~n17417 ;
  assign y3889 = n17426 ;
  assign y3890 = ~n17428 ;
  assign y3891 = ~1'b0 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = ~n17432 ;
  assign y3894 = n17433 ;
  assign y3895 = ~n17434 ;
  assign y3896 = n17435 ;
  assign y3897 = ~n17439 ;
  assign y3898 = ~n17441 ;
  assign y3899 = ~n17445 ;
  assign y3900 = n17447 ;
  assign y3901 = ~n17453 ;
  assign y3902 = ~n17464 ;
  assign y3903 = ~n17468 ;
  assign y3904 = n17473 ;
  assign y3905 = ~n17481 ;
  assign y3906 = n17486 ;
  assign y3907 = n17487 ;
  assign y3908 = ~n17493 ;
  assign y3909 = n17501 ;
  assign y3910 = n17503 ;
  assign y3911 = ~n17506 ;
  assign y3912 = ~n17511 ;
  assign y3913 = n17515 ;
  assign y3914 = ~n17521 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = ~n17524 ;
  assign y3917 = ~n17527 ;
  assign y3918 = ~n17531 ;
  assign y3919 = n17535 ;
  assign y3920 = ~n17537 ;
  assign y3921 = ~1'b0 ;
  assign y3922 = ~n17538 ;
  assign y3923 = ~n17539 ;
  assign y3924 = n17544 ;
  assign y3925 = n17546 ;
  assign y3926 = ~1'b0 ;
  assign y3927 = ~1'b0 ;
  assign y3928 = n17548 ;
  assign y3929 = ~n17554 ;
  assign y3930 = n17571 ;
  assign y3931 = ~n17572 ;
  assign y3932 = ~n17575 ;
  assign y3933 = n17586 ;
  assign y3934 = n17589 ;
  assign y3935 = n17592 ;
  assign y3936 = n17597 ;
  assign y3937 = ~n17603 ;
  assign y3938 = n17616 ;
  assign y3939 = ~n17618 ;
  assign y3940 = ~n17619 ;
  assign y3941 = ~n17625 ;
  assign y3942 = ~n17629 ;
  assign y3943 = ~n17633 ;
  assign y3944 = ~n17634 ;
  assign y3945 = n17636 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = n17637 ;
  assign y3948 = ~n17639 ;
  assign y3949 = n17646 ;
  assign y3950 = ~n17650 ;
  assign y3951 = ~n17654 ;
  assign y3952 = n17658 ;
  assign y3953 = n17661 ;
  assign y3954 = n17663 ;
  assign y3955 = ~x163 ;
  assign y3956 = n17667 ;
  assign y3957 = n17671 ;
  assign y3958 = ~1'b0 ;
  assign y3959 = ~n17672 ;
  assign y3960 = ~n17673 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = ~n17676 ;
  assign y3963 = n17679 ;
  assign y3964 = n17685 ;
  assign y3965 = n17703 ;
  assign y3966 = ~n17705 ;
  assign y3967 = n17706 ;
  assign y3968 = n17708 ;
  assign y3969 = ~n17709 ;
  assign y3970 = ~1'b0 ;
  assign y3971 = ~n17712 ;
  assign y3972 = ~n17715 ;
  assign y3973 = ~n17717 ;
  assign y3974 = n17718 ;
  assign y3975 = ~n17719 ;
  assign y3976 = n17720 ;
  assign y3977 = ~n17721 ;
  assign y3978 = n17723 ;
  assign y3979 = ~n17746 ;
  assign y3980 = ~n17750 ;
  assign y3981 = n17755 ;
  assign y3982 = n17756 ;
  assign y3983 = n17762 ;
  assign y3984 = ~1'b0 ;
  assign y3985 = ~n17774 ;
  assign y3986 = n14507 ;
  assign y3987 = ~n17778 ;
  assign y3988 = n17779 ;
  assign y3989 = n17781 ;
  assign y3990 = ~n17782 ;
  assign y3991 = n17786 ;
  assign y3992 = n17787 ;
  assign y3993 = n17796 ;
  assign y3994 = n17804 ;
  assign y3995 = n17805 ;
  assign y3996 = ~n17806 ;
  assign y3997 = n17808 ;
  assign y3998 = ~n17811 ;
  assign y3999 = n17813 ;
  assign y4000 = ~1'b0 ;
  assign y4001 = ~n17818 ;
  assign y4002 = n17821 ;
  assign y4003 = ~n17823 ;
  assign y4004 = n17828 ;
  assign y4005 = ~n17833 ;
  assign y4006 = ~n17836 ;
  assign y4007 = ~1'b0 ;
  assign y4008 = ~n17842 ;
  assign y4009 = ~n17846 ;
  assign y4010 = ~n17848 ;
  assign y4011 = ~1'b0 ;
  assign y4012 = ~n17850 ;
  assign y4013 = ~n17854 ;
  assign y4014 = n17859 ;
  assign y4015 = ~n17860 ;
  assign y4016 = ~n17862 ;
  assign y4017 = ~n17865 ;
  assign y4018 = n17866 ;
  assign y4019 = ~n17874 ;
  assign y4020 = ~n17875 ;
  assign y4021 = ~1'b0 ;
  assign y4022 = n17879 ;
  assign y4023 = n17881 ;
  assign y4024 = ~n17885 ;
  assign y4025 = ~n17891 ;
  assign y4026 = n17895 ;
  assign y4027 = ~1'b0 ;
  assign y4028 = ~n17898 ;
  assign y4029 = n17904 ;
  assign y4030 = ~n17905 ;
  assign y4031 = n17911 ;
  assign y4032 = n5185 ;
  assign y4033 = n17920 ;
  assign y4034 = ~n17921 ;
  assign y4035 = n17924 ;
  assign y4036 = n17927 ;
  assign y4037 = ~n17937 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = ~n17939 ;
  assign y4040 = ~n17943 ;
  assign y4041 = ~n17949 ;
  assign y4042 = ~n17953 ;
  assign y4043 = ~1'b0 ;
  assign y4044 = ~n17959 ;
  assign y4045 = n17963 ;
  assign y4046 = ~n17971 ;
  assign y4047 = ~1'b0 ;
  assign y4048 = n6601 ;
  assign y4049 = n17980 ;
  assign y4050 = n17984 ;
  assign y4051 = ~n17987 ;
  assign y4052 = ~n17988 ;
  assign y4053 = n17989 ;
  assign y4054 = ~n17994 ;
  assign y4055 = ~1'b0 ;
  assign y4056 = ~n17995 ;
  assign y4057 = n17996 ;
  assign y4058 = ~n17997 ;
  assign y4059 = ~1'b0 ;
  assign y4060 = n18002 ;
  assign y4061 = ~n18003 ;
  assign y4062 = n18006 ;
  assign y4063 = ~n18008 ;
  assign y4064 = ~1'b0 ;
  assign y4065 = n18017 ;
  assign y4066 = ~n18018 ;
  assign y4067 = n18020 ;
  assign y4068 = n18024 ;
  assign y4069 = n18028 ;
  assign y4070 = ~n18034 ;
  assign y4071 = n18040 ;
  assign y4072 = n18043 ;
  assign y4073 = ~n18046 ;
  assign y4074 = n18047 ;
  assign y4075 = n18057 ;
  assign y4076 = n18059 ;
  assign y4077 = n18062 ;
  assign y4078 = ~n18066 ;
  assign y4079 = n18070 ;
  assign y4080 = n18071 ;
  assign y4081 = ~n18074 ;
  assign y4082 = n18081 ;
  assign y4083 = ~n18086 ;
  assign y4084 = ~n18089 ;
  assign y4085 = n18093 ;
  assign y4086 = n18095 ;
  assign y4087 = n18096 ;
  assign y4088 = n18097 ;
  assign y4089 = ~n18099 ;
  assign y4090 = ~n18105 ;
  assign y4091 = ~n18106 ;
  assign y4092 = n18109 ;
  assign y4093 = n18113 ;
  assign y4094 = n18122 ;
  assign y4095 = ~n18128 ;
  assign y4096 = ~n18134 ;
  assign y4097 = ~n18137 ;
  assign y4098 = n18140 ;
  assign y4099 = n18142 ;
  assign y4100 = n18144 ;
  assign y4101 = n18146 ;
  assign y4102 = ~n18147 ;
  assign y4103 = ~n18151 ;
  assign y4104 = n18153 ;
  assign y4105 = ~n18154 ;
  assign y4106 = ~1'b0 ;
  assign y4107 = n18175 ;
  assign y4108 = ~n18180 ;
  assign y4109 = n18185 ;
  assign y4110 = n18187 ;
  assign y4111 = n18201 ;
  assign y4112 = ~n18204 ;
  assign y4113 = n18213 ;
  assign y4114 = n18214 ;
  assign y4115 = ~n18218 ;
  assign y4116 = n18225 ;
  assign y4117 = n18226 ;
  assign y4118 = ~n18230 ;
  assign y4119 = ~n18234 ;
  assign y4120 = ~n18236 ;
  assign y4121 = n18248 ;
  assign y4122 = n18252 ;
  assign y4123 = ~1'b0 ;
  assign y4124 = ~n18254 ;
  assign y4125 = n18255 ;
  assign y4126 = n18261 ;
  assign y4127 = n18262 ;
  assign y4128 = n18263 ;
  assign y4129 = ~n18264 ;
  assign y4130 = ~n18267 ;
  assign y4131 = n18269 ;
  assign y4132 = n18272 ;
  assign y4133 = ~n18276 ;
  assign y4134 = n18278 ;
  assign y4135 = ~n18281 ;
  assign y4136 = ~n18287 ;
  assign y4137 = n18290 ;
  assign y4138 = ~n18294 ;
  assign y4139 = n18297 ;
  assign y4140 = n18301 ;
  assign y4141 = ~n18302 ;
  assign y4142 = n18304 ;
  assign y4143 = n18305 ;
  assign y4144 = ~1'b0 ;
  assign y4145 = ~n18310 ;
  assign y4146 = ~n18311 ;
  assign y4147 = ~n18314 ;
  assign y4148 = n18320 ;
  assign y4149 = ~1'b0 ;
  assign y4150 = n18326 ;
  assign y4151 = ~n18327 ;
  assign y4152 = ~1'b0 ;
  assign y4153 = ~n18328 ;
  assign y4154 = n18333 ;
  assign y4155 = n18334 ;
  assign y4156 = ~1'b0 ;
  assign y4157 = n18337 ;
  assign y4158 = ~n18342 ;
  assign y4159 = n18346 ;
  assign y4160 = n18349 ;
  assign y4161 = ~n18354 ;
  assign y4162 = ~1'b0 ;
  assign y4163 = n18359 ;
  assign y4164 = n18362 ;
  assign y4165 = ~n18366 ;
  assign y4166 = ~n18367 ;
  assign y4167 = n18368 ;
  assign y4168 = ~n18380 ;
  assign y4169 = ~n18387 ;
  assign y4170 = n18389 ;
  assign y4171 = 1'b0 ;
  assign y4172 = ~n18390 ;
  assign y4173 = ~n18393 ;
  assign y4174 = ~n1926 ;
  assign y4175 = ~n18396 ;
  assign y4176 = n18406 ;
  assign y4177 = n18407 ;
  assign y4178 = ~1'b0 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = ~n18410 ;
  assign y4181 = n18411 ;
  assign y4182 = n18413 ;
  assign y4183 = ~n18418 ;
  assign y4184 = ~n18420 ;
  assign y4185 = n18426 ;
  assign y4186 = ~n18434 ;
  assign y4187 = n18444 ;
  assign y4188 = ~n18445 ;
  assign y4189 = ~n18447 ;
  assign y4190 = n18450 ;
  assign y4191 = ~n18455 ;
  assign y4192 = ~n18460 ;
  assign y4193 = n18461 ;
  assign y4194 = n18463 ;
  assign y4195 = n18465 ;
  assign y4196 = ~1'b0 ;
  assign y4197 = ~1'b0 ;
  assign y4198 = n18467 ;
  assign y4199 = ~n18473 ;
  assign y4200 = ~n18474 ;
  assign y4201 = ~n18478 ;
  assign y4202 = ~n18485 ;
  assign y4203 = ~n18492 ;
  assign y4204 = ~n18494 ;
  assign y4205 = ~n18496 ;
  assign y4206 = ~1'b0 ;
  assign y4207 = n18498 ;
  assign y4208 = n18503 ;
  assign y4209 = ~n18504 ;
  assign y4210 = ~n18505 ;
  assign y4211 = ~n18508 ;
  assign y4212 = ~n18512 ;
  assign y4213 = 1'b0 ;
  assign y4214 = n18514 ;
  assign y4215 = ~n18516 ;
  assign y4216 = ~1'b0 ;
  assign y4217 = ~n18520 ;
  assign y4218 = n18523 ;
  assign y4219 = n18534 ;
  assign y4220 = n18536 ;
  assign y4221 = ~1'b0 ;
  assign y4222 = n18537 ;
  assign y4223 = ~n18542 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~n18546 ;
  assign y4226 = n18548 ;
  assign y4227 = n18553 ;
  assign y4228 = n18555 ;
  assign y4229 = n18557 ;
  assign y4230 = ~1'b0 ;
  assign y4231 = n18560 ;
  assign y4232 = ~n18563 ;
  assign y4233 = n18564 ;
  assign y4234 = n18567 ;
  assign y4235 = ~n18571 ;
  assign y4236 = n18584 ;
  assign y4237 = ~n18587 ;
  assign y4238 = ~n18590 ;
  assign y4239 = ~n18593 ;
  assign y4240 = n18597 ;
  assign y4241 = ~n18600 ;
  assign y4242 = ~n18606 ;
  assign y4243 = ~n18610 ;
  assign y4244 = ~n18611 ;
  assign y4245 = n18612 ;
  assign y4246 = ~n18622 ;
  assign y4247 = n18623 ;
  assign y4248 = ~n18627 ;
  assign y4249 = ~n18628 ;
  assign y4250 = ~n18632 ;
  assign y4251 = n18647 ;
  assign y4252 = ~n18669 ;
  assign y4253 = ~n18675 ;
  assign y4254 = n18677 ;
  assign y4255 = ~n18683 ;
  assign y4256 = ~n18686 ;
  assign y4257 = n18692 ;
  assign y4258 = n18693 ;
  assign y4259 = ~n18695 ;
  assign y4260 = ~n18696 ;
  assign y4261 = n18700 ;
  assign y4262 = ~n18702 ;
  assign y4263 = ~n18703 ;
  assign y4264 = ~n18705 ;
  assign y4265 = n18711 ;
  assign y4266 = n18713 ;
  assign y4267 = ~n18715 ;
  assign y4268 = ~n18716 ;
  assign y4269 = n18719 ;
  assign y4270 = ~n18721 ;
  assign y4271 = ~n18728 ;
  assign y4272 = ~n18731 ;
  assign y4273 = ~n18741 ;
  assign y4274 = n18742 ;
  assign y4275 = n18743 ;
  assign y4276 = n18744 ;
  assign y4277 = ~n18748 ;
  assign y4278 = ~n18756 ;
  assign y4279 = n18758 ;
  assign y4280 = ~1'b0 ;
  assign y4281 = ~n18771 ;
  assign y4282 = ~n18774 ;
  assign y4283 = ~n18776 ;
  assign y4284 = ~n18781 ;
  assign y4285 = n18787 ;
  assign y4286 = ~n18793 ;
  assign y4287 = ~n18795 ;
  assign y4288 = ~n18796 ;
  assign y4289 = n18799 ;
  assign y4290 = n18800 ;
  assign y4291 = ~n18803 ;
  assign y4292 = n18806 ;
  assign y4293 = ~n18808 ;
  assign y4294 = n18815 ;
  assign y4295 = n18816 ;
  assign y4296 = n18817 ;
  assign y4297 = ~n18818 ;
  assign y4298 = ~n18824 ;
  assign y4299 = ~n18827 ;
  assign y4300 = n18829 ;
  assign y4301 = n18833 ;
  assign y4302 = ~1'b0 ;
  assign y4303 = n18843 ;
  assign y4304 = n18845 ;
  assign y4305 = n18849 ;
  assign y4306 = n18852 ;
  assign y4307 = ~n18853 ;
  assign y4308 = n18855 ;
  assign y4309 = ~n11745 ;
  assign y4310 = n18862 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = ~n18864 ;
  assign y4313 = ~1'b0 ;
  assign y4314 = ~n18871 ;
  assign y4315 = ~1'b0 ;
  assign y4316 = n18876 ;
  assign y4317 = ~n18878 ;
  assign y4318 = ~n18879 ;
  assign y4319 = n18885 ;
  assign y4320 = n18887 ;
  assign y4321 = ~1'b0 ;
  assign y4322 = ~n18892 ;
  assign y4323 = ~1'b0 ;
  assign y4324 = n18893 ;
  assign y4325 = ~n18900 ;
  assign y4326 = ~n18903 ;
  assign y4327 = n18907 ;
  assign y4328 = ~n18913 ;
  assign y4329 = n18914 ;
  assign y4330 = n18915 ;
  assign y4331 = n18916 ;
  assign y4332 = ~n18918 ;
  assign y4333 = n18923 ;
  assign y4334 = n18925 ;
  assign y4335 = n18927 ;
  assign y4336 = n18928 ;
  assign y4337 = n18933 ;
  assign y4338 = ~n18943 ;
  assign y4339 = ~n18945 ;
  assign y4340 = ~n18964 ;
  assign y4341 = n18970 ;
  assign y4342 = ~1'b0 ;
  assign y4343 = n18979 ;
  assign y4344 = ~n18980 ;
  assign y4345 = ~n18984 ;
  assign y4346 = n18988 ;
  assign y4347 = ~n18999 ;
  assign y4348 = n19000 ;
  assign y4349 = ~n19001 ;
  assign y4350 = n19003 ;
  assign y4351 = n19006 ;
  assign y4352 = n19007 ;
  assign y4353 = ~n19009 ;
  assign y4354 = ~n19012 ;
  assign y4355 = n19018 ;
  assign y4356 = n19021 ;
  assign y4357 = ~n19022 ;
  assign y4358 = ~n19025 ;
  assign y4359 = n19026 ;
  assign y4360 = n19035 ;
  assign y4361 = ~n19039 ;
  assign y4362 = n2864 ;
  assign y4363 = n19051 ;
  assign y4364 = ~n19057 ;
  assign y4365 = ~1'b0 ;
  assign y4366 = ~n19058 ;
  assign y4367 = ~n19059 ;
  assign y4368 = ~n19060 ;
  assign y4369 = n19062 ;
  assign y4370 = n19069 ;
  assign y4371 = n19075 ;
  assign y4372 = n19079 ;
  assign y4373 = ~n19083 ;
  assign y4374 = ~n19084 ;
  assign y4375 = n19085 ;
  assign y4376 = n19087 ;
  assign y4377 = ~n19090 ;
  assign y4378 = ~n19096 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = ~1'b0 ;
  assign y4381 = n19105 ;
  assign y4382 = ~n19111 ;
  assign y4383 = n19112 ;
  assign y4384 = n19124 ;
  assign y4385 = n13484 ;
  assign y4386 = ~n19126 ;
  assign y4387 = ~n19129 ;
  assign y4388 = ~n19132 ;
  assign y4389 = ~n19133 ;
  assign y4390 = ~n19135 ;
  assign y4391 = ~n19137 ;
  assign y4392 = n19151 ;
  assign y4393 = ~n19153 ;
  assign y4394 = n19154 ;
  assign y4395 = n19164 ;
  assign y4396 = n19166 ;
  assign y4397 = ~n19177 ;
  assign y4398 = n19178 ;
  assign y4399 = ~n19181 ;
  assign y4400 = ~n19183 ;
  assign y4401 = ~n19184 ;
  assign y4402 = ~n19185 ;
  assign y4403 = ~n19189 ;
  assign y4404 = n19196 ;
  assign y4405 = n19198 ;
  assign y4406 = n19199 ;
  assign y4407 = ~n19209 ;
  assign y4408 = n19214 ;
  assign y4409 = n19223 ;
  assign y4410 = n19225 ;
  assign y4411 = n19229 ;
  assign y4412 = n19230 ;
  assign y4413 = ~n19236 ;
  assign y4414 = ~n19240 ;
  assign y4415 = n19243 ;
  assign y4416 = ~n19247 ;
  assign y4417 = ~n19251 ;
  assign y4418 = n19253 ;
  assign y4419 = n19261 ;
  assign y4420 = ~n19264 ;
  assign y4421 = n19270 ;
  assign y4422 = n19272 ;
  assign y4423 = ~n19276 ;
  assign y4424 = n19277 ;
  assign y4425 = n19286 ;
  assign y4426 = n19287 ;
  assign y4427 = ~n19295 ;
  assign y4428 = ~n19301 ;
  assign y4429 = n19305 ;
  assign y4430 = n19307 ;
  assign y4431 = ~n19308 ;
  assign y4432 = ~n19311 ;
  assign y4433 = n19313 ;
  assign y4434 = ~n19318 ;
  assign y4435 = n19321 ;
  assign y4436 = n19323 ;
  assign y4437 = n19325 ;
  assign y4438 = ~n19331 ;
  assign y4439 = ~n19333 ;
  assign y4440 = n19339 ;
  assign y4441 = n19344 ;
  assign y4442 = n19348 ;
  assign y4443 = ~n19360 ;
  assign y4444 = ~n19361 ;
  assign y4445 = ~n19362 ;
  assign y4446 = ~n19366 ;
  assign y4447 = n19371 ;
  assign y4448 = ~n19375 ;
  assign y4449 = ~n19376 ;
  assign y4450 = ~n19379 ;
  assign y4451 = n19380 ;
  assign y4452 = n19386 ;
  assign y4453 = ~1'b0 ;
  assign y4454 = ~n19392 ;
  assign y4455 = ~n19397 ;
  assign y4456 = n19407 ;
  assign y4457 = ~n19414 ;
  assign y4458 = n19416 ;
  assign y4459 = ~n19418 ;
  assign y4460 = ~n16632 ;
  assign y4461 = n19423 ;
  assign y4462 = ~n19427 ;
  assign y4463 = n19428 ;
  assign y4464 = ~1'b0 ;
  assign y4465 = n19439 ;
  assign y4466 = n19440 ;
  assign y4467 = ~1'b0 ;
  assign y4468 = ~1'b0 ;
  assign y4469 = n19444 ;
  assign y4470 = ~n19449 ;
  assign y4471 = ~n19453 ;
  assign y4472 = n19458 ;
  assign y4473 = n19462 ;
  assign y4474 = ~n19466 ;
  assign y4475 = n19470 ;
  assign y4476 = n19481 ;
  assign y4477 = ~n19485 ;
  assign y4478 = n19488 ;
  assign y4479 = ~n19490 ;
  assign y4480 = ~n19492 ;
  assign y4481 = ~n19499 ;
  assign y4482 = ~n19502 ;
  assign y4483 = n19507 ;
  assign y4484 = ~n19510 ;
  assign y4485 = ~n19514 ;
  assign y4486 = ~n19522 ;
  assign y4487 = ~n19523 ;
  assign y4488 = n19533 ;
  assign y4489 = ~n19541 ;
  assign y4490 = n19545 ;
  assign y4491 = ~n19551 ;
  assign y4492 = n19554 ;
  assign y4493 = ~n19562 ;
  assign y4494 = ~n19565 ;
  assign y4495 = n19566 ;
  assign y4496 = ~n19571 ;
  assign y4497 = ~n19577 ;
  assign y4498 = n19578 ;
  assign y4499 = ~n19583 ;
  assign y4500 = n19585 ;
  assign y4501 = ~n19592 ;
  assign y4502 = n19593 ;
  assign y4503 = ~n19595 ;
  assign y4504 = ~n19597 ;
  assign y4505 = n19598 ;
  assign y4506 = n19602 ;
  assign y4507 = ~n19612 ;
  assign y4508 = ~n19615 ;
  assign y4509 = ~n19622 ;
  assign y4510 = n19623 ;
  assign y4511 = ~n19627 ;
  assign y4512 = n19628 ;
  assign y4513 = ~n19637 ;
  assign y4514 = n19641 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~n19644 ;
  assign y4517 = ~1'b0 ;
  assign y4518 = n19650 ;
  assign y4519 = n19652 ;
  assign y4520 = n19655 ;
  assign y4521 = n19659 ;
  assign y4522 = ~n19661 ;
  assign y4523 = n19663 ;
  assign y4524 = ~n19665 ;
  assign y4525 = n19678 ;
  assign y4526 = n19681 ;
  assign y4527 = ~n19686 ;
  assign y4528 = ~n19689 ;
  assign y4529 = ~1'b0 ;
  assign y4530 = n19690 ;
  assign y4531 = ~n19691 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = n19692 ;
  assign y4534 = n19696 ;
  assign y4535 = ~n19707 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = n19708 ;
  assign y4538 = n19714 ;
  assign y4539 = ~n19720 ;
  assign y4540 = ~n19722 ;
  assign y4541 = ~n19726 ;
  assign y4542 = ~n19727 ;
  assign y4543 = ~1'b0 ;
  assign y4544 = ~n19735 ;
  assign y4545 = ~n19744 ;
  assign y4546 = ~n19747 ;
  assign y4547 = ~n19749 ;
  assign y4548 = n19753 ;
  assign y4549 = ~n19769 ;
  assign y4550 = n19775 ;
  assign y4551 = ~n19783 ;
  assign y4552 = ~n19784 ;
  assign y4553 = ~1'b0 ;
  assign y4554 = ~1'b0 ;
  assign y4555 = n19786 ;
  assign y4556 = ~n19787 ;
  assign y4557 = ~n19789 ;
  assign y4558 = n19797 ;
  assign y4559 = n19799 ;
  assign y4560 = n19801 ;
  assign y4561 = n19812 ;
  assign y4562 = ~1'b0 ;
  assign y4563 = ~n19824 ;
  assign y4564 = ~n19830 ;
  assign y4565 = n19837 ;
  assign y4566 = ~1'b0 ;
  assign y4567 = ~1'b0 ;
  assign y4568 = ~n19839 ;
  assign y4569 = ~n19841 ;
  assign y4570 = ~n19847 ;
  assign y4571 = ~n19849 ;
  assign y4572 = ~n19851 ;
  assign y4573 = ~n19860 ;
  assign y4574 = n19864 ;
  assign y4575 = ~n19865 ;
  assign y4576 = n19866 ;
  assign y4577 = n19867 ;
  assign y4578 = ~n19872 ;
  assign y4579 = ~1'b0 ;
  assign y4580 = ~n19874 ;
  assign y4581 = ~n19876 ;
  assign y4582 = n19880 ;
  assign y4583 = ~n19887 ;
  assign y4584 = ~1'b0 ;
  assign y4585 = ~n19895 ;
  assign y4586 = n19898 ;
  assign y4587 = ~n19900 ;
  assign y4588 = n19905 ;
  assign y4589 = n19909 ;
  assign y4590 = ~n19910 ;
  assign y4591 = ~n19912 ;
  assign y4592 = ~n19913 ;
  assign y4593 = ~1'b0 ;
  assign y4594 = ~n19923 ;
  assign y4595 = ~n19924 ;
  assign y4596 = ~n19926 ;
  assign y4597 = ~n19928 ;
  assign y4598 = ~n19931 ;
  assign y4599 = ~n19940 ;
  assign y4600 = n19965 ;
  assign y4601 = ~n19973 ;
  assign y4602 = ~n19974 ;
  assign y4603 = n19976 ;
  assign y4604 = ~n19982 ;
  assign y4605 = ~n19989 ;
  assign y4606 = n19991 ;
  assign y4607 = ~n19994 ;
  assign y4608 = ~n19996 ;
  assign y4609 = ~1'b0 ;
  assign y4610 = n20001 ;
  assign y4611 = ~n20005 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = ~n20008 ;
  assign y4614 = ~n20018 ;
  assign y4615 = n20020 ;
  assign y4616 = ~n20021 ;
  assign y4617 = n20024 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = n20027 ;
  assign y4620 = n20034 ;
  assign y4621 = ~1'b0 ;
  assign y4622 = n20037 ;
  assign y4623 = ~n20039 ;
  assign y4624 = n20061 ;
  assign y4625 = ~n20065 ;
  assign y4626 = n20070 ;
  assign y4627 = n20072 ;
  assign y4628 = ~n20073 ;
  assign y4629 = ~n20085 ;
  assign y4630 = ~n20088 ;
  assign y4631 = ~n771 ;
  assign y4632 = ~n20089 ;
  assign y4633 = ~n20093 ;
  assign y4634 = ~n20098 ;
  assign y4635 = ~n20100 ;
  assign y4636 = n20107 ;
  assign y4637 = n20117 ;
  assign y4638 = ~n20118 ;
  assign y4639 = n20121 ;
  assign y4640 = ~n20125 ;
  assign y4641 = n20129 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = n20133 ;
  assign y4644 = ~n20135 ;
  assign y4645 = ~n20136 ;
  assign y4646 = ~n20137 ;
  assign y4647 = n20141 ;
  assign y4648 = ~n20142 ;
  assign y4649 = ~n20143 ;
  assign y4650 = ~n20146 ;
  assign y4651 = ~n20151 ;
  assign y4652 = ~1'b0 ;
  assign y4653 = n20155 ;
  assign y4654 = ~n20161 ;
  assign y4655 = ~n20166 ;
  assign y4656 = ~n20168 ;
  assign y4657 = ~n20176 ;
  assign y4658 = ~1'b0 ;
  assign y4659 = n20179 ;
  assign y4660 = ~n20182 ;
  assign y4661 = n20185 ;
  assign y4662 = n20194 ;
  assign y4663 = ~1'b0 ;
  assign y4664 = ~n20196 ;
  assign y4665 = n20197 ;
  assign y4666 = n20203 ;
  assign y4667 = ~n20204 ;
  assign y4668 = ~n20213 ;
  assign y4669 = ~n20217 ;
  assign y4670 = n20219 ;
  assign y4671 = n20224 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = ~n20225 ;
  assign y4674 = n20230 ;
  assign y4675 = n20235 ;
  assign y4676 = ~n20240 ;
  assign y4677 = n20241 ;
  assign y4678 = n20247 ;
  assign y4679 = n20250 ;
  assign y4680 = ~n20252 ;
  assign y4681 = n20263 ;
  assign y4682 = ~n20264 ;
  assign y4683 = n20275 ;
  assign y4684 = ~n20278 ;
  assign y4685 = n20280 ;
  assign y4686 = ~1'b0 ;
  assign y4687 = n20282 ;
  assign y4688 = ~n20287 ;
  assign y4689 = ~n20297 ;
  assign y4690 = n20299 ;
  assign y4691 = ~n20301 ;
  assign y4692 = ~n20302 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = n20303 ;
  assign y4695 = ~n20311 ;
  assign y4696 = n20313 ;
  assign y4697 = n20315 ;
  assign y4698 = ~1'b0 ;
  assign y4699 = n20316 ;
  assign y4700 = n20326 ;
  assign y4701 = ~n20335 ;
  assign y4702 = ~n20344 ;
  assign y4703 = ~n20346 ;
  assign y4704 = ~n20350 ;
  assign y4705 = n20363 ;
  assign y4706 = n6280 ;
  assign y4707 = ~n20366 ;
  assign y4708 = ~n20372 ;
  assign y4709 = n20381 ;
  assign y4710 = n20382 ;
  assign y4711 = n20387 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = n20388 ;
  assign y4714 = n20394 ;
  assign y4715 = n20401 ;
  assign y4716 = ~n20402 ;
  assign y4717 = ~n20420 ;
  assign y4718 = ~n20424 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = n20429 ;
  assign y4721 = ~1'b0 ;
  assign y4722 = ~n20430 ;
  assign y4723 = n20431 ;
  assign y4724 = ~n20453 ;
  assign y4725 = ~n20455 ;
  assign y4726 = ~n20457 ;
  assign y4727 = ~n20460 ;
  assign y4728 = ~1'b0 ;
  assign y4729 = ~n20464 ;
  assign y4730 = ~n20465 ;
  assign y4731 = ~n20468 ;
  assign y4732 = n20473 ;
  assign y4733 = ~n20474 ;
  assign y4734 = n20478 ;
  assign y4735 = n20481 ;
  assign y4736 = n20483 ;
  assign y4737 = n20492 ;
  assign y4738 = n20494 ;
  assign y4739 = ~n20500 ;
  assign y4740 = ~1'b0 ;
  assign y4741 = ~n20501 ;
  assign y4742 = n17332 ;
  assign y4743 = n20505 ;
  assign y4744 = n20507 ;
  assign y4745 = n20509 ;
  assign y4746 = n20520 ;
  assign y4747 = ~n20522 ;
  assign y4748 = n20529 ;
  assign y4749 = n20530 ;
  assign y4750 = n20538 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = n20544 ;
  assign y4753 = ~n20547 ;
  assign y4754 = ~n20548 ;
  assign y4755 = n20549 ;
  assign y4756 = n20551 ;
  assign y4757 = n20563 ;
  assign y4758 = ~n20574 ;
  assign y4759 = ~1'b0 ;
  assign y4760 = ~n20579 ;
  assign y4761 = ~n20583 ;
  assign y4762 = ~n20592 ;
  assign y4763 = ~n20602 ;
  assign y4764 = n20604 ;
  assign y4765 = ~n20605 ;
  assign y4766 = ~n20608 ;
  assign y4767 = n20609 ;
  assign y4768 = ~n20615 ;
  assign y4769 = n20617 ;
  assign y4770 = n20618 ;
  assign y4771 = n20621 ;
  assign y4772 = ~n20622 ;
  assign y4773 = ~n20625 ;
  assign y4774 = n20628 ;
  assign y4775 = ~n20632 ;
  assign y4776 = ~n20634 ;
  assign y4777 = n20639 ;
  assign y4778 = ~1'b0 ;
  assign y4779 = ~n20640 ;
  assign y4780 = n20643 ;
  assign y4781 = ~n20654 ;
  assign y4782 = ~1'b0 ;
  assign y4783 = ~n20659 ;
  assign y4784 = ~n20662 ;
  assign y4785 = n20665 ;
  assign y4786 = n20667 ;
  assign y4787 = ~n20670 ;
  assign y4788 = n20672 ;
  assign y4789 = ~n20681 ;
  assign y4790 = ~n20683 ;
  assign y4791 = n20684 ;
  assign y4792 = n20689 ;
  assign y4793 = ~n20691 ;
  assign y4794 = ~n20694 ;
  assign y4795 = n20699 ;
  assign y4796 = n20701 ;
  assign y4797 = ~n20705 ;
  assign y4798 = ~n20713 ;
  assign y4799 = n20714 ;
  assign y4800 = ~n20716 ;
  assign y4801 = ~n20720 ;
  assign y4802 = ~n20722 ;
  assign y4803 = n20723 ;
  assign y4804 = n20733 ;
  assign y4805 = n20734 ;
  assign y4806 = n20738 ;
  assign y4807 = n20743 ;
  assign y4808 = n20745 ;
  assign y4809 = ~n20749 ;
  assign y4810 = ~1'b0 ;
  assign y4811 = n20753 ;
  assign y4812 = ~n20760 ;
  assign y4813 = n20764 ;
  assign y4814 = ~n20768 ;
  assign y4815 = n20769 ;
  assign y4816 = n20771 ;
  assign y4817 = n20773 ;
  assign y4818 = ~n20775 ;
  assign y4819 = ~n20786 ;
  assign y4820 = ~n20791 ;
  assign y4821 = n20797 ;
  assign y4822 = n20799 ;
  assign y4823 = ~n20803 ;
  assign y4824 = ~n20805 ;
  assign y4825 = n20810 ;
  assign y4826 = n20812 ;
  assign y4827 = n20814 ;
  assign y4828 = n20816 ;
  assign y4829 = n20818 ;
  assign y4830 = n20825 ;
  assign y4831 = ~n20831 ;
  assign y4832 = ~1'b0 ;
  assign y4833 = n20836 ;
  assign y4834 = n20837 ;
  assign y4835 = n20843 ;
  assign y4836 = n20850 ;
  assign y4837 = n20854 ;
  assign y4838 = n20859 ;
  assign y4839 = n20862 ;
  assign y4840 = ~n20863 ;
  assign y4841 = n20867 ;
  assign y4842 = ~1'b0 ;
  assign y4843 = ~n20871 ;
  assign y4844 = ~n20879 ;
  assign y4845 = n20882 ;
  assign y4846 = ~n20883 ;
  assign y4847 = ~n20886 ;
  assign y4848 = ~n20888 ;
  assign y4849 = n20892 ;
  assign y4850 = n20897 ;
  assign y4851 = ~n20898 ;
  assign y4852 = ~1'b0 ;
  assign y4853 = n20900 ;
  assign y4854 = n20901 ;
  assign y4855 = n20906 ;
  assign y4856 = n20909 ;
  assign y4857 = n20914 ;
  assign y4858 = ~1'b0 ;
  assign y4859 = n20919 ;
  assign y4860 = ~n20920 ;
  assign y4861 = n20923 ;
  assign y4862 = n20926 ;
  assign y4863 = n20930 ;
  assign y4864 = ~n20936 ;
  assign y4865 = ~1'b0 ;
  assign y4866 = n20937 ;
  assign y4867 = ~n20938 ;
  assign y4868 = n20948 ;
  assign y4869 = n20951 ;
  assign y4870 = n20963 ;
  assign y4871 = n20967 ;
  assign y4872 = ~n20971 ;
  assign y4873 = n20975 ;
  assign y4874 = ~n20976 ;
  assign y4875 = n20977 ;
  assign y4876 = ~n20980 ;
  assign y4877 = ~n20982 ;
  assign y4878 = ~n20988 ;
  assign y4879 = ~n20993 ;
  assign y4880 = n21000 ;
  assign y4881 = ~n21007 ;
  assign y4882 = ~n21009 ;
  assign y4883 = ~n21012 ;
  assign y4884 = ~n21013 ;
  assign y4885 = n21014 ;
  assign y4886 = ~n21016 ;
  assign y4887 = ~n21017 ;
  assign y4888 = ~n21019 ;
  assign y4889 = ~n21021 ;
  assign y4890 = n21027 ;
  assign y4891 = n21028 ;
  assign y4892 = n21035 ;
  assign y4893 = n21037 ;
  assign y4894 = n21044 ;
  assign y4895 = ~n21047 ;
  assign y4896 = n21049 ;
  assign y4897 = n21051 ;
  assign y4898 = n21062 ;
  assign y4899 = ~n21064 ;
  assign y4900 = ~n21067 ;
  assign y4901 = n21072 ;
  assign y4902 = ~n21078 ;
  assign y4903 = n21081 ;
  assign y4904 = ~n21082 ;
  assign y4905 = ~n21089 ;
  assign y4906 = ~n21092 ;
  assign y4907 = n21094 ;
  assign y4908 = ~n21097 ;
  assign y4909 = ~n21098 ;
  assign y4910 = n21100 ;
  assign y4911 = ~n21103 ;
  assign y4912 = ~1'b0 ;
  assign y4913 = ~n21122 ;
  assign y4914 = n21124 ;
  assign y4915 = ~n21125 ;
  assign y4916 = ~1'b0 ;
  assign y4917 = n21127 ;
  assign y4918 = n21131 ;
  assign y4919 = ~n21132 ;
  assign y4920 = ~n21136 ;
  assign y4921 = ~n21147 ;
  assign y4922 = ~n21152 ;
  assign y4923 = n21153 ;
  assign y4924 = n21155 ;
  assign y4925 = n21176 ;
  assign y4926 = ~n21179 ;
  assign y4927 = n21180 ;
  assign y4928 = ~n21182 ;
  assign y4929 = ~1'b0 ;
  assign y4930 = ~1'b0 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = n21192 ;
  assign y4933 = n21193 ;
  assign y4934 = n21197 ;
  assign y4935 = n21202 ;
  assign y4936 = n21207 ;
  assign y4937 = n21213 ;
  assign y4938 = ~n21215 ;
  assign y4939 = n21221 ;
  assign y4940 = n21224 ;
  assign y4941 = n21234 ;
  assign y4942 = ~n21241 ;
  assign y4943 = ~n21244 ;
  assign y4944 = ~n21258 ;
  assign y4945 = ~n21266 ;
  assign y4946 = ~n21267 ;
  assign y4947 = ~n21270 ;
  assign y4948 = ~n21276 ;
  assign y4949 = ~n21279 ;
  assign y4950 = ~n21280 ;
  assign y4951 = ~n21285 ;
  assign y4952 = n21287 ;
  assign y4953 = ~1'b0 ;
  assign y4954 = n21293 ;
  assign y4955 = n21294 ;
  assign y4956 = ~n21295 ;
  assign y4957 = ~n21297 ;
  assign y4958 = ~n21302 ;
  assign y4959 = n21305 ;
  assign y4960 = n21311 ;
  assign y4961 = ~n21314 ;
  assign y4962 = ~n21317 ;
  assign y4963 = n6769 ;
  assign y4964 = ~1'b0 ;
  assign y4965 = n21326 ;
  assign y4966 = ~n21330 ;
  assign y4967 = n21331 ;
  assign y4968 = n21335 ;
  assign y4969 = ~n21340 ;
  assign y4970 = ~n21343 ;
  assign y4971 = n21347 ;
  assign y4972 = ~n21349 ;
  assign y4973 = ~n21352 ;
  assign y4974 = ~n21358 ;
  assign y4975 = n21362 ;
  assign y4976 = ~n21364 ;
  assign y4977 = n21370 ;
  assign y4978 = ~n21374 ;
  assign y4979 = ~n21375 ;
  assign y4980 = ~n21378 ;
  assign y4981 = n21379 ;
  assign y4982 = n21384 ;
  assign y4983 = n21387 ;
  assign y4984 = n21390 ;
  assign y4985 = ~n21391 ;
  assign y4986 = n21392 ;
  assign y4987 = n21396 ;
  assign y4988 = ~n21399 ;
  assign y4989 = n21400 ;
  assign y4990 = n21404 ;
  assign y4991 = ~n21408 ;
  assign y4992 = ~n21409 ;
  assign y4993 = ~n21412 ;
  assign y4994 = ~n21413 ;
  assign y4995 = ~n21415 ;
  assign y4996 = n21417 ;
  assign y4997 = n21422 ;
  assign y4998 = ~n21427 ;
  assign y4999 = n21428 ;
  assign y5000 = n21431 ;
  assign y5001 = ~1'b0 ;
  assign y5002 = ~n21433 ;
  assign y5003 = ~n21436 ;
  assign y5004 = ~n21437 ;
  assign y5005 = ~1'b0 ;
  assign y5006 = n21441 ;
  assign y5007 = n21445 ;
  assign y5008 = ~n21446 ;
  assign y5009 = n21454 ;
  assign y5010 = n21459 ;
  assign y5011 = ~n21463 ;
  assign y5012 = ~1'b0 ;
  assign y5013 = ~1'b0 ;
  assign y5014 = n21464 ;
  assign y5015 = n21465 ;
  assign y5016 = n21468 ;
  assign y5017 = n21470 ;
  assign y5018 = n21472 ;
  assign y5019 = n21476 ;
  assign y5020 = ~1'b0 ;
  assign y5021 = ~n21481 ;
  assign y5022 = n21493 ;
  assign y5023 = ~n21496 ;
  assign y5024 = ~n21499 ;
  assign y5025 = ~n21501 ;
  assign y5026 = n21504 ;
  assign y5027 = ~n21507 ;
  assign y5028 = ~n21509 ;
  assign y5029 = ~1'b0 ;
  assign y5030 = ~n21513 ;
  assign y5031 = n21514 ;
  assign y5032 = n21515 ;
  assign y5033 = ~n21517 ;
  assign y5034 = ~n21519 ;
  assign y5035 = n21520 ;
  assign y5036 = n21521 ;
  assign y5037 = n21522 ;
  assign y5038 = ~n21527 ;
  assign y5039 = n21528 ;
  assign y5040 = n21531 ;
  assign y5041 = ~n21542 ;
  assign y5042 = ~1'b0 ;
  assign y5043 = ~n21544 ;
  assign y5044 = ~n21547 ;
  assign y5045 = ~n21548 ;
  assign y5046 = ~1'b0 ;
  assign y5047 = ~1'b0 ;
  assign y5048 = n21551 ;
  assign y5049 = ~n21554 ;
  assign y5050 = n21556 ;
  assign y5051 = n21561 ;
  assign y5052 = n21564 ;
  assign y5053 = ~n21567 ;
  assign y5054 = ~n21572 ;
  assign y5055 = n21574 ;
  assign y5056 = ~1'b0 ;
  assign y5057 = ~n21578 ;
  assign y5058 = ~n21580 ;
  assign y5059 = n21586 ;
  assign y5060 = n21591 ;
  assign y5061 = ~n21593 ;
  assign y5062 = ~n21602 ;
  assign y5063 = ~n4680 ;
  assign y5064 = ~n21605 ;
  assign y5065 = ~n21611 ;
  assign y5066 = n21612 ;
  assign y5067 = ~n21614 ;
  assign y5068 = n21616 ;
  assign y5069 = ~n21625 ;
  assign y5070 = ~n21631 ;
  assign y5071 = n21633 ;
  assign y5072 = ~1'b0 ;
  assign y5073 = n21635 ;
  assign y5074 = ~n21637 ;
  assign y5075 = ~n21641 ;
  assign y5076 = n21645 ;
  assign y5077 = ~1'b0 ;
  assign y5078 = ~n21647 ;
  assign y5079 = n21649 ;
  assign y5080 = n21654 ;
  assign y5081 = ~n21655 ;
  assign y5082 = ~n21660 ;
  assign y5083 = n21663 ;
  assign y5084 = n21669 ;
  assign y5085 = n21670 ;
  assign y5086 = ~n21673 ;
  assign y5087 = ~n21676 ;
  assign y5088 = ~1'b0 ;
  assign y5089 = ~n21682 ;
  assign y5090 = ~n21683 ;
  assign y5091 = ~n21686 ;
  assign y5092 = ~n21689 ;
  assign y5093 = n21690 ;
  assign y5094 = n21692 ;
  assign y5095 = ~n21696 ;
  assign y5096 = 1'b0 ;
  assign y5097 = ~1'b0 ;
  assign y5098 = ~n21701 ;
  assign y5099 = n21704 ;
  assign y5100 = 1'b0 ;
  assign y5101 = n21706 ;
  assign y5102 = n21709 ;
  assign y5103 = n21714 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = n21715 ;
  assign y5106 = ~n21716 ;
  assign y5107 = ~n21721 ;
  assign y5108 = ~n21724 ;
  assign y5109 = n21728 ;
  assign y5110 = ~n21735 ;
  assign y5111 = ~n21743 ;
  assign y5112 = ~n21744 ;
  assign y5113 = ~1'b0 ;
  assign y5114 = ~n21746 ;
  assign y5115 = ~n21750 ;
  assign y5116 = ~n21755 ;
  assign y5117 = ~n21758 ;
  assign y5118 = ~n21764 ;
  assign y5119 = n21766 ;
  assign y5120 = n21775 ;
  assign y5121 = n21778 ;
  assign y5122 = n21784 ;
  assign y5123 = n21788 ;
  assign y5124 = ~n21794 ;
  assign y5125 = n21796 ;
  assign y5126 = ~n21797 ;
  assign y5127 = n21803 ;
  assign y5128 = ~1'b0 ;
  assign y5129 = n21805 ;
  assign y5130 = n21813 ;
  assign y5131 = ~1'b0 ;
  assign y5132 = ~1'b0 ;
  assign y5133 = ~n21814 ;
  assign y5134 = n21817 ;
  assign y5135 = n21824 ;
  assign y5136 = ~n21827 ;
  assign y5137 = ~n21834 ;
  assign y5138 = n21838 ;
  assign y5139 = n21843 ;
  assign y5140 = ~1'b0 ;
  assign y5141 = n21844 ;
  assign y5142 = ~1'b0 ;
  assign y5143 = ~n21845 ;
  assign y5144 = ~n21849 ;
  assign y5145 = n21856 ;
  assign y5146 = ~n11110 ;
  assign y5147 = n21859 ;
  assign y5148 = ~1'b0 ;
  assign y5149 = n21860 ;
  assign y5150 = n21861 ;
  assign y5151 = n21863 ;
  assign y5152 = n21864 ;
  assign y5153 = n21868 ;
  assign y5154 = n21873 ;
  assign y5155 = n21876 ;
  assign y5156 = n21877 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = n21879 ;
  assign y5159 = ~n21881 ;
  assign y5160 = n21891 ;
  assign y5161 = n21893 ;
  assign y5162 = n21896 ;
  assign y5163 = ~n21899 ;
  assign y5164 = n21901 ;
  assign y5165 = n21904 ;
  assign y5166 = n21907 ;
  assign y5167 = ~n21913 ;
  assign y5168 = n21915 ;
  assign y5169 = ~n21922 ;
  assign y5170 = n21925 ;
  assign y5171 = ~n21926 ;
  assign y5172 = n21928 ;
  assign y5173 = ~n21932 ;
  assign y5174 = ~n21933 ;
  assign y5175 = ~n21938 ;
  assign y5176 = n21939 ;
  assign y5177 = n21940 ;
  assign y5178 = n21942 ;
  assign y5179 = ~n21947 ;
  assign y5180 = ~n21949 ;
  assign y5181 = n21953 ;
  assign y5182 = ~n21955 ;
  assign y5183 = n21959 ;
  assign y5184 = n21961 ;
  assign y5185 = ~n21963 ;
  assign y5186 = ~n21964 ;
  assign y5187 = ~n21965 ;
  assign y5188 = n21968 ;
  assign y5189 = n21977 ;
  assign y5190 = n21978 ;
  assign y5191 = n21984 ;
  assign y5192 = n21990 ;
  assign y5193 = n21999 ;
  assign y5194 = n22001 ;
  assign y5195 = ~1'b0 ;
  assign y5196 = n22005 ;
  assign y5197 = n22006 ;
  assign y5198 = n22008 ;
  assign y5199 = ~n22011 ;
  assign y5200 = n22016 ;
  assign y5201 = n22018 ;
  assign y5202 = n22021 ;
  assign y5203 = ~n22032 ;
  assign y5204 = ~n22037 ;
  assign y5205 = n22040 ;
  assign y5206 = n22045 ;
  assign y5207 = n22048 ;
  assign y5208 = ~n22051 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = ~n22053 ;
  assign y5211 = n22054 ;
  assign y5212 = ~n22056 ;
  assign y5213 = ~n22059 ;
  assign y5214 = ~1'b0 ;
  assign y5215 = ~1'b0 ;
  assign y5216 = ~n22060 ;
  assign y5217 = ~n22065 ;
  assign y5218 = ~1'b0 ;
  assign y5219 = ~1'b0 ;
  assign y5220 = ~n22071 ;
  assign y5221 = n22074 ;
  assign y5222 = ~1'b0 ;
  assign y5223 = n22079 ;
  assign y5224 = ~n22082 ;
  assign y5225 = n2401 ;
  assign y5226 = n17589 ;
  assign y5227 = ~n22084 ;
  assign y5228 = ~n22086 ;
  assign y5229 = ~n22090 ;
  assign y5230 = n22098 ;
  assign y5231 = n22104 ;
  assign y5232 = n22106 ;
  assign y5233 = ~n22110 ;
  assign y5234 = ~n22120 ;
  assign y5235 = ~n22124 ;
  assign y5236 = ~n22126 ;
  assign y5237 = n22129 ;
  assign y5238 = ~1'b0 ;
  assign y5239 = ~n22134 ;
  assign y5240 = n22143 ;
  assign y5241 = n22146 ;
  assign y5242 = n22147 ;
  assign y5243 = ~1'b0 ;
  assign y5244 = n22151 ;
  assign y5245 = n22153 ;
  assign y5246 = n22161 ;
  assign y5247 = ~n22162 ;
  assign y5248 = n22166 ;
  assign y5249 = ~n22183 ;
  assign y5250 = n22189 ;
  assign y5251 = ~n22194 ;
  assign y5252 = ~n22206 ;
  assign y5253 = ~n22207 ;
  assign y5254 = ~n22210 ;
  assign y5255 = ~1'b0 ;
  assign y5256 = n22212 ;
  assign y5257 = n22216 ;
  assign y5258 = n22220 ;
  assign y5259 = n22225 ;
  assign y5260 = n22229 ;
  assign y5261 = n22231 ;
  assign y5262 = n22232 ;
  assign y5263 = n22238 ;
  assign y5264 = ~n22246 ;
  assign y5265 = n22255 ;
  assign y5266 = ~n22258 ;
  assign y5267 = ~n16404 ;
  assign y5268 = ~1'b0 ;
  assign y5269 = ~n22264 ;
  assign y5270 = ~n21737 ;
  assign y5271 = ~n22267 ;
  assign y5272 = n22274 ;
  assign y5273 = ~n22277 ;
  assign y5274 = n22281 ;
  assign y5275 = n22283 ;
  assign y5276 = n22284 ;
  assign y5277 = ~n22289 ;
  assign y5278 = n22291 ;
  assign y5279 = ~n22292 ;
  assign y5280 = ~n22295 ;
  assign y5281 = ~n22298 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = ~n22301 ;
  assign y5284 = n22303 ;
  assign y5285 = ~n22306 ;
  assign y5286 = n22309 ;
  assign y5287 = ~n22315 ;
  assign y5288 = ~n22321 ;
  assign y5289 = ~n22331 ;
  assign y5290 = n22340 ;
  assign y5291 = ~n22341 ;
  assign y5292 = n22342 ;
  assign y5293 = ~n22345 ;
  assign y5294 = n22347 ;
  assign y5295 = ~n22349 ;
  assign y5296 = n22350 ;
  assign y5297 = n22353 ;
  assign y5298 = ~n22359 ;
  assign y5299 = ~n22361 ;
  assign y5300 = n22365 ;
  assign y5301 = n22368 ;
  assign y5302 = n22370 ;
  assign y5303 = n22374 ;
  assign y5304 = n22375 ;
  assign y5305 = n22111 ;
  assign y5306 = ~n22377 ;
  assign y5307 = ~n22381 ;
  assign y5308 = n22383 ;
  assign y5309 = ~n22389 ;
  assign y5310 = n22395 ;
  assign y5311 = n22399 ;
  assign y5312 = ~1'b0 ;
  assign y5313 = n22405 ;
  assign y5314 = n22406 ;
  assign y5315 = ~1'b0 ;
  assign y5316 = ~n22419 ;
  assign y5317 = n22420 ;
  assign y5318 = n22423 ;
  assign y5319 = ~n22430 ;
  assign y5320 = ~n22437 ;
  assign y5321 = ~n22439 ;
  assign y5322 = n22443 ;
  assign y5323 = ~n22444 ;
  assign y5324 = n22445 ;
  assign y5325 = n22447 ;
  assign y5326 = ~n22451 ;
  assign y5327 = ~n22455 ;
  assign y5328 = n7505 ;
  assign y5329 = ~n22459 ;
  assign y5330 = n22460 ;
  assign y5331 = n22471 ;
  assign y5332 = ~n22475 ;
  assign y5333 = ~n22477 ;
  assign y5334 = ~n22479 ;
  assign y5335 = n22480 ;
  assign y5336 = ~n22481 ;
  assign y5337 = n22483 ;
  assign y5338 = n22492 ;
  assign y5339 = ~n22495 ;
  assign y5340 = ~n22503 ;
  assign y5341 = ~n22511 ;
  assign y5342 = n22513 ;
  assign y5343 = n22514 ;
  assign y5344 = n22531 ;
  assign y5345 = n22538 ;
  assign y5346 = ~n22542 ;
  assign y5347 = n22546 ;
  assign y5348 = n22548 ;
  assign y5349 = ~n22550 ;
  assign y5350 = ~n22559 ;
  assign y5351 = n22565 ;
  assign y5352 = ~1'b0 ;
  assign y5353 = n22570 ;
  assign y5354 = n22574 ;
  assign y5355 = n22577 ;
  assign y5356 = ~1'b0 ;
  assign y5357 = ~n22580 ;
  assign y5358 = ~n22581 ;
  assign y5359 = n22583 ;
  assign y5360 = ~n22586 ;
  assign y5361 = ~n22587 ;
  assign y5362 = n22588 ;
  assign y5363 = n22596 ;
  assign y5364 = ~n22607 ;
  assign y5365 = ~n22608 ;
  assign y5366 = n22620 ;
  assign y5367 = ~n22633 ;
  assign y5368 = n22634 ;
  assign y5369 = ~n22639 ;
  assign y5370 = ~n22641 ;
  assign y5371 = ~n22645 ;
  assign y5372 = n22649 ;
  assign y5373 = n22652 ;
  assign y5374 = ~n22656 ;
  assign y5375 = n22657 ;
  assign y5376 = ~n22659 ;
  assign y5377 = n22660 ;
  assign y5378 = ~n22661 ;
  assign y5379 = ~1'b0 ;
  assign y5380 = n22662 ;
  assign y5381 = ~n22663 ;
  assign y5382 = ~n22668 ;
  assign y5383 = ~n22669 ;
  assign y5384 = n22674 ;
  assign y5385 = n22678 ;
  assign y5386 = n22680 ;
  assign y5387 = ~n22684 ;
  assign y5388 = ~n22689 ;
  assign y5389 = n22691 ;
  assign y5390 = ~n22693 ;
  assign y5391 = n22695 ;
  assign y5392 = ~n22696 ;
  assign y5393 = ~n22698 ;
  assign y5394 = ~n22699 ;
  assign y5395 = ~n22703 ;
  assign y5396 = n22707 ;
  assign y5397 = ~n22709 ;
  assign y5398 = ~n22711 ;
  assign y5399 = ~1'b0 ;
  assign y5400 = ~n22722 ;
  assign y5401 = ~n22723 ;
  assign y5402 = ~n22729 ;
  assign y5403 = ~1'b0 ;
  assign y5404 = n22731 ;
  assign y5405 = ~n22736 ;
  assign y5406 = ~n22738 ;
  assign y5407 = n22741 ;
  assign y5408 = n22746 ;
  assign y5409 = n22749 ;
  assign y5410 = ~n22753 ;
  assign y5411 = n22757 ;
  assign y5412 = ~n22758 ;
  assign y5413 = n22764 ;
  assign y5414 = n22771 ;
  assign y5415 = n22773 ;
  assign y5416 = n22775 ;
  assign y5417 = n22782 ;
  assign y5418 = n22789 ;
  assign y5419 = ~n22791 ;
  assign y5420 = n22793 ;
  assign y5421 = n22794 ;
  assign y5422 = ~n22798 ;
  assign y5423 = n22799 ;
  assign y5424 = ~n22805 ;
  assign y5425 = n22808 ;
  assign y5426 = ~n12880 ;
  assign y5427 = n22810 ;
  assign y5428 = ~1'b0 ;
  assign y5429 = ~n22814 ;
  assign y5430 = n22815 ;
  assign y5431 = ~n22821 ;
  assign y5432 = n22827 ;
  assign y5433 = n22828 ;
  assign y5434 = ~n22829 ;
  assign y5435 = ~n22838 ;
  assign y5436 = n22839 ;
  assign y5437 = n22845 ;
  assign y5438 = n22847 ;
  assign y5439 = ~n22849 ;
  assign y5440 = ~n22851 ;
  assign y5441 = n22864 ;
  assign y5442 = ~n22866 ;
  assign y5443 = ~n22871 ;
  assign y5444 = n22873 ;
  assign y5445 = ~n22876 ;
  assign y5446 = n22878 ;
  assign y5447 = n22880 ;
  assign y5448 = n22886 ;
  assign y5449 = ~n22889 ;
  assign y5450 = ~n22892 ;
  assign y5451 = ~n22893 ;
  assign y5452 = ~n22895 ;
  assign y5453 = n22896 ;
  assign y5454 = n22902 ;
  assign y5455 = n22906 ;
  assign y5456 = ~1'b0 ;
  assign y5457 = n22908 ;
  assign y5458 = n22911 ;
  assign y5459 = ~1'b0 ;
  assign y5460 = ~n22912 ;
  assign y5461 = n22914 ;
  assign y5462 = n22918 ;
  assign y5463 = ~1'b0 ;
  assign y5464 = n22929 ;
  assign y5465 = ~n22936 ;
  assign y5466 = ~n22939 ;
  assign y5467 = ~n22944 ;
  assign y5468 = ~n22945 ;
  assign y5469 = n22950 ;
  assign y5470 = ~n22954 ;
  assign y5471 = ~1'b0 ;
  assign y5472 = ~n22956 ;
  assign y5473 = n22958 ;
  assign y5474 = n22963 ;
  assign y5475 = ~1'b0 ;
  assign y5476 = n22966 ;
  assign y5477 = n22968 ;
  assign y5478 = n22970 ;
  assign y5479 = n22974 ;
  assign y5480 = ~n22977 ;
  assign y5481 = ~n22980 ;
  assign y5482 = ~n22984 ;
  assign y5483 = n22988 ;
  assign y5484 = ~n22990 ;
  assign y5485 = ~n22994 ;
  assign y5486 = ~n22998 ;
  assign y5487 = ~n22999 ;
  assign y5488 = n23005 ;
  assign y5489 = ~n19685 ;
  assign y5490 = n23006 ;
  assign y5491 = n23008 ;
  assign y5492 = ~n23009 ;
  assign y5493 = n23014 ;
  assign y5494 = ~n23015 ;
  assign y5495 = ~n23025 ;
  assign y5496 = ~n23027 ;
  assign y5497 = n23029 ;
  assign y5498 = ~1'b0 ;
  assign y5499 = ~n23035 ;
  assign y5500 = ~n23039 ;
  assign y5501 = ~n23042 ;
  assign y5502 = ~n23044 ;
  assign y5503 = ~n23045 ;
  assign y5504 = ~n23054 ;
  assign y5505 = n23059 ;
  assign y5506 = n23060 ;
  assign y5507 = n23063 ;
  assign y5508 = ~1'b0 ;
  assign y5509 = ~n23064 ;
  assign y5510 = n23071 ;
  assign y5511 = n23073 ;
  assign y5512 = ~1'b0 ;
  assign y5513 = ~1'b0 ;
  assign y5514 = n23078 ;
  assign y5515 = ~n23086 ;
  assign y5516 = n23094 ;
  assign y5517 = n23097 ;
  assign y5518 = ~n23100 ;
  assign y5519 = ~n23101 ;
  assign y5520 = n23104 ;
  assign y5521 = ~n23105 ;
  assign y5522 = n23108 ;
  assign y5523 = ~n23110 ;
  assign y5524 = ~n23112 ;
  assign y5525 = n23117 ;
  assign y5526 = ~n23128 ;
  assign y5527 = ~n23131 ;
  assign y5528 = n23137 ;
  assign y5529 = n23139 ;
  assign y5530 = ~n23140 ;
  assign y5531 = ~n23145 ;
  assign y5532 = n23146 ;
  assign y5533 = n23154 ;
  assign y5534 = ~n2130 ;
  assign y5535 = n23155 ;
  assign y5536 = n23158 ;
  assign y5537 = ~n23160 ;
  assign y5538 = ~n23164 ;
  assign y5539 = ~n23176 ;
  assign y5540 = ~n23180 ;
  assign y5541 = ~1'b0 ;
  assign y5542 = ~n23195 ;
  assign y5543 = n23198 ;
  assign y5544 = ~1'b0 ;
  assign y5545 = n23202 ;
  assign y5546 = n23203 ;
  assign y5547 = ~n23206 ;
  assign y5548 = n23207 ;
  assign y5549 = n23218 ;
  assign y5550 = n23224 ;
  assign y5551 = 1'b0 ;
  assign y5552 = ~n23227 ;
  assign y5553 = n23228 ;
  assign y5554 = ~n23230 ;
  assign y5555 = ~n23236 ;
  assign y5556 = n23238 ;
  assign y5557 = n23239 ;
  assign y5558 = ~n23243 ;
  assign y5559 = ~n23257 ;
  assign y5560 = ~n23258 ;
  assign y5561 = n23261 ;
  assign y5562 = ~n23263 ;
  assign y5563 = ~1'b0 ;
  assign y5564 = n23267 ;
  assign y5565 = ~n23269 ;
  assign y5566 = n23273 ;
  assign y5567 = n14267 ;
  assign y5568 = ~n23279 ;
  assign y5569 = n23283 ;
  assign y5570 = n23284 ;
  assign y5571 = ~n23285 ;
  assign y5572 = n23299 ;
  assign y5573 = ~n23303 ;
  assign y5574 = ~1'b0 ;
  assign y5575 = ~n23305 ;
  assign y5576 = n14047 ;
  assign y5577 = ~n23306 ;
  assign y5578 = n23311 ;
  assign y5579 = n23313 ;
  assign y5580 = ~1'b0 ;
  assign y5581 = n23316 ;
  assign y5582 = ~n23320 ;
  assign y5583 = n23323 ;
  assign y5584 = n23324 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = ~n23326 ;
  assign y5587 = n23329 ;
  assign y5588 = n23334 ;
  assign y5589 = n23337 ;
  assign y5590 = n23339 ;
  assign y5591 = n23344 ;
  assign y5592 = ~n23346 ;
  assign y5593 = n23347 ;
  assign y5594 = n23350 ;
  assign y5595 = n23358 ;
  assign y5596 = n23362 ;
  assign y5597 = ~n23367 ;
  assign y5598 = ~n23373 ;
  assign y5599 = ~n23377 ;
  assign y5600 = ~n23379 ;
  assign y5601 = ~1'b0 ;
  assign y5602 = n23382 ;
  assign y5603 = n23384 ;
  assign y5604 = ~n23385 ;
  assign y5605 = n23389 ;
  assign y5606 = n23392 ;
  assign y5607 = n23400 ;
  assign y5608 = n23401 ;
  assign y5609 = ~n23404 ;
  assign y5610 = ~n23405 ;
  assign y5611 = ~n23406 ;
  assign y5612 = n23408 ;
  assign y5613 = n23417 ;
  assign y5614 = n23422 ;
  assign y5615 = n23424 ;
  assign y5616 = n23427 ;
  assign y5617 = n23432 ;
  assign y5618 = ~n23434 ;
  assign y5619 = ~n23437 ;
  assign y5620 = ~n23443 ;
  assign y5621 = ~n23445 ;
  assign y5622 = n23458 ;
  assign y5623 = n23462 ;
  assign y5624 = ~n23468 ;
  assign y5625 = n23470 ;
  assign y5626 = n23474 ;
  assign y5627 = n23476 ;
  assign y5628 = ~n23482 ;
  assign y5629 = ~1'b0 ;
  assign y5630 = ~n23484 ;
  assign y5631 = n23485 ;
  assign y5632 = ~n23489 ;
  assign y5633 = n23491 ;
  assign y5634 = ~1'b0 ;
  assign y5635 = ~1'b0 ;
  assign y5636 = ~n23499 ;
  assign y5637 = n23508 ;
  assign y5638 = ~1'b0 ;
  assign y5639 = ~n23513 ;
  assign y5640 = ~1'b0 ;
  assign y5641 = n23514 ;
  assign y5642 = ~n23515 ;
  assign y5643 = ~n23519 ;
  assign y5644 = n23520 ;
  assign y5645 = n23525 ;
  assign y5646 = ~n23527 ;
  assign y5647 = ~n23529 ;
  assign y5648 = n23534 ;
  assign y5649 = n23536 ;
  assign y5650 = n23545 ;
  assign y5651 = ~1'b0 ;
  assign y5652 = n23548 ;
  assign y5653 = n23550 ;
  assign y5654 = ~n23551 ;
  assign y5655 = ~n23554 ;
  assign y5656 = ~1'b0 ;
  assign y5657 = n23556 ;
  assign y5658 = n23559 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = ~n23563 ;
  assign y5661 = ~n23572 ;
  assign y5662 = ~n23575 ;
  assign y5663 = ~n23580 ;
  assign y5664 = ~n1515 ;
  assign y5665 = n23581 ;
  assign y5666 = n23583 ;
  assign y5667 = ~n23585 ;
  assign y5668 = ~n23586 ;
  assign y5669 = n23588 ;
  assign y5670 = ~n23590 ;
  assign y5671 = n18892 ;
  assign y5672 = ~n23595 ;
  assign y5673 = n23600 ;
  assign y5674 = n23602 ;
  assign y5675 = n23606 ;
  assign y5676 = ~n23609 ;
  assign y5677 = n23616 ;
  assign y5678 = n23617 ;
  assign y5679 = ~n23618 ;
  assign y5680 = ~n23625 ;
  assign y5681 = ~n23629 ;
  assign y5682 = ~n23638 ;
  assign y5683 = ~n23643 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = ~1'b0 ;
  assign y5686 = n23646 ;
  assign y5687 = ~n23647 ;
  assign y5688 = ~1'b0 ;
  assign y5689 = ~n23655 ;
  assign y5690 = n23656 ;
  assign y5691 = n23658 ;
  assign y5692 = n23668 ;
  assign y5693 = n23670 ;
  assign y5694 = ~n23675 ;
  assign y5695 = ~n23677 ;
  assign y5696 = n23683 ;
  assign y5697 = n23689 ;
  assign y5698 = n23692 ;
  assign y5699 = n23693 ;
  assign y5700 = ~n23696 ;
  assign y5701 = n23703 ;
  assign y5702 = ~1'b0 ;
  assign y5703 = n23711 ;
  assign y5704 = ~1'b0 ;
  assign y5705 = ~n23714 ;
  assign y5706 = ~n23719 ;
  assign y5707 = n23720 ;
  assign y5708 = n23723 ;
  assign y5709 = n23725 ;
  assign y5710 = n23728 ;
  assign y5711 = ~1'b0 ;
  assign y5712 = n23729 ;
  assign y5713 = n23732 ;
  assign y5714 = ~n23733 ;
  assign y5715 = n23743 ;
  assign y5716 = n23745 ;
  assign y5717 = n23750 ;
  assign y5718 = n23751 ;
  assign y5719 = n23764 ;
  assign y5720 = n23767 ;
  assign y5721 = ~n23769 ;
  assign y5722 = ~n23770 ;
  assign y5723 = ~n23775 ;
  assign y5724 = ~1'b0 ;
  assign y5725 = n23778 ;
  assign y5726 = n23779 ;
  assign y5727 = ~n23788 ;
  assign y5728 = ~n23789 ;
  assign y5729 = ~n23792 ;
  assign y5730 = ~n23794 ;
  assign y5731 = n23796 ;
  assign y5732 = ~n23800 ;
  assign y5733 = ~n23807 ;
  assign y5734 = n23808 ;
  assign y5735 = ~n23811 ;
  assign y5736 = n23812 ;
  assign y5737 = ~n23817 ;
  assign y5738 = n23819 ;
  assign y5739 = n23826 ;
  assign y5740 = n23841 ;
  assign y5741 = n23844 ;
  assign y5742 = ~n23847 ;
  assign y5743 = n23852 ;
  assign y5744 = ~n23855 ;
  assign y5745 = n23857 ;
  assign y5746 = n23858 ;
  assign y5747 = n23864 ;
  assign y5748 = n23866 ;
  assign y5749 = n23869 ;
  assign y5750 = ~n23880 ;
  assign y5751 = n23883 ;
  assign y5752 = n1133 ;
  assign y5753 = ~1'b0 ;
  assign y5754 = ~n23884 ;
  assign y5755 = ~1'b0 ;
  assign y5756 = ~n23885 ;
  assign y5757 = ~n23890 ;
  assign y5758 = n23891 ;
  assign y5759 = n23892 ;
  assign y5760 = ~n23900 ;
  assign y5761 = n23906 ;
  assign y5762 = n23909 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = ~n23911 ;
  assign y5765 = ~n23912 ;
  assign y5766 = n2979 ;
  assign y5767 = n23917 ;
  assign y5768 = ~n23918 ;
  assign y5769 = ~1'b0 ;
  assign y5770 = n23920 ;
  assign y5771 = n23921 ;
  assign y5772 = ~1'b0 ;
  assign y5773 = ~n23927 ;
  assign y5774 = ~1'b0 ;
  assign y5775 = n23930 ;
  assign y5776 = ~n23936 ;
  assign y5777 = ~1'b0 ;
  assign y5778 = n23937 ;
  assign y5779 = n23938 ;
  assign y5780 = n23940 ;
  assign y5781 = n23941 ;
  assign y5782 = n23945 ;
  assign y5783 = n23946 ;
  assign y5784 = ~1'b0 ;
  assign y5785 = ~n23954 ;
  assign y5786 = ~n23958 ;
  assign y5787 = ~n11553 ;
  assign y5788 = n23959 ;
  assign y5789 = n23971 ;
  assign y5790 = ~n23972 ;
  assign y5791 = ~n23976 ;
  assign y5792 = ~n23977 ;
  assign y5793 = n23981 ;
  assign y5794 = ~1'b0 ;
  assign y5795 = n23996 ;
  assign y5796 = n24001 ;
  assign y5797 = ~n24004 ;
  assign y5798 = n24009 ;
  assign y5799 = ~n24014 ;
  assign y5800 = ~n24022 ;
  assign y5801 = n24037 ;
  assign y5802 = n24041 ;
  assign y5803 = n24043 ;
  assign y5804 = ~n24047 ;
  assign y5805 = n24049 ;
  assign y5806 = ~n24058 ;
  assign y5807 = n24059 ;
  assign y5808 = ~n24064 ;
  assign y5809 = ~n24066 ;
  assign y5810 = ~n24071 ;
  assign y5811 = ~n24073 ;
  assign y5812 = ~n24079 ;
  assign y5813 = ~n24081 ;
  assign y5814 = ~n24090 ;
  assign y5815 = ~1'b0 ;
  assign y5816 = ~n24095 ;
  assign y5817 = n18010 ;
  assign y5818 = ~n24096 ;
  assign y5819 = ~n24101 ;
  assign y5820 = n24102 ;
  assign y5821 = ~n24104 ;
  assign y5822 = ~n24108 ;
  assign y5823 = n24109 ;
  assign y5824 = ~1'b0 ;
  assign y5825 = ~n24113 ;
  assign y5826 = n24119 ;
  assign y5827 = n24120 ;
  assign y5828 = ~n24121 ;
  assign y5829 = ~1'b0 ;
  assign y5830 = ~n24124 ;
  assign y5831 = n24129 ;
  assign y5832 = n24130 ;
  assign y5833 = ~n24131 ;
  assign y5834 = ~n24133 ;
  assign y5835 = n24146 ;
  assign y5836 = n24153 ;
  assign y5837 = ~n24158 ;
  assign y5838 = n24164 ;
  assign y5839 = ~n24165 ;
  assign y5840 = n24172 ;
  assign y5841 = ~n24174 ;
  assign y5842 = ~n24177 ;
  assign y5843 = n24182 ;
  assign y5844 = ~n24188 ;
  assign y5845 = n24191 ;
  assign y5846 = n24195 ;
  assign y5847 = ~1'b0 ;
  assign y5848 = n24199 ;
  assign y5849 = ~n24200 ;
  assign y5850 = n24216 ;
  assign y5851 = ~1'b0 ;
  assign y5852 = ~n24223 ;
  assign y5853 = ~n24225 ;
  assign y5854 = ~n24226 ;
  assign y5855 = n24237 ;
  assign y5856 = ~n24243 ;
  assign y5857 = n24250 ;
  assign y5858 = ~1'b0 ;
  assign y5859 = ~n24253 ;
  assign y5860 = ~n24254 ;
  assign y5861 = ~n24255 ;
  assign y5862 = ~1'b0 ;
  assign y5863 = ~n24258 ;
  assign y5864 = ~n24262 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = ~n24263 ;
  assign y5867 = n24268 ;
  assign y5868 = ~n24274 ;
  assign y5869 = ~n24277 ;
  assign y5870 = ~n24282 ;
  assign y5871 = ~n24285 ;
  assign y5872 = ~1'b0 ;
  assign y5873 = ~n24287 ;
  assign y5874 = n24289 ;
  assign y5875 = ~n24293 ;
  assign y5876 = ~1'b0 ;
  assign y5877 = n24296 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = n24300 ;
  assign y5880 = ~n24302 ;
  assign y5881 = ~n24308 ;
  assign y5882 = ~n24309 ;
  assign y5883 = ~n24314 ;
  assign y5884 = ~n24322 ;
  assign y5885 = n24324 ;
  assign y5886 = ~n24326 ;
  assign y5887 = ~n24328 ;
  assign y5888 = ~n24330 ;
  assign y5889 = ~n24331 ;
  assign y5890 = n24336 ;
  assign y5891 = n24339 ;
  assign y5892 = ~1'b0 ;
  assign y5893 = ~n24340 ;
  assign y5894 = ~n24353 ;
  assign y5895 = n24356 ;
  assign y5896 = ~1'b0 ;
  assign y5897 = ~n24360 ;
  assign y5898 = ~n24364 ;
  assign y5899 = ~n24365 ;
  assign y5900 = n24368 ;
  assign y5901 = ~n24370 ;
  assign y5902 = ~n24373 ;
  assign y5903 = ~n24379 ;
  assign y5904 = n24397 ;
  assign y5905 = 1'b0 ;
  assign y5906 = ~n24398 ;
  assign y5907 = n24399 ;
  assign y5908 = ~n24400 ;
  assign y5909 = ~n24401 ;
  assign y5910 = ~1'b0 ;
  assign y5911 = ~1'b0 ;
  assign y5912 = n24404 ;
  assign y5913 = n24405 ;
  assign y5914 = ~n24410 ;
  assign y5915 = n24419 ;
  assign y5916 = ~1'b0 ;
  assign y5917 = ~n24434 ;
  assign y5918 = ~n24436 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = n24438 ;
  assign y5921 = n24441 ;
  assign y5922 = n24445 ;
  assign y5923 = n24449 ;
  assign y5924 = n24450 ;
  assign y5925 = ~n24453 ;
  assign y5926 = ~n24455 ;
  assign y5927 = ~n24457 ;
  assign y5928 = ~n24462 ;
  assign y5929 = ~n24465 ;
  assign y5930 = ~n24469 ;
  assign y5931 = ~n24470 ;
  assign y5932 = ~n24471 ;
  assign y5933 = ~n24472 ;
  assign y5934 = n24473 ;
  assign y5935 = n24480 ;
  assign y5936 = ~n24481 ;
  assign y5937 = ~1'b0 ;
  assign y5938 = n24482 ;
  assign y5939 = n24489 ;
  assign y5940 = ~n24494 ;
  assign y5941 = n21483 ;
  assign y5942 = ~n24495 ;
  assign y5943 = ~n24501 ;
  assign y5944 = ~n24504 ;
  assign y5945 = n24510 ;
  assign y5946 = ~n24512 ;
  assign y5947 = n24517 ;
  assign y5948 = ~n24529 ;
  assign y5949 = ~n24532 ;
  assign y5950 = ~1'b0 ;
  assign y5951 = ~n24534 ;
  assign y5952 = n24538 ;
  assign y5953 = ~n24539 ;
  assign y5954 = ~n24545 ;
  assign y5955 = n24553 ;
  assign y5956 = ~n24557 ;
  assign y5957 = ~n24566 ;
  assign y5958 = ~1'b0 ;
  assign y5959 = ~n24568 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = n24570 ;
  assign y5962 = ~n24577 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = n24579 ;
  assign y5965 = n24590 ;
  assign y5966 = ~n24591 ;
  assign y5967 = ~n24598 ;
  assign y5968 = n24602 ;
  assign y5969 = ~n24607 ;
  assign y5970 = ~n24609 ;
  assign y5971 = ~n24612 ;
  assign y5972 = ~n24614 ;
  assign y5973 = ~n24616 ;
  assign y5974 = ~n24623 ;
  assign y5975 = ~n24629 ;
  assign y5976 = ~n24630 ;
  assign y5977 = ~n24634 ;
  assign y5978 = ~n24651 ;
  assign y5979 = n24654 ;
  assign y5980 = ~1'b0 ;
  assign y5981 = n24658 ;
  assign y5982 = ~1'b0 ;
  assign y5983 = ~n24663 ;
  assign y5984 = ~n24669 ;
  assign y5985 = ~1'b0 ;
  assign y5986 = ~n24674 ;
  assign y5987 = ~x76 ;
  assign y5988 = ~n24677 ;
  assign y5989 = ~n24679 ;
  assign y5990 = n24683 ;
  assign y5991 = n24688 ;
  assign y5992 = n24689 ;
  assign y5993 = n24690 ;
  assign y5994 = ~n24695 ;
  assign y5995 = n24696 ;
  assign y5996 = ~n24710 ;
  assign y5997 = n24713 ;
  assign y5998 = ~n24714 ;
  assign y5999 = ~n24720 ;
  assign y6000 = n24721 ;
  assign y6001 = n24727 ;
  assign y6002 = n24729 ;
  assign y6003 = ~n24732 ;
  assign y6004 = ~n24734 ;
  assign y6005 = n24739 ;
  assign y6006 = n24749 ;
  assign y6007 = ~1'b0 ;
  assign y6008 = n24750 ;
  assign y6009 = ~n24753 ;
  assign y6010 = ~1'b0 ;
  assign y6011 = ~n24755 ;
  assign y6012 = n24757 ;
  assign y6013 = ~n24766 ;
  assign y6014 = n24773 ;
  assign y6015 = ~n24775 ;
  assign y6016 = ~n24776 ;
  assign y6017 = ~n24778 ;
  assign y6018 = ~n24783 ;
  assign y6019 = n24784 ;
  assign y6020 = ~n24785 ;
  assign y6021 = ~n24786 ;
  assign y6022 = n24788 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = ~n24790 ;
  assign y6025 = ~n24793 ;
  assign y6026 = n24797 ;
  assign y6027 = ~n24800 ;
  assign y6028 = ~n24804 ;
  assign y6029 = ~n24805 ;
  assign y6030 = n24817 ;
  assign y6031 = ~n24819 ;
  assign y6032 = n24820 ;
  assign y6033 = n24826 ;
  assign y6034 = ~n24831 ;
  assign y6035 = n24833 ;
  assign y6036 = ~n1773 ;
  assign y6037 = ~n24834 ;
  assign y6038 = n24835 ;
  assign y6039 = ~n24837 ;
  assign y6040 = ~n24843 ;
  assign y6041 = ~n24846 ;
  assign y6042 = ~n24849 ;
  assign y6043 = ~n24853 ;
  assign y6044 = n24860 ;
  assign y6045 = ~1'b0 ;
  assign y6046 = ~n24866 ;
  assign y6047 = ~n24868 ;
  assign y6048 = ~n24869 ;
  assign y6049 = n24870 ;
  assign y6050 = n24875 ;
  assign y6051 = ~n24878 ;
  assign y6052 = n24886 ;
  assign y6053 = ~1'b0 ;
  assign y6054 = ~n24888 ;
  assign y6055 = n24890 ;
  assign y6056 = ~n24899 ;
  assign y6057 = ~n24900 ;
  assign y6058 = ~n24901 ;
  assign y6059 = ~n24902 ;
  assign y6060 = ~n24905 ;
  assign y6061 = ~n24906 ;
  assign y6062 = ~n24909 ;
  assign y6063 = n24917 ;
  assign y6064 = n24919 ;
  assign y6065 = n24923 ;
  assign y6066 = ~1'b0 ;
  assign y6067 = ~1'b0 ;
  assign y6068 = n24929 ;
  assign y6069 = n24933 ;
  assign y6070 = ~n24934 ;
  assign y6071 = ~n24937 ;
  assign y6072 = ~n24938 ;
  assign y6073 = ~n24940 ;
  assign y6074 = n24947 ;
  assign y6075 = n24948 ;
  assign y6076 = n24949 ;
  assign y6077 = n24951 ;
  assign y6078 = ~n24953 ;
  assign y6079 = ~1'b0 ;
  assign y6080 = ~n24958 ;
  assign y6081 = n24962 ;
  assign y6082 = n24964 ;
  assign y6083 = n24969 ;
  assign y6084 = ~n24970 ;
  assign y6085 = n24973 ;
  assign y6086 = n24978 ;
  assign y6087 = n24979 ;
  assign y6088 = n24986 ;
  assign y6089 = ~n24989 ;
  assign y6090 = ~n24990 ;
  assign y6091 = ~n24992 ;
  assign y6092 = ~n24994 ;
  assign y6093 = ~n24998 ;
  assign y6094 = ~n24999 ;
  assign y6095 = ~n25002 ;
  assign y6096 = n25006 ;
  assign y6097 = n25009 ;
  assign y6098 = ~n25011 ;
  assign y6099 = n25013 ;
  assign y6100 = ~n25015 ;
  assign y6101 = ~1'b0 ;
  assign y6102 = n25016 ;
  assign y6103 = n25020 ;
  assign y6104 = n25033 ;
  assign y6105 = ~n25037 ;
  assign y6106 = n25047 ;
  assign y6107 = n25048 ;
  assign y6108 = n25052 ;
  assign y6109 = n25054 ;
  assign y6110 = ~1'b0 ;
  assign y6111 = ~n25061 ;
  assign y6112 = ~n25065 ;
  assign y6113 = n25066 ;
  assign y6114 = ~n25068 ;
  assign y6115 = n25070 ;
  assign y6116 = ~n25072 ;
  assign y6117 = ~n25073 ;
  assign y6118 = n25081 ;
  assign y6119 = ~n25084 ;
  assign y6120 = ~n25085 ;
  assign y6121 = n25086 ;
  assign y6122 = n25087 ;
  assign y6123 = ~n25093 ;
  assign y6124 = ~n25100 ;
  assign y6125 = n25102 ;
  assign y6126 = ~n25104 ;
  assign y6127 = ~n25106 ;
  assign y6128 = n25108 ;
  assign y6129 = n25115 ;
  assign y6130 = n25124 ;
  assign y6131 = ~n25125 ;
  assign y6132 = ~1'b0 ;
  assign y6133 = ~n25126 ;
  assign y6134 = ~n25133 ;
  assign y6135 = n25143 ;
  assign y6136 = ~n25144 ;
  assign y6137 = ~n25146 ;
  assign y6138 = ~n25155 ;
  assign y6139 = ~n25159 ;
  assign y6140 = n25165 ;
  assign y6141 = ~n25169 ;
  assign y6142 = n25172 ;
  assign y6143 = n25181 ;
  assign y6144 = ~1'b0 ;
  assign y6145 = ~1'b0 ;
  assign y6146 = ~n25184 ;
  assign y6147 = n25185 ;
  assign y6148 = n13962 ;
  assign y6149 = ~n25189 ;
  assign y6150 = n25190 ;
  assign y6151 = ~n25191 ;
  assign y6152 = ~n25195 ;
  assign y6153 = n25202 ;
  assign y6154 = n25204 ;
  assign y6155 = ~1'b0 ;
  assign y6156 = ~n25210 ;
  assign y6157 = ~n25216 ;
  assign y6158 = ~n25224 ;
  assign y6159 = n25230 ;
  assign y6160 = n25237 ;
  assign y6161 = ~n25253 ;
  assign y6162 = n25254 ;
  assign y6163 = ~n25255 ;
  assign y6164 = n25260 ;
  assign y6165 = n25262 ;
  assign y6166 = n25266 ;
  assign y6167 = ~n25268 ;
  assign y6168 = ~1'b0 ;
  assign y6169 = ~n25269 ;
  assign y6170 = n25271 ;
  assign y6171 = ~1'b0 ;
  assign y6172 = ~1'b0 ;
  assign y6173 = n25276 ;
  assign y6174 = ~n25278 ;
  assign y6175 = n25280 ;
  assign y6176 = ~n25285 ;
  assign y6177 = n25286 ;
  assign y6178 = n25293 ;
  assign y6179 = ~n25294 ;
  assign y6180 = n25295 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = ~n25298 ;
  assign y6183 = n25299 ;
  assign y6184 = ~n25300 ;
  assign y6185 = n25302 ;
  assign y6186 = ~n25307 ;
  assign y6187 = n25315 ;
  assign y6188 = n25317 ;
  assign y6189 = ~n25323 ;
  assign y6190 = n25325 ;
  assign y6191 = n25327 ;
  assign y6192 = ~n25330 ;
  assign y6193 = n25333 ;
  assign y6194 = ~n25338 ;
  assign y6195 = ~n25345 ;
  assign y6196 = ~1'b0 ;
  assign y6197 = ~n25348 ;
  assign y6198 = n25353 ;
  assign y6199 = 1'b0 ;
  assign y6200 = n25361 ;
  assign y6201 = n25363 ;
  assign y6202 = ~n25367 ;
  assign y6203 = ~n25373 ;
  assign y6204 = ~n25386 ;
  assign y6205 = ~n25389 ;
  assign y6206 = ~n25394 ;
  assign y6207 = n25401 ;
  assign y6208 = n25406 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = n25412 ;
  assign y6211 = ~n25417 ;
  assign y6212 = ~n25418 ;
  assign y6213 = n25424 ;
  assign y6214 = ~n25427 ;
  assign y6215 = ~n25434 ;
  assign y6216 = ~n25437 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = ~n25438 ;
  assign y6219 = n25440 ;
  assign y6220 = ~n25441 ;
  assign y6221 = ~n25443 ;
  assign y6222 = ~n25448 ;
  assign y6223 = ~n25454 ;
  assign y6224 = ~n25463 ;
  assign y6225 = ~n25469 ;
  assign y6226 = ~n25471 ;
  assign y6227 = ~n25472 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = ~n25473 ;
  assign y6230 = n25474 ;
  assign y6231 = n25485 ;
  assign y6232 = n25491 ;
  assign y6233 = n25494 ;
  assign y6234 = ~n25496 ;
  assign y6235 = ~n25498 ;
  assign y6236 = n25501 ;
  assign y6237 = ~1'b0 ;
  assign y6238 = ~n25502 ;
  assign y6239 = n25504 ;
  assign y6240 = n25511 ;
  assign y6241 = n25513 ;
  assign y6242 = ~n25517 ;
  assign y6243 = ~1'b0 ;
  assign y6244 = ~1'b0 ;
  assign y6245 = ~n25524 ;
  assign y6246 = n25528 ;
  assign y6247 = ~n25529 ;
  assign y6248 = ~n25530 ;
  assign y6249 = n25531 ;
  assign y6250 = ~1'b0 ;
  assign y6251 = n25537 ;
  assign y6252 = ~n25540 ;
  assign y6253 = n25545 ;
  assign y6254 = n25547 ;
  assign y6255 = ~n25552 ;
  assign y6256 = ~n25553 ;
  assign y6257 = ~n25557 ;
  assign y6258 = ~n25561 ;
  assign y6259 = ~n25566 ;
  assign y6260 = ~n25567 ;
  assign y6261 = ~1'b0 ;
  assign y6262 = ~1'b0 ;
  assign y6263 = n25572 ;
  assign y6264 = ~n25576 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = n25577 ;
  assign y6267 = n25578 ;
  assign y6268 = ~1'b0 ;
  assign y6269 = ~n25581 ;
  assign y6270 = n25585 ;
  assign y6271 = n25591 ;
  assign y6272 = n25603 ;
  assign y6273 = ~n25605 ;
  assign y6274 = ~n25607 ;
  assign y6275 = ~n25611 ;
  assign y6276 = n25612 ;
  assign y6277 = n25613 ;
  assign y6278 = n25617 ;
  assign y6279 = n25618 ;
  assign y6280 = n25625 ;
  assign y6281 = n25626 ;
  assign y6282 = n25627 ;
  assign y6283 = ~n25634 ;
  assign y6284 = ~n25643 ;
  assign y6285 = ~n25644 ;
  assign y6286 = ~n25648 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = n25651 ;
  assign y6289 = n25656 ;
  assign y6290 = n25658 ;
  assign y6291 = n25664 ;
  assign y6292 = ~n25666 ;
  assign y6293 = n25668 ;
  assign y6294 = 1'b0 ;
  assign y6295 = ~1'b0 ;
  assign y6296 = n25670 ;
  assign y6297 = n25672 ;
  assign y6298 = n25679 ;
  assign y6299 = ~n25680 ;
  assign y6300 = ~1'b0 ;
  assign y6301 = ~n25684 ;
  assign y6302 = ~n25688 ;
  assign y6303 = n25691 ;
  assign y6304 = n25692 ;
  assign y6305 = n25696 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = n25702 ;
  assign y6308 = ~1'b0 ;
  assign y6309 = ~n25705 ;
  assign y6310 = n25707 ;
  assign y6311 = ~n25715 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = ~n25717 ;
  assign y6314 = n25718 ;
  assign y6315 = ~1'b0 ;
  assign y6316 = ~1'b0 ;
  assign y6317 = ~n25723 ;
  assign y6318 = ~n25724 ;
  assign y6319 = n25725 ;
  assign y6320 = ~n25731 ;
  assign y6321 = ~1'b0 ;
  assign y6322 = n25737 ;
  assign y6323 = n25742 ;
  assign y6324 = n25747 ;
  assign y6325 = ~n25748 ;
  assign y6326 = n25750 ;
  assign y6327 = n25758 ;
  assign y6328 = n25759 ;
  assign y6329 = n25760 ;
  assign y6330 = ~n25762 ;
  assign y6331 = ~n25768 ;
  assign y6332 = ~n25770 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = n25771 ;
  assign y6335 = ~n25776 ;
  assign y6336 = n25777 ;
  assign y6337 = ~n25779 ;
  assign y6338 = ~n25781 ;
  assign y6339 = ~n25782 ;
  assign y6340 = n25783 ;
  assign y6341 = ~n25786 ;
  assign y6342 = n25790 ;
  assign y6343 = ~n25793 ;
  assign y6344 = ~n25794 ;
  assign y6345 = ~n25796 ;
  assign y6346 = ~n25799 ;
  assign y6347 = ~n25804 ;
  assign y6348 = n25808 ;
  assign y6349 = ~1'b0 ;
  assign y6350 = ~n25817 ;
  assign y6351 = n25824 ;
  assign y6352 = ~1'b0 ;
  assign y6353 = ~1'b0 ;
  assign y6354 = n25826 ;
  assign y6355 = n25837 ;
  assign y6356 = ~n25840 ;
  assign y6357 = ~n25842 ;
  assign y6358 = ~n25843 ;
  assign y6359 = ~n8588 ;
  assign y6360 = ~n25850 ;
  assign y6361 = n25851 ;
  assign y6362 = ~1'b0 ;
  assign y6363 = ~1'b0 ;
  assign y6364 = ~n25856 ;
  assign y6365 = n25857 ;
  assign y6366 = ~n25859 ;
  assign y6367 = n25865 ;
  assign y6368 = n25866 ;
  assign y6369 = n25868 ;
  assign y6370 = n25874 ;
  assign y6371 = n25881 ;
  assign y6372 = ~n25885 ;
  assign y6373 = ~1'b0 ;
  assign y6374 = n25893 ;
  assign y6375 = ~n25895 ;
  assign y6376 = ~n25898 ;
  assign y6377 = ~n25899 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = ~n25903 ;
  assign y6380 = n25907 ;
  assign y6381 = n25909 ;
  assign y6382 = n25910 ;
  assign y6383 = n25911 ;
  assign y6384 = ~1'b0 ;
  assign y6385 = ~n25913 ;
  assign y6386 = ~n25919 ;
  assign y6387 = n25922 ;
  assign y6388 = n25924 ;
  assign y6389 = ~n25927 ;
  assign y6390 = n25932 ;
  assign y6391 = n25934 ;
  assign y6392 = n25938 ;
  assign y6393 = ~n25951 ;
  assign y6394 = n25953 ;
  assign y6395 = n25958 ;
  assign y6396 = n25968 ;
  assign y6397 = n25970 ;
  assign y6398 = ~n25971 ;
  assign y6399 = ~n25973 ;
  assign y6400 = ~n25977 ;
  assign y6401 = ~n25979 ;
  assign y6402 = n25982 ;
  assign y6403 = n25987 ;
  assign y6404 = ~1'b0 ;
  assign y6405 = ~n25990 ;
  assign y6406 = ~n25997 ;
  assign y6407 = n25999 ;
  assign y6408 = ~n26006 ;
  assign y6409 = ~n26016 ;
  assign y6410 = ~n26019 ;
  assign y6411 = n26024 ;
  assign y6412 = ~1'b0 ;
  assign y6413 = n26028 ;
  assign y6414 = ~n26029 ;
  assign y6415 = n26033 ;
  assign y6416 = ~n26039 ;
  assign y6417 = n26040 ;
  assign y6418 = ~n26045 ;
  assign y6419 = ~n26049 ;
  assign y6420 = ~n26053 ;
  assign y6421 = ~n26061 ;
  assign y6422 = n26065 ;
  assign y6423 = ~n26068 ;
  assign y6424 = n26075 ;
  assign y6425 = ~n26080 ;
  assign y6426 = ~n26090 ;
  assign y6427 = ~n26091 ;
  assign y6428 = n26094 ;
  assign y6429 = ~n26099 ;
  assign y6430 = ~n26107 ;
  assign y6431 = n26113 ;
  assign y6432 = ~n26120 ;
  assign y6433 = ~n26124 ;
  assign y6434 = ~n26126 ;
  assign y6435 = ~n26135 ;
  assign y6436 = ~n26140 ;
  assign y6437 = n26144 ;
  assign y6438 = n26147 ;
  assign y6439 = n26148 ;
  assign y6440 = ~n26153 ;
  assign y6441 = ~n26154 ;
  assign y6442 = ~1'b0 ;
  assign y6443 = ~n26157 ;
  assign y6444 = n26162 ;
  assign y6445 = n26164 ;
  assign y6446 = n26166 ;
  assign y6447 = n26170 ;
  assign y6448 = n26175 ;
  assign y6449 = ~n26181 ;
  assign y6450 = n26183 ;
  assign y6451 = ~n26202 ;
  assign y6452 = ~n26204 ;
  assign y6453 = n26208 ;
  assign y6454 = n26214 ;
  assign y6455 = ~n26215 ;
  assign y6456 = n26221 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = n26223 ;
  assign y6459 = ~n26224 ;
  assign y6460 = ~1'b0 ;
  assign y6461 = ~n26226 ;
  assign y6462 = ~n26227 ;
  assign y6463 = ~n26232 ;
  assign y6464 = ~1'b0 ;
  assign y6465 = ~n26235 ;
  assign y6466 = ~n26238 ;
  assign y6467 = n26239 ;
  assign y6468 = n26243 ;
  assign y6469 = ~1'b0 ;
  assign y6470 = ~n26247 ;
  assign y6471 = ~1'b0 ;
  assign y6472 = ~n26249 ;
  assign y6473 = ~n26250 ;
  assign y6474 = n26256 ;
  assign y6475 = ~n26257 ;
  assign y6476 = n26262 ;
  assign y6477 = n26263 ;
  assign y6478 = n26264 ;
  assign y6479 = n26265 ;
  assign y6480 = ~n26270 ;
  assign y6481 = ~n26271 ;
  assign y6482 = n26276 ;
  assign y6483 = ~n26277 ;
  assign y6484 = ~1'b0 ;
  assign y6485 = n26278 ;
  assign y6486 = ~n26280 ;
  assign y6487 = n26282 ;
  assign y6488 = n26289 ;
  assign y6489 = ~1'b0 ;
  assign y6490 = ~n26294 ;
  assign y6491 = n26295 ;
  assign y6492 = ~1'b0 ;
  assign y6493 = ~n26300 ;
  assign y6494 = n26302 ;
  assign y6495 = n26303 ;
  assign y6496 = ~n26305 ;
  assign y6497 = n26314 ;
  assign y6498 = n26315 ;
  assign y6499 = ~1'b0 ;
  assign y6500 = ~n26323 ;
  assign y6501 = n26324 ;
  assign y6502 = ~n26325 ;
  assign y6503 = n26326 ;
  assign y6504 = ~1'b0 ;
  assign y6505 = ~1'b0 ;
  assign y6506 = ~n26330 ;
  assign y6507 = n26334 ;
  assign y6508 = n26339 ;
  assign y6509 = n26340 ;
  assign y6510 = n26346 ;
  assign y6511 = ~1'b0 ;
  assign y6512 = n26354 ;
  assign y6513 = n26360 ;
  assign y6514 = ~n26368 ;
  assign y6515 = ~n26378 ;
  assign y6516 = ~n26382 ;
  assign y6517 = n26385 ;
  assign y6518 = n26386 ;
  assign y6519 = n26387 ;
  assign y6520 = ~n26390 ;
  assign y6521 = ~n26391 ;
  assign y6522 = n26392 ;
  assign y6523 = ~n26396 ;
  assign y6524 = ~1'b0 ;
  assign y6525 = ~n26397 ;
  assign y6526 = n26398 ;
  assign y6527 = n26400 ;
  assign y6528 = ~n26402 ;
  assign y6529 = ~1'b0 ;
  assign y6530 = n26405 ;
  assign y6531 = ~n26410 ;
  assign y6532 = ~1'b0 ;
  assign y6533 = n26414 ;
  assign y6534 = ~n26415 ;
  assign y6535 = n26418 ;
  assign y6536 = ~n26420 ;
  assign y6537 = ~n26423 ;
  assign y6538 = ~n26428 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = n26433 ;
  assign y6541 = n26435 ;
  assign y6542 = n26439 ;
  assign y6543 = ~n26440 ;
  assign y6544 = ~1'b0 ;
  assign y6545 = ~1'b0 ;
  assign y6546 = n26441 ;
  assign y6547 = ~n26445 ;
  assign y6548 = ~n26446 ;
  assign y6549 = n26448 ;
  assign y6550 = ~n26464 ;
  assign y6551 = ~n26466 ;
  assign y6552 = ~1'b0 ;
  assign y6553 = n26470 ;
  assign y6554 = ~n26476 ;
  assign y6555 = n26481 ;
  assign y6556 = ~n26483 ;
  assign y6557 = n2356 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = ~n26491 ;
  assign y6560 = n26493 ;
  assign y6561 = ~n26495 ;
  assign y6562 = n26496 ;
  assign y6563 = n26498 ;
  assign y6564 = ~n26500 ;
  assign y6565 = n26504 ;
  assign y6566 = n26507 ;
  assign y6567 = ~n26516 ;
  assign y6568 = n26521 ;
  assign y6569 = ~1'b0 ;
  assign y6570 = ~n26523 ;
  assign y6571 = n26526 ;
  assign y6572 = n26528 ;
  assign y6573 = n26533 ;
  assign y6574 = ~1'b0 ;
  assign y6575 = ~n26537 ;
  assign y6576 = ~n26538 ;
  assign y6577 = ~1'b0 ;
  assign y6578 = n26539 ;
  assign y6579 = ~n26541 ;
  assign y6580 = ~n26546 ;
  assign y6581 = n26552 ;
  assign y6582 = n26558 ;
  assign y6583 = ~n26563 ;
  assign y6584 = n26564 ;
  assign y6585 = n26569 ;
  assign y6586 = ~n26576 ;
  assign y6587 = ~n26577 ;
  assign y6588 = n26583 ;
  assign y6589 = ~n26584 ;
  assign y6590 = n26585 ;
  assign y6591 = ~n26588 ;
  assign y6592 = n26592 ;
  assign y6593 = n26598 ;
  assign y6594 = n26600 ;
  assign y6595 = ~n26603 ;
  assign y6596 = ~1'b0 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = ~1'b0 ;
  assign y6599 = ~n26604 ;
  assign y6600 = ~1'b0 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = ~n26608 ;
  assign y6604 = n26611 ;
  assign y6605 = ~n26615 ;
  assign y6606 = ~n26616 ;
  assign y6607 = n26618 ;
  assign y6608 = ~1'b0 ;
  assign y6609 = ~n26619 ;
  assign y6610 = ~n26623 ;
  assign y6611 = ~n26626 ;
  assign y6612 = n26630 ;
  assign y6613 = n26632 ;
  assign y6614 = ~n26634 ;
  assign y6615 = ~n26636 ;
  assign y6616 = ~n26648 ;
  assign y6617 = n26655 ;
  assign y6618 = ~n26657 ;
  assign y6619 = ~n26659 ;
  assign y6620 = ~n26664 ;
  assign y6621 = n26666 ;
  assign y6622 = n26667 ;
  assign y6623 = ~1'b0 ;
  assign y6624 = n26671 ;
  assign y6625 = ~n26674 ;
  assign y6626 = n26683 ;
  assign y6627 = ~n26685 ;
  assign y6628 = n24329 ;
  assign y6629 = ~n26686 ;
  assign y6630 = ~n26687 ;
  assign y6631 = ~n26689 ;
  assign y6632 = ~n26692 ;
  assign y6633 = ~n26699 ;
  assign y6634 = n26706 ;
  assign y6635 = n26707 ;
  assign y6636 = ~n26709 ;
  assign y6637 = ~n26712 ;
  assign y6638 = n26714 ;
  assign y6639 = n26715 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = n20902 ;
  assign y6642 = n26719 ;
  assign y6643 = ~n26722 ;
  assign y6644 = ~1'b0 ;
  assign y6645 = ~n26724 ;
  assign y6646 = ~n26725 ;
  assign y6647 = n26732 ;
  assign y6648 = ~n26736 ;
  assign y6649 = ~1'b0 ;
  assign y6650 = n26740 ;
  assign y6651 = ~1'b0 ;
  assign y6652 = ~n26746 ;
  assign y6653 = ~n26749 ;
  assign y6654 = n26754 ;
  assign y6655 = n26757 ;
  assign y6656 = ~n26760 ;
  assign y6657 = ~1'b0 ;
  assign y6658 = n26761 ;
  assign y6659 = n26762 ;
  assign y6660 = ~n26764 ;
  assign y6661 = ~n26768 ;
  assign y6662 = ~1'b0 ;
  assign y6663 = ~n26777 ;
  assign y6664 = n26780 ;
  assign y6665 = ~n26783 ;
  assign y6666 = n26785 ;
  assign y6667 = ~n26792 ;
  assign y6668 = ~n26795 ;
  assign y6669 = ~n26799 ;
  assign y6670 = n26802 ;
  assign y6671 = n26804 ;
  assign y6672 = ~n26806 ;
  assign y6673 = n26808 ;
  assign y6674 = ~n26809 ;
  assign y6675 = ~n26810 ;
  assign y6676 = ~n26811 ;
  assign y6677 = n26812 ;
  assign y6678 = ~n26813 ;
  assign y6679 = n26822 ;
  assign y6680 = ~n26830 ;
  assign y6681 = n26831 ;
  assign y6682 = ~n26833 ;
  assign y6683 = n26836 ;
  assign y6684 = n26837 ;
  assign y6685 = n26839 ;
  assign y6686 = ~n26840 ;
  assign y6687 = ~n26841 ;
  assign y6688 = ~n26843 ;
  assign y6689 = n26848 ;
  assign y6690 = ~n26850 ;
  assign y6691 = ~n26851 ;
  assign y6692 = n26854 ;
  assign y6693 = ~1'b0 ;
  assign y6694 = ~n26855 ;
  assign y6695 = n26858 ;
  assign y6696 = ~n26860 ;
  assign y6697 = ~1'b0 ;
  assign y6698 = ~n26862 ;
  assign y6699 = ~n26869 ;
  assign y6700 = n26871 ;
  assign y6701 = ~n26872 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = n26882 ;
  assign y6704 = n26885 ;
  assign y6705 = n26893 ;
  assign y6706 = ~n26899 ;
  assign y6707 = n26904 ;
  assign y6708 = n26906 ;
  assign y6709 = n26909 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~n26915 ;
  assign y6712 = ~n26916 ;
  assign y6713 = ~n26917 ;
  assign y6714 = n26918 ;
  assign y6715 = n26921 ;
  assign y6716 = ~n26929 ;
  assign y6717 = n26930 ;
  assign y6718 = n26932 ;
  assign y6719 = ~n26935 ;
  assign y6720 = n26939 ;
  assign y6721 = n26942 ;
  assign y6722 = ~n26943 ;
  assign y6723 = n26945 ;
  assign y6724 = ~n26948 ;
  assign y6725 = ~n26963 ;
  assign y6726 = n26966 ;
  assign y6727 = n26971 ;
  assign y6728 = ~1'b0 ;
  assign y6729 = ~n26972 ;
  assign y6730 = ~n26973 ;
  assign y6731 = n26975 ;
  assign y6732 = n26978 ;
  assign y6733 = ~1'b0 ;
  assign y6734 = ~n26981 ;
  assign y6735 = n26986 ;
  assign y6736 = n26991 ;
  assign y6737 = ~n26995 ;
  assign y6738 = ~n26997 ;
  assign y6739 = ~1'b0 ;
  assign y6740 = ~n27000 ;
  assign y6741 = n27001 ;
  assign y6742 = n27005 ;
  assign y6743 = n27007 ;
  assign y6744 = n27009 ;
  assign y6745 = ~1'b0 ;
  assign y6746 = n27011 ;
  assign y6747 = ~n27015 ;
  assign y6748 = n27016 ;
  assign y6749 = ~n16209 ;
  assign y6750 = ~n27018 ;
  assign y6751 = ~n27020 ;
  assign y6752 = ~n27022 ;
  assign y6753 = ~n27026 ;
  assign y6754 = n27029 ;
  assign y6755 = n27031 ;
  assign y6756 = ~n27032 ;
  assign y6757 = ~1'b0 ;
  assign y6758 = ~1'b0 ;
  assign y6759 = ~n27040 ;
  assign y6760 = n27050 ;
  assign y6761 = ~n27051 ;
  assign y6762 = ~n27053 ;
  assign y6763 = n27055 ;
  assign y6764 = ~1'b0 ;
  assign y6765 = n27062 ;
  assign y6766 = n27069 ;
  assign y6767 = n27075 ;
  assign y6768 = n27077 ;
  assign y6769 = ~n27078 ;
  assign y6770 = n27081 ;
  assign y6771 = n27082 ;
  assign y6772 = ~n27085 ;
  assign y6773 = ~n27087 ;
  assign y6774 = n27093 ;
  assign y6775 = ~1'b0 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~n27097 ;
  assign y6778 = n27101 ;
  assign y6779 = n27102 ;
  assign y6780 = n27105 ;
  assign y6781 = n27107 ;
  assign y6782 = ~n27109 ;
  assign y6783 = ~n27111 ;
  assign y6784 = n27116 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = ~n27123 ;
  assign y6787 = ~n27124 ;
  assign y6788 = ~n27126 ;
  assign y6789 = n27131 ;
  assign y6790 = n27133 ;
  assign y6791 = ~1'b0 ;
  assign y6792 = n27138 ;
  assign y6793 = n27144 ;
  assign y6794 = ~n27145 ;
  assign y6795 = ~n27148 ;
  assign y6796 = n27152 ;
  assign y6797 = n27154 ;
  assign y6798 = ~n27158 ;
  assign y6799 = ~1'b0 ;
  assign y6800 = n27162 ;
  assign y6801 = n27167 ;
  assign y6802 = ~n27177 ;
  assign y6803 = ~n27181 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = n27184 ;
  assign y6806 = n27185 ;
  assign y6807 = n27187 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = n27189 ;
  assign y6810 = n27190 ;
  assign y6811 = ~n27194 ;
  assign y6812 = ~n27201 ;
  assign y6813 = ~1'b0 ;
  assign y6814 = ~1'b0 ;
  assign y6815 = ~n27202 ;
  assign y6816 = ~n27210 ;
  assign y6817 = ~n27211 ;
  assign y6818 = ~n27213 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = n27217 ;
  assign y6821 = ~n27219 ;
  assign y6822 = ~n27222 ;
  assign y6823 = ~n27223 ;
  assign y6824 = n27224 ;
  assign y6825 = ~n27228 ;
  assign y6826 = n27230 ;
  assign y6827 = n27233 ;
  assign y6828 = n27236 ;
  assign y6829 = n27238 ;
  assign y6830 = n27240 ;
  assign y6831 = n27247 ;
  assign y6832 = ~n27249 ;
  assign y6833 = ~1'b0 ;
  assign y6834 = ~n27253 ;
  assign y6835 = ~n27258 ;
  assign y6836 = n27265 ;
  assign y6837 = n27270 ;
  assign y6838 = n27273 ;
  assign y6839 = ~n27281 ;
  assign y6840 = ~n27282 ;
  assign y6841 = n27287 ;
  assign y6842 = n27291 ;
  assign y6843 = ~1'b0 ;
  assign y6844 = ~n27295 ;
  assign y6845 = ~n27306 ;
  assign y6846 = ~n27307 ;
  assign y6847 = ~n27309 ;
  assign y6848 = ~n27311 ;
  assign y6849 = n27313 ;
  assign y6850 = n27315 ;
  assign y6851 = ~1'b0 ;
  assign y6852 = ~n27318 ;
  assign y6853 = n27319 ;
  assign y6854 = n27327 ;
  assign y6855 = ~n27329 ;
  assign y6856 = n27332 ;
  assign y6857 = ~n27336 ;
  assign y6858 = ~n27337 ;
  assign y6859 = ~n27340 ;
  assign y6860 = n27344 ;
  assign y6861 = n27346 ;
  assign y6862 = n27357 ;
  assign y6863 = ~n27359 ;
  assign y6864 = ~n27360 ;
  assign y6865 = n27368 ;
  assign y6866 = ~n27370 ;
  assign y6867 = n27372 ;
  assign y6868 = ~1'b0 ;
  assign y6869 = ~1'b0 ;
  assign y6870 = ~n27383 ;
  assign y6871 = ~n27384 ;
  assign y6872 = n27386 ;
  assign y6873 = n27387 ;
  assign y6874 = n27398 ;
  assign y6875 = ~n27403 ;
  assign y6876 = n27409 ;
  assign y6877 = ~n27410 ;
  assign y6878 = ~1'b0 ;
  assign y6879 = ~n27418 ;
  assign y6880 = ~n27420 ;
  assign y6881 = ~n27429 ;
  assign y6882 = ~n27433 ;
  assign y6883 = n27437 ;
  assign y6884 = ~1'b0 ;
  assign y6885 = n27441 ;
  assign y6886 = ~n27449 ;
  assign y6887 = ~n27452 ;
  assign y6888 = n27459 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = ~n27461 ;
  assign y6891 = ~n27463 ;
  assign y6892 = ~n27465 ;
  assign y6893 = n27467 ;
  assign y6894 = ~1'b0 ;
  assign y6895 = ~n27470 ;
  assign y6896 = ~1'b0 ;
  assign y6897 = ~n27472 ;
  assign y6898 = ~n27477 ;
  assign y6899 = ~n27479 ;
  assign y6900 = ~n27483 ;
  assign y6901 = ~n27488 ;
  assign y6902 = ~1'b0 ;
  assign y6903 = n27490 ;
  assign y6904 = ~n27492 ;
  assign y6905 = n27500 ;
  assign y6906 = n27502 ;
  assign y6907 = ~n27510 ;
  assign y6908 = ~n27514 ;
  assign y6909 = n27516 ;
  assign y6910 = ~n27524 ;
  assign y6911 = ~n27525 ;
  assign y6912 = n5628 ;
  assign y6913 = n27529 ;
  assign y6914 = ~n27530 ;
  assign y6915 = ~n27532 ;
  assign y6916 = n27534 ;
  assign y6917 = ~n27536 ;
  assign y6918 = n27537 ;
  assign y6919 = ~n27544 ;
  assign y6920 = n27549 ;
  assign y6921 = n27556 ;
  assign y6922 = ~1'b0 ;
  assign y6923 = ~n27562 ;
  assign y6924 = n27565 ;
  assign y6925 = ~n27569 ;
  assign y6926 = ~n27573 ;
  assign y6927 = n27579 ;
  assign y6928 = n27580 ;
  assign y6929 = n27589 ;
  assign y6930 = ~1'b0 ;
  assign y6931 = ~n27594 ;
  assign y6932 = ~n27596 ;
  assign y6933 = n27605 ;
  assign y6934 = ~n27609 ;
  assign y6935 = n27611 ;
  assign y6936 = ~1'b0 ;
  assign y6937 = ~n27613 ;
  assign y6938 = n27615 ;
  assign y6939 = ~n27616 ;
  assign y6940 = ~n27624 ;
  assign y6941 = ~n27628 ;
  assign y6942 = ~n27629 ;
  assign y6943 = ~n27639 ;
  assign y6944 = n27641 ;
  assign y6945 = n27642 ;
  assign y6946 = ~n27647 ;
  assign y6947 = ~n27648 ;
  assign y6948 = n27649 ;
  assign y6949 = ~n27657 ;
  assign y6950 = n27661 ;
  assign y6951 = ~n27665 ;
  assign y6952 = ~n27666 ;
  assign y6953 = ~1'b0 ;
  assign y6954 = n27668 ;
  assign y6955 = ~n27674 ;
  assign y6956 = n27675 ;
  assign y6957 = n27679 ;
  assign y6958 = ~n27681 ;
  assign y6959 = ~n27686 ;
  assign y6960 = n27693 ;
  assign y6961 = n27698 ;
  assign y6962 = n27701 ;
  assign y6963 = n27710 ;
  assign y6964 = n27712 ;
  assign y6965 = n27713 ;
  assign y6966 = n27717 ;
  assign y6967 = ~n27722 ;
  assign y6968 = n27727 ;
  assign y6969 = n27735 ;
  assign y6970 = ~n27738 ;
  assign y6971 = ~n27743 ;
  assign y6972 = ~n27744 ;
  assign y6973 = ~n27749 ;
  assign y6974 = n27754 ;
  assign y6975 = n27757 ;
  assign y6976 = n27760 ;
  assign y6977 = ~n27763 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = ~1'b0 ;
  assign y6980 = n27766 ;
  assign y6981 = ~n27773 ;
  assign y6982 = n27782 ;
  assign y6983 = n27784 ;
  assign y6984 = n27786 ;
  assign y6985 = n27796 ;
  assign y6986 = n27803 ;
  assign y6987 = ~1'b0 ;
  assign y6988 = n27804 ;
  assign y6989 = ~n27806 ;
  assign y6990 = n27808 ;
  assign y6991 = n27811 ;
  assign y6992 = n27815 ;
  assign y6993 = n27817 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = ~n27820 ;
  assign y6996 = ~n27821 ;
  assign y6997 = n27823 ;
  assign y6998 = 1'b0 ;
  assign y6999 = n27827 ;
  assign y7000 = ~n27829 ;
  assign y7001 = ~n27831 ;
  assign y7002 = ~n27837 ;
  assign y7003 = n27838 ;
  assign y7004 = ~1'b0 ;
  assign y7005 = n27843 ;
  assign y7006 = n27847 ;
  assign y7007 = n27850 ;
  assign y7008 = n27853 ;
  assign y7009 = ~1'b0 ;
  assign y7010 = n27854 ;
  assign y7011 = ~n27862 ;
  assign y7012 = ~n27863 ;
  assign y7013 = ~n24779 ;
  assign y7014 = ~1'b0 ;
  assign y7015 = n27868 ;
  assign y7016 = ~n27871 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = ~n27875 ;
  assign y7019 = n27880 ;
  assign y7020 = ~n27883 ;
  assign y7021 = n27891 ;
  assign y7022 = ~n27892 ;
  assign y7023 = n27895 ;
  assign y7024 = n27897 ;
  assign y7025 = ~n27899 ;
  assign y7026 = ~n27902 ;
  assign y7027 = ~n27903 ;
  assign y7028 = n27904 ;
  assign y7029 = ~n27907 ;
  assign y7030 = ~n27910 ;
  assign y7031 = ~n27912 ;
  assign y7032 = n27919 ;
  assign y7033 = ~n27930 ;
  assign y7034 = ~n27939 ;
  assign y7035 = ~n27943 ;
  assign y7036 = n27948 ;
  assign y7037 = ~n27952 ;
  assign y7038 = n27957 ;
  assign y7039 = n27961 ;
  assign y7040 = ~1'b0 ;
  assign y7041 = ~n27967 ;
  assign y7042 = ~n27969 ;
  assign y7043 = n27972 ;
  assign y7044 = n27975 ;
  assign y7045 = n27977 ;
  assign y7046 = n27982 ;
  assign y7047 = ~1'b0 ;
  assign y7048 = ~n27986 ;
  assign y7049 = n27991 ;
  assign y7050 = n27994 ;
  assign y7051 = n27999 ;
  assign y7052 = n28000 ;
  assign y7053 = n28002 ;
  assign y7054 = ~n28004 ;
  assign y7055 = n28007 ;
  assign y7056 = n28010 ;
  assign y7057 = ~n28019 ;
  assign y7058 = n28023 ;
  assign y7059 = ~n28027 ;
  assign y7060 = ~n28033 ;
  assign y7061 = ~n28045 ;
  assign y7062 = ~n28047 ;
  assign y7063 = n28057 ;
  assign y7064 = n28059 ;
  assign y7065 = ~n28060 ;
  assign y7066 = ~n28064 ;
  assign y7067 = ~n28068 ;
  assign y7068 = ~n28070 ;
  assign y7069 = ~1'b0 ;
  assign y7070 = n28072 ;
  assign y7071 = ~n28084 ;
  assign y7072 = n28085 ;
  assign y7073 = n28086 ;
  assign y7074 = ~n28089 ;
  assign y7075 = ~n28092 ;
  assign y7076 = ~1'b0 ;
  assign y7077 = ~n28096 ;
  assign y7078 = ~n28100 ;
  assign y7079 = ~n28101 ;
  assign y7080 = ~n28103 ;
  assign y7081 = ~n28107 ;
  assign y7082 = ~1'b0 ;
  assign y7083 = ~n28110 ;
  assign y7084 = n28111 ;
  assign y7085 = ~n28114 ;
  assign y7086 = n28116 ;
  assign y7087 = ~n28117 ;
  assign y7088 = n28118 ;
  assign y7089 = ~n28122 ;
  assign y7090 = n28123 ;
  assign y7091 = ~n28125 ;
  assign y7092 = ~n28130 ;
  assign y7093 = n28134 ;
  assign y7094 = n28142 ;
  assign y7095 = ~n28144 ;
  assign y7096 = ~1'b0 ;
  assign y7097 = n28146 ;
  assign y7098 = ~n28147 ;
  assign y7099 = ~n28158 ;
  assign y7100 = ~n28159 ;
  assign y7101 = ~1'b0 ;
  assign y7102 = ~n28167 ;
  assign y7103 = n28171 ;
  assign y7104 = ~n28172 ;
  assign y7105 = ~n28174 ;
  assign y7106 = ~n28178 ;
  assign y7107 = ~1'b0 ;
  assign y7108 = ~n28179 ;
  assign y7109 = ~n28182 ;
  assign y7110 = ~n28183 ;
  assign y7111 = ~1'b0 ;
  assign y7112 = ~n28185 ;
  assign y7113 = ~1'b0 ;
  assign y7114 = ~n28188 ;
  assign y7115 = n28190 ;
  assign y7116 = ~n28196 ;
  assign y7117 = ~n28201 ;
  assign y7118 = ~n28209 ;
  assign y7119 = ~n28215 ;
  assign y7120 = n28216 ;
  assign y7121 = ~n28217 ;
  assign y7122 = ~n28220 ;
  assign y7123 = ~n28222 ;
  assign y7124 = n28223 ;
  assign y7125 = ~n28224 ;
  assign y7126 = ~n28228 ;
  assign y7127 = ~1'b0 ;
  assign y7128 = ~1'b0 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = ~n28229 ;
  assign y7131 = ~n28232 ;
  assign y7132 = n28233 ;
  assign y7133 = ~n28236 ;
  assign y7134 = n28241 ;
  assign y7135 = ~n28254 ;
  assign y7136 = n28258 ;
  assign y7137 = n28270 ;
  assign y7138 = ~n28271 ;
  assign y7139 = n28272 ;
  assign y7140 = ~n28273 ;
  assign y7141 = n28276 ;
  assign y7142 = ~n28283 ;
  assign y7143 = ~1'b0 ;
  assign y7144 = n28286 ;
  assign y7145 = ~n28288 ;
  assign y7146 = n28296 ;
  assign y7147 = ~n28301 ;
  assign y7148 = ~n28306 ;
  assign y7149 = ~1'b0 ;
  assign y7150 = ~n28312 ;
  assign y7151 = ~n28313 ;
  assign y7152 = n28321 ;
  assign y7153 = ~n28323 ;
  assign y7154 = ~n28329 ;
  assign y7155 = ~n28337 ;
  assign y7156 = ~1'b0 ;
  assign y7157 = n28344 ;
  assign y7158 = n28345 ;
  assign y7159 = ~n28347 ;
  assign y7160 = ~n28349 ;
  assign y7161 = ~n28350 ;
  assign y7162 = ~1'b0 ;
  assign y7163 = ~n28353 ;
  assign y7164 = n28358 ;
  assign y7165 = ~n28361 ;
  assign y7166 = n28363 ;
  assign y7167 = ~1'b0 ;
  assign y7168 = n28364 ;
  assign y7169 = n28369 ;
  assign y7170 = ~n28370 ;
  assign y7171 = n28378 ;
  assign y7172 = ~n28381 ;
  assign y7173 = ~n28385 ;
  assign y7174 = n28388 ;
  assign y7175 = n28389 ;
  assign y7176 = n28390 ;
  assign y7177 = n28391 ;
  assign y7178 = ~1'b0 ;
  assign y7179 = ~n28392 ;
  assign y7180 = n28393 ;
  assign y7181 = ~n28396 ;
  assign y7182 = ~n28400 ;
  assign y7183 = n28403 ;
  assign y7184 = n28404 ;
  assign y7185 = n28409 ;
  assign y7186 = ~n28414 ;
  assign y7187 = n28423 ;
  assign y7188 = n28428 ;
  assign y7189 = ~n28430 ;
  assign y7190 = ~n28431 ;
  assign y7191 = n28434 ;
  assign y7192 = n28435 ;
  assign y7193 = ~n28441 ;
  assign y7194 = ~n28451 ;
  assign y7195 = n28459 ;
  assign y7196 = ~n28460 ;
  assign y7197 = ~n28461 ;
  assign y7198 = ~1'b0 ;
  assign y7199 = ~n28464 ;
  assign y7200 = ~1'b0 ;
  assign y7201 = ~n28466 ;
  assign y7202 = ~n28467 ;
  assign y7203 = ~n28468 ;
  assign y7204 = n28469 ;
  assign y7205 = n28476 ;
  assign y7206 = n28479 ;
  assign y7207 = n28480 ;
  assign y7208 = n28484 ;
  assign y7209 = ~n28488 ;
  assign y7210 = n28490 ;
  assign y7211 = ~n28491 ;
  assign y7212 = ~n28493 ;
  assign y7213 = n28495 ;
  assign y7214 = n28496 ;
  assign y7215 = n28499 ;
  assign y7216 = n28502 ;
  assign y7217 = n28506 ;
  assign y7218 = n28509 ;
  assign y7219 = ~n28512 ;
  assign y7220 = n28515 ;
  assign y7221 = ~1'b0 ;
  assign y7222 = n28526 ;
  assign y7223 = ~n28528 ;
  assign y7224 = ~n28532 ;
  assign y7225 = n28533 ;
  assign y7226 = ~n28541 ;
  assign y7227 = n28542 ;
  assign y7228 = n28545 ;
  assign y7229 = ~n28551 ;
  assign y7230 = n28553 ;
  assign y7231 = ~n28557 ;
  assign y7232 = ~n28563 ;
  assign y7233 = ~n28570 ;
  assign y7234 = n28578 ;
  assign y7235 = ~n28582 ;
  assign y7236 = ~n28583 ;
  assign y7237 = n28589 ;
  assign y7238 = n16683 ;
  assign y7239 = ~n28595 ;
  assign y7240 = ~n28596 ;
  assign y7241 = n28597 ;
  assign y7242 = n28601 ;
  assign y7243 = n28605 ;
  assign y7244 = ~n28607 ;
  assign y7245 = n28609 ;
  assign y7246 = ~1'b0 ;
  assign y7247 = ~n28610 ;
  assign y7248 = ~n28611 ;
  assign y7249 = n28612 ;
  assign y7250 = ~n28613 ;
  assign y7251 = ~n28616 ;
  assign y7252 = n28619 ;
  assign y7253 = n28622 ;
  assign y7254 = ~n28624 ;
  assign y7255 = ~n28631 ;
  assign y7256 = ~n28633 ;
  assign y7257 = ~1'b0 ;
  assign y7258 = n28641 ;
  assign y7259 = ~n28644 ;
  assign y7260 = 1'b0 ;
  assign y7261 = ~n28646 ;
  assign y7262 = ~n28648 ;
  assign y7263 = ~n28655 ;
  assign y7264 = ~n28657 ;
  assign y7265 = n28659 ;
  assign y7266 = n28663 ;
  assign y7267 = ~1'b0 ;
  assign y7268 = ~n28668 ;
  assign y7269 = n28676 ;
  assign y7270 = ~n28679 ;
  assign y7271 = ~n28681 ;
  assign y7272 = ~n28682 ;
  assign y7273 = n28686 ;
  assign y7274 = ~n28697 ;
  assign y7275 = n12238 ;
  assign y7276 = ~1'b0 ;
  assign y7277 = ~1'b0 ;
  assign y7278 = n28701 ;
  assign y7279 = ~n28702 ;
  assign y7280 = ~n28705 ;
  assign y7281 = n28708 ;
  assign y7282 = n28717 ;
  assign y7283 = ~n28726 ;
  assign y7284 = ~1'b0 ;
  assign y7285 = n28730 ;
  assign y7286 = n28731 ;
  assign y7287 = n28732 ;
  assign y7288 = ~1'b0 ;
  assign y7289 = ~n28735 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~n28737 ;
  assign y7292 = ~n28739 ;
  assign y7293 = ~n28740 ;
  assign y7294 = n28741 ;
  assign y7295 = n28742 ;
  assign y7296 = n28746 ;
  assign y7297 = ~1'b0 ;
  assign y7298 = n28747 ;
  assign y7299 = n28748 ;
  assign y7300 = ~n28751 ;
  assign y7301 = ~n28757 ;
  assign y7302 = n28758 ;
  assign y7303 = ~n28759 ;
  assign y7304 = ~1'b0 ;
  assign y7305 = n28761 ;
  assign y7306 = ~n28762 ;
  assign y7307 = ~n28766 ;
  assign y7308 = ~n28767 ;
  assign y7309 = n28768 ;
  assign y7310 = ~n28769 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = ~1'b0 ;
  assign y7313 = ~n28773 ;
  assign y7314 = ~n28775 ;
  assign y7315 = ~n28778 ;
  assign y7316 = ~n28780 ;
  assign y7317 = ~n28782 ;
  assign y7318 = n28784 ;
  assign y7319 = n28788 ;
  assign y7320 = ~n28796 ;
  assign y7321 = n28803 ;
  assign y7322 = ~n28804 ;
  assign y7323 = ~n28809 ;
  assign y7324 = ~n28811 ;
  assign y7325 = ~n28818 ;
  assign y7326 = ~n28819 ;
  assign y7327 = n28822 ;
  assign y7328 = ~n28824 ;
  assign y7329 = ~n28826 ;
  assign y7330 = n28827 ;
  assign y7331 = ~1'b0 ;
  assign y7332 = n28829 ;
  assign y7333 = ~n28832 ;
  assign y7334 = n28841 ;
  assign y7335 = ~n28843 ;
  assign y7336 = ~n28845 ;
  assign y7337 = ~1'b0 ;
  assign y7338 = n28852 ;
  assign y7339 = ~1'b0 ;
  assign y7340 = n28853 ;
  assign y7341 = ~n28866 ;
  assign y7342 = ~1'b0 ;
  assign y7343 = ~n28867 ;
  assign y7344 = n28868 ;
  assign y7345 = n28869 ;
  assign y7346 = n28872 ;
  assign y7347 = n28876 ;
  assign y7348 = ~n28877 ;
  assign y7349 = ~n28885 ;
  assign y7350 = n28891 ;
  assign y7351 = ~n28894 ;
  assign y7352 = ~n28896 ;
  assign y7353 = ~n28898 ;
  assign y7354 = ~n28907 ;
  assign y7355 = ~n28920 ;
  assign y7356 = n28922 ;
  assign y7357 = ~n28927 ;
  assign y7358 = n28928 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = ~n28930 ;
  assign y7361 = ~n28932 ;
  assign y7362 = n21634 ;
  assign y7363 = ~n28934 ;
  assign y7364 = ~n28937 ;
  assign y7365 = ~n28940 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = n28944 ;
  assign y7368 = ~n28946 ;
  assign y7369 = ~n28949 ;
  assign y7370 = n28950 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = n28952 ;
  assign y7373 = ~n28956 ;
  assign y7374 = ~1'b0 ;
  assign y7375 = n28961 ;
  assign y7376 = ~n28964 ;
  assign y7377 = ~n28970 ;
  assign y7378 = ~n28977 ;
  assign y7379 = n28981 ;
  assign y7380 = n28982 ;
  assign y7381 = n28984 ;
  assign y7382 = ~n28986 ;
  assign y7383 = ~n28989 ;
  assign y7384 = n28990 ;
  assign y7385 = ~n28991 ;
  assign y7386 = n28993 ;
  assign y7387 = n28998 ;
  assign y7388 = n29009 ;
  assign y7389 = ~n29010 ;
  assign y7390 = ~n29013 ;
  assign y7391 = ~n29014 ;
  assign y7392 = n29015 ;
  assign y7393 = n29017 ;
  assign y7394 = ~n29018 ;
  assign y7395 = ~n29023 ;
  assign y7396 = ~n29025 ;
  assign y7397 = ~n29026 ;
  assign y7398 = ~n29034 ;
  assign y7399 = n29036 ;
  assign y7400 = ~1'b0 ;
  assign y7401 = n29039 ;
  assign y7402 = ~n29044 ;
  assign y7403 = ~n29045 ;
  assign y7404 = n29047 ;
  assign y7405 = ~n29051 ;
  assign y7406 = ~n29055 ;
  assign y7407 = n29056 ;
  assign y7408 = ~n29064 ;
  assign y7409 = n29066 ;
  assign y7410 = ~n29071 ;
  assign y7411 = n29073 ;
  assign y7412 = ~n29074 ;
  assign y7413 = ~n29075 ;
  assign y7414 = ~n29081 ;
  assign y7415 = ~n29083 ;
  assign y7416 = ~n29089 ;
  assign y7417 = n29090 ;
  assign y7418 = n29093 ;
  assign y7419 = ~n29098 ;
  assign y7420 = n29100 ;
  assign y7421 = ~1'b0 ;
  assign y7422 = ~n29102 ;
  assign y7423 = n29108 ;
  assign y7424 = n29110 ;
  assign y7425 = n29113 ;
  assign y7426 = ~n29114 ;
  assign y7427 = ~n29119 ;
  assign y7428 = n29129 ;
  assign y7429 = n29134 ;
  assign y7430 = ~n29146 ;
  assign y7431 = n29147 ;
  assign y7432 = n29149 ;
  assign y7433 = ~n29153 ;
  assign y7434 = ~n29156 ;
  assign y7435 = ~1'b0 ;
  assign y7436 = n29158 ;
  assign y7437 = ~n29164 ;
  assign y7438 = ~n29166 ;
  assign y7439 = ~n29167 ;
  assign y7440 = ~n29172 ;
  assign y7441 = ~n29173 ;
  assign y7442 = n29177 ;
  assign y7443 = ~n29180 ;
  assign y7444 = ~n29181 ;
  assign y7445 = ~n29190 ;
  assign y7446 = ~n29194 ;
  assign y7447 = ~n29197 ;
  assign y7448 = ~n29198 ;
  assign y7449 = ~n29207 ;
  assign y7450 = ~1'b0 ;
  assign y7451 = n29213 ;
  assign y7452 = n29216 ;
  assign y7453 = ~n29218 ;
  assign y7454 = n29220 ;
  assign y7455 = ~1'b0 ;
  assign y7456 = ~n29223 ;
  assign y7457 = ~n29231 ;
  assign y7458 = ~1'b0 ;
  assign y7459 = n29232 ;
  assign y7460 = n17227 ;
  assign y7461 = ~n29233 ;
  assign y7462 = ~n29236 ;
  assign y7463 = n29238 ;
  assign y7464 = ~n29243 ;
  assign y7465 = n29244 ;
  assign y7466 = ~n29263 ;
  assign y7467 = n29267 ;
  assign y7468 = ~n29277 ;
  assign y7469 = n29282 ;
  assign y7470 = n29284 ;
  assign y7471 = n29286 ;
  assign y7472 = ~n29287 ;
  assign y7473 = ~n29290 ;
  assign y7474 = ~1'b0 ;
  assign y7475 = ~n29292 ;
  assign y7476 = n29296 ;
  assign y7477 = n29308 ;
  assign y7478 = n29309 ;
  assign y7479 = ~1'b0 ;
  assign y7480 = ~n29313 ;
  assign y7481 = ~n29318 ;
  assign y7482 = ~n29324 ;
  assign y7483 = n29328 ;
  assign y7484 = n29331 ;
  assign y7485 = n29334 ;
  assign y7486 = ~n29337 ;
  assign y7487 = n29338 ;
  assign y7488 = ~n29339 ;
  assign y7489 = n29346 ;
  assign y7490 = n29351 ;
  assign y7491 = n29353 ;
  assign y7492 = n29361 ;
  assign y7493 = n29363 ;
  assign y7494 = ~n29367 ;
  assign y7495 = n29370 ;
  assign y7496 = n29391 ;
  assign y7497 = ~n29392 ;
  assign y7498 = ~n16976 ;
  assign y7499 = ~n29399 ;
  assign y7500 = ~n29402 ;
  assign y7501 = n29404 ;
  assign y7502 = ~n29410 ;
  assign y7503 = ~n29414 ;
  assign y7504 = n29415 ;
  assign y7505 = ~n29419 ;
  assign y7506 = ~n29420 ;
  assign y7507 = n29423 ;
  assign y7508 = n29432 ;
  assign y7509 = ~n29441 ;
  assign y7510 = ~n29442 ;
  assign y7511 = n29445 ;
  assign y7512 = n29448 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = n29453 ;
  assign y7515 = n29454 ;
  assign y7516 = ~n10589 ;
  assign y7517 = ~1'b0 ;
  assign y7518 = ~n29458 ;
  assign y7519 = ~n29461 ;
  assign y7520 = n29462 ;
  assign y7521 = ~n29463 ;
  assign y7522 = n29465 ;
  assign y7523 = ~1'b0 ;
  assign y7524 = n29467 ;
  assign y7525 = ~1'b0 ;
  assign y7526 = ~n29469 ;
  assign y7527 = n29471 ;
  assign y7528 = ~n29475 ;
  assign y7529 = n29477 ;
  assign y7530 = n29484 ;
  assign y7531 = ~n29485 ;
  assign y7532 = n29488 ;
  assign y7533 = ~n29489 ;
  assign y7534 = n29495 ;
  assign y7535 = ~n29501 ;
  assign y7536 = ~n29507 ;
  assign y7537 = ~n29514 ;
  assign y7538 = 1'b0 ;
  assign y7539 = n29515 ;
  assign y7540 = n834 ;
  assign y7541 = n29516 ;
  assign y7542 = ~n29520 ;
  assign y7543 = n29521 ;
  assign y7544 = n29522 ;
  assign y7545 = ~n29524 ;
  assign y7546 = n29527 ;
  assign y7547 = n29532 ;
  assign y7548 = ~n29534 ;
  assign y7549 = n29543 ;
  assign y7550 = n29545 ;
  assign y7551 = n29549 ;
  assign y7552 = n29551 ;
  assign y7553 = ~n29555 ;
  assign y7554 = n29557 ;
  assign y7555 = n29558 ;
  assign y7556 = n29562 ;
  assign y7557 = n29566 ;
  assign y7558 = ~n29568 ;
  assign y7559 = ~n29570 ;
  assign y7560 = ~n29577 ;
  assign y7561 = ~n29579 ;
  assign y7562 = n29589 ;
  assign y7563 = n29590 ;
  assign y7564 = ~n29592 ;
  assign y7565 = ~n29599 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = n29600 ;
  assign y7568 = ~n29603 ;
  assign y7569 = ~n29609 ;
  assign y7570 = ~n29610 ;
  assign y7571 = n29611 ;
  assign y7572 = ~n29620 ;
  assign y7573 = n29622 ;
  assign y7574 = ~n27451 ;
  assign y7575 = ~n29626 ;
  assign y7576 = ~1'b0 ;
  assign y7577 = n29641 ;
  assign y7578 = ~n29642 ;
  assign y7579 = ~n29647 ;
  assign y7580 = ~n29648 ;
  assign y7581 = ~n29650 ;
  assign y7582 = ~n29652 ;
  assign y7583 = n29654 ;
  assign y7584 = n29655 ;
  assign y7585 = n29657 ;
  assign y7586 = n29660 ;
  assign y7587 = n29665 ;
  assign y7588 = n29666 ;
  assign y7589 = ~n29670 ;
  assign y7590 = ~n29671 ;
  assign y7591 = ~n29673 ;
  assign y7592 = ~n29675 ;
  assign y7593 = n29678 ;
  assign y7594 = n29689 ;
  assign y7595 = ~1'b0 ;
  assign y7596 = ~n29693 ;
  assign y7597 = n29700 ;
  assign y7598 = ~n29702 ;
  assign y7599 = ~n29715 ;
  assign y7600 = n29717 ;
  assign y7601 = n29720 ;
  assign y7602 = ~n29724 ;
  assign y7603 = n29725 ;
  assign y7604 = ~n29726 ;
  assign y7605 = 1'b0 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = ~1'b0 ;
  assign y7608 = ~n29728 ;
  assign y7609 = ~n29729 ;
  assign y7610 = ~n29732 ;
  assign y7611 = n29735 ;
  assign y7612 = ~n29738 ;
  assign y7613 = ~1'b0 ;
  assign y7614 = ~n29739 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = ~n29742 ;
  assign y7617 = ~n29743 ;
  assign y7618 = n29745 ;
  assign y7619 = ~n29749 ;
  assign y7620 = ~n29754 ;
  assign y7621 = n29755 ;
  assign y7622 = ~n29758 ;
  assign y7623 = n29762 ;
  assign y7624 = n29764 ;
  assign y7625 = ~n29765 ;
  assign y7626 = ~n29766 ;
  assign y7627 = n29767 ;
  assign y7628 = n29780 ;
  assign y7629 = ~n29781 ;
  assign y7630 = n29784 ;
  assign y7631 = n29788 ;
  assign y7632 = ~n29798 ;
  assign y7633 = n29799 ;
  assign y7634 = n29804 ;
  assign y7635 = ~n29808 ;
  assign y7636 = ~n29812 ;
  assign y7637 = ~n29813 ;
  assign y7638 = ~1'b0 ;
  assign y7639 = ~n29816 ;
  assign y7640 = n29818 ;
  assign y7641 = n29819 ;
  assign y7642 = ~n29820 ;
  assign y7643 = ~n29823 ;
  assign y7644 = n29828 ;
  assign y7645 = n29832 ;
  assign y7646 = ~1'b0 ;
  assign y7647 = n29833 ;
  assign y7648 = ~n29834 ;
  assign y7649 = n29837 ;
  assign y7650 = n29838 ;
  assign y7651 = n29840 ;
  assign y7652 = n29841 ;
  assign y7653 = ~1'b0 ;
  assign y7654 = n29843 ;
  assign y7655 = ~n29844 ;
  assign y7656 = ~n29845 ;
  assign y7657 = ~n29850 ;
  assign y7658 = ~n29853 ;
  assign y7659 = n29862 ;
  assign y7660 = ~n29870 ;
  assign y7661 = n29874 ;
  assign y7662 = ~n29877 ;
  assign y7663 = ~n29879 ;
  assign y7664 = n29883 ;
  assign y7665 = ~n29884 ;
  assign y7666 = ~n29887 ;
  assign y7667 = n29892 ;
  assign y7668 = ~1'b0 ;
  assign y7669 = ~n29895 ;
  assign y7670 = ~n29896 ;
  assign y7671 = n29906 ;
  assign y7672 = ~1'b0 ;
  assign y7673 = n29909 ;
  assign y7674 = n29912 ;
  assign y7675 = ~n29913 ;
  assign y7676 = ~n29915 ;
  assign y7677 = n29922 ;
  assign y7678 = ~n29923 ;
  assign y7679 = ~1'b0 ;
  assign y7680 = ~n29926 ;
  assign y7681 = n29928 ;
  assign y7682 = ~n29929 ;
  assign y7683 = n29932 ;
  assign y7684 = n29941 ;
  assign y7685 = ~n29943 ;
  assign y7686 = n29944 ;
  assign y7687 = ~n29945 ;
  assign y7688 = n29947 ;
  assign y7689 = ~n29949 ;
  assign y7690 = ~n29952 ;
  assign y7691 = ~n29953 ;
  assign y7692 = ~n29956 ;
  assign y7693 = ~n29963 ;
  assign y7694 = n29971 ;
  assign y7695 = n29976 ;
  assign y7696 = ~n29977 ;
  assign y7697 = n29978 ;
  assign y7698 = ~n29979 ;
  assign y7699 = ~n29986 ;
  assign y7700 = ~n29997 ;
  assign y7701 = ~n30000 ;
  assign y7702 = ~1'b0 ;
  assign y7703 = ~n30001 ;
  assign y7704 = ~n30005 ;
  assign y7705 = ~1'b0 ;
  assign y7706 = ~n30013 ;
  assign y7707 = ~1'b0 ;
  assign y7708 = ~1'b0 ;
  assign y7709 = ~n30014 ;
  assign y7710 = ~n30016 ;
  assign y7711 = ~n30028 ;
  assign y7712 = ~n30029 ;
  assign y7713 = ~n30030 ;
  assign y7714 = n30038 ;
  assign y7715 = ~n30041 ;
  assign y7716 = ~n30046 ;
  assign y7717 = ~1'b0 ;
  assign y7718 = ~n30047 ;
  assign y7719 = n30060 ;
  assign y7720 = n30063 ;
  assign y7721 = n30066 ;
  assign y7722 = ~n30068 ;
  assign y7723 = n30072 ;
  assign y7724 = ~n30078 ;
  assign y7725 = n30079 ;
  assign y7726 = n30084 ;
  assign y7727 = n30087 ;
  assign y7728 = ~n30088 ;
  assign y7729 = n30091 ;
  assign y7730 = ~n30092 ;
  assign y7731 = n30093 ;
  assign y7732 = ~n30094 ;
  assign y7733 = ~n30098 ;
  assign y7734 = n30100 ;
  assign y7735 = n30102 ;
  assign y7736 = n30105 ;
  assign y7737 = n30108 ;
  assign y7738 = ~1'b0 ;
  assign y7739 = n30109 ;
  assign y7740 = ~n30110 ;
  assign y7741 = ~1'b0 ;
  assign y7742 = ~n30111 ;
  assign y7743 = ~n30118 ;
  assign y7744 = ~n30119 ;
  assign y7745 = ~n30126 ;
  assign y7746 = n30129 ;
  assign y7747 = n30132 ;
  assign y7748 = ~n30135 ;
  assign y7749 = n30138 ;
  assign y7750 = ~n30140 ;
  assign y7751 = ~n30145 ;
  assign y7752 = n30146 ;
  assign y7753 = ~n30150 ;
  assign y7754 = ~n30151 ;
  assign y7755 = n30161 ;
  assign y7756 = ~n30162 ;
  assign y7757 = n30164 ;
  assign y7758 = n30169 ;
  assign y7759 = ~n30175 ;
  assign y7760 = ~n30181 ;
  assign y7761 = n30184 ;
  assign y7762 = n30188 ;
  assign y7763 = n30191 ;
  assign y7764 = ~n30194 ;
  assign y7765 = ~n30196 ;
  assign y7766 = ~n30197 ;
  assign y7767 = ~n30202 ;
  assign y7768 = ~n30205 ;
  assign y7769 = n30207 ;
  assign y7770 = ~n30209 ;
  assign y7771 = n30211 ;
  assign y7772 = n30214 ;
  assign y7773 = ~1'b0 ;
  assign y7774 = n30221 ;
  assign y7775 = n30222 ;
  assign y7776 = n30224 ;
  assign y7777 = ~1'b0 ;
  assign y7778 = n30226 ;
  assign y7779 = n30230 ;
  assign y7780 = n30232 ;
  assign y7781 = n30235 ;
  assign y7782 = ~1'b0 ;
  assign y7783 = ~n30240 ;
  assign y7784 = n30241 ;
  assign y7785 = ~n30244 ;
  assign y7786 = n30245 ;
  assign y7787 = ~n30252 ;
  assign y7788 = ~n30253 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = n30255 ;
  assign y7791 = ~n30256 ;
  assign y7792 = ~n30258 ;
  assign y7793 = n30262 ;
  assign y7794 = n30266 ;
  assign y7795 = ~n30269 ;
  assign y7796 = ~n30270 ;
  assign y7797 = ~n30271 ;
  assign y7798 = ~n30272 ;
  assign y7799 = ~n30278 ;
  assign y7800 = ~1'b0 ;
  assign y7801 = ~1'b0 ;
  assign y7802 = ~n30279 ;
  assign y7803 = n30282 ;
  assign y7804 = n30286 ;
  assign y7805 = ~n30289 ;
  assign y7806 = ~n30291 ;
  assign y7807 = ~1'b0 ;
  assign y7808 = n30293 ;
  assign y7809 = ~n30295 ;
  assign y7810 = ~n30301 ;
  assign y7811 = ~n30304 ;
  assign y7812 = n30308 ;
  assign y7813 = ~n30313 ;
  assign y7814 = ~n30315 ;
  assign y7815 = ~n30321 ;
  assign y7816 = ~n30324 ;
  assign y7817 = ~1'b0 ;
  assign y7818 = ~1'b0 ;
  assign y7819 = n30325 ;
  assign y7820 = n30331 ;
  assign y7821 = n30333 ;
  assign y7822 = ~n30334 ;
  assign y7823 = n30336 ;
  assign y7824 = ~1'b0 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = n30338 ;
  assign y7827 = n30339 ;
  assign y7828 = n30342 ;
  assign y7829 = ~n30349 ;
  assign y7830 = ~n30357 ;
  assign y7831 = ~n30362 ;
  assign y7832 = n30363 ;
  assign y7833 = ~n30364 ;
  assign y7834 = n30368 ;
  assign y7835 = n30373 ;
  assign y7836 = n30382 ;
  assign y7837 = ~n30395 ;
  assign y7838 = ~n30397 ;
  assign y7839 = ~n30399 ;
  assign y7840 = ~n30400 ;
  assign y7841 = n12090 ;
  assign y7842 = n30412 ;
  assign y7843 = ~n30416 ;
  assign y7844 = ~n30422 ;
  assign y7845 = n30427 ;
  assign y7846 = ~n30429 ;
  assign y7847 = ~n19599 ;
  assign y7848 = ~n30432 ;
  assign y7849 = ~1'b0 ;
  assign y7850 = ~1'b0 ;
  assign y7851 = ~n30433 ;
  assign y7852 = ~n30434 ;
  assign y7853 = n30439 ;
  assign y7854 = ~n30441 ;
  assign y7855 = ~n30442 ;
  assign y7856 = n30443 ;
  assign y7857 = n30448 ;
  assign y7858 = n30452 ;
  assign y7859 = ~n30453 ;
  assign y7860 = n30455 ;
  assign y7861 = ~n30458 ;
  assign y7862 = ~n30462 ;
  assign y7863 = ~n30466 ;
  assign y7864 = ~n30472 ;
  assign y7865 = n30474 ;
  assign y7866 = ~n30482 ;
  assign y7867 = ~n30484 ;
  assign y7868 = ~n30487 ;
  assign y7869 = ~n30489 ;
  assign y7870 = ~n30498 ;
  assign y7871 = ~n30506 ;
  assign y7872 = ~n30514 ;
  assign y7873 = n30517 ;
  assign y7874 = ~n30519 ;
  assign y7875 = ~n30523 ;
  assign y7876 = n30524 ;
  assign y7877 = ~n30536 ;
  assign y7878 = ~1'b0 ;
  assign y7879 = n30539 ;
  assign y7880 = ~n30540 ;
  assign y7881 = n30543 ;
  assign y7882 = ~n30544 ;
  assign y7883 = ~n30545 ;
  assign y7884 = ~n30549 ;
  assign y7885 = n30554 ;
  assign y7886 = ~n30555 ;
  assign y7887 = ~n30560 ;
  assign y7888 = n30562 ;
  assign y7889 = ~1'b0 ;
  assign y7890 = n30566 ;
  assign y7891 = n30567 ;
  assign y7892 = n30575 ;
  assign y7893 = n30580 ;
  assign y7894 = ~1'b0 ;
  assign y7895 = n30582 ;
  assign y7896 = n30583 ;
  assign y7897 = ~n30584 ;
  assign y7898 = ~n30588 ;
  assign y7899 = ~n30592 ;
  assign y7900 = n30593 ;
  assign y7901 = ~n30595 ;
  assign y7902 = ~n30599 ;
  assign y7903 = ~1'b0 ;
  assign y7904 = ~n30605 ;
  assign y7905 = n30617 ;
  assign y7906 = ~n30619 ;
  assign y7907 = ~n30623 ;
  assign y7908 = ~n30629 ;
  assign y7909 = n30634 ;
  assign y7910 = ~1'b0 ;
  assign y7911 = ~n30635 ;
  assign y7912 = n30637 ;
  assign y7913 = ~n30638 ;
  assign y7914 = n30640 ;
  assign y7915 = ~n30645 ;
  assign y7916 = ~n30646 ;
  assign y7917 = ~n30648 ;
  assign y7918 = ~n30652 ;
  assign y7919 = n30653 ;
  assign y7920 = ~n30655 ;
  assign y7921 = ~n30658 ;
  assign y7922 = ~n30664 ;
  assign y7923 = ~n30673 ;
  assign y7924 = ~1'b0 ;
  assign y7925 = n30679 ;
  assign y7926 = ~n30684 ;
  assign y7927 = ~n30685 ;
  assign y7928 = ~n30687 ;
  assign y7929 = n30690 ;
  assign y7930 = ~n30693 ;
  assign y7931 = ~1'b0 ;
  assign y7932 = n30697 ;
  assign y7933 = n30699 ;
  assign y7934 = n30703 ;
  assign y7935 = n30708 ;
  assign y7936 = ~n30716 ;
  assign y7937 = n30719 ;
  assign y7938 = ~n30721 ;
  assign y7939 = n30722 ;
  assign y7940 = n30723 ;
  assign y7941 = ~n30725 ;
  assign y7942 = n30726 ;
  assign y7943 = n30731 ;
  assign y7944 = ~n30738 ;
  assign y7945 = ~n30741 ;
  assign y7946 = n30746 ;
  assign y7947 = n30747 ;
  assign y7948 = n30754 ;
  assign y7949 = n30755 ;
  assign y7950 = n30758 ;
  assign y7951 = n30759 ;
  assign y7952 = ~n30764 ;
  assign y7953 = ~n30767 ;
  assign y7954 = ~1'b0 ;
  assign y7955 = ~1'b0 ;
  assign y7956 = n30771 ;
  assign y7957 = ~n30776 ;
  assign y7958 = ~n30777 ;
  assign y7959 = n30779 ;
  assign y7960 = n30781 ;
  assign y7961 = n30782 ;
  assign y7962 = n30783 ;
  assign y7963 = n30785 ;
  assign y7964 = n30789 ;
  assign y7965 = n30791 ;
  assign y7966 = ~n30794 ;
  assign y7967 = n30795 ;
  assign y7968 = ~1'b0 ;
  assign y7969 = n30800 ;
  assign y7970 = ~n30802 ;
  assign y7971 = n30806 ;
  assign y7972 = n30812 ;
  assign y7973 = n30816 ;
  assign y7974 = n30819 ;
  assign y7975 = n30824 ;
  assign y7976 = ~n30825 ;
  assign y7977 = ~n30829 ;
  assign y7978 = ~n30832 ;
  assign y7979 = n30833 ;
  assign y7980 = n30835 ;
  assign y7981 = n30837 ;
  assign y7982 = n30840 ;
  assign y7983 = n30850 ;
  assign y7984 = ~n30852 ;
  assign y7985 = ~n30854 ;
  assign y7986 = n30857 ;
  assign y7987 = ~n30865 ;
  assign y7988 = n30870 ;
  assign y7989 = ~1'b0 ;
  assign y7990 = n30879 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = n30881 ;
  assign y7993 = n30882 ;
  assign y7994 = ~1'b0 ;
  assign y7995 = ~n30888 ;
  assign y7996 = ~n30890 ;
  assign y7997 = n30901 ;
  assign y7998 = n30905 ;
  assign y7999 = n30907 ;
  assign y8000 = n30909 ;
  assign y8001 = n30910 ;
  assign y8002 = ~n30912 ;
  assign y8003 = n30927 ;
  assign y8004 = n18917 ;
  assign y8005 = n30930 ;
  assign y8006 = ~n30935 ;
  assign y8007 = n30939 ;
  assign y8008 = n30945 ;
  assign y8009 = ~n30947 ;
  assign y8010 = ~n30948 ;
  assign y8011 = n30950 ;
  assign y8012 = n30958 ;
  assign y8013 = ~n30964 ;
  assign y8014 = n30967 ;
  assign y8015 = n30968 ;
  assign y8016 = n30969 ;
  assign y8017 = n30976 ;
  assign y8018 = ~n30979 ;
  assign y8019 = n30981 ;
  assign y8020 = ~n30983 ;
  assign y8021 = n30988 ;
  assign y8022 = ~n30989 ;
  assign y8023 = n30990 ;
  assign y8024 = n30993 ;
  assign y8025 = ~n30994 ;
  assign y8026 = n30995 ;
  assign y8027 = ~n30999 ;
  assign y8028 = ~1'b0 ;
  assign y8029 = n31001 ;
  assign y8030 = n31003 ;
  assign y8031 = n31005 ;
  assign y8032 = ~n31009 ;
  assign y8033 = ~n31012 ;
  assign y8034 = ~1'b0 ;
  assign y8035 = ~n31014 ;
  assign y8036 = n31021 ;
  assign y8037 = n31022 ;
  assign y8038 = ~n31025 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = ~n31027 ;
  assign y8041 = n31031 ;
  assign y8042 = n31035 ;
  assign y8043 = n31037 ;
  assign y8044 = ~1'b0 ;
  assign y8045 = n31038 ;
  assign y8046 = ~n31039 ;
  assign y8047 = n31040 ;
  assign y8048 = n31041 ;
  assign y8049 = n31050 ;
  assign y8050 = ~1'b0 ;
  assign y8051 = ~n31051 ;
  assign y8052 = n31054 ;
  assign y8053 = n31057 ;
  assign y8054 = ~n31059 ;
  assign y8055 = ~n31060 ;
  assign y8056 = ~n31064 ;
  assign y8057 = ~n31066 ;
  assign y8058 = n31067 ;
  assign y8059 = n31069 ;
  assign y8060 = ~n31070 ;
  assign y8061 = ~n31071 ;
  assign y8062 = n31084 ;
  assign y8063 = ~n31088 ;
  assign y8064 = n31092 ;
  assign y8065 = n31093 ;
  assign y8066 = ~n31095 ;
  assign y8067 = n31096 ;
  assign y8068 = n31104 ;
  assign y8069 = n31105 ;
  assign y8070 = n31106 ;
  assign y8071 = n31108 ;
  assign y8072 = ~1'b0 ;
  assign y8073 = n31115 ;
  assign y8074 = n31116 ;
  assign y8075 = ~n31117 ;
  assign y8076 = n31119 ;
  assign y8077 = ~n31121 ;
  assign y8078 = n31122 ;
  assign y8079 = ~n31125 ;
  assign y8080 = n31128 ;
  assign y8081 = ~n31129 ;
  assign y8082 = n31131 ;
  assign y8083 = ~n31134 ;
  assign y8084 = n31138 ;
  assign y8085 = ~n31140 ;
  assign y8086 = ~n31142 ;
  assign y8087 = ~n31143 ;
  assign y8088 = ~n31146 ;
  assign y8089 = n31149 ;
  assign y8090 = n31151 ;
  assign y8091 = n31155 ;
  assign y8092 = n31161 ;
  assign y8093 = ~n31164 ;
  assign y8094 = ~n31166 ;
  assign y8095 = n31168 ;
  assign y8096 = ~n31176 ;
  assign y8097 = n31179 ;
  assign y8098 = ~n31180 ;
  assign y8099 = ~n31182 ;
  assign y8100 = ~n31183 ;
  assign y8101 = n31185 ;
  assign y8102 = ~n31188 ;
  assign y8103 = ~n31190 ;
  assign y8104 = ~n31196 ;
  assign y8105 = ~n31199 ;
  assign y8106 = ~n31203 ;
  assign y8107 = ~n31204 ;
  assign y8108 = n31206 ;
  assign y8109 = n31208 ;
  assign y8110 = ~n31210 ;
  assign y8111 = ~n31212 ;
  assign y8112 = n31216 ;
  assign y8113 = n31219 ;
  assign y8114 = ~1'b0 ;
  assign y8115 = ~n31226 ;
  assign y8116 = n31228 ;
  assign y8117 = n31230 ;
  assign y8118 = ~n31234 ;
  assign y8119 = ~n31243 ;
  assign y8120 = ~n31247 ;
  assign y8121 = ~n31249 ;
  assign y8122 = n31251 ;
  assign y8123 = n31252 ;
  assign y8124 = ~n31261 ;
  assign y8125 = ~n31264 ;
  assign y8126 = n31266 ;
  assign y8127 = ~n31268 ;
  assign y8128 = n31279 ;
  assign y8129 = ~n31282 ;
  assign y8130 = n31285 ;
  assign y8131 = ~1'b0 ;
  assign y8132 = ~n31286 ;
  assign y8133 = ~n31289 ;
  assign y8134 = n31292 ;
  assign y8135 = n31294 ;
  assign y8136 = n31295 ;
  assign y8137 = n31299 ;
  assign y8138 = ~n31304 ;
  assign y8139 = ~n31306 ;
  assign y8140 = ~n31308 ;
  assign y8141 = n31309 ;
  assign y8142 = n31312 ;
  assign y8143 = n31314 ;
  assign y8144 = ~n31317 ;
  assign y8145 = n31321 ;
  assign y8146 = ~n31325 ;
  assign y8147 = ~n31331 ;
  assign y8148 = n31333 ;
  assign y8149 = n31335 ;
  assign y8150 = ~n31351 ;
  assign y8151 = n31352 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = ~1'b0 ;
  assign y8154 = ~n31353 ;
  assign y8155 = n31358 ;
  assign y8156 = n31361 ;
  assign y8157 = n31364 ;
  assign y8158 = n31369 ;
  assign y8159 = ~1'b0 ;
  assign y8160 = ~n31370 ;
  assign y8161 = ~n31371 ;
  assign y8162 = ~n31373 ;
  assign y8163 = ~n31375 ;
  assign y8164 = ~n31377 ;
  assign y8165 = ~n31379 ;
  assign y8166 = ~n31380 ;
  assign y8167 = ~n31381 ;
  assign y8168 = n31391 ;
  assign y8169 = ~n31392 ;
  assign y8170 = n31395 ;
  assign y8171 = n31398 ;
  assign y8172 = ~n31403 ;
  assign y8173 = ~n31408 ;
  assign y8174 = n31411 ;
  assign y8175 = n31412 ;
  assign y8176 = ~1'b0 ;
  assign y8177 = ~n31418 ;
  assign y8178 = n31420 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = n31421 ;
  assign y8181 = ~n31425 ;
  assign y8182 = n31431 ;
  assign y8183 = ~n31437 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~n31438 ;
  assign y8186 = ~n31443 ;
  assign y8187 = n31447 ;
  assign y8188 = ~n31449 ;
  assign y8189 = ~n31450 ;
  assign y8190 = ~n31454 ;
  assign y8191 = ~n31457 ;
  assign y8192 = ~1'b0 ;
  assign y8193 = ~n31459 ;
  assign y8194 = ~n31461 ;
  assign y8195 = n31463 ;
  assign y8196 = ~n31466 ;
  assign y8197 = ~n31469 ;
  assign y8198 = ~1'b0 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = ~n31473 ;
  assign y8201 = ~n31474 ;
  assign y8202 = n31475 ;
  assign y8203 = ~n31478 ;
  assign y8204 = ~n31481 ;
  assign y8205 = n31488 ;
  assign y8206 = n31490 ;
  assign y8207 = n31491 ;
  assign y8208 = ~n31493 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = n31497 ;
  assign y8211 = n31500 ;
  assign y8212 = n31513 ;
  assign y8213 = ~n31514 ;
  assign y8214 = ~n31515 ;
  assign y8215 = n31517 ;
  assign y8216 = n31519 ;
  assign y8217 = n31525 ;
  assign y8218 = ~n31526 ;
  assign y8219 = n31531 ;
  assign y8220 = ~n31533 ;
  assign y8221 = n31544 ;
  assign y8222 = ~1'b0 ;
  assign y8223 = ~n31555 ;
  assign y8224 = ~n31558 ;
  assign y8225 = ~n31560 ;
  assign y8226 = n31563 ;
  assign y8227 = n31565 ;
  assign y8228 = n31576 ;
  assign y8229 = n31582 ;
  assign y8230 = ~n31583 ;
  assign y8231 = n31584 ;
  assign y8232 = n31585 ;
  assign y8233 = ~n31596 ;
  assign y8234 = n31600 ;
  assign y8235 = ~n31601 ;
  assign y8236 = ~n31608 ;
  assign y8237 = n31609 ;
  assign y8238 = n31617 ;
  assign y8239 = n31619 ;
  assign y8240 = ~n31623 ;
  assign y8241 = n31624 ;
  assign y8242 = ~n31626 ;
  assign y8243 = ~n31631 ;
  assign y8244 = ~n31634 ;
  assign y8245 = n31641 ;
  assign y8246 = n31642 ;
  assign y8247 = n31644 ;
  assign y8248 = ~n31652 ;
  assign y8249 = ~n31653 ;
  assign y8250 = n31659 ;
  assign y8251 = ~1'b0 ;
  assign y8252 = ~1'b0 ;
  assign y8253 = n31661 ;
  assign y8254 = n31663 ;
  assign y8255 = ~n31666 ;
  assign y8256 = n21866 ;
  assign y8257 = ~n31667 ;
  assign y8258 = n31670 ;
  assign y8259 = ~n31673 ;
  assign y8260 = n31682 ;
  assign y8261 = ~n31683 ;
  assign y8262 = ~n31684 ;
  assign y8263 = n31686 ;
  assign y8264 = ~1'b0 ;
  assign y8265 = n31688 ;
  assign y8266 = n31690 ;
  assign y8267 = ~n31691 ;
  assign y8268 = ~n31693 ;
  assign y8269 = ~n31695 ;
  assign y8270 = ~1'b0 ;
  assign y8271 = n31696 ;
  assign y8272 = ~n31699 ;
  assign y8273 = n31709 ;
  assign y8274 = ~1'b0 ;
  assign y8275 = ~n31713 ;
  assign y8276 = ~n31715 ;
  assign y8277 = n31717 ;
  assign y8278 = ~n31719 ;
  assign y8279 = n31726 ;
  assign y8280 = ~n31729 ;
  assign y8281 = n31731 ;
  assign y8282 = ~n31732 ;
  assign y8283 = n31734 ;
  assign y8284 = ~1'b0 ;
  assign y8285 = n31741 ;
  assign y8286 = n31743 ;
  assign y8287 = n31749 ;
  assign y8288 = ~n31752 ;
  assign y8289 = ~n31754 ;
  assign y8290 = n31756 ;
  assign y8291 = ~n31758 ;
  assign y8292 = ~n31761 ;
  assign y8293 = ~n31763 ;
  assign y8294 = n31766 ;
  assign y8295 = n31767 ;
  assign y8296 = ~n31770 ;
  assign y8297 = n31775 ;
  assign y8298 = n31779 ;
  assign y8299 = ~n31788 ;
  assign y8300 = n31793 ;
  assign y8301 = ~n31795 ;
  assign y8302 = ~n31796 ;
  assign y8303 = ~1'b0 ;
  assign y8304 = ~1'b0 ;
  assign y8305 = ~n31797 ;
  assign y8306 = n31798 ;
  assign y8307 = n31799 ;
  assign y8308 = ~n31805 ;
  assign y8309 = ~n31807 ;
  assign y8310 = n31811 ;
  assign y8311 = n31814 ;
  assign y8312 = ~n31815 ;
  assign y8313 = ~1'b0 ;
  assign y8314 = n31816 ;
  assign y8315 = n31818 ;
  assign y8316 = ~n31819 ;
  assign y8317 = ~n31823 ;
  assign y8318 = ~n31826 ;
  assign y8319 = ~n31828 ;
  assign y8320 = n31833 ;
  assign y8321 = ~n31837 ;
  assign y8322 = ~n31838 ;
  assign y8323 = ~n31842 ;
  assign y8324 = ~n31845 ;
  assign y8325 = ~n31848 ;
  assign y8326 = ~n31852 ;
  assign y8327 = ~1'b0 ;
  assign y8328 = n31853 ;
  assign y8329 = n31854 ;
  assign y8330 = n31859 ;
  assign y8331 = ~n31862 ;
  assign y8332 = ~n31866 ;
  assign y8333 = ~n31867 ;
  assign y8334 = n31870 ;
  assign y8335 = n31873 ;
  assign y8336 = n31875 ;
  assign y8337 = ~1'b0 ;
  assign y8338 = ~n31879 ;
  assign y8339 = ~n31880 ;
  assign y8340 = ~n31883 ;
  assign y8341 = ~n31885 ;
  assign y8342 = n31889 ;
  assign y8343 = ~n31895 ;
  assign y8344 = n31898 ;
  assign y8345 = ~n31904 ;
  assign y8346 = n31905 ;
  assign y8347 = n31906 ;
  assign y8348 = ~n31908 ;
  assign y8349 = n31911 ;
  assign y8350 = n31914 ;
  assign y8351 = ~n31916 ;
  assign y8352 = ~n31917 ;
  assign y8353 = ~n31918 ;
  assign y8354 = n31920 ;
  assign y8355 = ~1'b0 ;
  assign y8356 = n31927 ;
  assign y8357 = n31932 ;
  assign y8358 = n31939 ;
  assign y8359 = ~n31941 ;
  assign y8360 = n31943 ;
  assign y8361 = n31944 ;
  assign y8362 = n31947 ;
  assign y8363 = ~1'b0 ;
  assign y8364 = ~1'b0 ;
  assign y8365 = n31949 ;
  assign y8366 = n31951 ;
  assign y8367 = n31952 ;
  assign y8368 = ~n31954 ;
  assign y8369 = ~n31959 ;
  assign y8370 = ~1'b0 ;
  assign y8371 = ~n31960 ;
  assign y8372 = ~n31964 ;
  assign y8373 = n23062 ;
  assign y8374 = ~n31966 ;
  assign y8375 = ~n31967 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = n31968 ;
  assign y8378 = n31975 ;
  assign y8379 = n31976 ;
  assign y8380 = ~n31981 ;
  assign y8381 = n31982 ;
  assign y8382 = n31985 ;
  assign y8383 = ~n31987 ;
  assign y8384 = n31990 ;
  assign y8385 = ~1'b0 ;
  assign y8386 = ~1'b0 ;
  assign y8387 = ~n31991 ;
  assign y8388 = n31992 ;
  assign y8389 = ~n31998 ;
  assign y8390 = ~1'b0 ;
  assign y8391 = ~n27649 ;
  assign y8392 = n31999 ;
  assign y8393 = n32006 ;
  assign y8394 = n32007 ;
  assign y8395 = ~n32015 ;
  assign y8396 = ~n32017 ;
  assign y8397 = n32021 ;
  assign y8398 = ~n32022 ;
  assign y8399 = ~n32023 ;
  assign y8400 = ~n32025 ;
  assign y8401 = ~n32028 ;
  assign y8402 = ~n32030 ;
  assign y8403 = ~n32034 ;
  assign y8404 = n32039 ;
  assign y8405 = ~1'b0 ;
  assign y8406 = ~n32041 ;
  assign y8407 = ~n32043 ;
  assign y8408 = n32048 ;
  assign y8409 = n32049 ;
  assign y8410 = ~n32052 ;
  assign y8411 = n32053 ;
  assign y8412 = ~n32056 ;
  assign y8413 = n32062 ;
  assign y8414 = ~n32063 ;
  assign y8415 = ~n32064 ;
  assign y8416 = n32069 ;
  assign y8417 = ~n32076 ;
  assign y8418 = n32080 ;
  assign y8419 = n32090 ;
  assign y8420 = n32091 ;
  assign y8421 = ~n32093 ;
  assign y8422 = ~1'b0 ;
  assign y8423 = n31049 ;
  assign y8424 = n32094 ;
  assign y8425 = n32102 ;
  assign y8426 = n32104 ;
  assign y8427 = n32109 ;
  assign y8428 = ~n32113 ;
  assign y8429 = ~n32115 ;
  assign y8430 = ~n32126 ;
  assign y8431 = n32129 ;
  assign y8432 = ~n32134 ;
  assign y8433 = ~n32136 ;
  assign y8434 = ~1'b0 ;
  assign y8435 = n32139 ;
  assign y8436 = n32140 ;
  assign y8437 = ~n32144 ;
  assign y8438 = ~n32145 ;
  assign y8439 = ~n32148 ;
  assign y8440 = n32152 ;
  assign y8441 = n32154 ;
  assign y8442 = n32155 ;
  assign y8443 = ~n32160 ;
  assign y8444 = ~n32164 ;
  assign y8445 = n32165 ;
  assign y8446 = ~1'b0 ;
  assign y8447 = n32166 ;
  assign y8448 = n32169 ;
  assign y8449 = n32170 ;
  assign y8450 = ~n32171 ;
  assign y8451 = ~1'b0 ;
  assign y8452 = n32172 ;
  assign y8453 = ~n32174 ;
  assign y8454 = n32178 ;
  assign y8455 = ~n32180 ;
  assign y8456 = ~n8194 ;
  assign y8457 = n32181 ;
  assign y8458 = ~n32183 ;
  assign y8459 = ~n32190 ;
  assign y8460 = ~n32191 ;
  assign y8461 = n32201 ;
  assign y8462 = ~n32203 ;
  assign y8463 = ~n32206 ;
  assign y8464 = ~n32209 ;
  assign y8465 = ~n32210 ;
  assign y8466 = n32213 ;
  assign y8467 = n32216 ;
  assign y8468 = n32220 ;
  assign y8469 = n32225 ;
  assign y8470 = 1'b0 ;
  assign y8471 = n32226 ;
  assign y8472 = ~n32228 ;
  assign y8473 = ~1'b0 ;
  assign y8474 = n32229 ;
  assign y8475 = ~n32233 ;
  assign y8476 = ~n32236 ;
  assign y8477 = n32239 ;
  assign y8478 = n32246 ;
  assign y8479 = n32247 ;
  assign y8480 = ~n32249 ;
  assign y8481 = ~n32252 ;
  assign y8482 = n32258 ;
  assign y8483 = n32260 ;
  assign y8484 = ~n32268 ;
  assign y8485 = ~n32272 ;
  assign y8486 = n32274 ;
  assign y8487 = ~n32276 ;
  assign y8488 = ~n32279 ;
  assign y8489 = n32283 ;
  assign y8490 = ~n32285 ;
  assign y8491 = ~n32297 ;
  assign y8492 = ~n32298 ;
  assign y8493 = ~n32299 ;
  assign y8494 = n32300 ;
  assign y8495 = n32306 ;
  assign y8496 = ~n32307 ;
  assign y8497 = ~n32309 ;
  assign y8498 = ~1'b0 ;
  assign y8499 = n32311 ;
  assign y8500 = ~n32313 ;
  assign y8501 = ~n32315 ;
  assign y8502 = n32322 ;
  assign y8503 = ~n32325 ;
  assign y8504 = n32326 ;
  assign y8505 = ~n32327 ;
  assign y8506 = ~n32329 ;
  assign y8507 = ~n32330 ;
  assign y8508 = ~n32335 ;
  assign y8509 = ~n32337 ;
  assign y8510 = n32338 ;
  assign y8511 = n32344 ;
  assign y8512 = ~n32346 ;
  assign y8513 = n32347 ;
  assign y8514 = n32348 ;
  assign y8515 = n32349 ;
  assign y8516 = ~n32352 ;
  assign y8517 = n32358 ;
  assign y8518 = ~1'b0 ;
  assign y8519 = ~n32360 ;
  assign y8520 = ~1'b0 ;
  assign y8521 = ~n32364 ;
  assign y8522 = ~1'b0 ;
  assign y8523 = n32371 ;
  assign y8524 = ~n32382 ;
  assign y8525 = n32383 ;
  assign y8526 = n32385 ;
  assign y8527 = ~n32388 ;
  assign y8528 = n32390 ;
  assign y8529 = ~n32394 ;
  assign y8530 = ~n32396 ;
  assign y8531 = n30804 ;
  assign y8532 = n32399 ;
  assign y8533 = n32400 ;
  assign y8534 = ~n32407 ;
  assign y8535 = n32408 ;
  assign y8536 = ~n32410 ;
  assign y8537 = n32412 ;
  assign y8538 = ~n32417 ;
  assign y8539 = n32418 ;
  assign y8540 = n32424 ;
  assign y8541 = ~n32427 ;
  assign y8542 = n32432 ;
  assign y8543 = n32437 ;
  assign y8544 = n32440 ;
  assign y8545 = ~n32447 ;
  assign y8546 = ~n32448 ;
  assign y8547 = n32449 ;
  assign y8548 = ~n32450 ;
  assign y8549 = ~n32452 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~n32455 ;
  assign y8552 = ~n32456 ;
  assign y8553 = ~n32457 ;
  assign y8554 = n32460 ;
  assign y8555 = ~n32462 ;
  assign y8556 = ~n32473 ;
  assign y8557 = ~n32480 ;
  assign y8558 = ~n32482 ;
  assign y8559 = ~n32486 ;
  assign y8560 = ~n32489 ;
  assign y8561 = ~n32492 ;
  assign y8562 = n32494 ;
  assign y8563 = n32496 ;
  assign y8564 = ~n32499 ;
  assign y8565 = ~n32506 ;
  assign y8566 = ~1'b0 ;
  assign y8567 = ~n32508 ;
  assign y8568 = ~n32509 ;
  assign y8569 = n32511 ;
  assign y8570 = ~n32512 ;
  assign y8571 = ~n32516 ;
  assign y8572 = ~n32519 ;
  assign y8573 = n32521 ;
  assign y8574 = n32522 ;
  assign y8575 = n32523 ;
  assign y8576 = ~n32526 ;
  assign y8577 = ~1'b0 ;
  assign y8578 = ~n32529 ;
  assign y8579 = ~n32531 ;
  assign y8580 = n32537 ;
  assign y8581 = ~n32542 ;
  assign y8582 = n32545 ;
  assign y8583 = n32548 ;
  assign y8584 = ~n32549 ;
  assign y8585 = n32553 ;
  assign y8586 = ~1'b0 ;
  assign y8587 = ~n32554 ;
  assign y8588 = n32558 ;
  assign y8589 = ~n32562 ;
  assign y8590 = n32563 ;
  assign y8591 = ~n32569 ;
  assign y8592 = ~1'b0 ;
  assign y8593 = ~1'b0 ;
  assign y8594 = ~n32576 ;
  assign y8595 = ~n32578 ;
  assign y8596 = ~n32583 ;
  assign y8597 = n32584 ;
  assign y8598 = ~n32589 ;
  assign y8599 = ~n32590 ;
  assign y8600 = n32596 ;
  assign y8601 = ~n32600 ;
  assign y8602 = n32601 ;
  assign y8603 = n32608 ;
  assign y8604 = ~1'b0 ;
  assign y8605 = n32609 ;
  assign y8606 = ~1'b0 ;
  assign y8607 = ~n32616 ;
  assign y8608 = ~n32619 ;
  assign y8609 = n32621 ;
  assign y8610 = n32625 ;
  assign y8611 = n32627 ;
  assign y8612 = ~1'b0 ;
  assign y8613 = ~1'b0 ;
  assign y8614 = n32628 ;
  assign y8615 = ~n32631 ;
  assign y8616 = n32644 ;
  assign y8617 = ~n32645 ;
  assign y8618 = n32646 ;
  assign y8619 = n32648 ;
  assign y8620 = n32652 ;
  assign y8621 = ~1'b0 ;
  assign y8622 = ~n32655 ;
  assign y8623 = ~n32657 ;
  assign y8624 = ~n32661 ;
  assign y8625 = n32665 ;
  assign y8626 = ~n32667 ;
  assign y8627 = n32672 ;
  assign y8628 = n32673 ;
  assign y8629 = ~1'b0 ;
  assign y8630 = ~n32675 ;
  assign y8631 = n32679 ;
  assign y8632 = ~n32680 ;
  assign y8633 = ~n32682 ;
  assign y8634 = n32684 ;
  assign y8635 = n32686 ;
  assign y8636 = ~n32691 ;
  assign y8637 = n32693 ;
  assign y8638 = ~n32694 ;
  assign y8639 = n32695 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = n32697 ;
  assign y8642 = ~1'b0 ;
  assign y8643 = n32701 ;
  assign y8644 = n32704 ;
  assign y8645 = n32709 ;
  assign y8646 = n32711 ;
  assign y8647 = n32715 ;
  assign y8648 = n32717 ;
  assign y8649 = n32718 ;
  assign y8650 = n32722 ;
  assign y8651 = n32725 ;
  assign y8652 = n32732 ;
  assign y8653 = ~n32733 ;
  assign y8654 = ~n32734 ;
  assign y8655 = ~n32735 ;
  assign y8656 = n32737 ;
  assign y8657 = ~n32738 ;
  assign y8658 = ~n32739 ;
  assign y8659 = ~n32742 ;
  assign y8660 = n32750 ;
  assign y8661 = n32757 ;
  assign y8662 = ~n32759 ;
  assign y8663 = n32760 ;
  assign y8664 = ~n32762 ;
  assign y8665 = n12473 ;
  assign y8666 = n32763 ;
  assign y8667 = ~n32768 ;
  assign y8668 = n32774 ;
  assign y8669 = ~n32776 ;
  assign y8670 = n32778 ;
  assign y8671 = ~n32780 ;
  assign y8672 = ~n32783 ;
  assign y8673 = ~n32784 ;
  assign y8674 = ~1'b0 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = n32786 ;
  assign y8677 = n32789 ;
  assign y8678 = n32791 ;
  assign y8679 = ~n7158 ;
  assign y8680 = ~n32792 ;
  assign y8681 = ~n32793 ;
  assign y8682 = n32795 ;
  assign y8683 = ~n32797 ;
  assign y8684 = ~n32799 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = ~n32803 ;
  assign y8687 = ~n32810 ;
  assign y8688 = ~n32812 ;
  assign y8689 = n32813 ;
  assign y8690 = ~n32814 ;
  assign y8691 = n32815 ;
  assign y8692 = ~n32817 ;
  assign y8693 = n32822 ;
  assign y8694 = n32830 ;
  assign y8695 = n32831 ;
  assign y8696 = ~n550 ;
  assign y8697 = ~n32836 ;
  assign y8698 = n32839 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = ~n32840 ;
  assign y8701 = n32841 ;
  assign y8702 = n32842 ;
  assign y8703 = n32844 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = ~n32849 ;
  assign y8706 = ~n32850 ;
  assign y8707 = ~n32854 ;
  assign y8708 = n32859 ;
  assign y8709 = n32863 ;
  assign y8710 = ~n32866 ;
  assign y8711 = ~n32870 ;
  assign y8712 = n32873 ;
  assign y8713 = ~n32876 ;
  assign y8714 = ~n32880 ;
  assign y8715 = ~n32884 ;
  assign y8716 = 1'b0 ;
  assign y8717 = n32887 ;
  assign y8718 = ~n32891 ;
  assign y8719 = ~n32894 ;
  assign y8720 = n32898 ;
  assign y8721 = ~n32903 ;
  assign y8722 = ~n32904 ;
  assign y8723 = n1527 ;
  assign y8724 = ~1'b0 ;
  assign y8725 = ~n32908 ;
  assign y8726 = ~n32910 ;
  assign y8727 = ~n32917 ;
  assign y8728 = n32920 ;
  assign y8729 = n32924 ;
  assign y8730 = ~n32925 ;
  assign y8731 = ~n32929 ;
  assign y8732 = ~n32931 ;
  assign y8733 = n32945 ;
  assign y8734 = ~n32947 ;
  assign y8735 = ~n32949 ;
  assign y8736 = ~n32950 ;
  assign y8737 = ~1'b0 ;
  assign y8738 = ~n32957 ;
  assign y8739 = ~n32959 ;
  assign y8740 = n32962 ;
  assign y8741 = ~n32963 ;
  assign y8742 = n32964 ;
  assign y8743 = ~n32968 ;
  assign y8744 = n32969 ;
  assign y8745 = ~n32970 ;
  assign y8746 = ~n32972 ;
  assign y8747 = n32975 ;
  assign y8748 = ~n32979 ;
  assign y8749 = n32983 ;
  assign y8750 = n32984 ;
  assign y8751 = n32987 ;
  assign y8752 = ~n32988 ;
  assign y8753 = ~1'b0 ;
  assign y8754 = n32992 ;
  assign y8755 = n32996 ;
  assign y8756 = ~n32997 ;
  assign y8757 = ~n33002 ;
  assign y8758 = n33006 ;
  assign y8759 = ~1'b0 ;
  assign y8760 = n33007 ;
  assign y8761 = ~n33010 ;
  assign y8762 = n33015 ;
  assign y8763 = ~n33021 ;
  assign y8764 = ~n33023 ;
  assign y8765 = n33025 ;
  assign y8766 = ~n33027 ;
  assign y8767 = ~n33030 ;
  assign y8768 = ~1'b0 ;
  assign y8769 = n33032 ;
  assign y8770 = n33034 ;
  assign y8771 = ~1'b0 ;
  assign y8772 = ~1'b0 ;
  assign y8773 = ~n33036 ;
  assign y8774 = n33048 ;
  assign y8775 = n33051 ;
  assign y8776 = ~n33052 ;
  assign y8777 = n33053 ;
  assign y8778 = ~1'b0 ;
  assign y8779 = ~1'b0 ;
  assign y8780 = n33055 ;
  assign y8781 = ~n33057 ;
  assign y8782 = n33058 ;
  assign y8783 = ~n33062 ;
  assign y8784 = n33065 ;
  assign y8785 = n33069 ;
  assign y8786 = ~n33071 ;
  assign y8787 = n33072 ;
  assign y8788 = ~n33075 ;
  assign y8789 = n33078 ;
  assign y8790 = ~1'b0 ;
  assign y8791 = n33081 ;
  assign y8792 = n33082 ;
  assign y8793 = n33087 ;
  assign y8794 = ~1'b0 ;
  assign y8795 = ~n33090 ;
  assign y8796 = n33091 ;
  assign y8797 = ~n33094 ;
  assign y8798 = n33096 ;
  assign y8799 = n33099 ;
  assign y8800 = n33105 ;
  assign y8801 = ~n33113 ;
  assign y8802 = n33121 ;
  assign y8803 = n33123 ;
  assign y8804 = n33129 ;
  assign y8805 = ~n33131 ;
  assign y8806 = ~n33135 ;
  assign y8807 = ~n33141 ;
  assign y8808 = ~n33147 ;
  assign y8809 = ~1'b0 ;
  assign y8810 = ~n33148 ;
  assign y8811 = ~n33149 ;
  assign y8812 = n33150 ;
  assign y8813 = ~n33151 ;
  assign y8814 = n33155 ;
  assign y8815 = ~n33157 ;
  assign y8816 = n33158 ;
  assign y8817 = ~1'b0 ;
  assign y8818 = ~n33160 ;
  assign y8819 = ~1'b0 ;
  assign y8820 = ~1'b0 ;
  assign y8821 = n33161 ;
  assign y8822 = ~n33162 ;
  assign y8823 = ~n33164 ;
  assign y8824 = n33167 ;
  assign y8825 = ~1'b0 ;
  assign y8826 = n33169 ;
  assign y8827 = ~n33170 ;
  assign y8828 = n33171 ;
  assign y8829 = ~1'b0 ;
  assign y8830 = ~n33182 ;
  assign y8831 = n33183 ;
  assign y8832 = ~n33186 ;
  assign y8833 = n33187 ;
  assign y8834 = ~n33195 ;
  assign y8835 = ~n33196 ;
  assign y8836 = ~n33199 ;
  assign y8837 = ~n33204 ;
  assign y8838 = n33206 ;
  assign y8839 = ~n33209 ;
  assign y8840 = ~n33212 ;
  assign y8841 = ~n33213 ;
  assign y8842 = ~n33215 ;
  assign y8843 = n33218 ;
  assign y8844 = ~n33221 ;
  assign y8845 = n33224 ;
  assign y8846 = ~n33226 ;
  assign y8847 = ~n33228 ;
  assign y8848 = n6318 ;
  assign y8849 = ~n33229 ;
  assign y8850 = ~n33231 ;
  assign y8851 = ~n33235 ;
  assign y8852 = ~n33239 ;
  assign y8853 = ~n33240 ;
  assign y8854 = n33249 ;
  assign y8855 = n33254 ;
  assign y8856 = n33258 ;
  assign y8857 = ~n33265 ;
  assign y8858 = ~n33266 ;
  assign y8859 = n33267 ;
  assign y8860 = 1'b0 ;
  assign y8861 = n33270 ;
  assign y8862 = ~n33275 ;
  assign y8863 = n33277 ;
  assign y8864 = ~n33278 ;
  assign y8865 = ~n33280 ;
  assign y8866 = n33281 ;
  assign y8867 = ~n33286 ;
  assign y8868 = ~n33289 ;
  assign y8869 = n33293 ;
  assign y8870 = ~n33295 ;
  assign y8871 = ~n33301 ;
  assign y8872 = n33302 ;
  assign y8873 = ~1'b0 ;
  assign y8874 = ~1'b0 ;
  assign y8875 = ~n33307 ;
  assign y8876 = ~1'b0 ;
  assign y8877 = ~n33310 ;
  assign y8878 = ~n33313 ;
  assign y8879 = ~n33315 ;
  assign y8880 = ~n33318 ;
  assign y8881 = n33319 ;
  assign y8882 = ~n33320 ;
  assign y8883 = n33322 ;
  assign y8884 = n33324 ;
  assign y8885 = n33329 ;
  assign y8886 = n33331 ;
  assign y8887 = n33333 ;
  assign y8888 = n33340 ;
  assign y8889 = n33341 ;
  assign y8890 = ~n33344 ;
  assign y8891 = ~n33347 ;
  assign y8892 = ~n33350 ;
  assign y8893 = ~n33355 ;
  assign y8894 = ~1'b0 ;
  assign y8895 = ~n33358 ;
  assign y8896 = ~n33363 ;
  assign y8897 = ~n33370 ;
  assign y8898 = ~n33374 ;
  assign y8899 = n33380 ;
  assign y8900 = n33384 ;
  assign y8901 = ~n33386 ;
  assign y8902 = n33392 ;
  assign y8903 = ~n33393 ;
  assign y8904 = ~n33394 ;
  assign y8905 = ~n33395 ;
  assign y8906 = ~n33399 ;
  assign y8907 = ~n33402 ;
  assign y8908 = ~n33404 ;
  assign y8909 = ~n33406 ;
  assign y8910 = ~n33407 ;
  assign y8911 = n33409 ;
  assign y8912 = ~n33415 ;
  assign y8913 = ~n33416 ;
  assign y8914 = ~n33417 ;
  assign y8915 = ~n33418 ;
  assign y8916 = n33420 ;
  assign y8917 = n33422 ;
  assign y8918 = ~n33423 ;
  assign y8919 = n33424 ;
  assign y8920 = n33427 ;
  assign y8921 = n33429 ;
  assign y8922 = n33431 ;
  assign y8923 = ~n18223 ;
  assign y8924 = ~n33443 ;
  assign y8925 = n33445 ;
  assign y8926 = n33450 ;
  assign y8927 = n33454 ;
  assign y8928 = ~n33455 ;
  assign y8929 = n33460 ;
  assign y8930 = n33465 ;
  assign y8931 = ~n33467 ;
  assign y8932 = ~n33469 ;
  assign y8933 = n33473 ;
  assign y8934 = n33482 ;
  assign y8935 = ~n33487 ;
  assign y8936 = n33488 ;
  assign y8937 = n33491 ;
  assign y8938 = ~n33494 ;
  assign y8939 = ~1'b0 ;
  assign y8940 = n33497 ;
  assign y8941 = ~n2909 ;
  assign y8942 = n33500 ;
  assign y8943 = ~n33502 ;
  assign y8944 = ~1'b0 ;
  assign y8945 = n33503 ;
  assign y8946 = n33505 ;
  assign y8947 = ~n33506 ;
  assign y8948 = ~n33507 ;
  assign y8949 = ~n33509 ;
  assign y8950 = ~n33511 ;
  assign y8951 = ~n33515 ;
  assign y8952 = ~n33517 ;
  assign y8953 = ~n33518 ;
  assign y8954 = ~n33520 ;
  assign y8955 = n33522 ;
  assign y8956 = ~n33527 ;
  assign y8957 = n33528 ;
  assign y8958 = n33530 ;
  assign y8959 = ~n33531 ;
  assign y8960 = ~n33533 ;
  assign y8961 = n33534 ;
  assign y8962 = ~n33542 ;
  assign y8963 = n33544 ;
  assign y8964 = ~n33548 ;
  assign y8965 = n33550 ;
  assign y8966 = ~n33554 ;
  assign y8967 = ~n33555 ;
  assign y8968 = n33560 ;
  assign y8969 = n33561 ;
  assign y8970 = n33572 ;
  assign y8971 = ~n33574 ;
  assign y8972 = n33577 ;
  assign y8973 = ~1'b0 ;
  assign y8974 = n33581 ;
  assign y8975 = n33582 ;
  assign y8976 = ~n33589 ;
  assign y8977 = n33594 ;
  assign y8978 = n33596 ;
  assign y8979 = n33599 ;
  assign y8980 = ~n23091 ;
  assign y8981 = ~n33606 ;
  assign y8982 = ~n33607 ;
  assign y8983 = ~n33609 ;
  assign y8984 = n33613 ;
  assign y8985 = ~n33617 ;
  assign y8986 = n33618 ;
  assign y8987 = ~n33623 ;
  assign y8988 = ~n33625 ;
  assign y8989 = n33626 ;
  assign y8990 = n23555 ;
  assign y8991 = n33631 ;
  assign y8992 = n33636 ;
  assign y8993 = ~1'b0 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = ~n33639 ;
  assign y8996 = n33643 ;
  assign y8997 = n33647 ;
  assign y8998 = n33648 ;
  assign y8999 = ~n33653 ;
  assign y9000 = n33657 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = n33658 ;
  assign y9003 = n33659 ;
  assign y9004 = n33660 ;
  assign y9005 = ~n33661 ;
  assign y9006 = ~n33666 ;
  assign y9007 = n33668 ;
  assign y9008 = n33670 ;
  assign y9009 = n33672 ;
  assign y9010 = n33674 ;
  assign y9011 = ~1'b0 ;
  assign y9012 = n33677 ;
  assign y9013 = n33678 ;
  assign y9014 = ~n33683 ;
  assign y9015 = ~n33685 ;
  assign y9016 = ~n33688 ;
  assign y9017 = n33700 ;
  assign y9018 = ~n33701 ;
  assign y9019 = ~n33702 ;
  assign y9020 = n33709 ;
  assign y9021 = ~1'b0 ;
  assign y9022 = ~n33711 ;
  assign y9023 = n33713 ;
  assign y9024 = n33715 ;
  assign y9025 = n33716 ;
  assign y9026 = ~n33718 ;
  assign y9027 = n33720 ;
  assign y9028 = n33721 ;
  assign y9029 = n33722 ;
  assign y9030 = n33726 ;
  assign y9031 = ~n33727 ;
  assign y9032 = ~n33733 ;
  assign y9033 = n33734 ;
  assign y9034 = ~n33737 ;
  assign y9035 = ~n33740 ;
  assign y9036 = n33748 ;
  assign y9037 = n33751 ;
  assign y9038 = ~n33756 ;
  assign y9039 = ~1'b0 ;
  assign y9040 = n33757 ;
  assign y9041 = ~n33759 ;
  assign y9042 = ~n33775 ;
  assign y9043 = n33779 ;
  assign y9044 = ~n33780 ;
  assign y9045 = ~n33782 ;
  assign y9046 = ~n33783 ;
  assign y9047 = ~n33784 ;
  assign y9048 = n33791 ;
  assign y9049 = n33794 ;
  assign y9050 = n33795 ;
  assign y9051 = ~n33796 ;
  assign y9052 = n33801 ;
  assign y9053 = ~n33802 ;
  assign y9054 = n33809 ;
  assign y9055 = n33811 ;
  assign y9056 = ~n33817 ;
  assign y9057 = n33819 ;
  assign y9058 = ~1'b0 ;
  assign y9059 = ~n33820 ;
  assign y9060 = n33825 ;
  assign y9061 = n33827 ;
  assign y9062 = ~n33831 ;
  assign y9063 = n33833 ;
  assign y9064 = ~n33840 ;
  assign y9065 = ~n33847 ;
  assign y9066 = n33855 ;
  assign y9067 = n33858 ;
  assign y9068 = ~n33861 ;
  assign y9069 = ~n33862 ;
  assign y9070 = ~1'b0 ;
  assign y9071 = n33863 ;
  assign y9072 = ~n1918 ;
  assign y9073 = ~n33864 ;
  assign y9074 = n33865 ;
  assign y9075 = ~n33867 ;
  assign y9076 = ~n33868 ;
  assign y9077 = ~1'b0 ;
  assign y9078 = n33869 ;
  assign y9079 = n33875 ;
  assign y9080 = ~n33879 ;
  assign y9081 = n33881 ;
  assign y9082 = ~n33884 ;
  assign y9083 = n33887 ;
  assign y9084 = n33891 ;
  assign y9085 = n33892 ;
  assign y9086 = ~n33893 ;
  assign y9087 = n33894 ;
  assign y9088 = ~n33900 ;
  assign y9089 = ~1'b0 ;
  assign y9090 = ~1'b0 ;
  assign y9091 = ~n33902 ;
  assign y9092 = ~n33904 ;
  assign y9093 = n33909 ;
  assign y9094 = n33913 ;
  assign y9095 = ~1'b0 ;
  assign y9096 = n33914 ;
  assign y9097 = ~n33918 ;
  assign y9098 = n33919 ;
  assign y9099 = n33921 ;
  assign y9100 = n33922 ;
  assign y9101 = n33924 ;
  assign y9102 = ~n33929 ;
  assign y9103 = ~n33934 ;
  assign y9104 = ~n33939 ;
  assign y9105 = ~n33942 ;
  assign y9106 = ~n33945 ;
  assign y9107 = ~1'b0 ;
  assign y9108 = ~1'b0 ;
  assign y9109 = n33947 ;
  assign y9110 = n33951 ;
  assign y9111 = ~n33958 ;
  assign y9112 = n33959 ;
  assign y9113 = ~n33968 ;
  assign y9114 = ~1'b0 ;
  assign y9115 = ~1'b0 ;
  assign y9116 = ~n33976 ;
  assign y9117 = ~n33977 ;
  assign y9118 = ~n33983 ;
  assign y9119 = ~n33987 ;
  assign y9120 = ~1'b0 ;
  assign y9121 = ~n33989 ;
  assign y9122 = n33990 ;
  assign y9123 = ~1'b0 ;
  assign y9124 = n33991 ;
  assign y9125 = n33994 ;
  assign y9126 = n34000 ;
  assign y9127 = ~1'b0 ;
  assign y9128 = n34002 ;
  assign y9129 = n34004 ;
  assign y9130 = ~n34007 ;
  assign y9131 = n34012 ;
  assign y9132 = ~n34013 ;
  assign y9133 = ~1'b0 ;
  assign y9134 = ~n34015 ;
  assign y9135 = n34019 ;
  assign y9136 = ~n34023 ;
  assign y9137 = ~n34026 ;
  assign y9138 = n34029 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = n34031 ;
  assign y9141 = ~n34035 ;
  assign y9142 = ~n34038 ;
  assign y9143 = n34042 ;
  assign y9144 = n34045 ;
  assign y9145 = n34052 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = ~1'b0 ;
  assign y9148 = ~n34053 ;
  assign y9149 = ~n34055 ;
  assign y9150 = n34059 ;
  assign y9151 = n34060 ;
  assign y9152 = ~n34064 ;
  assign y9153 = ~1'b0 ;
  assign y9154 = n34067 ;
  assign y9155 = n34068 ;
  assign y9156 = ~n34069 ;
  assign y9157 = n34070 ;
  assign y9158 = n34077 ;
  assign y9159 = ~n34080 ;
  assign y9160 = ~n34086 ;
  assign y9161 = n34092 ;
  assign y9162 = ~n34094 ;
  assign y9163 = ~n34096 ;
  assign y9164 = ~n34106 ;
  assign y9165 = n34108 ;
  assign y9166 = ~1'b0 ;
  assign y9167 = ~n34113 ;
  assign y9168 = n34114 ;
  assign y9169 = n34116 ;
  assign y9170 = ~n34122 ;
  assign y9171 = n34123 ;
  assign y9172 = n34125 ;
  assign y9173 = ~n34130 ;
  assign y9174 = n34131 ;
  assign y9175 = ~n34139 ;
  assign y9176 = n34142 ;
  assign y9177 = n26200 ;
  assign y9178 = ~n34143 ;
  assign y9179 = n34149 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = n34151 ;
  assign y9182 = ~n34152 ;
  assign y9183 = ~n34153 ;
  assign y9184 = n34157 ;
  assign y9185 = ~1'b0 ;
  assign y9186 = n34159 ;
  assign y9187 = n34160 ;
  assign y9188 = n34168 ;
  assign y9189 = ~n34170 ;
  assign y9190 = ~n34173 ;
  assign y9191 = ~n34177 ;
  assign y9192 = n34181 ;
  assign y9193 = n34185 ;
  assign y9194 = n34196 ;
  assign y9195 = n34197 ;
  assign y9196 = n34209 ;
  assign y9197 = ~n8144 ;
  assign y9198 = ~n34211 ;
  assign y9199 = ~n34212 ;
  assign y9200 = n34213 ;
  assign y9201 = n34216 ;
  assign y9202 = n34219 ;
  assign y9203 = n34221 ;
  assign y9204 = n34224 ;
  assign y9205 = ~n34231 ;
  assign y9206 = ~n34234 ;
  assign y9207 = n34237 ;
  assign y9208 = n34238 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = n34241 ;
  assign y9211 = n34245 ;
  assign y9212 = n34246 ;
  assign y9213 = n34249 ;
  assign y9214 = ~n34256 ;
  assign y9215 = ~n34258 ;
  assign y9216 = ~n34263 ;
  assign y9217 = n34265 ;
  assign y9218 = ~n34267 ;
  assign y9219 = n34269 ;
  assign y9220 = ~n34270 ;
  assign y9221 = ~n34272 ;
  assign y9222 = ~n34273 ;
  assign y9223 = ~n34278 ;
  assign y9224 = ~n34281 ;
  assign y9225 = n34285 ;
  assign y9226 = ~n34287 ;
  assign y9227 = n34295 ;
  assign y9228 = n34298 ;
  assign y9229 = ~1'b0 ;
  assign y9230 = ~n34299 ;
  assign y9231 = ~n34305 ;
  assign y9232 = ~1'b0 ;
  assign y9233 = n34307 ;
  assign y9234 = ~n34314 ;
  assign y9235 = ~n34318 ;
  assign y9236 = ~n34321 ;
  assign y9237 = ~n34328 ;
  assign y9238 = ~n34333 ;
  assign y9239 = n34338 ;
  assign y9240 = ~n34339 ;
  assign y9241 = n34340 ;
  assign y9242 = ~1'b0 ;
  assign y9243 = ~1'b0 ;
  assign y9244 = ~n34343 ;
  assign y9245 = ~n34349 ;
  assign y9246 = n34351 ;
  assign y9247 = ~n34354 ;
  assign y9248 = n34360 ;
  assign y9249 = n34361 ;
  assign y9250 = ~1'b0 ;
  assign y9251 = n34366 ;
  assign y9252 = ~n34368 ;
  assign y9253 = n34371 ;
  assign y9254 = ~n34373 ;
  assign y9255 = ~n34374 ;
  assign y9256 = ~n34375 ;
  assign y9257 = ~1'b0 ;
  assign y9258 = ~n34377 ;
  assign y9259 = ~1'b0 ;
  assign y9260 = n34384 ;
  assign y9261 = ~n34390 ;
  assign y9262 = n34392 ;
  assign y9263 = ~1'b0 ;
  assign y9264 = ~1'b0 ;
  assign y9265 = ~1'b0 ;
  assign y9266 = ~n34393 ;
  assign y9267 = n34396 ;
  assign y9268 = n34398 ;
  assign y9269 = ~n34399 ;
  assign y9270 = ~n34407 ;
  assign y9271 = n34409 ;
  assign y9272 = ~n34410 ;
  assign y9273 = n34414 ;
  assign y9274 = ~n34415 ;
  assign y9275 = ~n34418 ;
  assign y9276 = ~n34421 ;
  assign y9277 = n34423 ;
  assign y9278 = ~1'b0 ;
  assign y9279 = ~n34425 ;
  assign y9280 = n34435 ;
  assign y9281 = n34436 ;
  assign y9282 = ~n34438 ;
  assign y9283 = ~1'b0 ;
  assign y9284 = ~1'b0 ;
  assign y9285 = ~n34442 ;
  assign y9286 = n34447 ;
  assign y9287 = ~n34450 ;
  assign y9288 = n34459 ;
  assign y9289 = ~n34464 ;
  assign y9290 = ~n34466 ;
  assign y9291 = ~n34472 ;
  assign y9292 = n34478 ;
  assign y9293 = n34479 ;
  assign y9294 = ~n34482 ;
  assign y9295 = n34483 ;
  assign y9296 = n34485 ;
  assign y9297 = ~n34488 ;
  assign y9298 = ~n34491 ;
  assign y9299 = n34497 ;
  assign y9300 = ~n34501 ;
  assign y9301 = ~n34503 ;
  assign y9302 = n34504 ;
  assign y9303 = ~n34506 ;
  assign y9304 = n34511 ;
  assign y9305 = n34513 ;
  assign y9306 = ~n34517 ;
  assign y9307 = ~1'b0 ;
  assign y9308 = n34518 ;
  assign y9309 = n34519 ;
  assign y9310 = n34520 ;
  assign y9311 = ~n34525 ;
  assign y9312 = n34528 ;
  assign y9313 = ~n34529 ;
  assign y9314 = ~n34533 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = n34535 ;
  assign y9317 = ~n34536 ;
  assign y9318 = ~n34537 ;
  assign y9319 = n34539 ;
  assign y9320 = n34540 ;
  assign y9321 = n34547 ;
  assign y9322 = n34549 ;
  assign y9323 = n34551 ;
  assign y9324 = ~n34552 ;
  assign y9325 = ~n34555 ;
  assign y9326 = n34559 ;
  assign y9327 = ~n34560 ;
  assign y9328 = ~1'b0 ;
  assign y9329 = ~n34562 ;
  assign y9330 = n34565 ;
  assign y9331 = ~n34567 ;
  assign y9332 = n34570 ;
  assign y9333 = ~n34574 ;
  assign y9334 = ~1'b0 ;
  assign y9335 = n34578 ;
  assign y9336 = ~n34579 ;
  assign y9337 = n34584 ;
  assign y9338 = ~n34585 ;
  assign y9339 = ~n34586 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = ~n34588 ;
  assign y9342 = n34589 ;
  assign y9343 = n34591 ;
  assign y9344 = ~n34592 ;
  assign y9345 = n34598 ;
  assign y9346 = ~n34604 ;
  assign y9347 = n34605 ;
  assign y9348 = n34606 ;
  assign y9349 = n34609 ;
  assign y9350 = ~n34611 ;
  assign y9351 = ~1'b0 ;
  assign y9352 = ~n34615 ;
  assign y9353 = ~n34628 ;
  assign y9354 = n34633 ;
  assign y9355 = ~n34635 ;
  assign y9356 = ~n34636 ;
  assign y9357 = ~n34640 ;
  assign y9358 = n34647 ;
  assign y9359 = ~n34650 ;
  assign y9360 = n34651 ;
  assign y9361 = ~n34652 ;
  assign y9362 = n34655 ;
  assign y9363 = ~n34657 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = ~n34659 ;
  assign y9366 = ~n34663 ;
  assign y9367 = ~n34664 ;
  assign y9368 = ~1'b0 ;
  assign y9369 = ~n34668 ;
  assign y9370 = n34671 ;
  assign y9371 = ~n34674 ;
  assign y9372 = n34675 ;
  assign y9373 = n34678 ;
  assign y9374 = n34682 ;
  assign y9375 = n34685 ;
  assign y9376 = ~n34686 ;
  assign y9377 = n34687 ;
  assign y9378 = n34688 ;
  assign y9379 = ~n34689 ;
  assign y9380 = ~n34691 ;
  assign y9381 = ~n34705 ;
  assign y9382 = n34706 ;
  assign y9383 = ~n34710 ;
  assign y9384 = n34713 ;
  assign y9385 = ~n34716 ;
  assign y9386 = ~1'b0 ;
  assign y9387 = n34717 ;
  assign y9388 = n34719 ;
  assign y9389 = ~n34721 ;
  assign y9390 = n14225 ;
  assign y9391 = n34722 ;
  assign y9392 = ~1'b0 ;
  assign y9393 = n34728 ;
  assign y9394 = n34730 ;
  assign y9395 = ~n34734 ;
  assign y9396 = n34735 ;
  assign y9397 = n34737 ;
  assign y9398 = ~n34739 ;
  assign y9399 = ~n24615 ;
  assign y9400 = ~n34744 ;
  assign y9401 = n34746 ;
  assign y9402 = n34748 ;
  assign y9403 = n34752 ;
  assign y9404 = ~n34755 ;
  assign y9405 = ~n34761 ;
  assign y9406 = ~n34764 ;
  assign y9407 = n34766 ;
  assign y9408 = ~n34768 ;
  assign y9409 = n34771 ;
  assign y9410 = n34772 ;
  assign y9411 = ~n34774 ;
  assign y9412 = n34778 ;
  assign y9413 = n34779 ;
  assign y9414 = ~n34783 ;
  assign y9415 = n34784 ;
  assign y9416 = n34789 ;
  assign y9417 = ~1'b0 ;
  assign y9418 = ~n34790 ;
  assign y9419 = ~n34791 ;
  assign y9420 = n34792 ;
  assign y9421 = n34794 ;
  assign y9422 = ~1'b0 ;
  assign y9423 = ~n34795 ;
  assign y9424 = n34796 ;
  assign y9425 = ~n34798 ;
  assign y9426 = ~n34801 ;
  assign y9427 = n34802 ;
  assign y9428 = ~n34803 ;
  assign y9429 = n34804 ;
  assign y9430 = n34811 ;
  assign y9431 = ~1'b0 ;
  assign y9432 = ~n34812 ;
  assign y9433 = ~n34827 ;
  assign y9434 = ~n34831 ;
  assign y9435 = ~n34832 ;
  assign y9436 = n34841 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = ~n34843 ;
  assign y9439 = ~n34844 ;
  assign y9440 = n34845 ;
  assign y9441 = n34850 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = n34852 ;
  assign y9444 = ~n34855 ;
  assign y9445 = ~n34858 ;
  assign y9446 = ~1'b0 ;
  assign y9447 = n34860 ;
  assign y9448 = ~n34868 ;
  assign y9449 = ~n34873 ;
  assign y9450 = n10990 ;
  assign y9451 = ~n34875 ;
  assign y9452 = ~n34879 ;
  assign y9453 = n34881 ;
  assign y9454 = ~n34882 ;
  assign y9455 = ~n34886 ;
  assign y9456 = ~n34888 ;
  assign y9457 = ~n34890 ;
  assign y9458 = ~n34895 ;
  assign y9459 = ~n34900 ;
  assign y9460 = ~n34901 ;
  assign y9461 = n34902 ;
  assign y9462 = ~n34904 ;
  assign y9463 = ~n34906 ;
  assign y9464 = ~n34911 ;
  assign y9465 = ~n34914 ;
  assign y9466 = ~n34921 ;
  assign y9467 = n34923 ;
  assign y9468 = ~n34926 ;
  assign y9469 = n34928 ;
  assign y9470 = n34932 ;
  assign y9471 = ~n34937 ;
  assign y9472 = n34938 ;
  assign y9473 = ~n34942 ;
  assign y9474 = ~n34943 ;
  assign y9475 = ~1'b0 ;
  assign y9476 = n34949 ;
  assign y9477 = n34950 ;
  assign y9478 = n34951 ;
  assign y9479 = ~n34955 ;
  assign y9480 = ~n34957 ;
  assign y9481 = ~1'b0 ;
  assign y9482 = n34959 ;
  assign y9483 = ~n34961 ;
  assign y9484 = ~n34962 ;
  assign y9485 = ~n34965 ;
  assign y9486 = ~n34967 ;
  assign y9487 = ~n34971 ;
  assign y9488 = ~n34981 ;
  assign y9489 = ~n34982 ;
  assign y9490 = n34989 ;
  assign y9491 = ~n34992 ;
  assign y9492 = n34993 ;
  assign y9493 = n34996 ;
  assign y9494 = n34997 ;
  assign y9495 = n34998 ;
  assign y9496 = ~1'b0 ;
  assign y9497 = n35005 ;
  assign y9498 = ~1'b0 ;
  assign y9499 = n35006 ;
  assign y9500 = n35009 ;
  assign y9501 = n35010 ;
  assign y9502 = ~n35012 ;
  assign y9503 = ~n35014 ;
  assign y9504 = ~n35015 ;
  assign y9505 = n35020 ;
  assign y9506 = n35026 ;
  assign y9507 = ~n35028 ;
  assign y9508 = n35030 ;
  assign y9509 = ~n35035 ;
  assign y9510 = n35038 ;
  assign y9511 = ~1'b0 ;
  assign y9512 = ~1'b0 ;
  assign y9513 = ~n35043 ;
  assign y9514 = ~n35047 ;
  assign y9515 = ~n35050 ;
  assign y9516 = ~n35051 ;
  assign y9517 = n35056 ;
  assign y9518 = n35058 ;
  assign y9519 = ~n35061 ;
  assign y9520 = n35066 ;
  assign y9521 = ~n35068 ;
  assign y9522 = n35073 ;
  assign y9523 = ~1'b0 ;
  assign y9524 = ~n35079 ;
  assign y9525 = n35080 ;
  assign y9526 = n35081 ;
  assign y9527 = ~n35085 ;
  assign y9528 = ~n35087 ;
  assign y9529 = ~n35089 ;
  assign y9530 = n35091 ;
  assign y9531 = n35096 ;
  assign y9532 = ~n35097 ;
  assign y9533 = ~n35098 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = ~n35101 ;
  assign y9536 = n35103 ;
  assign y9537 = ~n35108 ;
  assign y9538 = ~n35110 ;
  assign y9539 = ~n35113 ;
  assign y9540 = ~n35121 ;
  assign y9541 = ~n35125 ;
  assign y9542 = ~n35126 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = n35127 ;
  assign y9545 = ~n35128 ;
  assign y9546 = n35129 ;
  assign y9547 = ~n35133 ;
  assign y9548 = n35140 ;
  assign y9549 = ~n35144 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = n35145 ;
  assign y9552 = n35146 ;
  assign y9553 = n35152 ;
  assign y9554 = n35157 ;
  assign y9555 = ~1'b0 ;
  assign y9556 = n35158 ;
  assign y9557 = n35166 ;
  assign y9558 = n35169 ;
  assign y9559 = ~n35172 ;
  assign y9560 = n35173 ;
  assign y9561 = ~n35175 ;
  assign y9562 = n35177 ;
  assign y9563 = ~n35179 ;
  assign y9564 = ~1'b0 ;
  assign y9565 = ~1'b0 ;
  assign y9566 = ~1'b0 ;
  assign y9567 = ~n35180 ;
  assign y9568 = n35182 ;
  assign y9569 = n35198 ;
  assign y9570 = ~n35202 ;
  assign y9571 = ~n35209 ;
  assign y9572 = ~n35210 ;
  assign y9573 = ~n35211 ;
  assign y9574 = n35213 ;
  assign y9575 = ~n1508 ;
  assign y9576 = n35218 ;
  assign y9577 = ~n35220 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = ~n35222 ;
  assign y9580 = n35226 ;
  assign y9581 = ~n35229 ;
  assign y9582 = ~n35235 ;
  assign y9583 = ~n35239 ;
  assign y9584 = ~n35241 ;
  assign y9585 = ~n35242 ;
  assign y9586 = ~n35243 ;
  assign y9587 = ~n35245 ;
  assign y9588 = n35256 ;
  assign y9589 = n35258 ;
  assign y9590 = ~n35260 ;
  assign y9591 = n35262 ;
  assign y9592 = ~n35265 ;
  assign y9593 = n35266 ;
  assign y9594 = n35271 ;
  assign y9595 = n35274 ;
  assign y9596 = ~n35275 ;
  assign y9597 = n35276 ;
  assign y9598 = ~1'b0 ;
  assign y9599 = ~n35279 ;
  assign y9600 = ~n35299 ;
  assign y9601 = n35302 ;
  assign y9602 = n35306 ;
  assign y9603 = ~n35311 ;
  assign y9604 = ~n35314 ;
  assign y9605 = n35318 ;
  assign y9606 = ~n35322 ;
  assign y9607 = ~n35323 ;
  assign y9608 = ~n35326 ;
  assign y9609 = n35327 ;
  assign y9610 = ~n35332 ;
  assign y9611 = ~1'b0 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = ~1'b0 ;
  assign y9614 = n35335 ;
  assign y9615 = ~n35336 ;
  assign y9616 = ~1'b0 ;
  assign y9617 = ~n29958 ;
  assign y9618 = n35339 ;
  assign y9619 = n35344 ;
  assign y9620 = n35345 ;
  assign y9621 = ~1'b0 ;
  assign y9622 = ~n35349 ;
  assign y9623 = n35351 ;
  assign y9624 = n35352 ;
  assign y9625 = ~n35354 ;
  assign y9626 = n35359 ;
  assign y9627 = ~n35365 ;
  assign y9628 = n35366 ;
  assign y9629 = ~n35374 ;
  assign y9630 = ~n35375 ;
  assign y9631 = ~n35376 ;
  assign y9632 = n35380 ;
  assign y9633 = ~n35385 ;
  assign y9634 = ~n35387 ;
  assign y9635 = ~n35391 ;
  assign y9636 = n35392 ;
  assign y9637 = ~n35394 ;
  assign y9638 = n35401 ;
  assign y9639 = ~n35405 ;
  assign y9640 = ~n35406 ;
  assign y9641 = n35407 ;
  assign y9642 = ~n35408 ;
  assign y9643 = ~n35409 ;
  assign y9644 = ~n35414 ;
  assign y9645 = ~n35418 ;
  assign y9646 = ~n35420 ;
  assign y9647 = ~1'b0 ;
  assign y9648 = ~n35423 ;
  assign y9649 = ~n35426 ;
  assign y9650 = ~n35427 ;
  assign y9651 = ~n35429 ;
  assign y9652 = ~n35431 ;
  assign y9653 = ~1'b0 ;
  assign y9654 = n35437 ;
  assign y9655 = ~n35439 ;
  assign y9656 = ~n35442 ;
  assign y9657 = ~n35444 ;
  assign y9658 = ~n35446 ;
  assign y9659 = ~n35450 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~n35451 ;
  assign y9662 = ~n35455 ;
  assign y9663 = n35456 ;
  assign y9664 = n35458 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~n35462 ;
  assign y9667 = ~n35465 ;
  assign y9668 = n35467 ;
  assign y9669 = ~n35470 ;
  assign y9670 = ~n35473 ;
  assign y9671 = n35474 ;
  assign y9672 = n35476 ;
  assign y9673 = ~n35482 ;
  assign y9674 = ~n35486 ;
  assign y9675 = n35490 ;
  assign y9676 = n35491 ;
  assign y9677 = n35493 ;
  assign y9678 = n35495 ;
  assign y9679 = ~n35496 ;
  assign y9680 = ~n35500 ;
  assign y9681 = ~n35505 ;
  assign y9682 = n35507 ;
  assign y9683 = ~n35508 ;
  assign y9684 = n35513 ;
  assign y9685 = ~n35516 ;
  assign y9686 = n35517 ;
  assign y9687 = ~1'b0 ;
  assign y9688 = n35523 ;
  assign y9689 = n35526 ;
  assign y9690 = ~1'b0 ;
  assign y9691 = ~n35528 ;
  assign y9692 = n35529 ;
  assign y9693 = ~n35535 ;
  assign y9694 = ~n35536 ;
  assign y9695 = n35538 ;
  assign y9696 = n35540 ;
  assign y9697 = ~n35541 ;
  assign y9698 = n35546 ;
  assign y9699 = n35548 ;
  assign y9700 = ~n35551 ;
  assign y9701 = ~n35553 ;
  assign y9702 = n35558 ;
  assign y9703 = ~n35559 ;
  assign y9704 = ~n35567 ;
  assign y9705 = ~1'b0 ;
  assign y9706 = ~n35569 ;
  assign y9707 = ~n35571 ;
  assign y9708 = ~n35574 ;
  assign y9709 = n35576 ;
  assign y9710 = n35578 ;
  assign y9711 = n35581 ;
  assign y9712 = ~1'b0 ;
  assign y9713 = ~1'b0 ;
  assign y9714 = ~n35583 ;
  assign y9715 = n35589 ;
  assign y9716 = n35591 ;
  assign y9717 = n35592 ;
  assign y9718 = ~1'b0 ;
  assign y9719 = ~1'b0 ;
  assign y9720 = n35594 ;
  assign y9721 = ~n35596 ;
  assign y9722 = n35597 ;
  assign y9723 = ~n35601 ;
  assign y9724 = ~n35607 ;
  assign y9725 = ~n35608 ;
  assign y9726 = n35609 ;
  assign y9727 = ~n35612 ;
  assign y9728 = n35613 ;
  assign y9729 = n35619 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = ~n35622 ;
  assign y9732 = n35623 ;
  assign y9733 = ~n35628 ;
  assign y9734 = ~n35629 ;
  assign y9735 = n35632 ;
  assign y9736 = n35635 ;
  assign y9737 = n35637 ;
  assign y9738 = ~n35640 ;
  assign y9739 = ~n35642 ;
  assign y9740 = n35654 ;
  assign y9741 = ~1'b0 ;
  assign y9742 = n35656 ;
  assign y9743 = n35658 ;
  assign y9744 = n35660 ;
  assign y9745 = ~n35662 ;
  assign y9746 = n35663 ;
  assign y9747 = ~n35667 ;
  assign y9748 = n35669 ;
  assign y9749 = ~n35673 ;
  assign y9750 = ~n35675 ;
  assign y9751 = n35676 ;
  assign y9752 = ~n35678 ;
  assign y9753 = ~1'b0 ;
  assign y9754 = ~n35684 ;
  assign y9755 = n35690 ;
  assign y9756 = n35692 ;
  assign y9757 = ~n35697 ;
  assign y9758 = ~n35702 ;
  assign y9759 = ~n35703 ;
  assign y9760 = ~n35704 ;
  assign y9761 = ~n35706 ;
  assign y9762 = ~n35707 ;
  assign y9763 = n35708 ;
  assign y9764 = ~n35709 ;
  assign y9765 = n35712 ;
  assign y9766 = ~1'b0 ;
  assign y9767 = ~n35713 ;
  assign y9768 = n35715 ;
  assign y9769 = ~n35722 ;
  assign y9770 = ~n35723 ;
  assign y9771 = n35726 ;
  assign y9772 = ~n35730 ;
  assign y9773 = ~1'b0 ;
  assign y9774 = n35095 ;
  assign y9775 = ~n35736 ;
  assign y9776 = n35739 ;
  assign y9777 = ~n35740 ;
  assign y9778 = n35742 ;
  assign y9779 = ~1'b0 ;
  assign y9780 = ~n35743 ;
  assign y9781 = n35744 ;
  assign y9782 = n35751 ;
  assign y9783 = ~1'b0 ;
  assign y9784 = n35752 ;
  assign y9785 = ~n35754 ;
  assign y9786 = n35760 ;
  assign y9787 = ~n35761 ;
  assign y9788 = ~1'b0 ;
  assign y9789 = ~n35766 ;
  assign y9790 = n35769 ;
  assign y9791 = ~1'b0 ;
  assign y9792 = n35771 ;
  assign y9793 = n35780 ;
  assign y9794 = n35781 ;
  assign y9795 = ~n35785 ;
  assign y9796 = ~n35788 ;
  assign y9797 = n35789 ;
  assign y9798 = ~n35791 ;
  assign y9799 = n35793 ;
  assign y9800 = ~n35795 ;
  assign y9801 = n35798 ;
  assign y9802 = n35805 ;
  assign y9803 = n35808 ;
  assign y9804 = ~n35809 ;
  assign y9805 = n35814 ;
  assign y9806 = n35818 ;
  assign y9807 = n35821 ;
  assign y9808 = ~n35826 ;
  assign y9809 = n35829 ;
  assign y9810 = n35830 ;
  assign y9811 = ~n35832 ;
  assign y9812 = ~n35836 ;
  assign y9813 = n35838 ;
  assign y9814 = n35839 ;
  assign y9815 = n35842 ;
  assign y9816 = ~n35848 ;
  assign y9817 = n35851 ;
  assign y9818 = ~n35855 ;
  assign y9819 = ~n35856 ;
  assign y9820 = n35857 ;
  assign y9821 = n35858 ;
  assign y9822 = n35867 ;
  assign y9823 = ~1'b0 ;
  assign y9824 = ~1'b0 ;
  assign y9825 = ~n35870 ;
  assign y9826 = n35871 ;
  assign y9827 = n35873 ;
  assign y9828 = ~n35876 ;
  assign y9829 = n35880 ;
  assign y9830 = n35882 ;
  assign y9831 = ~n35884 ;
  assign y9832 = ~n35888 ;
  assign y9833 = n35890 ;
  assign y9834 = n35892 ;
  assign y9835 = n35899 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = ~n35906 ;
  assign y9838 = ~n35908 ;
  assign y9839 = n35911 ;
  assign y9840 = n35912 ;
  assign y9841 = n35913 ;
  assign y9842 = ~n35920 ;
  assign y9843 = ~1'b0 ;
  assign y9844 = ~n35922 ;
  assign y9845 = n35924 ;
  assign y9846 = ~n35929 ;
  assign y9847 = ~n35933 ;
  assign y9848 = ~n35934 ;
  assign y9849 = ~n35940 ;
  assign y9850 = ~1'b0 ;
  assign y9851 = ~n35942 ;
  assign y9852 = ~1'b0 ;
  assign y9853 = n35944 ;
  assign y9854 = n35951 ;
  assign y9855 = ~n35952 ;
  assign y9856 = n35957 ;
  assign y9857 = n35958 ;
  assign y9858 = ~n35964 ;
  assign y9859 = ~n35966 ;
  assign y9860 = ~1'b0 ;
  assign y9861 = ~1'b0 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = ~n35967 ;
  assign y9864 = n35968 ;
  assign y9865 = ~1'b0 ;
  assign y9866 = n35972 ;
  assign y9867 = n35974 ;
  assign y9868 = n35978 ;
  assign y9869 = ~1'b0 ;
  assign y9870 = ~1'b0 ;
  assign y9871 = ~n35982 ;
  assign y9872 = n35983 ;
  assign y9873 = ~n35989 ;
  assign y9874 = ~n35992 ;
  assign y9875 = n35996 ;
  assign y9876 = n35997 ;
  assign y9877 = n35998 ;
  assign y9878 = ~n35999 ;
  assign y9879 = ~n36004 ;
  assign y9880 = ~n36006 ;
  assign y9881 = n36009 ;
  assign y9882 = ~n36011 ;
  assign y9883 = ~n36012 ;
  assign y9884 = ~n36013 ;
  assign y9885 = n36016 ;
  assign y9886 = n15825 ;
  assign y9887 = ~n36018 ;
  assign y9888 = n36020 ;
  assign y9889 = ~n36021 ;
  assign y9890 = n36024 ;
  assign y9891 = n36031 ;
  assign y9892 = ~n36034 ;
  assign y9893 = ~1'b0 ;
  assign y9894 = ~n36042 ;
  assign y9895 = n36044 ;
  assign y9896 = ~n36046 ;
  assign y9897 = ~n36048 ;
  assign y9898 = ~1'b0 ;
  assign y9899 = n36049 ;
  assign y9900 = n36055 ;
  assign y9901 = n36058 ;
  assign y9902 = n36060 ;
  assign y9903 = ~n36064 ;
  assign y9904 = ~n36071 ;
  assign y9905 = n36072 ;
  assign y9906 = n36074 ;
  assign y9907 = n36087 ;
  assign y9908 = n36089 ;
  assign y9909 = ~n36093 ;
  assign y9910 = ~n36096 ;
  assign y9911 = ~1'b0 ;
  assign y9912 = ~n36098 ;
  assign y9913 = ~n36100 ;
  assign y9914 = n36103 ;
  assign y9915 = ~n36112 ;
  assign y9916 = n36113 ;
  assign y9917 = n36114 ;
  assign y9918 = ~n36119 ;
  assign y9919 = n36123 ;
  assign y9920 = n36129 ;
  assign y9921 = n36136 ;
  assign y9922 = n36137 ;
  assign y9923 = ~n36138 ;
  assign y9924 = n36141 ;
  assign y9925 = ~n36142 ;
  assign y9926 = n36144 ;
  assign y9927 = ~n36153 ;
  assign y9928 = n36154 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = n36157 ;
  assign y9931 = ~n36158 ;
  assign y9932 = n36160 ;
  assign y9933 = n36162 ;
  assign y9934 = ~n36165 ;
  assign y9935 = n36169 ;
  assign y9936 = n36170 ;
  assign y9937 = ~1'b0 ;
  assign y9938 = n36172 ;
  assign y9939 = n36173 ;
  assign y9940 = ~n36175 ;
  assign y9941 = n36177 ;
  assign y9942 = n36178 ;
  assign y9943 = n36180 ;
  assign y9944 = ~n36183 ;
  assign y9945 = ~n36185 ;
  assign y9946 = n36190 ;
  assign y9947 = n36193 ;
  assign y9948 = ~n36194 ;
  assign y9949 = n36195 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = n36198 ;
  assign y9952 = n36199 ;
  assign y9953 = ~n36200 ;
  assign y9954 = ~n36201 ;
  assign y9955 = n36203 ;
  assign y9956 = n36204 ;
  assign y9957 = ~n36206 ;
  assign y9958 = n36207 ;
  assign y9959 = ~1'b0 ;
  assign y9960 = ~1'b0 ;
  assign y9961 = n36210 ;
  assign y9962 = n25347 ;
  assign y9963 = n36211 ;
  assign y9964 = ~1'b0 ;
  assign y9965 = ~n36214 ;
  assign y9966 = ~n36216 ;
  assign y9967 = n36217 ;
  assign y9968 = ~n36219 ;
  assign y9969 = n36221 ;
  assign y9970 = n36222 ;
  assign y9971 = n36225 ;
  assign y9972 = n36226 ;
  assign y9973 = ~n36227 ;
  assign y9974 = n36230 ;
  assign y9975 = ~n36231 ;
  assign y9976 = ~n36235 ;
  assign y9977 = n36241 ;
  assign y9978 = ~n36243 ;
  assign y9979 = ~n36251 ;
  assign y9980 = ~n36253 ;
  assign y9981 = ~n36256 ;
  assign y9982 = n36263 ;
  assign y9983 = n36264 ;
  assign y9984 = n36266 ;
  assign y9985 = n36270 ;
  assign y9986 = ~1'b0 ;
  assign y9987 = ~n36272 ;
  assign y9988 = ~n36275 ;
  assign y9989 = n36276 ;
  assign y9990 = ~1'b0 ;
  assign y9991 = n36279 ;
  assign y9992 = ~n36280 ;
  assign y9993 = n36282 ;
  assign y9994 = ~n36283 ;
  assign y9995 = ~n36285 ;
  assign y9996 = n36286 ;
  assign y9997 = ~n36290 ;
  assign y9998 = ~n36292 ;
  assign y9999 = ~1'b0 ;
  assign y10000 = n36298 ;
  assign y10001 = n36307 ;
  assign y10002 = ~n36309 ;
  assign y10003 = n36314 ;
  assign y10004 = ~n36320 ;
  assign y10005 = n36324 ;
  assign y10006 = n36328 ;
  assign y10007 = n36331 ;
  assign y10008 = ~n36332 ;
  assign y10009 = n36338 ;
  assign y10010 = ~n36342 ;
  assign y10011 = ~n36344 ;
  assign y10012 = ~n36346 ;
  assign y10013 = ~n36347 ;
  assign y10014 = n36350 ;
  assign y10015 = ~n36351 ;
  assign y10016 = ~n36354 ;
  assign y10017 = ~n36355 ;
  assign y10018 = n36359 ;
  assign y10019 = ~n36364 ;
  assign y10020 = n36367 ;
  assign y10021 = n36372 ;
  assign y10022 = n36377 ;
  assign y10023 = n36381 ;
  assign y10024 = ~n36382 ;
  assign y10025 = ~1'b0 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = n36384 ;
  assign y10028 = n36385 ;
  assign y10029 = ~n36386 ;
  assign y10030 = ~n36388 ;
  assign y10031 = n36389 ;
  assign y10032 = ~n36390 ;
  assign y10033 = ~1'b0 ;
  assign y10034 = n36394 ;
  assign y10035 = n36396 ;
  assign y10036 = n36397 ;
  assign y10037 = ~n36400 ;
  assign y10038 = ~1'b0 ;
  assign y10039 = ~n36406 ;
  assign y10040 = n36407 ;
  assign y10041 = n36408 ;
  assign y10042 = ~n36409 ;
  assign y10043 = ~n36410 ;
  assign y10044 = n36419 ;
  assign y10045 = n36421 ;
  assign y10046 = n36424 ;
  assign y10047 = ~n36427 ;
  assign y10048 = ~n36432 ;
  assign y10049 = ~n36434 ;
  assign y10050 = n36435 ;
  assign y10051 = ~n36436 ;
  assign y10052 = ~n36437 ;
  assign y10053 = ~1'b0 ;
  assign y10054 = ~n36438 ;
  assign y10055 = ~n36439 ;
  assign y10056 = n36441 ;
  assign y10057 = n36443 ;
  assign y10058 = ~n36449 ;
  assign y10059 = ~n36450 ;
  assign y10060 = ~n36453 ;
  assign y10061 = n36456 ;
  assign y10062 = ~n11158 ;
  assign y10063 = n36458 ;
  assign y10064 = ~n36464 ;
  assign y10065 = ~n36466 ;
  assign y10066 = n36467 ;
  assign y10067 = n36468 ;
  assign y10068 = ~n36472 ;
  assign y10069 = n36473 ;
  assign y10070 = ~n36475 ;
  assign y10071 = ~n36476 ;
  assign y10072 = ~n36477 ;
  assign y10073 = n36478 ;
  assign y10074 = ~1'b0 ;
  assign y10075 = ~1'b0 ;
  assign y10076 = ~n36479 ;
  assign y10077 = n36482 ;
  assign y10078 = ~n36483 ;
  assign y10079 = n36484 ;
  assign y10080 = ~n36489 ;
  assign y10081 = ~n36494 ;
  assign y10082 = ~n36498 ;
  assign y10083 = ~n36502 ;
  assign y10084 = n36506 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = ~n36508 ;
  assign y10087 = ~n36516 ;
  assign y10088 = n36518 ;
  assign y10089 = ~n36523 ;
  assign y10090 = n36526 ;
  assign y10091 = n36534 ;
  assign y10092 = ~n36535 ;
  assign y10093 = ~n36537 ;
  assign y10094 = n36541 ;
  assign y10095 = n36543 ;
  assign y10096 = n36544 ;
  assign y10097 = n36551 ;
  assign y10098 = ~n36554 ;
  assign y10099 = ~1'b0 ;
  assign y10100 = n36558 ;
  assign y10101 = ~1'b0 ;
  assign y10102 = n36563 ;
  assign y10103 = n36564 ;
  assign y10104 = n36565 ;
  assign y10105 = n36566 ;
  assign y10106 = ~1'b0 ;
  assign y10107 = n36568 ;
  assign y10108 = ~n36569 ;
  assign y10109 = ~n36572 ;
  assign y10110 = n36576 ;
  assign y10111 = n36577 ;
  assign y10112 = n36580 ;
  assign y10113 = n36586 ;
  assign y10114 = ~n36589 ;
  assign y10115 = ~n36597 ;
  assign y10116 = n36599 ;
  assign y10117 = ~n36602 ;
  assign y10118 = n36605 ;
  assign y10119 = ~1'b0 ;
  assign y10120 = ~n36607 ;
  assign y10121 = ~1'b0 ;
  assign y10122 = n36609 ;
  assign y10123 = n36610 ;
  assign y10124 = n36612 ;
  assign y10125 = n36613 ;
  assign y10126 = n36616 ;
  assign y10127 = ~n36617 ;
  assign y10128 = ~n36619 ;
  assign y10129 = n36627 ;
  assign y10130 = n36628 ;
  assign y10131 = ~n36629 ;
  assign y10132 = n26194 ;
  assign y10133 = n36630 ;
  assign y10134 = ~n36631 ;
  assign y10135 = n36635 ;
  assign y10136 = n36636 ;
  assign y10137 = ~n36638 ;
  assign y10138 = ~n36640 ;
  assign y10139 = n36641 ;
  assign y10140 = n36643 ;
  assign y10141 = n36654 ;
  assign y10142 = ~n36655 ;
  assign y10143 = ~n36659 ;
  assign y10144 = ~n36662 ;
  assign y10145 = n36666 ;
  assign y10146 = ~n36667 ;
  assign y10147 = ~n36671 ;
  assign y10148 = ~n36672 ;
  assign y10149 = ~n36674 ;
  assign y10150 = ~1'b0 ;
  assign y10151 = ~n36679 ;
  assign y10152 = n36686 ;
  assign y10153 = ~n36694 ;
  assign y10154 = ~n36696 ;
  assign y10155 = n36697 ;
  assign y10156 = n36698 ;
  assign y10157 = ~n36701 ;
  assign y10158 = n36707 ;
  assign y10159 = ~n36708 ;
  assign y10160 = n36709 ;
  assign y10161 = n36712 ;
  assign y10162 = n36718 ;
  assign y10163 = ~n36720 ;
  assign y10164 = n36721 ;
  assign y10165 = ~n36723 ;
  assign y10166 = n36726 ;
  assign y10167 = ~1'b0 ;
  assign y10168 = ~1'b0 ;
  assign y10169 = n36731 ;
  assign y10170 = n36732 ;
  assign y10171 = n36735 ;
  assign y10172 = n36740 ;
  assign y10173 = n36741 ;
  assign y10174 = ~n36743 ;
  assign y10175 = ~n36745 ;
  assign y10176 = n36748 ;
  assign y10177 = n36749 ;
  assign y10178 = n36752 ;
  assign y10179 = n36754 ;
  assign y10180 = ~n36755 ;
  assign y10181 = n36756 ;
  assign y10182 = ~n36761 ;
  assign y10183 = n36763 ;
  assign y10184 = ~n36767 ;
  assign y10185 = ~n36770 ;
  assign y10186 = ~1'b0 ;
  assign y10187 = n36775 ;
  assign y10188 = n36777 ;
  assign y10189 = n36779 ;
  assign y10190 = ~n36782 ;
  assign y10191 = n36785 ;
  assign y10192 = n36791 ;
  assign y10193 = n36792 ;
  assign y10194 = ~n36795 ;
  assign y10195 = ~n36796 ;
  assign y10196 = n36800 ;
  assign y10197 = n36803 ;
  assign y10198 = ~n36807 ;
  assign y10199 = ~n36810 ;
  assign y10200 = ~1'b0 ;
  assign y10201 = n36811 ;
  assign y10202 = n36813 ;
  assign y10203 = n36815 ;
  assign y10204 = n36816 ;
  assign y10205 = ~n36818 ;
  assign y10206 = ~n36820 ;
  assign y10207 = n36822 ;
  assign y10208 = n36824 ;
  assign y10209 = ~n36825 ;
  assign y10210 = n36829 ;
  assign y10211 = ~n36831 ;
  assign y10212 = n36833 ;
  assign y10213 = n36837 ;
  assign y10214 = ~n36841 ;
  assign y10215 = n36842 ;
  assign y10216 = n36843 ;
  assign y10217 = ~n36844 ;
  assign y10218 = n36845 ;
  assign y10219 = n36852 ;
  assign y10220 = ~1'b0 ;
  assign y10221 = ~n36854 ;
  assign y10222 = n36856 ;
  assign y10223 = ~n36858 ;
  assign y10224 = ~n36861 ;
  assign y10225 = ~n36862 ;
  assign y10226 = ~n36864 ;
  assign y10227 = ~n36869 ;
  assign y10228 = n36873 ;
  assign y10229 = ~n36880 ;
  assign y10230 = n36881 ;
  assign y10231 = n36884 ;
  assign y10232 = ~n36893 ;
  assign y10233 = ~n36894 ;
  assign y10234 = ~n36895 ;
  assign y10235 = ~n36897 ;
  assign y10236 = n36899 ;
  assign y10237 = n36901 ;
  assign y10238 = n36903 ;
  assign y10239 = n36905 ;
  assign y10240 = n16111 ;
  assign y10241 = n36907 ;
  assign y10242 = ~1'b0 ;
  assign y10243 = ~n36908 ;
  assign y10244 = n36909 ;
  assign y10245 = ~n36910 ;
  assign y10246 = ~1'b0 ;
  assign y10247 = ~1'b0 ;
  assign y10248 = n32499 ;
  assign y10249 = n36913 ;
  assign y10250 = n36914 ;
  assign y10251 = n36917 ;
  assign y10252 = n36921 ;
  assign y10253 = ~n36923 ;
  assign y10254 = ~n36925 ;
  assign y10255 = ~n36930 ;
  assign y10256 = ~n36933 ;
  assign y10257 = ~1'b0 ;
  assign y10258 = ~1'b0 ;
  assign y10259 = n36935 ;
  assign y10260 = n36938 ;
  assign y10261 = n36939 ;
  assign y10262 = ~n36940 ;
  assign y10263 = n36941 ;
  assign y10264 = ~n36942 ;
  assign y10265 = n36944 ;
  assign y10266 = ~n36948 ;
  assign y10267 = n36949 ;
  assign y10268 = n36953 ;
  assign y10269 = ~n36958 ;
  assign y10270 = ~n36959 ;
  assign y10271 = n36962 ;
  assign y10272 = n36965 ;
  assign y10273 = ~n36966 ;
  assign y10274 = ~n36969 ;
  assign y10275 = ~n36972 ;
  assign y10276 = n36973 ;
  assign y10277 = n36976 ;
  assign y10278 = ~n36980 ;
  assign y10279 = ~n36983 ;
  assign y10280 = n36986 ;
  assign y10281 = n36989 ;
  assign y10282 = ~n36997 ;
  assign y10283 = ~n37003 ;
  assign y10284 = n37009 ;
  assign y10285 = ~1'b0 ;
  assign y10286 = n37014 ;
  assign y10287 = n37015 ;
  assign y10288 = ~n37016 ;
  assign y10289 = n37021 ;
  assign y10290 = ~n37026 ;
  assign y10291 = ~n37028 ;
  assign y10292 = ~n37029 ;
  assign y10293 = ~n37030 ;
  assign y10294 = n37033 ;
  assign y10295 = ~n37035 ;
  assign y10296 = n37045 ;
  assign y10297 = ~n37047 ;
  assign y10298 = ~1'b0 ;
  assign y10299 = ~n37054 ;
  assign y10300 = n37056 ;
  assign y10301 = ~n37059 ;
  assign y10302 = n37068 ;
  assign y10303 = ~n37070 ;
  assign y10304 = n37072 ;
  assign y10305 = ~n37077 ;
  assign y10306 = n37078 ;
  assign y10307 = n37081 ;
  assign y10308 = ~n37084 ;
  assign y10309 = ~n37085 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = ~n37087 ;
  assign y10312 = ~n37091 ;
  assign y10313 = n37095 ;
  assign y10314 = n37097 ;
  assign y10315 = ~n37098 ;
  assign y10316 = ~n37099 ;
  assign y10317 = ~n37100 ;
  assign y10318 = ~n37101 ;
  assign y10319 = n37105 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = ~1'b0 ;
  assign y10322 = ~n37109 ;
  assign y10323 = ~n37110 ;
  assign y10324 = ~n37114 ;
  assign y10325 = n37115 ;
  assign y10326 = n37117 ;
  assign y10327 = ~1'b0 ;
  assign y10328 = ~n37119 ;
  assign y10329 = ~n37126 ;
  assign y10330 = n37127 ;
  assign y10331 = ~n37130 ;
  assign y10332 = n37132 ;
  assign y10333 = ~n37133 ;
  assign y10334 = ~1'b0 ;
  assign y10335 = ~n37134 ;
  assign y10336 = ~n37135 ;
  assign y10337 = n32921 ;
  assign y10338 = n37139 ;
  assign y10339 = n37145 ;
  assign y10340 = n37149 ;
  assign y10341 = n37159 ;
  assign y10342 = n37161 ;
  assign y10343 = n37162 ;
  assign y10344 = n37164 ;
  assign y10345 = ~1'b0 ;
  assign y10346 = n37169 ;
  assign y10347 = n37170 ;
  assign y10348 = n37174 ;
  assign y10349 = n37177 ;
  assign y10350 = ~n37178 ;
  assign y10351 = ~n37181 ;
  assign y10352 = ~n37185 ;
  assign y10353 = ~n37187 ;
  assign y10354 = n37188 ;
  assign y10355 = n37189 ;
  assign y10356 = ~n37190 ;
  assign y10357 = ~n37193 ;
  assign y10358 = ~n37198 ;
  assign y10359 = ~n37206 ;
  assign y10360 = ~n37209 ;
  assign y10361 = ~n16567 ;
  assign y10362 = n37210 ;
  assign y10363 = n37211 ;
  assign y10364 = ~n37214 ;
  assign y10365 = ~1'b0 ;
  assign y10366 = n37216 ;
  assign y10367 = ~n37217 ;
  assign y10368 = ~n37221 ;
  assign y10369 = ~n37222 ;
  assign y10370 = ~n37223 ;
  assign y10371 = ~n37224 ;
  assign y10372 = ~1'b0 ;
  assign y10373 = ~n37225 ;
  assign y10374 = ~n37229 ;
  assign y10375 = n37234 ;
  assign y10376 = ~n37235 ;
  assign y10377 = ~n37237 ;
  assign y10378 = n37239 ;
  assign y10379 = n37240 ;
  assign y10380 = ~n37241 ;
  assign y10381 = ~n37244 ;
  assign y10382 = ~n37251 ;
  assign y10383 = n37257 ;
  assign y10384 = n37260 ;
  assign y10385 = ~n37270 ;
  assign y10386 = n37272 ;
  assign y10387 = ~n37274 ;
  assign y10388 = ~n37281 ;
  assign y10389 = ~n37282 ;
  assign y10390 = n37283 ;
  assign y10391 = n37286 ;
  assign y10392 = n37287 ;
  assign y10393 = ~n37289 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = n37294 ;
  assign y10396 = n37297 ;
  assign y10397 = n37300 ;
  assign y10398 = n37301 ;
  assign y10399 = ~n37312 ;
  assign y10400 = n37314 ;
  assign y10401 = n37318 ;
  assign y10402 = n37322 ;
  assign y10403 = ~n37328 ;
  assign y10404 = ~n37329 ;
  assign y10405 = ~n37331 ;
  assign y10406 = n37333 ;
  assign y10407 = ~n37336 ;
  assign y10408 = ~n37338 ;
  assign y10409 = n37339 ;
  assign y10410 = n37340 ;
  assign y10411 = ~n37345 ;
  assign y10412 = n37346 ;
  assign y10413 = n37348 ;
  assign y10414 = ~1'b0 ;
  assign y10415 = ~n37352 ;
  assign y10416 = ~n37354 ;
  assign y10417 = ~1'b0 ;
  assign y10418 = n37355 ;
  assign y10419 = ~n37361 ;
  assign y10420 = n37363 ;
  assign y10421 = n37366 ;
  assign y10422 = n37368 ;
  assign y10423 = ~1'b0 ;
  assign y10424 = ~n37375 ;
  assign y10425 = n37383 ;
  assign y10426 = n37389 ;
  assign y10427 = n37390 ;
  assign y10428 = ~n37393 ;
  assign y10429 = ~n37395 ;
  assign y10430 = ~1'b0 ;
  assign y10431 = n37398 ;
  assign y10432 = ~n37399 ;
  assign y10433 = ~n37400 ;
  assign y10434 = ~n37404 ;
  assign y10435 = n37405 ;
  assign y10436 = ~n37408 ;
  assign y10437 = ~n37409 ;
  assign y10438 = ~n37411 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = ~n37412 ;
  assign y10441 = ~n37413 ;
  assign y10442 = ~n37416 ;
  assign y10443 = n37417 ;
  assign y10444 = ~n37420 ;
  assign y10445 = ~n37425 ;
  assign y10446 = n37427 ;
  assign y10447 = ~n37429 ;
  assign y10448 = ~n37431 ;
  assign y10449 = ~n37433 ;
  assign y10450 = n37434 ;
  assign y10451 = ~1'b0 ;
  assign y10452 = ~n37440 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = n37441 ;
  assign y10455 = ~n37442 ;
  assign y10456 = ~n37448 ;
  assign y10457 = n37450 ;
  assign y10458 = ~n37451 ;
  assign y10459 = ~n37452 ;
  assign y10460 = ~n37453 ;
  assign y10461 = n37454 ;
  assign y10462 = n37456 ;
  assign y10463 = ~1'b0 ;
  assign y10464 = ~n37457 ;
  assign y10465 = ~n37460 ;
  assign y10466 = ~n37463 ;
  assign y10467 = n37464 ;
  assign y10468 = n37467 ;
  assign y10469 = ~n37468 ;
  assign y10470 = ~n37469 ;
  assign y10471 = ~n37471 ;
  assign y10472 = ~n37473 ;
  assign y10473 = ~1'b0 ;
  assign y10474 = n37477 ;
  assign y10475 = n37479 ;
  assign y10476 = n37487 ;
  assign y10477 = ~n37490 ;
  assign y10478 = ~n37491 ;
  assign y10479 = ~n37493 ;
  assign y10480 = n37494 ;
  assign y10481 = ~1'b0 ;
  assign y10482 = ~n37500 ;
  assign y10483 = ~n37501 ;
  assign y10484 = n37503 ;
  assign y10485 = ~n37504 ;
  assign y10486 = ~1'b0 ;
  assign y10487 = ~n37506 ;
  assign y10488 = ~1'b0 ;
  assign y10489 = ~n37507 ;
  assign y10490 = ~n37510 ;
  assign y10491 = n37512 ;
  assign y10492 = n37516 ;
  assign y10493 = n37520 ;
  assign y10494 = ~1'b0 ;
  assign y10495 = ~n37523 ;
  assign y10496 = ~n37525 ;
  assign y10497 = n37528 ;
  assign y10498 = ~n37531 ;
  assign y10499 = n37532 ;
  assign y10500 = n37535 ;
  assign y10501 = n37537 ;
  assign y10502 = ~n37539 ;
  assign y10503 = ~1'b0 ;
  assign y10504 = ~n37546 ;
  assign y10505 = ~1'b0 ;
  assign y10506 = n37554 ;
  assign y10507 = n37555 ;
  assign y10508 = ~n37564 ;
  assign y10509 = n37565 ;
  assign y10510 = n37567 ;
  assign y10511 = ~n37576 ;
  assign y10512 = ~n37581 ;
  assign y10513 = ~n37586 ;
  assign y10514 = n37588 ;
  assign y10515 = n37591 ;
  assign y10516 = ~n37593 ;
  assign y10517 = ~n37594 ;
  assign y10518 = n37599 ;
  assign y10519 = ~n37601 ;
  assign y10520 = n37602 ;
  assign y10521 = n37603 ;
  assign y10522 = n37604 ;
  assign y10523 = ~n37606 ;
  assign y10524 = n37608 ;
  assign y10525 = n37617 ;
  assign y10526 = ~1'b0 ;
  assign y10527 = ~1'b0 ;
  assign y10528 = ~n37619 ;
  assign y10529 = n37625 ;
  assign y10530 = n37627 ;
  assign y10531 = ~n13761 ;
  assign y10532 = ~n37628 ;
  assign y10533 = n37629 ;
  assign y10534 = n37630 ;
  assign y10535 = ~n37631 ;
  assign y10536 = n37632 ;
  assign y10537 = ~n37633 ;
  assign y10538 = ~n37634 ;
  assign y10539 = ~n37651 ;
  assign y10540 = ~n37654 ;
  assign y10541 = ~n37655 ;
  assign y10542 = n37659 ;
  assign y10543 = ~n37662 ;
  assign y10544 = ~n37663 ;
  assign y10545 = n37664 ;
  assign y10546 = n37665 ;
  assign y10547 = ~n37674 ;
  assign y10548 = ~n37676 ;
  assign y10549 = n37680 ;
  assign y10550 = ~n37682 ;
  assign y10551 = ~1'b0 ;
  assign y10552 = ~n37684 ;
  assign y10553 = n37689 ;
  assign y10554 = ~n37694 ;
  assign y10555 = ~n37697 ;
  assign y10556 = ~n37699 ;
  assign y10557 = ~n37700 ;
  assign y10558 = n37702 ;
  assign y10559 = ~1'b0 ;
  assign y10560 = n37711 ;
  assign y10561 = n37713 ;
  assign y10562 = ~n37714 ;
  assign y10563 = n37716 ;
  assign y10564 = ~n37720 ;
  assign y10565 = n37721 ;
  assign y10566 = n37728 ;
  assign y10567 = n37729 ;
  assign y10568 = ~n37733 ;
  assign y10569 = n37735 ;
  assign y10570 = n37741 ;
  assign y10571 = n37742 ;
  assign y10572 = ~n37744 ;
  assign y10573 = ~n37749 ;
  assign y10574 = ~1'b0 ;
  assign y10575 = ~n37751 ;
  assign y10576 = n37752 ;
  assign y10577 = ~n37754 ;
  assign y10578 = ~n37756 ;
  assign y10579 = ~n37757 ;
  assign y10580 = n37764 ;
  assign y10581 = ~1'b0 ;
  assign y10582 = ~n37774 ;
  assign y10583 = n37775 ;
  assign y10584 = ~n37778 ;
  assign y10585 = ~n37780 ;
  assign y10586 = ~n37782 ;
  assign y10587 = ~1'b0 ;
  assign y10588 = ~n37783 ;
  assign y10589 = n37787 ;
  assign y10590 = ~n37792 ;
  assign y10591 = ~n37796 ;
  assign y10592 = n37801 ;
  assign y10593 = n37812 ;
  assign y10594 = n37813 ;
  assign y10595 = ~n37815 ;
  assign y10596 = n37819 ;
  assign y10597 = ~1'b0 ;
  assign y10598 = ~n37823 ;
  assign y10599 = n6589 ;
  assign y10600 = ~n37825 ;
  assign y10601 = ~n37826 ;
  assign y10602 = n37829 ;
  assign y10603 = ~n37834 ;
  assign y10604 = ~n37835 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = ~1'b0 ;
  assign y10607 = ~n37837 ;
  assign y10608 = n37840 ;
  assign y10609 = ~n37842 ;
  assign y10610 = ~n37843 ;
  assign y10611 = ~n37846 ;
  assign y10612 = n1827 ;
  assign y10613 = n37848 ;
  assign y10614 = ~n37854 ;
  assign y10615 = n37865 ;
  assign y10616 = ~n37866 ;
  assign y10617 = n37869 ;
  assign y10618 = ~n37870 ;
  assign y10619 = ~n37873 ;
  assign y10620 = n37880 ;
  assign y10621 = n3804 ;
  assign y10622 = n37882 ;
  assign y10623 = n37886 ;
  assign y10624 = ~n37891 ;
  assign y10625 = n37893 ;
  assign y10626 = n37898 ;
  assign y10627 = n37902 ;
  assign y10628 = n37903 ;
  assign y10629 = ~1'b0 ;
  assign y10630 = n37915 ;
  assign y10631 = ~n37918 ;
  assign y10632 = n37928 ;
  assign y10633 = ~n37934 ;
  assign y10634 = ~1'b0 ;
  assign y10635 = ~n37936 ;
  assign y10636 = n37937 ;
  assign y10637 = n37940 ;
  assign y10638 = ~n37944 ;
  assign y10639 = ~n37945 ;
  assign y10640 = ~n37947 ;
  assign y10641 = ~n37948 ;
  assign y10642 = n37950 ;
  assign y10643 = n37951 ;
  assign y10644 = ~n37956 ;
  assign y10645 = n37958 ;
  assign y10646 = n37959 ;
  assign y10647 = ~n37960 ;
  assign y10648 = n37964 ;
  assign y10649 = ~n37967 ;
  assign y10650 = n37968 ;
  assign y10651 = ~n37971 ;
  assign y10652 = n37973 ;
  assign y10653 = ~n37976 ;
  assign y10654 = ~n37981 ;
  assign y10655 = ~n37982 ;
  assign y10656 = n37985 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = ~n37990 ;
  assign y10659 = ~n37992 ;
  assign y10660 = ~n37994 ;
  assign y10661 = n37996 ;
  assign y10662 = n37997 ;
  assign y10663 = n38002 ;
  assign y10664 = ~n38003 ;
  assign y10665 = ~n38007 ;
  assign y10666 = ~1'b0 ;
  assign y10667 = n38009 ;
  assign y10668 = n38010 ;
  assign y10669 = ~n38011 ;
  assign y10670 = ~1'b0 ;
  assign y10671 = n38013 ;
  assign y10672 = n38016 ;
  assign y10673 = ~n38019 ;
  assign y10674 = n38021 ;
  assign y10675 = ~n38024 ;
  assign y10676 = ~n38029 ;
  assign y10677 = ~1'b0 ;
  assign y10678 = ~n38032 ;
  assign y10679 = n38033 ;
  assign y10680 = n38039 ;
  assign y10681 = ~n38040 ;
  assign y10682 = ~n38041 ;
  assign y10683 = ~n38044 ;
  assign y10684 = n38048 ;
  assign y10685 = n38049 ;
  assign y10686 = ~n38050 ;
  assign y10687 = ~1'b0 ;
  assign y10688 = ~n11983 ;
  assign y10689 = ~1'b0 ;
  assign y10690 = ~1'b0 ;
  assign y10691 = ~n38052 ;
  assign y10692 = n38054 ;
  assign y10693 = n38055 ;
  assign y10694 = ~n38058 ;
  assign y10695 = ~n38060 ;
  assign y10696 = n38064 ;
  assign y10697 = ~n38065 ;
  assign y10698 = ~n38067 ;
  assign y10699 = ~1'b0 ;
  assign y10700 = n38070 ;
  assign y10701 = n38071 ;
  assign y10702 = ~n38073 ;
  assign y10703 = n38079 ;
  assign y10704 = ~n38081 ;
  assign y10705 = ~n38082 ;
  assign y10706 = ~n38083 ;
  assign y10707 = n38084 ;
  assign y10708 = ~n38091 ;
  assign y10709 = ~n38093 ;
  assign y10710 = ~n38097 ;
  assign y10711 = ~n38099 ;
  assign y10712 = ~n38103 ;
  assign y10713 = ~n38105 ;
  assign y10714 = ~1'b0 ;
  assign y10715 = ~n38106 ;
  assign y10716 = ~n38110 ;
  assign y10717 = ~n38113 ;
  assign y10718 = ~n38116 ;
  assign y10719 = ~n38121 ;
  assign y10720 = n9355 ;
  assign y10721 = n38123 ;
  assign y10722 = ~1'b0 ;
  assign y10723 = ~1'b0 ;
  assign y10724 = ~1'b0 ;
  assign y10725 = ~n38124 ;
  assign y10726 = ~n38125 ;
  assign y10727 = ~n38127 ;
  assign y10728 = n38134 ;
  assign y10729 = ~1'b0 ;
  assign y10730 = n38139 ;
  assign y10731 = ~n38140 ;
  assign y10732 = n38142 ;
  assign y10733 = n38147 ;
  assign y10734 = ~1'b0 ;
  assign y10735 = n38151 ;
  assign y10736 = ~n38152 ;
  assign y10737 = ~n38156 ;
  assign y10738 = ~n38157 ;
  assign y10739 = ~n38161 ;
  assign y10740 = n38163 ;
  assign y10741 = n38164 ;
  assign y10742 = n38167 ;
  assign y10743 = ~n38168 ;
  assign y10744 = ~n38173 ;
  assign y10745 = ~n38177 ;
  assign y10746 = n38178 ;
  assign y10747 = n38182 ;
  assign y10748 = ~n38184 ;
  assign y10749 = n38186 ;
  assign y10750 = ~n38188 ;
  assign y10751 = ~n38190 ;
  assign y10752 = ~1'b0 ;
  assign y10753 = n38191 ;
  assign y10754 = n38192 ;
  assign y10755 = n38203 ;
  assign y10756 = n38205 ;
  assign y10757 = n38206 ;
  assign y10758 = n38207 ;
  assign y10759 = n38210 ;
  assign y10760 = ~n38211 ;
  assign y10761 = n38214 ;
  assign y10762 = ~n38223 ;
  assign y10763 = n38231 ;
  assign y10764 = ~1'b0 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = n38233 ;
  assign y10767 = ~n38235 ;
  assign y10768 = n38237 ;
  assign y10769 = ~n38240 ;
  assign y10770 = ~n38243 ;
  assign y10771 = n38244 ;
  assign y10772 = ~n38246 ;
  assign y10773 = ~n38249 ;
  assign y10774 = n38250 ;
  assign y10775 = ~n38251 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = n38253 ;
  assign y10778 = n38254 ;
  assign y10779 = n38256 ;
  assign y10780 = ~n38258 ;
  assign y10781 = ~n38263 ;
  assign y10782 = n38265 ;
  assign y10783 = ~1'b0 ;
  assign y10784 = ~n38268 ;
  assign y10785 = ~n38271 ;
  assign y10786 = n38273 ;
  assign y10787 = n38278 ;
  assign y10788 = ~n38280 ;
  assign y10789 = ~n38285 ;
  assign y10790 = n38288 ;
  assign y10791 = ~n38291 ;
  assign y10792 = ~n38296 ;
  assign y10793 = ~n38300 ;
  assign y10794 = ~n38301 ;
  assign y10795 = n38303 ;
  assign y10796 = ~n630 ;
  assign y10797 = n38305 ;
  assign y10798 = ~n38313 ;
  assign y10799 = n38315 ;
  assign y10800 = 1'b0 ;
  assign y10801 = ~n38316 ;
  assign y10802 = n38319 ;
  assign y10803 = ~1'b0 ;
  assign y10804 = n38323 ;
  assign y10805 = n38324 ;
  assign y10806 = n38325 ;
  assign y10807 = ~n38328 ;
  assign y10808 = ~n38331 ;
  assign y10809 = ~n38333 ;
  assign y10810 = n38334 ;
  assign y10811 = n38335 ;
  assign y10812 = n38338 ;
  assign y10813 = ~n38339 ;
  assign y10814 = n38342 ;
  assign y10815 = n38343 ;
  assign y10816 = ~1'b0 ;
  assign y10817 = ~n38346 ;
  assign y10818 = ~1'b0 ;
  assign y10819 = ~n38352 ;
  assign y10820 = ~n38354 ;
  assign y10821 = n38357 ;
  assign y10822 = ~n38364 ;
  assign y10823 = n38366 ;
  assign y10824 = ~n38367 ;
  assign y10825 = n38368 ;
  assign y10826 = n38369 ;
  assign y10827 = n38372 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = n38374 ;
  assign y10830 = n38378 ;
  assign y10831 = n38379 ;
  assign y10832 = n38385 ;
  assign y10833 = n38389 ;
  assign y10834 = ~n38393 ;
  assign y10835 = ~n38396 ;
  assign y10836 = n38398 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = ~n38399 ;
  assign y10840 = n38403 ;
  assign y10841 = ~n38404 ;
  assign y10842 = ~n38405 ;
  assign y10843 = ~n38406 ;
  assign y10844 = ~1'b0 ;
  assign y10845 = ~n38409 ;
  assign y10846 = ~n38410 ;
  assign y10847 = n38411 ;
  assign y10848 = ~n38420 ;
  assign y10849 = ~n38421 ;
  assign y10850 = n38424 ;
  assign y10851 = ~n38425 ;
  assign y10852 = ~1'b0 ;
  assign y10853 = ~n38427 ;
  assign y10854 = n38431 ;
  assign y10855 = n38438 ;
  assign y10856 = n38439 ;
  assign y10857 = ~n38447 ;
  assign y10858 = ~n38453 ;
  assign y10859 = ~1'b0 ;
  assign y10860 = n38458 ;
  assign y10861 = ~n38459 ;
  assign y10862 = n38462 ;
  assign y10863 = n38470 ;
  assign y10864 = ~n38472 ;
  assign y10865 = ~n38478 ;
  assign y10866 = ~1'b0 ;
  assign y10867 = n38483 ;
  assign y10868 = n38484 ;
  assign y10869 = n38486 ;
  assign y10870 = ~n38487 ;
  assign y10871 = n38491 ;
  assign y10872 = ~n38494 ;
  assign y10873 = n38497 ;
  assign y10874 = ~n38499 ;
  assign y10875 = ~n38500 ;
  assign y10876 = ~n38504 ;
  assign y10877 = ~n38506 ;
  assign y10878 = ~n38507 ;
  assign y10879 = ~n38512 ;
  assign y10880 = n38513 ;
  assign y10881 = ~n38516 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = ~n38517 ;
  assign y10884 = ~n38518 ;
  assign y10885 = ~n38519 ;
  assign y10886 = ~n38520 ;
  assign y10887 = ~n38522 ;
  assign y10888 = ~n38523 ;
  assign y10889 = ~n38528 ;
  assign y10890 = ~n38530 ;
  assign y10891 = n38532 ;
  assign y10892 = ~1'b0 ;
  assign y10893 = ~n38534 ;
  assign y10894 = ~n38537 ;
  assign y10895 = ~n38546 ;
  assign y10896 = n38547 ;
  assign y10897 = ~n38554 ;
  assign y10898 = n38556 ;
  assign y10899 = n38557 ;
  assign y10900 = ~n38561 ;
  assign y10901 = ~n38565 ;
  assign y10902 = n38566 ;
  assign y10903 = n38568 ;
  assign y10904 = n38571 ;
  assign y10905 = ~n38575 ;
  assign y10906 = ~n38578 ;
  assign y10907 = n38583 ;
  assign y10908 = ~n38586 ;
  assign y10909 = n38588 ;
  assign y10910 = n38596 ;
  assign y10911 = ~n38601 ;
  assign y10912 = n38602 ;
  assign y10913 = n38603 ;
  assign y10914 = ~1'b0 ;
  assign y10915 = ~n38608 ;
  assign y10916 = n38610 ;
  assign y10917 = ~n38611 ;
  assign y10918 = n38612 ;
  assign y10919 = ~n38616 ;
  assign y10920 = ~n38618 ;
  assign y10921 = ~n38619 ;
  assign y10922 = ~n38620 ;
  assign y10923 = n38624 ;
  assign y10924 = ~n38628 ;
  assign y10925 = ~1'b0 ;
  assign y10926 = ~1'b0 ;
  assign y10927 = n38635 ;
  assign y10928 = ~n38637 ;
  assign y10929 = ~n31066 ;
  assign y10930 = n38638 ;
  assign y10931 = ~1'b0 ;
  assign y10932 = n38640 ;
  assign y10933 = n38643 ;
  assign y10934 = n38649 ;
  assign y10935 = n38653 ;
  assign y10936 = n38655 ;
  assign y10937 = ~n38659 ;
  assign y10938 = n38661 ;
  assign y10939 = n38663 ;
  assign y10940 = ~n38665 ;
  assign y10941 = ~n38668 ;
  assign y10942 = ~1'b0 ;
  assign y10943 = n38670 ;
  assign y10944 = ~n38674 ;
  assign y10945 = n38679 ;
  assign y10946 = n38682 ;
  assign y10947 = ~1'b0 ;
  assign y10948 = ~n38690 ;
  assign y10949 = ~n38692 ;
  assign y10950 = ~n38693 ;
  assign y10951 = ~1'b0 ;
  assign y10952 = n38694 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~n38696 ;
  assign y10955 = ~n38700 ;
  assign y10956 = n38705 ;
  assign y10957 = n38707 ;
  assign y10958 = n38708 ;
  assign y10959 = ~n38709 ;
  assign y10960 = ~n38711 ;
  assign y10961 = ~n38716 ;
  assign y10962 = n38717 ;
  assign y10963 = n38729 ;
  assign y10964 = ~n38731 ;
  assign y10965 = ~n38732 ;
  assign y10966 = ~n38734 ;
  assign y10967 = n38737 ;
  assign y10968 = n38738 ;
  assign y10969 = ~n38740 ;
  assign y10970 = ~n38743 ;
  assign y10971 = n38749 ;
  assign y10972 = n38752 ;
  assign y10973 = ~n38754 ;
  assign y10974 = n38755 ;
  assign y10975 = ~n38758 ;
  assign y10976 = ~1'b0 ;
  assign y10977 = ~n38760 ;
  assign y10978 = ~1'b0 ;
  assign y10979 = ~n38761 ;
  assign y10980 = ~n38764 ;
  assign y10981 = n38769 ;
  assign y10982 = n38770 ;
  assign y10983 = ~n38775 ;
  assign y10984 = ~n38777 ;
  assign y10985 = n38784 ;
  assign y10986 = n38787 ;
  assign y10987 = n38788 ;
  assign y10988 = ~n38791 ;
  assign y10989 = ~n38793 ;
  assign y10990 = ~n38796 ;
  assign y10991 = n38797 ;
  assign y10992 = n38799 ;
  assign y10993 = n38801 ;
  assign y10994 = n38806 ;
  assign y10995 = n38808 ;
  assign y10996 = ~n38811 ;
  assign y10997 = n38812 ;
  assign y10998 = n38815 ;
  assign y10999 = ~n38816 ;
  assign y11000 = ~n38817 ;
  assign y11001 = n38818 ;
  assign y11002 = ~n38819 ;
  assign y11003 = n38824 ;
  assign y11004 = ~1'b0 ;
  assign y11005 = ~n38829 ;
  assign y11006 = n38835 ;
  assign y11007 = n38836 ;
  assign y11008 = ~n38837 ;
  assign y11009 = n38841 ;
  assign y11010 = n38846 ;
  assign y11011 = n38855 ;
  assign y11012 = n38857 ;
  assign y11013 = ~n38859 ;
  assign y11014 = n38866 ;
  assign y11015 = n38869 ;
  assign y11016 = ~n21506 ;
  assign y11017 = ~n38872 ;
  assign y11018 = n38875 ;
  assign y11019 = ~1'b0 ;
  assign y11020 = n38876 ;
  assign y11021 = ~n38879 ;
  assign y11022 = n38880 ;
  assign y11023 = ~n38882 ;
  assign y11024 = ~n38891 ;
  assign y11025 = ~n38896 ;
  assign y11026 = ~n38897 ;
  assign y11027 = ~1'b0 ;
  assign y11028 = n38898 ;
  assign y11029 = n38901 ;
  assign y11030 = n38903 ;
  assign y11031 = ~n38912 ;
  assign y11032 = n38916 ;
  assign y11033 = n38918 ;
  assign y11034 = n38920 ;
  assign y11035 = n38929 ;
  assign y11036 = ~n38934 ;
  assign y11037 = ~n38936 ;
  assign y11038 = ~1'b0 ;
  assign y11039 = ~n38938 ;
  assign y11040 = ~n38940 ;
  assign y11041 = ~n38944 ;
  assign y11042 = ~n38946 ;
  assign y11043 = ~n38955 ;
  assign y11044 = ~1'b0 ;
  assign y11045 = ~n38958 ;
  assign y11046 = n38962 ;
  assign y11047 = ~n38964 ;
  assign y11048 = ~n38965 ;
  assign y11049 = ~n38969 ;
  assign y11050 = ~n38974 ;
  assign y11051 = n38976 ;
  assign y11052 = n38977 ;
  assign y11053 = n38978 ;
  assign y11054 = ~1'b0 ;
  assign y11055 = ~1'b0 ;
  assign y11056 = ~n38979 ;
  assign y11057 = ~n38981 ;
  assign y11058 = ~n38986 ;
  assign y11059 = n38988 ;
  assign y11060 = ~n38989 ;
  assign y11061 = n38992 ;
  assign y11062 = n38994 ;
  assign y11063 = ~n38999 ;
  assign y11064 = ~n39000 ;
  assign y11065 = ~n39006 ;
  assign y11066 = ~n39010 ;
  assign y11067 = n39013 ;
  assign y11068 = n39016 ;
  assign y11069 = n39018 ;
  assign y11070 = n39021 ;
  assign y11071 = n39024 ;
  assign y11072 = n39025 ;
  assign y11073 = n39027 ;
  assign y11074 = n39028 ;
  assign y11075 = ~n39030 ;
  assign y11076 = ~n39031 ;
  assign y11077 = ~n39034 ;
  assign y11078 = n39037 ;
  assign y11079 = ~n39039 ;
  assign y11080 = n39040 ;
  assign y11081 = n39041 ;
  assign y11082 = n39045 ;
  assign y11083 = ~n39057 ;
  assign y11084 = ~n39059 ;
  assign y11085 = ~1'b0 ;
  assign y11086 = ~n39065 ;
  assign y11087 = ~n39068 ;
  assign y11088 = ~n39070 ;
  assign y11089 = n39071 ;
  assign y11090 = n39073 ;
  assign y11091 = n39076 ;
  assign y11092 = n39077 ;
  assign y11093 = ~n39080 ;
  assign y11094 = ~n39082 ;
  assign y11095 = ~n39088 ;
  assign y11096 = n39090 ;
  assign y11097 = ~n39096 ;
  assign y11098 = ~n39100 ;
  assign y11099 = n39101 ;
  assign y11100 = n39102 ;
  assign y11101 = n39106 ;
  assign y11102 = n39108 ;
  assign y11103 = n39110 ;
  assign y11104 = ~n39114 ;
  assign y11105 = n39117 ;
  assign y11106 = ~n39122 ;
  assign y11107 = n39123 ;
  assign y11108 = n39124 ;
  assign y11109 = n39125 ;
  assign y11110 = ~n39129 ;
  assign y11111 = n39130 ;
  assign y11112 = ~n39132 ;
  assign y11113 = ~n39134 ;
  assign y11114 = ~n39140 ;
  assign y11115 = ~n39142 ;
  assign y11116 = n39143 ;
  assign y11117 = ~1'b0 ;
  assign y11118 = n39145 ;
  assign y11119 = n39148 ;
  assign y11120 = ~n39151 ;
  assign y11121 = ~n39156 ;
  assign y11122 = ~n39163 ;
  assign y11123 = ~n39167 ;
  assign y11124 = ~n39170 ;
  assign y11125 = n39171 ;
  assign y11126 = ~n39173 ;
  assign y11127 = ~n39176 ;
  assign y11128 = n39177 ;
  assign y11129 = n39178 ;
  assign y11130 = ~n39180 ;
  assign y11131 = ~1'b0 ;
  assign y11132 = ~n39182 ;
  assign y11133 = ~n39185 ;
  assign y11134 = n39187 ;
  assign y11135 = n39188 ;
  assign y11136 = ~1'b0 ;
  assign y11137 = n39195 ;
  assign y11138 = n39203 ;
  assign y11139 = ~n39210 ;
  assign y11140 = n39216 ;
  assign y11141 = ~n39219 ;
  assign y11142 = n39220 ;
  assign y11143 = ~n39231 ;
  assign y11144 = ~n39232 ;
  assign y11145 = ~n39234 ;
  assign y11146 = ~n39238 ;
  assign y11147 = n39239 ;
  assign y11148 = ~n39245 ;
  assign y11149 = n39248 ;
  assign y11150 = n39251 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~1'b0 ;
  assign y11153 = ~n39257 ;
  assign y11154 = ~n39261 ;
  assign y11155 = n39263 ;
  assign y11156 = ~n39265 ;
  assign y11157 = ~n39268 ;
  assign y11158 = ~1'b0 ;
  assign y11159 = n39270 ;
  assign y11160 = ~n39271 ;
  assign y11161 = ~n39275 ;
  assign y11162 = n39277 ;
  assign y11163 = n39281 ;
  assign y11164 = n39284 ;
  assign y11165 = n39286 ;
  assign y11166 = ~1'b0 ;
  assign y11167 = n39288 ;
  assign y11168 = n39289 ;
  assign y11169 = n39290 ;
  assign y11170 = ~n39292 ;
  assign y11171 = ~n39294 ;
  assign y11172 = ~n39296 ;
  assign y11173 = ~1'b0 ;
  assign y11174 = n39299 ;
  assign y11175 = n39300 ;
  assign y11176 = ~n39306 ;
  assign y11177 = ~n39307 ;
  assign y11178 = n39312 ;
  assign y11179 = n39316 ;
  assign y11180 = ~n39317 ;
  assign y11181 = ~1'b0 ;
  assign y11182 = ~1'b0 ;
  assign y11183 = n39319 ;
  assign y11184 = n39320 ;
  assign y11185 = ~n39321 ;
  assign y11186 = n39325 ;
  assign y11187 = n39327 ;
  assign y11188 = n39329 ;
  assign y11189 = n39331 ;
  assign y11190 = n39335 ;
  assign y11191 = ~1'b0 ;
  assign y11192 = n39337 ;
  assign y11193 = ~1'b0 ;
  assign y11194 = ~n39341 ;
  assign y11195 = ~n39345 ;
  assign y11196 = ~n39346 ;
  assign y11197 = n39347 ;
  assign y11198 = ~n39349 ;
  assign y11199 = n39355 ;
  assign y11200 = ~1'b0 ;
  assign y11201 = n39357 ;
  assign y11202 = ~n39363 ;
  assign y11203 = ~n39364 ;
  assign y11204 = n39365 ;
  assign y11205 = ~n39369 ;
  assign y11206 = ~n39375 ;
  assign y11207 = ~n39378 ;
  assign y11208 = n39380 ;
  assign y11209 = ~1'b0 ;
  assign y11210 = ~n39384 ;
  assign y11211 = ~n39387 ;
  assign y11212 = n39388 ;
  assign y11213 = n39390 ;
  assign y11214 = ~n39393 ;
  assign y11215 = n39395 ;
  assign y11216 = ~n39399 ;
  assign y11217 = n39400 ;
  assign y11218 = ~1'b0 ;
  assign y11219 = ~1'b0 ;
  assign y11220 = ~n39402 ;
  assign y11221 = ~n39404 ;
  assign y11222 = ~n39408 ;
  assign y11223 = n39409 ;
  assign y11224 = ~1'b0 ;
  assign y11225 = ~n39416 ;
  assign y11226 = ~n39419 ;
  assign y11227 = ~n39422 ;
  assign y11228 = ~n39424 ;
  assign y11229 = ~n39425 ;
  assign y11230 = ~n39428 ;
  assign y11231 = ~1'b0 ;
  assign y11232 = n39429 ;
  assign y11233 = n39433 ;
  assign y11234 = n39435 ;
  assign y11235 = n39436 ;
  assign y11236 = ~n39440 ;
  assign y11237 = n39443 ;
  assign y11238 = ~n39447 ;
  assign y11239 = n39451 ;
  assign y11240 = n39454 ;
  assign y11241 = ~1'b0 ;
  assign y11242 = ~n39461 ;
  assign y11243 = n39469 ;
  assign y11244 = n39470 ;
  assign y11245 = n39471 ;
  assign y11246 = ~n39474 ;
  assign y11247 = ~n39479 ;
  assign y11248 = ~n39481 ;
  assign y11249 = ~n39485 ;
  assign y11250 = n39488 ;
  assign y11251 = ~n39489 ;
  assign y11252 = ~n39490 ;
  assign y11253 = n39491 ;
  assign y11254 = ~n39501 ;
  assign y11255 = ~n39503 ;
  assign y11256 = n39506 ;
  assign y11257 = ~n39510 ;
  assign y11258 = n39512 ;
  assign y11259 = ~1'b0 ;
  assign y11260 = ~n39518 ;
  assign y11261 = ~1'b0 ;
  assign y11262 = ~n39519 ;
  assign y11263 = ~n39522 ;
  assign y11264 = n39523 ;
  assign y11265 = ~n39524 ;
  assign y11266 = ~n39529 ;
  assign y11267 = ~1'b0 ;
  assign y11268 = ~n39538 ;
  assign y11269 = n39540 ;
  assign y11270 = ~n39541 ;
  assign y11271 = ~n39542 ;
  assign y11272 = ~n39543 ;
  assign y11273 = n39545 ;
  assign y11274 = ~n39549 ;
  assign y11275 = ~n39552 ;
  assign y11276 = ~n39553 ;
  assign y11277 = ~n39558 ;
  assign y11278 = n39560 ;
  assign y11279 = n39563 ;
  assign y11280 = ~n39566 ;
  assign y11281 = ~n39568 ;
  assign y11282 = n39578 ;
  assign y11283 = n39579 ;
  assign y11284 = n39583 ;
  assign y11285 = n39589 ;
  assign y11286 = n39593 ;
  assign y11287 = n39597 ;
  assign y11288 = n39601 ;
  assign y11289 = ~n39604 ;
  assign y11290 = ~n39606 ;
  assign y11291 = ~n39607 ;
  assign y11292 = ~n39609 ;
  assign y11293 = n39611 ;
  assign y11294 = n39613 ;
  assign y11295 = n39615 ;
  assign y11296 = n39616 ;
  assign y11297 = ~n39618 ;
  assign y11298 = n39620 ;
  assign y11299 = ~n39623 ;
  assign y11300 = ~n39624 ;
  assign y11301 = n39625 ;
  assign y11302 = ~1'b0 ;
  assign y11303 = ~n39628 ;
  assign y11304 = ~n39630 ;
  assign y11305 = n39631 ;
  assign y11306 = ~n39635 ;
  assign y11307 = n39638 ;
  assign y11308 = n39640 ;
  assign y11309 = ~n39645 ;
  assign y11310 = n39646 ;
  assign y11311 = n39653 ;
  assign y11312 = ~n39654 ;
  assign y11313 = n39657 ;
  assign y11314 = n39662 ;
  assign y11315 = ~1'b0 ;
  assign y11316 = n39664 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = n39666 ;
  assign y11319 = ~n39668 ;
  assign y11320 = n39672 ;
  assign y11321 = n39674 ;
  assign y11322 = ~n39675 ;
  assign y11323 = n39676 ;
  assign y11324 = ~1'b0 ;
  assign y11325 = ~1'b0 ;
  assign y11326 = ~n39679 ;
  assign y11327 = ~n39681 ;
  assign y11328 = ~n39682 ;
  assign y11329 = n39683 ;
  assign y11330 = ~n39684 ;
  assign y11331 = ~1'b0 ;
  assign y11332 = ~n39691 ;
  assign y11333 = n39692 ;
  assign y11334 = n39206 ;
  assign y11335 = n39694 ;
  assign y11336 = n39697 ;
  assign y11337 = ~n39699 ;
  assign y11338 = n39701 ;
  assign y11339 = ~n39704 ;
  assign y11340 = ~n39707 ;
  assign y11341 = ~n39708 ;
  assign y11342 = n39709 ;
  assign y11343 = ~1'b0 ;
  assign y11344 = ~n39712 ;
  assign y11345 = ~1'b0 ;
  assign y11346 = n39713 ;
  assign y11347 = n39715 ;
  assign y11348 = n39718 ;
  assign y11349 = n39719 ;
  assign y11350 = n39726 ;
  assign y11351 = ~1'b0 ;
  assign y11352 = ~n39728 ;
  assign y11353 = ~n39730 ;
  assign y11354 = ~n39733 ;
  assign y11355 = ~n39734 ;
  assign y11356 = ~n39735 ;
  assign y11357 = ~n39739 ;
  assign y11358 = n39741 ;
  assign y11359 = ~1'b0 ;
  assign y11360 = ~1'b0 ;
  assign y11361 = n39746 ;
  assign y11362 = n39381 ;
  assign y11363 = n11238 ;
  assign y11364 = n39751 ;
  assign y11365 = ~n39752 ;
  assign y11366 = n39753 ;
  assign y11367 = ~1'b0 ;
  assign y11368 = n39756 ;
  assign y11369 = n39764 ;
  assign y11370 = n39765 ;
  assign y11371 = n39767 ;
  assign y11372 = ~n39771 ;
  assign y11373 = ~n39776 ;
  assign y11374 = ~n39779 ;
  assign y11375 = n39783 ;
  assign y11376 = n39784 ;
  assign y11377 = n39785 ;
  assign y11378 = n39787 ;
  assign y11379 = ~n39790 ;
  assign y11380 = ~n39795 ;
  assign y11381 = ~n39798 ;
  assign y11382 = n39801 ;
  assign y11383 = ~n39804 ;
  assign y11384 = ~n39807 ;
  assign y11385 = n39809 ;
  assign y11386 = ~n39814 ;
  assign y11387 = ~n39817 ;
  assign y11388 = ~n39819 ;
  assign y11389 = ~n39821 ;
  assign y11390 = ~n39822 ;
  assign y11391 = n39825 ;
  assign y11392 = n39828 ;
  assign y11393 = n39832 ;
  assign y11394 = n39833 ;
  assign y11395 = n39835 ;
  assign y11396 = n39839 ;
  assign y11397 = n39840 ;
  assign y11398 = ~n39843 ;
  assign y11399 = n39844 ;
  assign y11400 = n39845 ;
  assign y11401 = n39846 ;
  assign y11402 = ~n39849 ;
  assign y11403 = ~1'b0 ;
  assign y11404 = n39850 ;
  assign y11405 = ~1'b0 ;
  assign y11406 = ~n39854 ;
  assign y11407 = ~n39856 ;
  assign y11408 = n39859 ;
  assign y11409 = n39861 ;
  assign y11410 = ~n39862 ;
  assign y11411 = n26641 ;
  assign y11412 = ~n39864 ;
  assign y11413 = ~n39866 ;
  assign y11414 = ~n39871 ;
  assign y11415 = n39875 ;
  assign y11416 = n39877 ;
  assign y11417 = n39878 ;
  assign y11418 = ~n39884 ;
  assign y11419 = n39888 ;
  assign y11420 = n39891 ;
  assign y11421 = ~n39895 ;
  assign y11422 = ~n39900 ;
  assign y11423 = n39903 ;
  assign y11424 = n34364 ;
  assign y11425 = n39906 ;
  assign y11426 = ~n39907 ;
  assign y11427 = n39908 ;
  assign y11428 = n39909 ;
  assign y11429 = n39913 ;
  assign y11430 = ~n39916 ;
  assign y11431 = ~n39918 ;
  assign y11432 = ~n39919 ;
  assign y11433 = ~n39921 ;
  assign y11434 = ~n39924 ;
  assign y11435 = n39928 ;
  assign y11436 = ~1'b0 ;
  assign y11437 = n39929 ;
  assign y11438 = ~n39942 ;
  assign y11439 = ~n39945 ;
  assign y11440 = ~n39946 ;
  assign y11441 = n39950 ;
  assign y11442 = n39954 ;
  assign y11443 = ~n39956 ;
  assign y11444 = n17534 ;
  assign y11445 = n39958 ;
  assign y11446 = n39962 ;
  assign y11447 = ~n39963 ;
  assign y11448 = n39964 ;
  assign y11449 = ~n39965 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = n39973 ;
  assign y11452 = n39974 ;
  assign y11453 = ~n39977 ;
  assign y11454 = n39981 ;
  assign y11455 = n39988 ;
  assign y11456 = n39989 ;
  assign y11457 = ~n39990 ;
  assign y11458 = ~n39991 ;
  assign y11459 = ~1'b0 ;
  assign y11460 = ~1'b0 ;
  assign y11461 = n39992 ;
  assign y11462 = ~n39994 ;
  assign y11463 = n39995 ;
  assign y11464 = n39996 ;
  assign y11465 = ~n40000 ;
  assign y11466 = ~n40010 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = ~n40011 ;
  assign y11469 = ~n40012 ;
  assign y11470 = ~n40013 ;
  assign y11471 = n40014 ;
  assign y11472 = ~n40016 ;
  assign y11473 = n40024 ;
  assign y11474 = n40027 ;
  assign y11475 = ~n5470 ;
  assign y11476 = n40029 ;
  assign y11477 = ~n40030 ;
  assign y11478 = ~n40031 ;
  assign y11479 = ~n40032 ;
  assign y11480 = ~n40034 ;
  assign y11481 = n40039 ;
  assign y11482 = ~n40040 ;
  assign y11483 = n40042 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = n40043 ;
  assign y11486 = n40048 ;
  assign y11487 = n40052 ;
  assign y11488 = n40053 ;
  assign y11489 = ~n40054 ;
  assign y11490 = ~n40060 ;
  assign y11491 = n40063 ;
  assign y11492 = ~1'b0 ;
  assign y11493 = ~n40068 ;
  assign y11494 = ~1'b0 ;
  assign y11495 = n40069 ;
  assign y11496 = ~n40072 ;
  assign y11497 = ~n40077 ;
  assign y11498 = ~n40087 ;
  assign y11499 = ~n40089 ;
  assign y11500 = n40092 ;
  assign y11501 = n40093 ;
  assign y11502 = n40094 ;
  assign y11503 = n40097 ;
  assign y11504 = ~n40098 ;
  assign y11505 = ~n40099 ;
  assign y11506 = n40103 ;
  assign y11507 = ~n40106 ;
  assign y11508 = n40111 ;
  assign y11509 = ~n40112 ;
  assign y11510 = n40115 ;
  assign y11511 = ~n40120 ;
  assign y11512 = n40121 ;
  assign y11513 = n40124 ;
  assign y11514 = n40126 ;
  assign y11515 = n40129 ;
  assign y11516 = ~n40130 ;
  assign y11517 = ~n40132 ;
  assign y11518 = n40135 ;
  assign y11519 = n40142 ;
  assign y11520 = n40145 ;
  assign y11521 = ~n40150 ;
  assign y11522 = ~n40153 ;
  assign y11523 = ~1'b0 ;
  assign y11524 = ~n40155 ;
  assign y11525 = n40156 ;
  assign y11526 = ~n40161 ;
  assign y11527 = ~n40162 ;
  assign y11528 = n40164 ;
  assign y11529 = ~n40169 ;
  assign y11530 = ~n40173 ;
  assign y11531 = ~1'b0 ;
  assign y11532 = ~n40174 ;
  assign y11533 = ~n40177 ;
  assign y11534 = ~n40181 ;
  assign y11535 = ~n40184 ;
  assign y11536 = ~n40188 ;
  assign y11537 = ~n40190 ;
  assign y11538 = ~n40191 ;
  assign y11539 = n40192 ;
  assign y11540 = ~n40196 ;
  assign y11541 = ~1'b0 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = ~n40201 ;
  assign y11544 = ~n40203 ;
  assign y11545 = ~1'b0 ;
  assign y11546 = ~n40206 ;
  assign y11547 = n40207 ;
  assign y11548 = ~n40208 ;
  assign y11549 = ~n40211 ;
  assign y11550 = n40212 ;
  assign y11551 = ~1'b0 ;
  assign y11552 = ~n40213 ;
  assign y11553 = n40216 ;
  assign y11554 = ~n40218 ;
  assign y11555 = ~n40219 ;
  assign y11556 = n40220 ;
  assign y11557 = n40222 ;
  assign y11558 = n40223 ;
  assign y11559 = n40227 ;
  assign y11560 = ~n40230 ;
  assign y11561 = ~1'b0 ;
  assign y11562 = n40234 ;
  assign y11563 = ~n40240 ;
  assign y11564 = ~n40246 ;
  assign y11565 = n40248 ;
  assign y11566 = ~n40250 ;
  assign y11567 = ~n40253 ;
  assign y11568 = ~n40264 ;
  assign y11569 = n16296 ;
  assign y11570 = n40267 ;
  assign y11571 = n40272 ;
  assign y11572 = ~n40275 ;
  assign y11573 = ~n40280 ;
  assign y11574 = ~n40283 ;
  assign y11575 = ~n40285 ;
  assign y11576 = ~n40286 ;
  assign y11577 = n40287 ;
  assign y11578 = ~n40290 ;
  assign y11579 = ~n40293 ;
  assign y11580 = n40299 ;
  assign y11581 = ~n40301 ;
  assign y11582 = n40302 ;
  assign y11583 = ~n40312 ;
  assign y11584 = ~n40313 ;
  assign y11585 = n40325 ;
  assign y11586 = ~n40326 ;
  assign y11587 = n40329 ;
  assign y11588 = ~n40333 ;
  assign y11589 = n40334 ;
  assign y11590 = ~n40335 ;
  assign y11591 = ~n40342 ;
  assign y11592 = ~n40344 ;
  assign y11593 = ~n40349 ;
  assign y11594 = n40354 ;
  assign y11595 = n40356 ;
  assign y11596 = ~1'b0 ;
  assign y11597 = n40358 ;
  assign y11598 = n40362 ;
  assign y11599 = ~n40364 ;
  assign y11600 = n40365 ;
  assign y11601 = n40368 ;
  assign y11602 = n40377 ;
  assign y11603 = ~n40380 ;
  assign y11604 = n40387 ;
  assign y11605 = ~1'b0 ;
  assign y11606 = ~n40390 ;
  assign y11607 = ~n40393 ;
  assign y11608 = ~n40394 ;
  assign y11609 = ~n40395 ;
  assign y11610 = n40396 ;
  assign y11611 = ~n40399 ;
  assign y11612 = ~n40401 ;
  assign y11613 = ~n40404 ;
  assign y11614 = ~n40410 ;
  assign y11615 = ~1'b0 ;
  assign y11616 = ~1'b0 ;
  assign y11617 = n40417 ;
  assign y11618 = ~n40418 ;
  assign y11619 = n40419 ;
  assign y11620 = ~n40420 ;
  assign y11621 = ~n40423 ;
  assign y11622 = ~1'b0 ;
  assign y11623 = n40425 ;
  assign y11624 = ~n40428 ;
  assign y11625 = n40429 ;
  assign y11626 = ~n40431 ;
  assign y11627 = n40433 ;
  assign y11628 = ~1'b0 ;
  assign y11629 = ~n40434 ;
  assign y11630 = ~1'b0 ;
  assign y11631 = n40436 ;
  assign y11632 = n40442 ;
  assign y11633 = n40445 ;
  assign y11634 = ~1'b0 ;
  assign y11635 = ~n40451 ;
  assign y11636 = n40458 ;
  assign y11637 = n40459 ;
  assign y11638 = n40461 ;
  assign y11639 = n40462 ;
  assign y11640 = ~n40465 ;
  assign y11641 = n40466 ;
  assign y11642 = n40467 ;
  assign y11643 = ~n40471 ;
  assign y11644 = n40475 ;
  assign y11645 = n40477 ;
  assign y11646 = ~n40481 ;
  assign y11647 = n40482 ;
  assign y11648 = ~n40483 ;
  assign y11649 = n40487 ;
  assign y11650 = ~1'b0 ;
  assign y11651 = ~1'b0 ;
  assign y11652 = n40491 ;
  assign y11653 = ~n40493 ;
  assign y11654 = n40497 ;
  assign y11655 = n40499 ;
  assign y11656 = ~n40509 ;
  assign y11657 = ~n40512 ;
  assign y11658 = n40523 ;
  assign y11659 = ~n40526 ;
  assign y11660 = ~1'b0 ;
  assign y11661 = ~n40528 ;
  assign y11662 = n40531 ;
  assign y11663 = n40535 ;
  assign y11664 = n40537 ;
  assign y11665 = n40542 ;
  assign y11666 = ~n40545 ;
  assign y11667 = n40559 ;
  assign y11668 = n40563 ;
  assign y11669 = ~n40567 ;
  assign y11670 = n40568 ;
  assign y11671 = ~1'b0 ;
  assign y11672 = ~1'b0 ;
  assign y11673 = ~n40573 ;
  assign y11674 = ~n40574 ;
  assign y11675 = n40576 ;
  assign y11676 = ~n40579 ;
  assign y11677 = n40582 ;
  assign y11678 = ~n40584 ;
  assign y11679 = n40587 ;
  assign y11680 = n40588 ;
  assign y11681 = n40591 ;
  assign y11682 = n40592 ;
  assign y11683 = ~n40601 ;
  assign y11684 = ~n40603 ;
  assign y11685 = n40607 ;
  assign y11686 = n40609 ;
  assign y11687 = n633 ;
  assign y11688 = n40613 ;
  assign y11689 = n40617 ;
  assign y11690 = ~n40620 ;
  assign y11691 = ~n40623 ;
  assign y11692 = n40627 ;
  assign y11693 = n40629 ;
  assign y11694 = ~1'b0 ;
  assign y11695 = n40632 ;
  assign y11696 = ~n40633 ;
  assign y11697 = n40635 ;
  assign y11698 = n40643 ;
  assign y11699 = n40645 ;
  assign y11700 = ~n40652 ;
  assign y11701 = n40657 ;
  assign y11702 = ~1'b0 ;
  assign y11703 = ~n40658 ;
  assign y11704 = ~n40661 ;
  assign y11705 = n40666 ;
  assign y11706 = n40670 ;
  assign y11707 = ~n40671 ;
  assign y11708 = n40677 ;
  assign y11709 = ~1'b0 ;
  assign y11710 = ~1'b0 ;
  assign y11711 = ~n40678 ;
  assign y11712 = ~n40684 ;
  assign y11713 = n40685 ;
  assign y11714 = n40688 ;
  assign y11715 = n40690 ;
  assign y11716 = n40691 ;
  assign y11717 = ~n40694 ;
  assign y11718 = ~n40699 ;
  assign y11719 = ~n40702 ;
  assign y11720 = n40705 ;
  assign y11721 = n40707 ;
  assign y11722 = ~n40711 ;
  assign y11723 = ~n40712 ;
  assign y11724 = ~1'b0 ;
  assign y11725 = ~n40714 ;
  assign y11726 = ~n40716 ;
  assign y11727 = ~n40717 ;
  assign y11728 = ~1'b0 ;
  assign y11729 = ~n40722 ;
  assign y11730 = n40723 ;
  assign y11731 = ~n40724 ;
  assign y11732 = ~n40730 ;
  assign y11733 = ~n40732 ;
  assign y11734 = n40735 ;
  assign y11735 = n40743 ;
  assign y11736 = ~1'b0 ;
  assign y11737 = ~n40745 ;
  assign y11738 = n40746 ;
  assign y11739 = n40747 ;
  assign y11740 = ~n40755 ;
  assign y11741 = n40757 ;
  assign y11742 = ~1'b0 ;
  assign y11743 = ~n40762 ;
  assign y11744 = ~1'b0 ;
  assign y11745 = n40768 ;
  assign y11746 = n40769 ;
  assign y11747 = n40771 ;
  assign y11748 = ~n40776 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = ~1'b0 ;
  assign y11751 = ~n40780 ;
  assign y11752 = ~n40781 ;
  assign y11753 = ~n40782 ;
  assign y11754 = ~n40787 ;
  assign y11755 = ~1'b0 ;
  assign y11756 = ~n40788 ;
  assign y11757 = n40794 ;
  assign y11758 = n40795 ;
  assign y11759 = ~n40797 ;
  assign y11760 = ~1'b0 ;
  assign y11761 = ~n40798 ;
  assign y11762 = n40802 ;
  assign y11763 = n40803 ;
  assign y11764 = n40805 ;
  assign y11765 = n40807 ;
  assign y11766 = ~n40814 ;
  assign y11767 = ~1'b0 ;
  assign y11768 = n40816 ;
  assign y11769 = n40817 ;
  assign y11770 = ~n40818 ;
  assign y11771 = n40827 ;
  assign y11772 = ~1'b0 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = ~1'b0 ;
  assign y11775 = ~n40831 ;
  assign y11776 = n40833 ;
  assign y11777 = n40834 ;
  assign y11778 = n40836 ;
  assign y11779 = n40837 ;
  assign y11780 = ~n40838 ;
  assign y11781 = n40839 ;
  assign y11782 = ~n40843 ;
  assign y11783 = ~n40844 ;
  assign y11784 = n40845 ;
  assign y11785 = n40847 ;
  assign y11786 = n40857 ;
  assign y11787 = n40860 ;
  assign y11788 = ~n40864 ;
  assign y11789 = n40867 ;
  assign y11790 = n40875 ;
  assign y11791 = ~n40877 ;
  assign y11792 = ~n40880 ;
  assign y11793 = ~1'b0 ;
  assign y11794 = ~n40881 ;
  assign y11795 = n40884 ;
  assign y11796 = ~n40888 ;
  assign y11797 = ~n40889 ;
  assign y11798 = ~n40894 ;
  assign y11799 = n40896 ;
  assign y11800 = ~n40899 ;
  assign y11801 = ~1'b0 ;
  assign y11802 = n40900 ;
  assign y11803 = n40903 ;
  assign y11804 = n40904 ;
  assign y11805 = ~1'b0 ;
  assign y11806 = ~1'b0 ;
  assign y11807 = ~n40907 ;
  assign y11808 = n40916 ;
  assign y11809 = ~n40917 ;
  assign y11810 = ~n40918 ;
  assign y11811 = n40920 ;
  assign y11812 = n40926 ;
  assign y11813 = ~n40928 ;
  assign y11814 = ~n40929 ;
  assign y11815 = ~n40931 ;
  assign y11816 = n40937 ;
  assign y11817 = n40938 ;
  assign y11818 = ~n40941 ;
  assign y11819 = n40942 ;
  assign y11820 = n40944 ;
  assign y11821 = ~n40945 ;
  assign y11822 = n40949 ;
  assign y11823 = ~n40950 ;
  assign y11824 = ~n40953 ;
  assign y11825 = ~n829 ;
  assign y11826 = n40959 ;
  assign y11827 = n40961 ;
  assign y11828 = n40962 ;
  assign y11829 = ~1'b0 ;
  assign y11830 = ~n40967 ;
  assign y11831 = ~n40969 ;
  assign y11832 = ~n40970 ;
  assign y11833 = n40976 ;
  assign y11834 = n40978 ;
  assign y11835 = ~n40984 ;
  assign y11836 = ~n40986 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = ~1'b0 ;
  assign y11839 = ~n40988 ;
  assign y11840 = ~n40989 ;
  assign y11841 = n40993 ;
  assign y11842 = n40996 ;
  assign y11843 = ~n41002 ;
  assign y11844 = n41006 ;
  assign y11845 = ~n41007 ;
  assign y11846 = ~1'b0 ;
  assign y11847 = n41009 ;
  assign y11848 = ~1'b0 ;
  assign y11849 = n41011 ;
  assign y11850 = n41015 ;
  assign y11851 = ~n41018 ;
  assign y11852 = ~n41021 ;
  assign y11853 = ~n41022 ;
  assign y11854 = ~n41024 ;
  assign y11855 = n41029 ;
  assign y11856 = ~n41033 ;
  assign y11857 = ~n41035 ;
  assign y11858 = ~n41038 ;
  assign y11859 = n41041 ;
  assign y11860 = ~n41043 ;
  assign y11861 = ~n41044 ;
  assign y11862 = ~n41048 ;
  assign y11863 = n41050 ;
  assign y11864 = n41052 ;
  assign y11865 = n41053 ;
  assign y11866 = n41062 ;
  assign y11867 = n41065 ;
  assign y11868 = ~1'b0 ;
  assign y11869 = n41068 ;
  assign y11870 = n41069 ;
  assign y11871 = ~n41071 ;
  assign y11872 = ~n41075 ;
  assign y11873 = ~n41077 ;
  assign y11874 = n41079 ;
  assign y11875 = ~n41082 ;
  assign y11876 = ~n41084 ;
  assign y11877 = ~n41086 ;
  assign y11878 = n41088 ;
  assign y11879 = ~1'b0 ;
  assign y11880 = ~n41090 ;
  assign y11881 = ~n41091 ;
  assign y11882 = ~n32046 ;
  assign y11883 = ~n41092 ;
  assign y11884 = n41095 ;
  assign y11885 = ~n41096 ;
  assign y11886 = n41097 ;
  assign y11887 = n41106 ;
  assign y11888 = ~n41107 ;
  assign y11889 = n41109 ;
  assign y11890 = ~n41110 ;
  assign y11891 = n41112 ;
  assign y11892 = n41115 ;
  assign y11893 = ~1'b0 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = ~n41125 ;
  assign y11896 = ~n41127 ;
  assign y11897 = n41128 ;
  assign y11898 = n41130 ;
  assign y11899 = n41133 ;
  assign y11900 = ~n41140 ;
  assign y11901 = ~n41141 ;
  assign y11902 = ~n41143 ;
  assign y11903 = n41144 ;
  assign y11904 = ~n41146 ;
  assign y11905 = n41147 ;
  assign y11906 = n41152 ;
  assign y11907 = ~n41154 ;
  assign y11908 = n41156 ;
  assign y11909 = ~n41157 ;
  assign y11910 = ~n41159 ;
  assign y11911 = ~1'b0 ;
  assign y11912 = ~1'b0 ;
  assign y11913 = ~1'b0 ;
  assign y11914 = n41160 ;
  assign y11915 = ~n41169 ;
  assign y11916 = n41171 ;
  assign y11917 = ~1'b0 ;
  assign y11918 = ~1'b0 ;
  assign y11919 = ~1'b0 ;
  assign y11920 = n41172 ;
  assign y11921 = n41175 ;
  assign y11922 = n41177 ;
  assign y11923 = n41178 ;
  assign y11924 = ~n41183 ;
  assign y11925 = ~n41185 ;
  assign y11926 = n41187 ;
  assign y11927 = ~1'b0 ;
  assign y11928 = ~n41189 ;
  assign y11929 = n41190 ;
  assign y11930 = n41191 ;
  assign y11931 = n41192 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~n41193 ;
  assign y11934 = n41196 ;
  assign y11935 = n41197 ;
  assign y11936 = n41204 ;
  assign y11937 = n41205 ;
  assign y11938 = n41206 ;
  assign y11939 = n41207 ;
  assign y11940 = ~1'b0 ;
  assign y11941 = ~n41210 ;
  assign y11942 = n41211 ;
  assign y11943 = ~n41214 ;
  assign y11944 = ~n41215 ;
  assign y11945 = ~n41218 ;
  assign y11946 = ~n41223 ;
  assign y11947 = n41227 ;
  assign y11948 = n41233 ;
  assign y11949 = ~n41234 ;
  assign y11950 = n41236 ;
  assign y11951 = n41237 ;
  assign y11952 = ~n41240 ;
  assign y11953 = ~n41241 ;
  assign y11954 = n41242 ;
  assign y11955 = n41247 ;
  assign y11956 = ~n41249 ;
  assign y11957 = ~n41250 ;
  assign y11958 = ~n41251 ;
  assign y11959 = n41252 ;
  assign y11960 = ~n41254 ;
  assign y11961 = ~n41255 ;
  assign y11962 = n41257 ;
  assign y11963 = n41259 ;
  assign y11964 = ~n41263 ;
  assign y11965 = n41264 ;
  assign y11966 = n41267 ;
  assign y11967 = ~n41268 ;
  assign y11968 = n41271 ;
  assign y11969 = n41272 ;
  assign y11970 = ~1'b0 ;
  assign y11971 = ~n41277 ;
  assign y11972 = ~n41285 ;
  assign y11973 = ~n41289 ;
  assign y11974 = n41295 ;
  assign y11975 = ~n41296 ;
  assign y11976 = n41299 ;
  assign y11977 = ~n41303 ;
  assign y11978 = ~n41306 ;
  assign y11979 = ~1'b0 ;
  assign y11980 = n41307 ;
  assign y11981 = n41309 ;
  assign y11982 = ~n41311 ;
  assign y11983 = ~n41315 ;
  assign y11984 = ~n41316 ;
  assign y11985 = ~n41327 ;
  assign y11986 = 1'b0 ;
  assign y11987 = n41329 ;
  assign y11988 = ~n41331 ;
  assign y11989 = ~n41332 ;
  assign y11990 = ~n41333 ;
  assign y11991 = n41336 ;
  assign y11992 = ~n41341 ;
  assign y11993 = n41347 ;
  assign y11994 = ~1'b0 ;
  assign y11995 = ~n41355 ;
  assign y11996 = ~n41357 ;
  assign y11997 = ~n41360 ;
  assign y11998 = ~n41361 ;
  assign y11999 = n41362 ;
  assign y12000 = ~n41368 ;
  assign y12001 = n41371 ;
  assign y12002 = ~n41373 ;
  assign y12003 = ~1'b0 ;
  assign y12004 = ~n41375 ;
  assign y12005 = 1'b0 ;
  assign y12006 = ~n41376 ;
  assign y12007 = n41377 ;
  assign y12008 = n41379 ;
  assign y12009 = ~n41380 ;
  assign y12010 = n41382 ;
  assign y12011 = ~1'b0 ;
  assign y12012 = ~1'b0 ;
  assign y12013 = n41383 ;
  assign y12014 = n41384 ;
  assign y12015 = n41386 ;
  assign y12016 = ~n41387 ;
  assign y12017 = n41388 ;
  assign y12018 = ~1'b0 ;
  assign y12019 = ~n41391 ;
  assign y12020 = n41392 ;
  assign y12021 = n41393 ;
  assign y12022 = n41398 ;
  assign y12023 = ~n41404 ;
  assign y12024 = ~n41409 ;
  assign y12025 = n41410 ;
  assign y12026 = ~1'b0 ;
  assign y12027 = n41411 ;
  assign y12028 = n41414 ;
  assign y12029 = ~n41415 ;
  assign y12030 = n41416 ;
  assign y12031 = n41417 ;
  assign y12032 = n41423 ;
  assign y12033 = ~n41429 ;
  assign y12034 = ~1'b0 ;
  assign y12035 = n41432 ;
  assign y12036 = ~n41433 ;
  assign y12037 = n41440 ;
  assign y12038 = n41442 ;
  assign y12039 = n41443 ;
  assign y12040 = ~1'b0 ;
  assign y12041 = ~n41450 ;
  assign y12042 = n41451 ;
  assign y12043 = n41457 ;
  assign y12044 = ~n41461 ;
  assign y12045 = ~n41463 ;
  assign y12046 = n41469 ;
  assign y12047 = ~n41472 ;
  assign y12048 = n41478 ;
  assign y12049 = ~n41479 ;
  assign y12050 = ~n41486 ;
  assign y12051 = n41487 ;
  assign y12052 = ~n41489 ;
  assign y12053 = n41490 ;
  assign y12054 = ~n41491 ;
  assign y12055 = n41492 ;
  assign y12056 = n41497 ;
  assign y12057 = n41499 ;
  assign y12058 = n41502 ;
  assign y12059 = n41503 ;
  assign y12060 = n41505 ;
  assign y12061 = ~n41508 ;
  assign y12062 = n41512 ;
  assign y12063 = ~n41517 ;
  assign y12064 = n41519 ;
  assign y12065 = ~n41523 ;
  assign y12066 = n41528 ;
  assign y12067 = ~n41533 ;
  assign y12068 = ~n41538 ;
  assign y12069 = ~n41543 ;
  assign y12070 = n41544 ;
  assign y12071 = n41546 ;
  assign y12072 = ~n41547 ;
  assign y12073 = ~n41550 ;
  assign y12074 = ~n41557 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = n41559 ;
  assign y12077 = ~n41561 ;
  assign y12078 = n41565 ;
  assign y12079 = n41566 ;
  assign y12080 = n41567 ;
  assign y12081 = n41569 ;
  assign y12082 = ~n41571 ;
  assign y12083 = ~n41573 ;
  assign y12084 = n41579 ;
  assign y12085 = n41581 ;
  assign y12086 = n41582 ;
  assign y12087 = n41584 ;
  assign y12088 = ~n41589 ;
  assign y12089 = n41594 ;
  assign y12090 = n41600 ;
  assign y12091 = ~n41602 ;
  assign y12092 = n41604 ;
  assign y12093 = ~n41607 ;
  assign y12094 = n41610 ;
  assign y12095 = ~n41616 ;
  assign y12096 = n41617 ;
  assign y12097 = ~n41620 ;
  assign y12098 = ~n41625 ;
  assign y12099 = n41628 ;
  assign y12100 = n41629 ;
  assign y12101 = n41634 ;
  assign y12102 = ~n41636 ;
  assign y12103 = n41637 ;
  assign y12104 = ~n41640 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = n41642 ;
  assign y12107 = ~n41644 ;
  assign y12108 = ~n41651 ;
  assign y12109 = n41654 ;
  assign y12110 = n41655 ;
  assign y12111 = ~n41657 ;
  assign y12112 = ~n41658 ;
  assign y12113 = n41664 ;
  assign y12114 = ~1'b0 ;
  assign y12115 = ~n41666 ;
  assign y12116 = n41668 ;
  assign y12117 = ~1'b0 ;
  assign y12118 = ~n41669 ;
  assign y12119 = ~n41671 ;
  assign y12120 = n41674 ;
  assign y12121 = ~n41679 ;
  assign y12122 = n41680 ;
  assign y12123 = ~n41684 ;
  assign y12124 = ~n41685 ;
  assign y12125 = n41687 ;
  assign y12126 = n41688 ;
  assign y12127 = n41689 ;
  assign y12128 = n41690 ;
  assign y12129 = ~n41691 ;
  assign y12130 = n41698 ;
  assign y12131 = n41702 ;
  assign y12132 = ~1'b0 ;
  assign y12133 = ~n41703 ;
  assign y12134 = ~1'b0 ;
  assign y12135 = n41704 ;
  assign y12136 = ~n41709 ;
  assign y12137 = ~n41710 ;
  assign y12138 = ~n41711 ;
  assign y12139 = n41712 ;
  assign y12140 = ~n41714 ;
  assign y12141 = n41715 ;
  assign y12142 = ~n41721 ;
  assign y12143 = n41724 ;
  assign y12144 = ~n41725 ;
  assign y12145 = ~n41730 ;
  assign y12146 = n41731 ;
  assign y12147 = ~n41732 ;
  assign y12148 = ~1'b0 ;
  assign y12149 = ~1'b0 ;
  assign y12150 = n41739 ;
  assign y12151 = n41742 ;
  assign y12152 = n41743 ;
  assign y12153 = n41747 ;
  assign y12154 = ~n41754 ;
  assign y12155 = ~n41759 ;
  assign y12156 = ~n41761 ;
  assign y12157 = ~n41765 ;
  assign y12158 = ~n41769 ;
  assign y12159 = ~1'b0 ;
  assign y12160 = ~n41773 ;
  assign y12161 = ~n41775 ;
  assign y12162 = n41777 ;
  assign y12163 = n41782 ;
  assign y12164 = ~n41783 ;
  assign y12165 = ~n41784 ;
  assign y12166 = n41789 ;
  assign y12167 = n41791 ;
  assign y12168 = ~n41795 ;
  assign y12169 = n41798 ;
  assign y12170 = ~1'b0 ;
  assign y12171 = ~n41801 ;
  assign y12172 = n41802 ;
  assign y12173 = n41805 ;
  assign y12174 = n41807 ;
  assign y12175 = ~n41808 ;
  assign y12176 = ~n41811 ;
  assign y12177 = n41812 ;
  assign y12178 = ~n41815 ;
  assign y12179 = ~n41816 ;
  assign y12180 = ~1'b0 ;
  assign y12181 = n41817 ;
  assign y12182 = ~n41818 ;
  assign y12183 = ~n41820 ;
  assign y12184 = n41828 ;
  assign y12185 = ~n41830 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = n41831 ;
  assign y12188 = ~n41833 ;
  assign y12189 = ~n41838 ;
  assign y12190 = ~n41839 ;
  assign y12191 = ~n41840 ;
  assign y12192 = n41841 ;
  assign y12193 = ~n41843 ;
  assign y12194 = n41848 ;
  assign y12195 = ~n6316 ;
  assign y12196 = n41849 ;
  assign y12197 = ~n41851 ;
  assign y12198 = ~n41854 ;
  assign y12199 = ~n41855 ;
  assign y12200 = n41860 ;
  assign y12201 = ~n41869 ;
  assign y12202 = ~n41874 ;
  assign y12203 = ~n41881 ;
  assign y12204 = n41886 ;
  assign y12205 = n41893 ;
  assign y12206 = ~n41894 ;
  assign y12207 = n41898 ;
  assign y12208 = n41899 ;
  assign y12209 = n41903 ;
  assign y12210 = ~n41908 ;
  assign y12211 = n41909 ;
  assign y12212 = ~n41910 ;
  assign y12213 = n41914 ;
  assign y12214 = n41915 ;
  assign y12215 = n41916 ;
  assign y12216 = n41918 ;
  assign y12217 = n41919 ;
  assign y12218 = ~1'b0 ;
  assign y12219 = ~n41922 ;
  assign y12220 = ~n41926 ;
  assign y12221 = ~1'b0 ;
  assign y12222 = n41929 ;
  assign y12223 = ~n41932 ;
  assign y12224 = n41933 ;
  assign y12225 = ~n41936 ;
  assign y12226 = n41939 ;
  assign y12227 = ~1'b0 ;
  assign y12228 = ~1'b0 ;
  assign y12229 = ~1'b0 ;
  assign y12230 = n41943 ;
  assign y12231 = n41946 ;
  assign y12232 = n41948 ;
  assign y12233 = ~n41950 ;
  assign y12234 = n41953 ;
  assign y12235 = n41955 ;
  assign y12236 = n41957 ;
  assign y12237 = ~n41958 ;
  assign y12238 = n41959 ;
  assign y12239 = n41960 ;
  assign y12240 = n41961 ;
  assign y12241 = ~n41962 ;
  assign y12242 = ~n26612 ;
  assign y12243 = ~n41964 ;
  assign y12244 = ~1'b0 ;
  assign y12245 = ~n41967 ;
  assign y12246 = ~1'b0 ;
  assign y12247 = n41970 ;
  assign y12248 = ~n41972 ;
  assign y12249 = ~n41973 ;
  assign y12250 = ~n41976 ;
  assign y12251 = n41984 ;
  assign y12252 = ~n41989 ;
  assign y12253 = ~1'b0 ;
  assign y12254 = ~n42000 ;
  assign y12255 = ~n42002 ;
  assign y12256 = n42003 ;
  assign y12257 = n42005 ;
  assign y12258 = ~n42009 ;
  assign y12259 = n42012 ;
  assign y12260 = ~1'b0 ;
  assign y12261 = ~n42014 ;
  assign y12262 = ~n42016 ;
  assign y12263 = n42027 ;
  assign y12264 = ~n42028 ;
  assign y12265 = ~n42030 ;
  assign y12266 = ~n42035 ;
  assign y12267 = ~n42040 ;
  assign y12268 = ~n42042 ;
  assign y12269 = ~n42048 ;
  assign y12270 = ~1'b0 ;
  assign y12271 = ~n42053 ;
  assign y12272 = ~n42054 ;
  assign y12273 = ~n42056 ;
  assign y12274 = ~n42063 ;
  assign y12275 = ~n42064 ;
  assign y12276 = ~1'b0 ;
  assign y12277 = ~1'b0 ;
  assign y12278 = ~n42065 ;
  assign y12279 = n42071 ;
  assign y12280 = ~n42073 ;
  assign y12281 = ~n42076 ;
  assign y12282 = n42081 ;
  assign y12283 = ~n42083 ;
  assign y12284 = n42086 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = ~n42087 ;
  assign y12288 = ~1'b0 ;
  assign y12289 = n42089 ;
  assign y12290 = n42090 ;
  assign y12291 = n42092 ;
  assign y12292 = n42095 ;
  assign y12293 = ~1'b0 ;
  assign y12294 = ~n42101 ;
  assign y12295 = n42105 ;
  assign y12296 = ~n42108 ;
  assign y12297 = ~n42109 ;
  assign y12298 = n42113 ;
  assign y12299 = n42116 ;
  assign y12300 = ~n42118 ;
  assign y12301 = ~n42120 ;
  assign y12302 = n42123 ;
  assign y12303 = n42126 ;
  assign y12304 = n42133 ;
  assign y12305 = n42135 ;
  assign y12306 = n42140 ;
  assign y12307 = ~n42144 ;
  assign y12308 = n42146 ;
  assign y12309 = ~n42148 ;
  assign y12310 = n42149 ;
  assign y12311 = ~n42154 ;
  assign y12312 = ~n42165 ;
  assign y12313 = ~n42166 ;
  assign y12314 = ~n42169 ;
  assign y12315 = ~n42171 ;
  assign y12316 = n42175 ;
  assign y12317 = ~1'b0 ;
  assign y12318 = n42176 ;
  assign y12319 = ~n42178 ;
  assign y12320 = ~n42181 ;
  assign y12321 = ~n42182 ;
  assign y12322 = n42185 ;
  assign y12323 = n42187 ;
  assign y12324 = ~n42192 ;
  assign y12325 = n42194 ;
  assign y12326 = n42196 ;
  assign y12327 = n42199 ;
  assign y12328 = n42200 ;
  assign y12329 = n24099 ;
  assign y12330 = n42201 ;
  assign y12331 = ~n42202 ;
  assign y12332 = n42205 ;
  assign y12333 = n42206 ;
  assign y12334 = ~1'b0 ;
  assign y12335 = n42207 ;
  assign y12336 = ~n42208 ;
  assign y12337 = ~n42209 ;
  assign y12338 = ~n42210 ;
  assign y12339 = ~n42212 ;
  assign y12340 = n42215 ;
  assign y12341 = ~1'b0 ;
  assign y12342 = ~1'b0 ;
  assign y12343 = ~n42216 ;
  assign y12344 = ~n42219 ;
  assign y12345 = ~n13484 ;
  assign y12346 = ~n42222 ;
  assign y12347 = n42224 ;
  assign y12348 = n42225 ;
  assign y12349 = ~n42228 ;
  assign y12350 = n42232 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = n42233 ;
  assign y12353 = n42234 ;
  assign y12354 = n42248 ;
  assign y12355 = n42253 ;
  assign y12356 = ~n42258 ;
  assign y12357 = ~n42263 ;
  assign y12358 = n42265 ;
  assign y12359 = ~n42266 ;
  assign y12360 = ~n42271 ;
  assign y12361 = n42275 ;
  assign y12362 = ~1'b0 ;
  assign y12363 = ~n42280 ;
  assign y12364 = n42281 ;
  assign y12365 = n42282 ;
  assign y12366 = n42288 ;
  assign y12367 = ~n42291 ;
  assign y12368 = n42292 ;
  assign y12369 = ~1'b0 ;
  assign y12370 = ~1'b0 ;
  assign y12371 = ~n42295 ;
  assign y12372 = ~n42298 ;
  assign y12373 = n42302 ;
  assign y12374 = n42307 ;
  assign y12375 = ~n42308 ;
  assign y12376 = ~n42310 ;
  assign y12377 = n42313 ;
  assign y12378 = ~n42314 ;
  assign y12379 = n42315 ;
  assign y12380 = ~n42317 ;
  assign y12381 = n42319 ;
  assign y12382 = n42331 ;
  assign y12383 = ~n42332 ;
  assign y12384 = n42333 ;
  assign y12385 = n42335 ;
  assign y12386 = ~1'b0 ;
  assign y12387 = ~1'b0 ;
  assign y12388 = n42336 ;
  assign y12389 = n42338 ;
  assign y12390 = n42339 ;
  assign y12391 = ~n42341 ;
  assign y12392 = n42349 ;
  assign y12393 = n42353 ;
  assign y12394 = n42354 ;
  assign y12395 = ~n42357 ;
  assign y12396 = ~n42358 ;
  assign y12397 = ~n42361 ;
  assign y12398 = ~n42364 ;
  assign y12399 = ~n42366 ;
  assign y12400 = ~n42369 ;
  assign y12401 = n42371 ;
  assign y12402 = n42377 ;
  assign y12403 = n42384 ;
  assign y12404 = n42386 ;
  assign y12405 = n42389 ;
  assign y12406 = ~n42391 ;
  assign y12407 = ~n42392 ;
  assign y12408 = ~n42393 ;
  assign y12409 = ~1'b0 ;
  assign y12410 = n42396 ;
  assign y12411 = ~1'b0 ;
  assign y12412 = n42398 ;
  assign y12413 = ~n42401 ;
  assign y12414 = n23237 ;
  assign y12415 = ~n42402 ;
  assign y12416 = ~n42408 ;
  assign y12417 = n42410 ;
  assign y12418 = ~n42411 ;
  assign y12419 = n42412 ;
  assign y12420 = ~n42413 ;
  assign y12421 = ~n42414 ;
  assign y12422 = ~n42415 ;
  assign y12423 = n42419 ;
  assign y12424 = ~n42421 ;
  assign y12425 = ~1'b0 ;
  assign y12426 = n42422 ;
  assign y12427 = n42424 ;
  assign y12428 = n42428 ;
  assign y12429 = n42432 ;
  assign y12430 = ~n42433 ;
  assign y12431 = ~n42434 ;
  assign y12432 = ~n42436 ;
  assign y12433 = ~n42442 ;
  assign y12434 = ~n42445 ;
  assign y12435 = n42455 ;
  assign y12436 = ~n42458 ;
  assign y12437 = ~1'b0 ;
  assign y12438 = ~n42465 ;
  assign y12439 = n42466 ;
  assign y12440 = ~1'b0 ;
  assign y12441 = ~n42467 ;
  assign y12442 = ~n42468 ;
  assign y12443 = ~n42469 ;
  assign y12444 = ~n42470 ;
  assign y12445 = ~1'b0 ;
  assign y12446 = ~n42471 ;
  assign y12447 = ~n42473 ;
  assign y12448 = n42475 ;
  assign y12449 = ~n42477 ;
  assign y12450 = ~n42478 ;
  assign y12451 = ~n42480 ;
  assign y12452 = ~n42484 ;
  assign y12453 = n42485 ;
  assign y12454 = ~n42489 ;
  assign y12455 = n42491 ;
  assign y12456 = n42492 ;
  assign y12457 = n42494 ;
  assign y12458 = ~1'b0 ;
  assign y12459 = ~n42495 ;
  assign y12460 = ~n42505 ;
  assign y12461 = n42507 ;
  assign y12462 = n42511 ;
  assign y12463 = n42517 ;
  assign y12464 = ~1'b0 ;
  assign y12465 = ~1'b0 ;
  assign y12466 = n42518 ;
  assign y12467 = n16047 ;
  assign y12468 = n42519 ;
  assign y12469 = ~n42522 ;
  assign y12470 = ~n42527 ;
  assign y12471 = n42528 ;
  assign y12472 = n42536 ;
  assign y12473 = ~n42538 ;
  assign y12474 = ~n42546 ;
  assign y12475 = n42547 ;
  assign y12476 = ~n42549 ;
  assign y12477 = ~n42550 ;
  assign y12478 = n14906 ;
  assign y12479 = ~1'b0 ;
  assign y12480 = ~n42551 ;
  assign y12481 = n42552 ;
  assign y12482 = ~n42556 ;
  assign y12483 = n42560 ;
  assign y12484 = n42563 ;
  assign y12485 = n42565 ;
  assign y12486 = n42569 ;
  assign y12487 = ~n42571 ;
  assign y12488 = ~n42578 ;
  assign y12489 = n42580 ;
  assign y12490 = ~n42588 ;
  assign y12491 = ~n42597 ;
  assign y12492 = n42603 ;
  assign y12493 = ~n42606 ;
  assign y12494 = ~n42610 ;
  assign y12495 = ~n42615 ;
  assign y12496 = n42618 ;
  assign y12497 = n42620 ;
  assign y12498 = n42623 ;
  assign y12499 = ~1'b0 ;
  assign y12500 = n42626 ;
  assign y12501 = n42627 ;
  assign y12502 = ~n42629 ;
  assign y12503 = n42631 ;
  assign y12504 = ~n42633 ;
  assign y12505 = n42634 ;
  assign y12506 = ~1'b0 ;
  assign y12507 = ~n42638 ;
  assign y12508 = ~n42639 ;
  assign y12509 = n42641 ;
  assign y12510 = ~n42643 ;
  assign y12511 = ~n42650 ;
  assign y12512 = n42651 ;
  assign y12513 = n42653 ;
  assign y12514 = ~n42656 ;
  assign y12515 = n42658 ;
  assign y12516 = n42660 ;
  assign y12517 = n42663 ;
  assign y12518 = n42670 ;
  assign y12519 = n42673 ;
  assign y12520 = ~n42675 ;
  assign y12521 = ~n42676 ;
  assign y12522 = n42678 ;
  assign y12523 = ~1'b0 ;
  assign y12524 = n42680 ;
  assign y12525 = n42683 ;
  assign y12526 = n42685 ;
  assign y12527 = ~n42688 ;
  assign y12528 = n42689 ;
  assign y12529 = ~n42690 ;
  assign y12530 = n42691 ;
  assign y12531 = ~1'b0 ;
  assign y12532 = ~n42699 ;
  assign y12533 = ~1'b0 ;
  assign y12534 = n42700 ;
  assign y12535 = ~n42701 ;
  assign y12536 = ~n42702 ;
  assign y12537 = n42706 ;
  assign y12538 = ~n42711 ;
  assign y12539 = ~n42713 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = n42716 ;
  assign y12542 = ~n42720 ;
  assign y12543 = n42723 ;
  assign y12544 = n42726 ;
  assign y12545 = ~n42727 ;
  assign y12546 = n42730 ;
  assign y12547 = ~n42732 ;
  assign y12548 = ~n42733 ;
  assign y12549 = n42740 ;
  assign y12550 = ~n42741 ;
  assign y12551 = n42744 ;
  assign y12552 = ~n42746 ;
  assign y12553 = n42749 ;
  assign y12554 = ~n42754 ;
  assign y12555 = ~n42755 ;
  assign y12556 = ~n42757 ;
  assign y12557 = n42762 ;
  assign y12558 = n25461 ;
  assign y12559 = ~n42767 ;
  assign y12560 = ~n42771 ;
  assign y12561 = ~1'b0 ;
  assign y12562 = ~1'b0 ;
  assign y12563 = n42774 ;
  assign y12564 = ~n42776 ;
  assign y12565 = n42782 ;
  assign y12566 = ~n42790 ;
  assign y12567 = n42794 ;
  assign y12568 = ~n42796 ;
  assign y12569 = ~n42797 ;
  assign y12570 = n42799 ;
  assign y12571 = ~n42804 ;
  assign y12572 = ~n42805 ;
  assign y12573 = ~n42810 ;
  assign y12574 = ~n42811 ;
  assign y12575 = n42813 ;
  assign y12576 = n42815 ;
  assign y12577 = n42817 ;
  assign y12578 = ~1'b0 ;
  assign y12579 = ~1'b0 ;
  assign y12580 = ~n42818 ;
  assign y12581 = ~n42821 ;
  assign y12582 = n42822 ;
  assign y12583 = n42823 ;
  assign y12584 = ~n42825 ;
  assign y12585 = ~1'b0 ;
  assign y12586 = n42828 ;
  assign y12587 = ~n42830 ;
  assign y12588 = ~n42832 ;
  assign y12589 = ~n42838 ;
  assign y12590 = n42840 ;
  assign y12591 = ~n42841 ;
  assign y12592 = ~n42844 ;
  assign y12593 = n42845 ;
  assign y12594 = n42853 ;
  assign y12595 = ~n42856 ;
  assign y12596 = n42860 ;
  assign y12597 = n42863 ;
  assign y12598 = ~n42867 ;
  assign y12599 = ~n42868 ;
  assign y12600 = n42869 ;
  assign y12601 = ~n42871 ;
  assign y12602 = n42877 ;
  assign y12603 = ~n42878 ;
  assign y12604 = n42879 ;
  assign y12605 = n42881 ;
  assign y12606 = ~1'b0 ;
  assign y12607 = ~n42883 ;
  assign y12608 = n42888 ;
  assign y12609 = n42890 ;
  assign y12610 = ~n42891 ;
  assign y12611 = ~n14314 ;
  assign y12612 = n42893 ;
  assign y12613 = ~n42896 ;
  assign y12614 = n42897 ;
  assign y12615 = n42898 ;
  assign y12616 = n42901 ;
  assign y12617 = ~n42902 ;
  assign y12618 = n42907 ;
  assign y12619 = n42908 ;
  assign y12620 = ~n42909 ;
  assign y12621 = n42911 ;
  assign y12622 = n42913 ;
  assign y12623 = ~n42915 ;
  assign y12624 = n42916 ;
  assign y12625 = n42922 ;
  assign y12626 = ~n42923 ;
  assign y12627 = n42924 ;
  assign y12628 = n42929 ;
  assign y12629 = ~n42930 ;
  assign y12630 = ~n42931 ;
  assign y12631 = n42935 ;
  assign y12632 = n42937 ;
  assign y12633 = n42938 ;
  assign y12634 = ~n42940 ;
  assign y12635 = ~1'b0 ;
  assign y12636 = ~n42943 ;
  assign y12637 = n42949 ;
  assign y12638 = n42952 ;
  assign y12639 = ~n42953 ;
  assign y12640 = ~n42956 ;
  assign y12641 = ~n42957 ;
  assign y12642 = n42958 ;
  assign y12643 = ~1'b0 ;
  assign y12644 = ~1'b0 ;
  assign y12645 = n42961 ;
  assign y12646 = ~n42965 ;
  assign y12647 = ~n42966 ;
  assign y12648 = ~n42967 ;
  assign y12649 = n42969 ;
  assign y12650 = ~n42970 ;
  assign y12651 = ~n42972 ;
  assign y12652 = n42974 ;
  assign y12653 = n27128 ;
  assign y12654 = n42976 ;
  assign y12655 = n42978 ;
  assign y12656 = ~n42979 ;
  assign y12657 = n42982 ;
  assign y12658 = ~1'b0 ;
  assign y12659 = n42983 ;
  assign y12660 = n42986 ;
  assign y12661 = ~n42987 ;
  assign y12662 = ~n12187 ;
  assign y12663 = n42988 ;
  assign y12664 = ~n42989 ;
  assign y12665 = n4724 ;
  assign y12666 = ~n42991 ;
  assign y12667 = n42998 ;
  assign y12668 = ~n43000 ;
  assign y12669 = ~n43005 ;
  assign y12670 = n43008 ;
  assign y12671 = ~n43010 ;
  assign y12672 = n43011 ;
  assign y12673 = n43012 ;
  assign y12674 = ~n43013 ;
  assign y12675 = ~n43015 ;
  assign y12676 = ~n43018 ;
  assign y12677 = n43025 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = n43026 ;
  assign y12680 = ~n43029 ;
  assign y12681 = ~n43033 ;
  assign y12682 = ~n43034 ;
  assign y12683 = ~n43036 ;
  assign y12684 = n43039 ;
  assign y12685 = n43046 ;
  assign y12686 = ~1'b0 ;
  assign y12687 = ~n43049 ;
  assign y12688 = n43056 ;
  assign y12689 = ~n43057 ;
  assign y12690 = n43061 ;
  assign y12691 = n43062 ;
  assign y12692 = ~n43068 ;
  assign y12693 = ~n43070 ;
  assign y12694 = n43071 ;
  assign y12695 = ~1'b0 ;
  assign y12696 = n43073 ;
  assign y12697 = n43077 ;
  assign y12698 = n43080 ;
  assign y12699 = ~n43083 ;
  assign y12700 = ~n43085 ;
  assign y12701 = n43088 ;
  assign y12702 = ~n43089 ;
  assign y12703 = n43092 ;
  assign y12704 = ~1'b0 ;
  assign y12705 = n43094 ;
  assign y12706 = ~n43101 ;
  assign y12707 = ~n43102 ;
  assign y12708 = n43103 ;
  assign y12709 = ~n43104 ;
  assign y12710 = n43105 ;
  assign y12711 = ~n43107 ;
  assign y12712 = ~n43110 ;
  assign y12713 = n43112 ;
  assign y12714 = ~n43113 ;
  assign y12715 = n43117 ;
  assign y12716 = n43120 ;
  assign y12717 = ~n43125 ;
  assign y12718 = ~n43127 ;
  assign y12719 = ~1'b0 ;
  assign y12720 = ~1'b0 ;
  assign y12721 = n43130 ;
  assign y12722 = n43131 ;
  assign y12723 = ~n43132 ;
  assign y12724 = n43134 ;
  assign y12725 = ~n43135 ;
  assign y12726 = n43138 ;
  assign y12727 = ~n43139 ;
  assign y12728 = ~n43141 ;
  assign y12729 = ~1'b0 ;
  assign y12730 = ~1'b0 ;
  assign y12731 = ~n43142 ;
  assign y12732 = n43144 ;
  assign y12733 = ~n43145 ;
  assign y12734 = n43148 ;
  assign y12735 = n43152 ;
  assign y12736 = n43153 ;
  assign y12737 = ~n43158 ;
  assign y12738 = ~n43161 ;
  assign y12739 = ~n43163 ;
  assign y12740 = n43166 ;
  assign y12741 = n43169 ;
  assign y12742 = ~n43173 ;
  assign y12743 = ~n43176 ;
  assign y12744 = n43182 ;
  assign y12745 = n43183 ;
  assign y12746 = ~n43186 ;
  assign y12747 = ~n43189 ;
  assign y12748 = ~n43190 ;
  assign y12749 = ~n43193 ;
  assign y12750 = n43194 ;
  assign y12751 = ~n43195 ;
  assign y12752 = ~n43199 ;
  assign y12753 = ~n43201 ;
  assign y12754 = n43202 ;
  assign y12755 = n43204 ;
  assign y12756 = n43206 ;
  assign y12757 = ~n43207 ;
  assign y12758 = n43211 ;
  assign y12759 = ~n43214 ;
  assign y12760 = ~n43220 ;
  assign y12761 = n43223 ;
  assign y12762 = n43228 ;
  assign y12763 = ~n43232 ;
  assign y12764 = n43234 ;
  assign y12765 = n43235 ;
  assign y12766 = n43236 ;
  assign y12767 = n43239 ;
  assign y12768 = ~n43245 ;
  assign y12769 = ~n43251 ;
  assign y12770 = ~n43258 ;
  assign y12771 = n43260 ;
  assign y12772 = ~n43262 ;
  assign y12773 = n43263 ;
  assign y12774 = n43266 ;
  assign y12775 = n43270 ;
  assign y12776 = ~1'b0 ;
  assign y12777 = ~n43274 ;
  assign y12778 = n43276 ;
  assign y12779 = ~n43277 ;
  assign y12780 = ~n5192 ;
  assign y12781 = n43281 ;
  assign y12782 = ~n43282 ;
  assign y12783 = n43285 ;
  assign y12784 = 1'b0 ;
  assign y12785 = n43287 ;
  assign y12786 = ~n43289 ;
  assign y12787 = n43294 ;
  assign y12788 = ~n43295 ;
  assign y12789 = n43300 ;
  assign y12790 = n43303 ;
  assign y12791 = n43307 ;
  assign y12792 = ~n43313 ;
  assign y12793 = ~n43318 ;
  assign y12794 = n43319 ;
  assign y12795 = n43320 ;
  assign y12796 = n43321 ;
  assign y12797 = n43322 ;
  assign y12798 = n43325 ;
  assign y12799 = n43327 ;
  assign y12800 = n43329 ;
  assign y12801 = ~n43332 ;
  assign y12802 = ~n43334 ;
  assign y12803 = ~n43338 ;
  assign y12804 = n43341 ;
  assign y12805 = ~n43346 ;
  assign y12806 = ~n43347 ;
  assign y12807 = ~n43350 ;
  assign y12808 = ~n43351 ;
  assign y12809 = n43353 ;
  assign y12810 = n43354 ;
  assign y12811 = n43359 ;
  assign y12812 = n43360 ;
  assign y12813 = ~n43361 ;
  assign y12814 = ~n43364 ;
  assign y12815 = ~n43367 ;
  assign y12816 = n43369 ;
  assign y12817 = ~n43371 ;
  assign y12818 = ~1'b0 ;
  assign y12819 = ~n43372 ;
  assign y12820 = n43374 ;
  assign y12821 = n43378 ;
  assign y12822 = n43379 ;
  assign y12823 = ~n43381 ;
  assign y12824 = ~n43384 ;
  assign y12825 = ~n43385 ;
  assign y12826 = ~n43386 ;
  assign y12827 = ~n43389 ;
  assign y12828 = ~n43391 ;
  assign y12829 = ~n43395 ;
  assign y12830 = n43397 ;
  assign y12831 = ~n43400 ;
  assign y12832 = n43404 ;
  assign y12833 = ~n43409 ;
  assign y12834 = n43416 ;
  assign y12835 = ~n43417 ;
  assign y12836 = n43424 ;
  assign y12837 = ~n43428 ;
  assign y12838 = ~n43429 ;
  assign y12839 = n43430 ;
  assign y12840 = ~n43431 ;
  assign y12841 = ~1'b0 ;
  assign y12842 = ~n43432 ;
  assign y12843 = ~n43435 ;
  assign y12844 = n43438 ;
  assign y12845 = ~n43448 ;
  assign y12846 = ~n43457 ;
  assign y12847 = ~n43462 ;
  assign y12848 = n43463 ;
  assign y12849 = ~n43466 ;
  assign y12850 = ~1'b0 ;
  assign y12851 = ~n43468 ;
  assign y12852 = n43471 ;
  assign y12853 = ~n43474 ;
  assign y12854 = ~n43477 ;
  assign y12855 = ~n43478 ;
  assign y12856 = ~n43482 ;
  assign y12857 = ~1'b0 ;
  assign y12858 = n43487 ;
  assign y12859 = ~n43488 ;
  assign y12860 = ~n17710 ;
  assign y12861 = ~n43491 ;
  assign y12862 = ~n43492 ;
  assign y12863 = ~n43494 ;
  assign y12864 = ~n43498 ;
  assign y12865 = n43500 ;
  assign y12866 = n43502 ;
  assign y12867 = ~n43504 ;
  assign y12868 = ~n43505 ;
  assign y12869 = ~n43510 ;
  assign y12870 = n43511 ;
  assign y12871 = n43517 ;
  assign y12872 = n43519 ;
  assign y12873 = n43524 ;
  assign y12874 = ~n43527 ;
  assign y12875 = ~n43533 ;
  assign y12876 = n43534 ;
  assign y12877 = n43536 ;
  assign y12878 = ~n43538 ;
  assign y12879 = n43539 ;
  assign y12880 = n43540 ;
  assign y12881 = n43541 ;
  assign y12882 = n43542 ;
  assign y12883 = ~n43548 ;
  assign y12884 = n43550 ;
  assign y12885 = ~n43553 ;
  assign y12886 = n43555 ;
  assign y12887 = n43556 ;
  assign y12888 = ~n43557 ;
  assign y12889 = n43561 ;
  assign y12890 = n43568 ;
  assign y12891 = ~1'b0 ;
  assign y12892 = n43570 ;
  assign y12893 = ~n43571 ;
  assign y12894 = n43572 ;
  assign y12895 = n43573 ;
  assign y12896 = ~n43575 ;
  assign y12897 = ~n43579 ;
  assign y12898 = n43582 ;
  assign y12899 = n43584 ;
  assign y12900 = n43586 ;
  assign y12901 = n43589 ;
  assign y12902 = ~n43597 ;
  assign y12903 = ~n43598 ;
  assign y12904 = n43602 ;
  assign y12905 = n43605 ;
  assign y12906 = n43608 ;
  assign y12907 = ~n43618 ;
  assign y12908 = n43621 ;
  assign y12909 = n43623 ;
  assign y12910 = ~n43624 ;
  assign y12911 = n43625 ;
  assign y12912 = ~n43626 ;
  assign y12913 = ~n43627 ;
  assign y12914 = ~n43628 ;
  assign y12915 = ~n43630 ;
  assign y12916 = ~n43632 ;
  assign y12917 = ~1'b0 ;
  assign y12918 = ~n43633 ;
  assign y12919 = n43634 ;
  assign y12920 = ~n43637 ;
  assign y12921 = ~1'b0 ;
  assign y12922 = ~1'b0 ;
  assign y12923 = n43640 ;
  assign y12924 = ~1'b0 ;
  assign y12925 = ~n43644 ;
  assign y12926 = ~n43646 ;
  assign y12927 = ~n43649 ;
  assign y12928 = ~1'b0 ;
  assign y12929 = ~n43651 ;
  assign y12930 = n43663 ;
  assign y12931 = ~n43668 ;
  assign y12932 = n43670 ;
  assign y12933 = n43672 ;
  assign y12934 = ~n43674 ;
  assign y12935 = n43676 ;
  assign y12936 = ~1'b0 ;
  assign y12937 = ~n43677 ;
  assign y12938 = ~n43681 ;
  assign y12939 = n43686 ;
  assign y12940 = ~n43687 ;
  assign y12941 = ~n43689 ;
  assign y12942 = ~1'b0 ;
  assign y12943 = ~n43692 ;
  assign y12944 = ~n43696 ;
  assign y12945 = ~n43703 ;
  assign y12946 = ~n43708 ;
  assign y12947 = ~n43711 ;
  assign y12948 = n43714 ;
  assign y12949 = n43716 ;
  assign y12950 = n43718 ;
  assign y12951 = n43720 ;
  assign y12952 = ~n43721 ;
  assign y12953 = ~n43722 ;
  assign y12954 = ~n11619 ;
  assign y12955 = n43726 ;
  assign y12956 = n43727 ;
  assign y12957 = ~n43728 ;
  assign y12958 = ~n43736 ;
  assign y12959 = ~1'b0 ;
  assign y12960 = ~n40167 ;
  assign y12961 = ~n43737 ;
  assign y12962 = n43741 ;
  assign y12963 = ~n43743 ;
  assign y12964 = n43744 ;
  assign y12965 = ~n43746 ;
  assign y12966 = n43753 ;
  assign y12967 = ~n43758 ;
  assign y12968 = n43759 ;
  assign y12969 = ~n43761 ;
  assign y12970 = n43764 ;
  assign y12971 = ~1'b0 ;
  assign y12972 = n43766 ;
  assign y12973 = ~n43768 ;
  assign y12974 = ~1'b0 ;
  assign y12975 = ~n43770 ;
  assign y12976 = n43771 ;
  assign y12977 = n43772 ;
  assign y12978 = n43777 ;
  assign y12979 = ~n43779 ;
  assign y12980 = ~1'b0 ;
  assign y12981 = n43781 ;
  assign y12982 = ~n43786 ;
  assign y12983 = ~n43790 ;
  assign y12984 = ~n43791 ;
  assign y12985 = ~n43795 ;
  assign y12986 = ~n43799 ;
  assign y12987 = n43801 ;
  assign y12988 = ~1'b0 ;
  assign y12989 = ~n43804 ;
  assign y12990 = ~n43807 ;
  assign y12991 = ~n43811 ;
  assign y12992 = ~n43812 ;
  assign y12993 = n43815 ;
  assign y12994 = ~n43818 ;
  assign y12995 = n43821 ;
  assign y12996 = n43823 ;
  assign y12997 = ~n43826 ;
  assign y12998 = n43828 ;
  assign y12999 = ~n43831 ;
  assign y13000 = n43833 ;
  assign y13001 = n43834 ;
  assign y13002 = n43837 ;
  assign y13003 = n43839 ;
  assign y13004 = ~1'b0 ;
  assign y13005 = ~n43842 ;
  assign y13006 = n43845 ;
  assign y13007 = ~n43846 ;
  assign y13008 = n43847 ;
  assign y13009 = n43849 ;
  assign y13010 = ~n43854 ;
  assign y13011 = ~n43857 ;
  assign y13012 = n43859 ;
  assign y13013 = n43860 ;
  assign y13014 = ~n43864 ;
  assign y13015 = ~n43866 ;
  assign y13016 = n43871 ;
  assign y13017 = n43875 ;
  assign y13018 = ~n43876 ;
  assign y13019 = n43878 ;
  assign y13020 = ~n43879 ;
  assign y13021 = ~n43880 ;
  assign y13022 = ~n43881 ;
  assign y13023 = n13547 ;
  assign y13024 = ~n43885 ;
  assign y13025 = n43887 ;
  assign y13026 = ~n43888 ;
  assign y13027 = ~n43890 ;
  assign y13028 = ~n43892 ;
  assign y13029 = ~1'b0 ;
  assign y13030 = ~n43894 ;
  assign y13031 = ~1'b0 ;
  assign y13032 = ~1'b0 ;
  assign y13033 = ~n43896 ;
  assign y13034 = ~n43901 ;
  assign y13035 = n43902 ;
  assign y13036 = ~n14930 ;
  assign y13037 = ~n43903 ;
  assign y13038 = ~n3336 ;
  assign y13039 = n43907 ;
  assign y13040 = ~n43911 ;
  assign y13041 = ~n43912 ;
  assign y13042 = ~n43913 ;
  assign y13043 = n43917 ;
  assign y13044 = n43918 ;
  assign y13045 = ~n43921 ;
  assign y13046 = ~n43924 ;
  assign y13047 = n43926 ;
  assign y13048 = 1'b0 ;
  assign y13049 = n43928 ;
  assign y13050 = n43929 ;
  assign y13051 = ~n43932 ;
  assign y13052 = ~n43933 ;
  assign y13053 = n43938 ;
  assign y13054 = ~n43940 ;
  assign y13055 = ~n43945 ;
  assign y13056 = ~n43948 ;
  assign y13057 = ~n43952 ;
  assign y13058 = n43955 ;
  assign y13059 = n43956 ;
  assign y13060 = n43959 ;
  assign y13061 = n43960 ;
  assign y13062 = ~n43963 ;
  assign y13063 = n43964 ;
  assign y13064 = n43968 ;
  assign y13065 = ~n43969 ;
  assign y13066 = n43970 ;
  assign y13067 = ~n43974 ;
  assign y13068 = ~n43976 ;
  assign y13069 = ~1'b0 ;
  assign y13070 = n43977 ;
  assign y13071 = ~n43978 ;
  assign y13072 = ~n43979 ;
  assign y13073 = ~n43980 ;
  assign y13074 = ~n43981 ;
  assign y13075 = ~n32853 ;
  assign y13076 = ~1'b0 ;
  assign y13077 = ~n43983 ;
  assign y13078 = n43986 ;
  assign y13079 = ~n43990 ;
  assign y13080 = ~n43993 ;
  assign y13081 = ~n43997 ;
  assign y13082 = n44000 ;
  assign y13083 = ~n44002 ;
  assign y13084 = n44004 ;
  assign y13085 = ~n44005 ;
  assign y13086 = ~n44008 ;
  assign y13087 = n44016 ;
  assign y13088 = ~n44018 ;
  assign y13089 = ~n44021 ;
  assign y13090 = ~n44026 ;
  assign y13091 = ~1'b0 ;
  assign y13092 = ~1'b0 ;
  assign y13093 = ~n44028 ;
  assign y13094 = ~n44030 ;
  assign y13095 = n44032 ;
  assign y13096 = n44035 ;
  assign y13097 = ~n44037 ;
  assign y13098 = ~n44039 ;
  assign y13099 = ~1'b0 ;
  assign y13100 = ~1'b0 ;
  assign y13101 = ~1'b0 ;
  assign y13102 = n44040 ;
  assign y13103 = ~n44042 ;
  assign y13104 = n44045 ;
  assign y13105 = ~n44046 ;
  assign y13106 = ~n44050 ;
  assign y13107 = n44052 ;
  assign y13108 = n44057 ;
  assign y13109 = ~n44059 ;
  assign y13110 = n44061 ;
  assign y13111 = n44062 ;
  assign y13112 = n44065 ;
  assign y13113 = n44066 ;
  assign y13114 = n44068 ;
  assign y13115 = ~n44069 ;
  assign y13116 = ~n44071 ;
  assign y13117 = n44075 ;
  assign y13118 = n44076 ;
  assign y13119 = ~1'b0 ;
  assign y13120 = ~n44084 ;
  assign y13121 = ~n38443 ;
  assign y13122 = ~n44085 ;
  assign y13123 = n44086 ;
  assign y13124 = ~n44089 ;
  assign y13125 = ~n44098 ;
  assign y13126 = ~n44099 ;
  assign y13127 = n44101 ;
  assign y13128 = n44103 ;
  assign y13129 = ~1'b0 ;
  assign y13130 = n44105 ;
  assign y13131 = ~n44107 ;
  assign y13132 = n44109 ;
  assign y13133 = n44111 ;
  assign y13134 = n44115 ;
  assign y13135 = ~n44117 ;
  assign y13136 = ~n44118 ;
  assign y13137 = n44122 ;
  assign y13138 = n44124 ;
  assign y13139 = n44126 ;
  assign y13140 = ~1'b0 ;
  assign y13141 = ~n44129 ;
  assign y13142 = n44132 ;
  assign y13143 = ~n44134 ;
  assign y13144 = n44139 ;
  assign y13145 = n44142 ;
  assign y13146 = n44145 ;
  assign y13147 = ~n44147 ;
  assign y13148 = ~1'b0 ;
  assign y13149 = n44149 ;
  assign y13150 = ~n44150 ;
  assign y13151 = n44151 ;
  assign y13152 = ~n44152 ;
  assign y13153 = n44155 ;
  assign y13154 = ~1'b0 ;
  assign y13155 = n44160 ;
  assign y13156 = n44164 ;
  assign y13157 = ~n44165 ;
  assign y13158 = n44167 ;
  assign y13159 = ~n44168 ;
  assign y13160 = n44170 ;
  assign y13161 = ~1'b0 ;
  assign y13162 = n44171 ;
  assign y13163 = ~n44173 ;
  assign y13164 = ~n44177 ;
  assign y13165 = n44178 ;
  assign y13166 = ~n44179 ;
  assign y13167 = n44180 ;
  assign y13168 = n44183 ;
  assign y13169 = ~n44191 ;
  assign y13170 = n44193 ;
  assign y13171 = ~n44195 ;
  assign y13172 = ~n44197 ;
  assign y13173 = ~n44200 ;
  assign y13174 = ~n44204 ;
  assign y13175 = n18768 ;
  assign y13176 = ~n44205 ;
  assign y13177 = n44207 ;
  assign y13178 = n44208 ;
  assign y13179 = ~1'b0 ;
  assign y13180 = ~1'b0 ;
  assign y13181 = ~n44211 ;
  assign y13182 = ~n44213 ;
  assign y13183 = n44214 ;
  assign y13184 = n44216 ;
  assign y13185 = n44217 ;
  assign y13186 = n44219 ;
  assign y13187 = n44229 ;
  assign y13188 = n44231 ;
  assign y13189 = ~n44238 ;
  assign y13190 = ~1'b0 ;
  assign y13191 = ~n44240 ;
  assign y13192 = ~n44241 ;
  assign y13193 = ~n44245 ;
  assign y13194 = n44248 ;
  assign y13195 = n44251 ;
  assign y13196 = n44255 ;
  assign y13197 = ~n44258 ;
  assign y13198 = ~1'b0 ;
  assign y13199 = ~n44260 ;
  assign y13200 = n44261 ;
  assign y13201 = n44263 ;
  assign y13202 = n44266 ;
  assign y13203 = ~n44267 ;
  assign y13204 = n44268 ;
  assign y13205 = n44277 ;
  assign y13206 = n44280 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = ~n44281 ;
  assign y13209 = n44282 ;
  assign y13210 = n44284 ;
  assign y13211 = ~n44286 ;
  assign y13212 = ~n44291 ;
  assign y13213 = ~n44294 ;
  assign y13214 = n44298 ;
  assign y13215 = ~n44300 ;
  assign y13216 = n44301 ;
  assign y13217 = n44302 ;
  assign y13218 = n44303 ;
  assign y13219 = ~n44304 ;
  assign y13220 = ~n44305 ;
  assign y13221 = ~n44307 ;
  assign y13222 = n44312 ;
  assign y13223 = ~1'b0 ;
  assign y13224 = ~n44314 ;
  assign y13225 = n44315 ;
  assign y13226 = ~n6933 ;
  assign y13227 = ~n44317 ;
  assign y13228 = n44321 ;
  assign y13229 = ~n44326 ;
  assign y13230 = ~n44328 ;
  assign y13231 = n44330 ;
  assign y13232 = ~1'b0 ;
  assign y13233 = ~1'b0 ;
  assign y13234 = n44332 ;
  assign y13235 = ~n44333 ;
  assign y13236 = n44335 ;
  assign y13237 = ~n44337 ;
  assign y13238 = ~n44339 ;
  assign y13239 = ~n44340 ;
  assign y13240 = n44344 ;
  assign y13241 = ~1'b0 ;
  assign y13242 = n44346 ;
  assign y13243 = ~n44348 ;
  assign y13244 = ~n44357 ;
  assign y13245 = n44358 ;
  assign y13246 = n44359 ;
  assign y13247 = n44362 ;
  assign y13248 = ~n44364 ;
  assign y13249 = ~1'b0 ;
  assign y13250 = ~1'b0 ;
  assign y13251 = ~n44368 ;
  assign y13252 = n44370 ;
  assign y13253 = ~n44371 ;
  assign y13254 = n44379 ;
  assign y13255 = ~n44380 ;
  assign y13256 = ~n44383 ;
  assign y13257 = ~1'b0 ;
  assign y13258 = n44388 ;
  assign y13259 = n44389 ;
  assign y13260 = ~n44392 ;
  assign y13261 = ~n44393 ;
  assign y13262 = n44401 ;
  assign y13263 = ~n44405 ;
  assign y13264 = ~n40906 ;
  assign y13265 = ~1'b0 ;
  assign y13266 = ~1'b0 ;
  assign y13267 = ~n44407 ;
  assign y13268 = ~n44408 ;
  assign y13269 = ~n44413 ;
  assign y13270 = ~n44418 ;
  assign y13271 = ~1'b0 ;
  assign y13272 = ~1'b0 ;
  assign y13273 = ~n44420 ;
  assign y13274 = ~n44422 ;
  assign y13275 = n44423 ;
  assign y13276 = ~n44427 ;
  assign y13277 = ~n44428 ;
  assign y13278 = ~n44431 ;
  assign y13279 = n44434 ;
  assign y13280 = n44436 ;
  assign y13281 = ~n44438 ;
  assign y13282 = ~1'b0 ;
  assign y13283 = n44440 ;
  assign y13284 = n44441 ;
  assign y13285 = n44443 ;
  assign y13286 = n44444 ;
  assign y13287 = n44447 ;
  assign y13288 = ~n44448 ;
  assign y13289 = ~n44452 ;
  assign y13290 = n44455 ;
  assign y13291 = ~1'b0 ;
  assign y13292 = n44458 ;
  assign y13293 = ~n44462 ;
  assign y13294 = n44468 ;
  assign y13295 = n44470 ;
  assign y13296 = n44471 ;
  assign y13297 = ~n44472 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~n44473 ;
  assign y13300 = ~n44474 ;
  assign y13301 = ~n44475 ;
  assign y13302 = ~n44478 ;
  assign y13303 = ~n44480 ;
  assign y13304 = ~n44481 ;
  assign y13305 = n44484 ;
  assign y13306 = ~n44486 ;
  assign y13307 = ~n44487 ;
  assign y13308 = n44488 ;
  assign y13309 = n44490 ;
  assign y13310 = n44491 ;
  assign y13311 = ~n44494 ;
  assign y13312 = ~n44495 ;
  assign y13313 = ~n44497 ;
  assign y13314 = ~1'b0 ;
  assign y13315 = ~n44498 ;
  assign y13316 = n44501 ;
  assign y13317 = n44503 ;
  assign y13318 = n44507 ;
  assign y13319 = n44510 ;
  assign y13320 = ~n44512 ;
  assign y13321 = ~1'b0 ;
  assign y13322 = n44517 ;
  assign y13323 = n44521 ;
  assign y13324 = n44524 ;
  assign y13325 = n44525 ;
  assign y13326 = n44526 ;
  assign y13327 = ~n44529 ;
  assign y13328 = n44531 ;
  assign y13329 = ~1'b0 ;
  assign y13330 = n44536 ;
  assign y13331 = n44537 ;
  assign y13332 = ~n44539 ;
  assign y13333 = n44540 ;
  assign y13334 = n44541 ;
  assign y13335 = ~n44543 ;
  assign y13336 = ~n44545 ;
  assign y13337 = ~n44549 ;
  assign y13338 = ~n44551 ;
  assign y13339 = ~n44554 ;
  assign y13340 = n44556 ;
  assign y13341 = ~n44559 ;
  assign y13342 = ~n44562 ;
  assign y13343 = n44564 ;
  assign y13344 = n44568 ;
  assign y13345 = n44574 ;
  assign y13346 = n44576 ;
  assign y13347 = ~1'b0 ;
  assign y13348 = ~1'b0 ;
  assign y13349 = ~1'b0 ;
  assign y13350 = n44580 ;
  assign y13351 = n44581 ;
  assign y13352 = n44583 ;
  assign y13353 = n44587 ;
  assign y13354 = ~n44588 ;
  assign y13355 = n44591 ;
  assign y13356 = ~1'b0 ;
  assign y13357 = ~1'b0 ;
  assign y13358 = n44595 ;
  assign y13359 = n44599 ;
  assign y13360 = n44601 ;
  assign y13361 = ~n44602 ;
  assign y13362 = n44604 ;
  assign y13363 = ~n44605 ;
  assign y13364 = n44607 ;
  assign y13365 = ~1'b0 ;
  assign y13366 = ~1'b0 ;
  assign y13367 = ~1'b0 ;
  assign y13368 = n44609 ;
  assign y13369 = ~n44610 ;
  assign y13370 = n44611 ;
  assign y13371 = n44612 ;
  assign y13372 = ~n44615 ;
  assign y13373 = n44619 ;
  assign y13374 = ~n44622 ;
  assign y13375 = n44626 ;
  assign y13376 = n44630 ;
  assign y13377 = ~n44633 ;
  assign y13378 = n44637 ;
  assign y13379 = ~n44643 ;
  assign y13380 = n44645 ;
  assign y13381 = ~n44651 ;
  assign y13382 = ~1'b0 ;
  assign y13383 = n44652 ;
  assign y13384 = n44660 ;
  assign y13385 = n44661 ;
  assign y13386 = n44664 ;
  assign y13387 = n44667 ;
  assign y13388 = n44668 ;
  assign y13389 = n44672 ;
  assign y13390 = n44674 ;
  assign y13391 = n44676 ;
  assign y13392 = ~n44678 ;
  assign y13393 = ~n44679 ;
  assign y13394 = ~n44684 ;
  assign y13395 = n44687 ;
  assign y13396 = ~n44690 ;
  assign y13397 = n44692 ;
  assign y13398 = ~n44694 ;
  assign y13399 = n44698 ;
  assign y13400 = ~n44699 ;
  assign y13401 = ~n44703 ;
  assign y13402 = ~n44708 ;
  assign y13403 = n44713 ;
  assign y13404 = ~n44714 ;
  assign y13405 = n44718 ;
  assign y13406 = ~1'b0 ;
  assign y13407 = ~n44719 ;
  assign y13408 = n44721 ;
  assign y13409 = n44722 ;
  assign y13410 = ~n44723 ;
  assign y13411 = n44724 ;
  assign y13412 = ~n44725 ;
  assign y13413 = ~n44727 ;
  assign y13414 = n44732 ;
  assign y13415 = ~1'b0 ;
  assign y13416 = ~n44734 ;
  assign y13417 = ~n44736 ;
  assign y13418 = ~n44738 ;
  assign y13419 = n44740 ;
  assign y13420 = n44745 ;
  assign y13421 = n44746 ;
  assign y13422 = n44749 ;
  assign y13423 = ~n44754 ;
  assign y13424 = ~n44756 ;
  assign y13425 = ~1'b0 ;
  assign y13426 = ~n44758 ;
  assign y13427 = ~1'b0 ;
  assign y13428 = ~n44762 ;
  assign y13429 = ~n44764 ;
  assign y13430 = n44765 ;
  assign y13431 = ~n44766 ;
  assign y13432 = n44767 ;
  assign y13433 = n44772 ;
  assign y13434 = ~n44775 ;
  assign y13435 = n44777 ;
  assign y13436 = n44780 ;
  assign y13437 = n44782 ;
  assign y13438 = ~n44785 ;
  assign y13439 = ~n44787 ;
  assign y13440 = ~n44788 ;
  assign y13441 = n44790 ;
  assign y13442 = ~n44791 ;
  assign y13443 = n44797 ;
  assign y13444 = ~1'b0 ;
  assign y13445 = n44798 ;
  assign y13446 = n44799 ;
  assign y13447 = n44804 ;
  assign y13448 = ~n44807 ;
  assign y13449 = n44808 ;
  assign y13450 = n44809 ;
  assign y13451 = n44810 ;
  assign y13452 = ~1'b0 ;
  assign y13453 = n44814 ;
  assign y13454 = n44820 ;
  assign y13455 = ~n44821 ;
  assign y13456 = n44822 ;
  assign y13457 = n44824 ;
  assign y13458 = ~n44828 ;
  assign y13459 = ~1'b0 ;
  assign y13460 = ~n44833 ;
  assign y13461 = n44835 ;
  assign y13462 = n44837 ;
  assign y13463 = ~n44839 ;
  assign y13464 = ~n44840 ;
  assign y13465 = n44841 ;
  assign y13466 = ~n44845 ;
  assign y13467 = ~n44848 ;
  assign y13468 = n44856 ;
  assign y13469 = ~n44859 ;
  assign y13470 = ~1'b0 ;
  assign y13471 = ~n44861 ;
  assign y13472 = ~n44866 ;
  assign y13473 = n44867 ;
  assign y13474 = ~n44868 ;
  assign y13475 = ~n44870 ;
  assign y13476 = n44873 ;
  assign y13477 = n44874 ;
  assign y13478 = n44875 ;
  assign y13479 = n44877 ;
  assign y13480 = n44884 ;
  assign y13481 = n44885 ;
  assign y13482 = n44887 ;
  assign y13483 = n44890 ;
  assign y13484 = ~n44891 ;
  assign y13485 = ~n44894 ;
  assign y13486 = ~n44895 ;
  assign y13487 = ~1'b0 ;
  assign y13488 = ~1'b0 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = n44897 ;
  assign y13491 = ~n44900 ;
  assign y13492 = ~n44903 ;
  assign y13493 = ~n44912 ;
  assign y13494 = ~n44915 ;
  assign y13495 = ~n44917 ;
  assign y13496 = ~n44919 ;
  assign y13497 = ~n44924 ;
  assign y13498 = ~n44926 ;
  assign y13499 = n44927 ;
  assign y13500 = ~n44932 ;
  assign y13501 = ~n44936 ;
  assign y13502 = n44937 ;
  assign y13503 = ~n44941 ;
  assign y13504 = ~1'b0 ;
  assign y13505 = ~n44943 ;
  assign y13506 = ~n44946 ;
  assign y13507 = ~n44947 ;
  assign y13508 = n44948 ;
  assign y13509 = n44950 ;
  assign y13510 = ~n44957 ;
  assign y13511 = ~n44958 ;
  assign y13512 = n44959 ;
  assign y13513 = n44961 ;
  assign y13514 = n44963 ;
  assign y13515 = ~n44967 ;
  assign y13516 = n44970 ;
  assign y13517 = ~n44973 ;
  assign y13518 = ~n44974 ;
  assign y13519 = ~n44977 ;
  assign y13520 = ~n44978 ;
  assign y13521 = ~1'b0 ;
  assign y13522 = n44983 ;
  assign y13523 = ~n44985 ;
  assign y13524 = n44992 ;
  assign y13525 = ~n44995 ;
  assign y13526 = ~n44996 ;
  assign y13527 = ~n44997 ;
  assign y13528 = n44998 ;
  assign y13529 = ~n45006 ;
  assign y13530 = ~n45007 ;
  assign y13531 = ~n45009 ;
  assign y13532 = n45013 ;
  assign y13533 = ~n45014 ;
  assign y13534 = ~n45021 ;
  assign y13535 = ~n45022 ;
  assign y13536 = n45023 ;
  assign y13537 = ~n45025 ;
  assign y13538 = ~n45026 ;
  assign y13539 = ~n45028 ;
  assign y13540 = ~n45029 ;
  assign y13541 = n45032 ;
  assign y13542 = n45034 ;
  assign y13543 = ~n45037 ;
  assign y13544 = n45038 ;
  assign y13545 = n45042 ;
  assign y13546 = n45043 ;
  assign y13547 = ~1'b0 ;
  assign y13548 = n45044 ;
  assign y13549 = ~n45046 ;
  assign y13550 = n45049 ;
  assign y13551 = n45052 ;
  assign y13552 = n45055 ;
  assign y13553 = ~1'b0 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = ~n45057 ;
  assign y13556 = ~n45058 ;
  assign y13557 = ~n45059 ;
  assign y13558 = ~n45060 ;
  assign y13559 = n45062 ;
  assign y13560 = n45063 ;
  assign y13561 = ~n45066 ;
  assign y13562 = ~n45070 ;
  assign y13563 = ~1'b0 ;
  assign y13564 = n45075 ;
  assign y13565 = ~1'b0 ;
  assign y13566 = ~n45077 ;
  assign y13567 = ~n45078 ;
  assign y13568 = n45080 ;
  assign y13569 = ~n45082 ;
  assign y13570 = n45085 ;
  assign y13571 = ~n45086 ;
  assign y13572 = n45088 ;
  assign y13573 = ~n45095 ;
  assign y13574 = ~n45097 ;
  assign y13575 = n45102 ;
  assign y13576 = n45116 ;
  assign y13577 = ~n45117 ;
  assign y13578 = n45118 ;
  assign y13579 = n45120 ;
  assign y13580 = ~n45121 ;
  assign y13581 = ~1'b0 ;
  assign y13582 = ~1'b0 ;
  assign y13583 = n45123 ;
  assign y13584 = ~n45124 ;
  assign y13585 = n45127 ;
  assign y13586 = n45130 ;
  assign y13587 = n45131 ;
  assign y13588 = n45132 ;
  assign y13589 = n45133 ;
  assign y13590 = n45136 ;
  assign y13591 = ~n45138 ;
  assign y13592 = n45142 ;
  assign y13593 = n45146 ;
  assign y13594 = n45149 ;
  assign y13595 = n45151 ;
  assign y13596 = n45152 ;
  assign y13597 = n45154 ;
  assign y13598 = ~n45156 ;
  assign y13599 = ~n45157 ;
  assign y13600 = n45162 ;
  assign y13601 = n45164 ;
  assign y13602 = ~n45166 ;
  assign y13603 = ~n45167 ;
  assign y13604 = ~n45172 ;
  assign y13605 = ~n45175 ;
  assign y13606 = n7310 ;
  assign y13607 = n45180 ;
  assign y13608 = ~n45183 ;
  assign y13609 = ~1'b0 ;
  assign y13610 = ~n45184 ;
  assign y13611 = n45190 ;
  assign y13612 = n45191 ;
  assign y13613 = ~n45192 ;
  assign y13614 = ~1'b0 ;
  assign y13615 = n45194 ;
  assign y13616 = ~1'b0 ;
  assign y13617 = ~n45195 ;
  assign y13618 = n45196 ;
  assign y13619 = n45197 ;
  assign y13620 = ~n45200 ;
  assign y13621 = ~n45201 ;
  assign y13622 = ~n45204 ;
  assign y13623 = ~n45205 ;
  assign y13624 = n45207 ;
  assign y13625 = ~n45214 ;
  assign y13626 = ~1'b0 ;
  assign y13627 = ~n45221 ;
  assign y13628 = ~n45225 ;
  assign y13629 = n45232 ;
  assign y13630 = n45233 ;
  assign y13631 = n45237 ;
  assign y13632 = ~1'b0 ;
  assign y13633 = n45238 ;
  assign y13634 = n45240 ;
  assign y13635 = n45246 ;
  assign y13636 = ~n45248 ;
  assign y13637 = ~n45249 ;
  assign y13638 = ~n45252 ;
  assign y13639 = n45255 ;
  assign y13640 = n45257 ;
  assign y13641 = ~n45258 ;
  assign y13642 = n45273 ;
  assign y13643 = n45276 ;
  assign y13644 = ~n45279 ;
  assign y13645 = n45280 ;
  assign y13646 = n45282 ;
  assign y13647 = n45286 ;
  assign y13648 = n45288 ;
  assign y13649 = n45290 ;
  assign y13650 = n45294 ;
  assign y13651 = ~n45296 ;
  assign y13652 = ~n45300 ;
  assign y13653 = ~n45302 ;
  assign y13654 = ~n45303 ;
  assign y13655 = ~n45304 ;
  assign y13656 = ~1'b0 ;
  assign y13657 = ~n45306 ;
  assign y13658 = ~n45309 ;
  assign y13659 = ~n45312 ;
  assign y13660 = ~1'b0 ;
  assign y13661 = n45316 ;
  assign y13662 = ~n45322 ;
  assign y13663 = ~n45324 ;
  assign y13664 = ~n45326 ;
  assign y13665 = n45329 ;
  assign y13666 = n45331 ;
  assign y13667 = ~1'b0 ;
  assign y13668 = ~1'b0 ;
  assign y13669 = ~n45333 ;
  assign y13670 = ~n45335 ;
  assign y13671 = ~n45336 ;
  assign y13672 = ~n45344 ;
  assign y13673 = ~n45345 ;
  assign y13674 = ~n45346 ;
  assign y13675 = n45348 ;
  assign y13676 = ~n45351 ;
  assign y13677 = ~1'b0 ;
  assign y13678 = ~n45353 ;
  assign y13679 = n45355 ;
  assign y13680 = ~n45358 ;
  assign y13681 = n45364 ;
  assign y13682 = ~n45366 ;
  assign y13683 = ~n45370 ;
  assign y13684 = n45376 ;
  assign y13685 = ~n45377 ;
  assign y13686 = ~n45379 ;
  assign y13687 = ~n45380 ;
  assign y13688 = n45381 ;
  assign y13689 = ~n45383 ;
  assign y13690 = ~n45387 ;
  assign y13691 = ~1'b0 ;
  assign y13692 = ~n45391 ;
  assign y13693 = n45396 ;
  assign y13694 = n45401 ;
  assign y13695 = ~n45402 ;
  assign y13696 = n45410 ;
  assign y13697 = ~n45415 ;
  assign y13698 = n22485 ;
  assign y13699 = n45418 ;
  assign y13700 = ~1'b0 ;
  assign y13701 = ~n45421 ;
  assign y13702 = n45423 ;
  assign y13703 = ~n45425 ;
  assign y13704 = ~n45427 ;
  assign y13705 = ~n45429 ;
  assign y13706 = ~n45431 ;
  assign y13707 = ~n45433 ;
  assign y13708 = ~n45435 ;
  assign y13709 = n45437 ;
  assign y13710 = n45439 ;
  assign y13711 = ~n45443 ;
  assign y13712 = n45446 ;
  assign y13713 = ~n45450 ;
  assign y13714 = ~n45456 ;
  assign y13715 = ~n45457 ;
  assign y13716 = ~n45458 ;
  assign y13717 = n45460 ;
  assign y13718 = n45461 ;
  assign y13719 = n45462 ;
  assign y13720 = ~1'b0 ;
  assign y13721 = ~1'b0 ;
  assign y13722 = n45463 ;
  assign y13723 = ~1'b0 ;
  assign y13724 = n45464 ;
  assign y13725 = n45465 ;
  assign y13726 = n45467 ;
  assign y13727 = n45469 ;
  assign y13728 = n45472 ;
  assign y13729 = ~1'b0 ;
  assign y13730 = ~n45476 ;
  assign y13731 = ~1'b0 ;
  assign y13732 = ~n45480 ;
  assign y13733 = n45481 ;
  assign y13734 = ~n45483 ;
  assign y13735 = n45486 ;
  assign y13736 = ~n45489 ;
  assign y13737 = n45490 ;
  assign y13738 = ~n45493 ;
  assign y13739 = ~n45495 ;
  assign y13740 = ~1'b0 ;
  assign y13741 = n45496 ;
  assign y13742 = ~n45497 ;
  assign y13743 = ~n45498 ;
  assign y13744 = ~n45500 ;
  assign y13745 = n45502 ;
  assign y13746 = ~1'b0 ;
  assign y13747 = ~1'b0 ;
  assign y13748 = n45506 ;
  assign y13749 = n45510 ;
  assign y13750 = n45513 ;
  assign y13751 = n45514 ;
  assign y13752 = ~n45515 ;
  assign y13753 = ~1'b0 ;
  assign y13754 = ~n45518 ;
  assign y13755 = ~n45519 ;
  assign y13756 = n45520 ;
  assign y13757 = n45523 ;
  assign y13758 = n28310 ;
  assign y13759 = ~n45524 ;
  assign y13760 = ~n45529 ;
  assign y13761 = ~n45531 ;
  assign y13762 = ~1'b0 ;
  assign y13763 = ~n45532 ;
  assign y13764 = n45533 ;
  assign y13765 = n45534 ;
  assign y13766 = ~n45539 ;
  assign y13767 = ~n45540 ;
  assign y13768 = ~n45544 ;
  assign y13769 = ~n45545 ;
  assign y13770 = n45546 ;
  assign y13771 = n45550 ;
  assign y13772 = ~n45551 ;
  assign y13773 = n45554 ;
  assign y13774 = ~1'b0 ;
  assign y13775 = n45555 ;
  assign y13776 = ~n45560 ;
  assign y13777 = n45563 ;
  assign y13778 = n45564 ;
  assign y13779 = ~n45565 ;
  assign y13780 = n45567 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = n45570 ;
  assign y13783 = ~1'b0 ;
  assign y13784 = ~n45574 ;
  assign y13785 = n45575 ;
  assign y13786 = ~n45579 ;
  assign y13787 = n45582 ;
  assign y13788 = n45584 ;
  assign y13789 = n45585 ;
  assign y13790 = ~n45587 ;
  assign y13791 = ~1'b0 ;
  assign y13792 = ~n45589 ;
  assign y13793 = n45592 ;
  assign y13794 = n45594 ;
  assign y13795 = ~n45599 ;
  assign y13796 = n45608 ;
  assign y13797 = n45611 ;
  assign y13798 = ~n45614 ;
  assign y13799 = n45617 ;
  assign y13800 = ~n45622 ;
  assign y13801 = n45625 ;
  assign y13802 = ~n45626 ;
  assign y13803 = ~n45628 ;
  assign y13804 = n45629 ;
  assign y13805 = ~n45630 ;
  assign y13806 = n45633 ;
  assign y13807 = n45638 ;
  assign y13808 = ~n45646 ;
  assign y13809 = ~n45648 ;
  assign y13810 = ~1'b0 ;
  assign y13811 = n45650 ;
  assign y13812 = ~n45651 ;
  assign y13813 = ~n45653 ;
  assign y13814 = ~n45656 ;
  assign y13815 = ~n45657 ;
  assign y13816 = n45659 ;
  assign y13817 = n45663 ;
  assign y13818 = ~1'b0 ;
  assign y13819 = n45666 ;
  assign y13820 = n45671 ;
  assign y13821 = n45674 ;
  assign y13822 = ~n45675 ;
  assign y13823 = ~n45677 ;
  assign y13824 = ~n45678 ;
  assign y13825 = ~n45679 ;
  assign y13826 = ~n45686 ;
  assign y13827 = ~n45689 ;
  assign y13828 = ~n45692 ;
  assign y13829 = ~n45695 ;
  assign y13830 = n45697 ;
  assign y13831 = n45701 ;
  assign y13832 = ~n45702 ;
  assign y13833 = ~n45707 ;
  assign y13834 = ~n45713 ;
  assign y13835 = ~n45723 ;
  assign y13836 = n45724 ;
  assign y13837 = ~1'b0 ;
  assign y13838 = ~1'b0 ;
  assign y13839 = ~1'b0 ;
  assign y13840 = ~n45725 ;
  assign y13841 = n45729 ;
  assign y13842 = n45730 ;
  assign y13843 = ~n45731 ;
  assign y13844 = ~n45734 ;
  assign y13845 = ~1'b0 ;
  assign y13846 = ~n45736 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = ~n45738 ;
  assign y13849 = n45750 ;
  assign y13850 = n45753 ;
  assign y13851 = ~n45756 ;
  assign y13852 = n45757 ;
  assign y13853 = ~n45758 ;
  assign y13854 = n45760 ;
  assign y13855 = ~n45762 ;
  assign y13856 = ~n45764 ;
  assign y13857 = ~n45765 ;
  assign y13858 = ~n45766 ;
  assign y13859 = n45767 ;
  assign y13860 = ~n45771 ;
  assign y13861 = ~n45772 ;
  assign y13862 = ~1'b0 ;
  assign y13863 = ~n45776 ;
  assign y13864 = n45778 ;
  assign y13865 = ~n45779 ;
  assign y13866 = n45780 ;
  assign y13867 = ~n42996 ;
  assign y13868 = ~n45784 ;
  assign y13869 = ~n45785 ;
  assign y13870 = ~n45791 ;
  assign y13871 = ~n45795 ;
  assign y13872 = ~1'b0 ;
  assign y13873 = n45797 ;
  assign y13874 = n45798 ;
  assign y13875 = n45799 ;
  assign y13876 = ~n45801 ;
  assign y13877 = n45803 ;
  assign y13878 = n45805 ;
  assign y13879 = n45806 ;
  assign y13880 = ~1'b0 ;
  assign y13881 = n45809 ;
  assign y13882 = n45811 ;
  assign y13883 = ~n45812 ;
  assign y13884 = ~n45813 ;
  assign y13885 = ~n45816 ;
  assign y13886 = n45818 ;
  assign y13887 = ~n45819 ;
  assign y13888 = ~n45827 ;
  assign y13889 = ~n45829 ;
  assign y13890 = n45830 ;
  assign y13891 = 1'b0 ;
  assign y13892 = ~n45833 ;
  assign y13893 = n45834 ;
  assign y13894 = n45839 ;
  assign y13895 = n45841 ;
  assign y13896 = n45842 ;
  assign y13897 = n45846 ;
  assign y13898 = ~n45851 ;
  assign y13899 = ~n45853 ;
  assign y13900 = ~n45858 ;
  assign y13901 = n45860 ;
  assign y13902 = ~n45864 ;
  assign y13903 = n45873 ;
  assign y13904 = ~n45878 ;
  assign y13905 = n45884 ;
  assign y13906 = ~1'b0 ;
  assign y13907 = ~1'b0 ;
  assign y13908 = ~n45887 ;
  assign y13909 = n45890 ;
  assign y13910 = n45893 ;
  assign y13911 = n45897 ;
  assign y13912 = ~n45898 ;
  assign y13913 = ~n45901 ;
  assign y13914 = n45902 ;
  assign y13915 = ~n45905 ;
  assign y13916 = ~n45907 ;
  assign y13917 = ~1'b0 ;
  assign y13918 = n45914 ;
  assign y13919 = ~n45918 ;
  assign y13920 = n45922 ;
  assign y13921 = ~n45924 ;
  assign y13922 = n45926 ;
  assign y13923 = n45930 ;
  assign y13924 = ~n45933 ;
  assign y13925 = n45937 ;
  assign y13926 = n45938 ;
  assign y13927 = ~n45942 ;
  assign y13928 = ~n45943 ;
  assign y13929 = ~n45944 ;
  assign y13930 = n45947 ;
  assign y13931 = ~1'b0 ;
  assign y13932 = n45948 ;
  assign y13933 = n45950 ;
  assign y13934 = n45951 ;
  assign y13935 = n45952 ;
  assign y13936 = ~n45958 ;
  assign y13937 = ~n45965 ;
  assign y13938 = n45969 ;
  assign y13939 = n45970 ;
  assign y13940 = n45971 ;
  assign y13941 = n45972 ;
  assign y13942 = n45976 ;
  assign y13943 = ~n45977 ;
  assign y13944 = ~1'b0 ;
  assign y13945 = ~1'b0 ;
  assign y13946 = n45979 ;
  assign y13947 = ~n45982 ;
  assign y13948 = n45991 ;
  assign y13949 = n45993 ;
  assign y13950 = ~n45994 ;
  assign y13951 = ~n45996 ;
  assign y13952 = ~n45998 ;
  assign y13953 = n46002 ;
  assign y13954 = ~n46003 ;
  assign y13955 = ~n46006 ;
  assign y13956 = ~n46007 ;
  assign y13957 = ~n46008 ;
  assign y13958 = n46009 ;
  assign y13959 = ~n46013 ;
  assign y13960 = ~n46015 ;
  assign y13961 = ~n46016 ;
  assign y13962 = ~n46019 ;
  assign y13963 = n46022 ;
  assign y13964 = ~n46023 ;
  assign y13965 = n46030 ;
  assign y13966 = n46035 ;
  assign y13967 = n46037 ;
  assign y13968 = ~n46040 ;
  assign y13969 = n46041 ;
  assign y13970 = ~n46043 ;
  assign y13971 = n46044 ;
  assign y13972 = n46047 ;
  assign y13973 = n46048 ;
  assign y13974 = n46052 ;
  assign y13975 = ~n46055 ;
  assign y13976 = n46058 ;
  assign y13977 = ~n46061 ;
  assign y13978 = n46064 ;
  assign y13979 = ~1'b0 ;
  assign y13980 = ~n46065 ;
  assign y13981 = n46069 ;
  assign y13982 = n46070 ;
  assign y13983 = ~n46072 ;
  assign y13984 = n46073 ;
  assign y13985 = n46074 ;
  assign y13986 = n46076 ;
  assign y13987 = n46080 ;
  assign y13988 = n46083 ;
  assign y13989 = ~n46084 ;
  assign y13990 = n46087 ;
  assign y13991 = ~n46090 ;
  assign y13992 = n46095 ;
  assign y13993 = ~n46096 ;
  assign y13994 = ~n46098 ;
  assign y13995 = ~n46101 ;
  assign y13996 = ~1'b0 ;
  assign y13997 = ~n46102 ;
  assign y13998 = ~n46103 ;
  assign y13999 = n46107 ;
  assign y14000 = n46111 ;
  assign y14001 = n46116 ;
  assign y14002 = ~1'b0 ;
  assign y14003 = ~1'b0 ;
  assign y14004 = ~n10272 ;
  assign y14005 = ~n46122 ;
  assign y14006 = ~n46127 ;
  assign y14007 = n46129 ;
  assign y14008 = n46130 ;
  assign y14009 = n46131 ;
  assign y14010 = n46138 ;
  assign y14011 = n46142 ;
  assign y14012 = ~n46143 ;
  assign y14013 = ~1'b0 ;
  assign y14014 = ~1'b0 ;
  assign y14015 = ~n46146 ;
  assign y14016 = ~n46149 ;
  assign y14017 = n46150 ;
  assign y14018 = ~n46152 ;
  assign y14019 = n46154 ;
  assign y14020 = n46156 ;
  assign y14021 = ~n46159 ;
  assign y14022 = ~n46162 ;
  assign y14023 = n46163 ;
  assign y14024 = n46165 ;
  assign y14025 = n46166 ;
  assign y14026 = ~n46168 ;
  assign y14027 = n46170 ;
  assign y14028 = ~n46173 ;
  assign y14029 = n46176 ;
  assign y14030 = ~n46180 ;
  assign y14031 = ~n46181 ;
  assign y14032 = n46185 ;
  assign y14033 = n46188 ;
  assign y14034 = n46191 ;
  assign y14035 = ~n46195 ;
  assign y14036 = n46201 ;
  assign y14037 = n46204 ;
  assign y14038 = ~n46206 ;
  assign y14039 = ~n46210 ;
  assign y14040 = n46211 ;
  assign y14041 = ~n46212 ;
  assign y14042 = ~n46213 ;
  assign y14043 = n46214 ;
  assign y14044 = n46220 ;
  assign y14045 = ~n46222 ;
  assign y14046 = n46226 ;
  assign y14047 = ~n46229 ;
  assign y14048 = ~1'b0 ;
  assign y14049 = ~n46232 ;
  assign y14050 = n46242 ;
  assign y14051 = ~n46246 ;
  assign y14052 = ~n46250 ;
  assign y14053 = ~n46251 ;
  assign y14054 = n46255 ;
  assign y14055 = ~n46257 ;
  assign y14056 = ~n46258 ;
  assign y14057 = ~n46263 ;
  assign y14058 = n46267 ;
  assign y14059 = ~n46268 ;
  assign y14060 = n46271 ;
  assign y14061 = ~n46272 ;
  assign y14062 = n46273 ;
  assign y14063 = ~n46275 ;
  assign y14064 = ~n46277 ;
  assign y14065 = ~n46280 ;
  assign y14066 = ~n46282 ;
  assign y14067 = ~n46283 ;
  assign y14068 = ~n46285 ;
  assign y14069 = ~n46286 ;
  assign y14070 = n46288 ;
  assign y14071 = n46290 ;
  assign y14072 = n46293 ;
  assign y14073 = ~1'b0 ;
  assign y14074 = ~n46294 ;
  assign y14075 = n46296 ;
  assign y14076 = n46297 ;
  assign y14077 = ~n46299 ;
  assign y14078 = ~n46302 ;
  assign y14079 = ~1'b0 ;
  assign y14080 = n46305 ;
  assign y14081 = ~n46308 ;
  assign y14082 = ~n46309 ;
  assign y14083 = ~n46311 ;
  assign y14084 = ~n46314 ;
  assign y14085 = ~n46316 ;
  assign y14086 = n46317 ;
  assign y14087 = ~1'b0 ;
  assign y14088 = n46320 ;
  assign y14089 = ~n46324 ;
  assign y14090 = n46327 ;
  assign y14091 = ~n46331 ;
  assign y14092 = ~n46332 ;
  assign y14093 = ~n46335 ;
  assign y14094 = n46338 ;
  assign y14095 = n46341 ;
  assign y14096 = ~n46342 ;
  assign y14097 = n46347 ;
  assign y14098 = ~n46349 ;
  assign y14099 = n46351 ;
  assign y14100 = n46353 ;
  assign y14101 = ~n46355 ;
  assign y14102 = ~n46356 ;
  assign y14103 = n46359 ;
  assign y14104 = ~n46360 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = n46361 ;
  assign y14107 = n46364 ;
  assign y14108 = n46368 ;
  assign y14109 = n46369 ;
  assign y14110 = n46373 ;
  assign y14111 = ~1'b0 ;
  assign y14112 = ~n46377 ;
  assign y14113 = n46383 ;
  assign y14114 = ~n46387 ;
  assign y14115 = ~n46388 ;
  assign y14116 = n46390 ;
  assign y14117 = ~n46391 ;
  assign y14118 = ~n46398 ;
  assign y14119 = ~n46399 ;
  assign y14120 = n46403 ;
  assign y14121 = n46406 ;
  assign y14122 = ~1'b0 ;
  assign y14123 = n46411 ;
  assign y14124 = ~n46413 ;
  assign y14125 = ~n46414 ;
  assign y14126 = ~n35269 ;
  assign y14127 = n46418 ;
  assign y14128 = ~n46419 ;
  assign y14129 = ~n46422 ;
  assign y14130 = ~n46425 ;
  assign y14131 = n46427 ;
  assign y14132 = ~1'b0 ;
  assign y14133 = ~1'b0 ;
  assign y14134 = n46429 ;
  assign y14135 = ~n46432 ;
  assign y14136 = n46434 ;
  assign y14137 = n46435 ;
  assign y14138 = ~n46437 ;
  assign y14139 = ~n46442 ;
  assign y14140 = ~n46444 ;
  assign y14141 = ~1'b0 ;
  assign y14142 = n46446 ;
  assign y14143 = n46449 ;
  assign y14144 = ~n46451 ;
  assign y14145 = ~n46452 ;
  assign y14146 = ~n46455 ;
  assign y14147 = ~n38443 ;
  assign y14148 = ~n46459 ;
  assign y14149 = ~n46462 ;
  assign y14150 = ~n46463 ;
  assign y14151 = n46465 ;
  assign y14152 = n46467 ;
  assign y14153 = n46470 ;
  assign y14154 = n46473 ;
  assign y14155 = ~n46476 ;
  assign y14156 = n46479 ;
  assign y14157 = n46484 ;
  assign y14158 = n30804 ;
  assign y14159 = ~1'b0 ;
  assign y14160 = ~1'b0 ;
  assign y14161 = ~n46488 ;
  assign y14162 = n46492 ;
  assign y14163 = ~n46493 ;
  assign y14164 = ~n46497 ;
  assign y14165 = ~n46499 ;
  assign y14166 = ~n46501 ;
  assign y14167 = ~n46502 ;
  assign y14168 = ~n46504 ;
  assign y14169 = ~n46506 ;
  assign y14170 = n46507 ;
  assign y14171 = n46510 ;
  assign y14172 = ~n46513 ;
  assign y14173 = ~n46514 ;
  assign y14174 = ~n46516 ;
  assign y14175 = ~n46519 ;
  assign y14176 = ~n46527 ;
  assign y14177 = ~n46532 ;
  assign y14178 = n46533 ;
  assign y14179 = ~n46537 ;
  assign y14180 = ~n46539 ;
  assign y14181 = n46540 ;
  assign y14182 = ~n46541 ;
  assign y14183 = ~n46544 ;
  assign y14184 = n46546 ;
  assign y14185 = n46548 ;
  assign y14186 = n46551 ;
  assign y14187 = ~n46552 ;
  assign y14188 = ~n46556 ;
  assign y14189 = n46557 ;
  assign y14190 = n46561 ;
  assign y14191 = n46562 ;
  assign y14192 = ~n46564 ;
  assign y14193 = n46567 ;
  assign y14194 = ~1'b0 ;
  assign y14195 = ~1'b0 ;
  assign y14196 = n46568 ;
  assign y14197 = ~n46571 ;
  assign y14198 = n46572 ;
  assign y14199 = ~n46575 ;
  assign y14200 = ~n46578 ;
  assign y14201 = n46582 ;
  assign y14202 = ~n46583 ;
  assign y14203 = n46585 ;
  assign y14204 = ~n46587 ;
  assign y14205 = n46589 ;
  assign y14206 = n46595 ;
  assign y14207 = ~n46603 ;
  assign y14208 = ~n46604 ;
  assign y14209 = ~n46606 ;
  assign y14210 = ~n46609 ;
  assign y14211 = ~n46610 ;
  assign y14212 = n46612 ;
  assign y14213 = ~n46613 ;
  assign y14214 = ~1'b0 ;
  assign y14215 = n46615 ;
  assign y14216 = ~1'b0 ;
  assign y14217 = ~n46618 ;
  assign y14218 = n46621 ;
  assign y14219 = ~n46624 ;
  assign y14220 = n46625 ;
  assign y14221 = n46626 ;
  assign y14222 = ~n46627 ;
  assign y14223 = n46629 ;
  assign y14224 = ~n46634 ;
  assign y14225 = n46636 ;
  assign y14226 = n46639 ;
  assign y14227 = n46643 ;
  assign y14228 = ~n46644 ;
  assign y14229 = n46650 ;
  assign y14230 = ~n46651 ;
  assign y14231 = n46652 ;
  assign y14232 = n46654 ;
  assign y14233 = ~n10700 ;
  assign y14234 = n46657 ;
  assign y14235 = ~1'b0 ;
  assign y14236 = n46660 ;
  assign y14237 = n46662 ;
  assign y14238 = n46663 ;
  assign y14239 = ~n46665 ;
  assign y14240 = n46666 ;
  assign y14241 = n46669 ;
  assign y14242 = n46670 ;
  assign y14243 = ~1'b0 ;
  assign y14244 = n46673 ;
  assign y14245 = ~n46684 ;
  assign y14246 = ~1'b0 ;
  assign y14247 = n46685 ;
  assign y14248 = ~n46689 ;
  assign y14249 = n46694 ;
  assign y14250 = ~n46696 ;
  assign y14251 = n46697 ;
  assign y14252 = n46702 ;
  assign y14253 = ~1'b0 ;
  assign y14254 = n46706 ;
  assign y14255 = ~1'b0 ;
  assign y14256 = n46710 ;
  assign y14257 = n46711 ;
  assign y14258 = ~n46716 ;
  assign y14259 = ~n46718 ;
  assign y14260 = ~n7580 ;
  assign y14261 = ~n46727 ;
  assign y14262 = ~n46729 ;
  assign y14263 = ~n46731 ;
  assign y14264 = n46734 ;
  assign y14265 = ~n46735 ;
  assign y14266 = ~n46737 ;
  assign y14267 = ~n46738 ;
  assign y14268 = n46740 ;
  assign y14269 = ~1'b0 ;
  assign y14270 = n46742 ;
  assign y14271 = n46743 ;
  assign y14272 = ~n46750 ;
  assign y14273 = ~n46751 ;
  assign y14274 = ~n46752 ;
  assign y14275 = n46753 ;
  assign y14276 = ~1'b0 ;
  assign y14277 = ~1'b0 ;
  assign y14278 = n46755 ;
  assign y14279 = n46762 ;
  assign y14280 = ~n46767 ;
  assign y14281 = n46773 ;
  assign y14282 = n46776 ;
  assign y14283 = ~n46779 ;
  assign y14284 = ~n46782 ;
  assign y14285 = ~n46786 ;
  assign y14286 = ~n46791 ;
  assign y14287 = ~1'b0 ;
  assign y14288 = n46795 ;
  assign y14289 = ~1'b0 ;
  assign y14290 = n46796 ;
  assign y14291 = n46797 ;
  assign y14292 = n46803 ;
  assign y14293 = n46804 ;
  assign y14294 = ~n46807 ;
  assign y14295 = ~n46812 ;
  assign y14296 = ~1'b0 ;
  assign y14297 = ~n46815 ;
  assign y14298 = n46817 ;
  assign y14299 = n46819 ;
  assign y14300 = n46822 ;
  assign y14301 = ~1'b0 ;
  assign y14302 = ~1'b0 ;
  assign y14303 = ~n46823 ;
  assign y14304 = n46826 ;
  assign y14305 = n46828 ;
  assign y14306 = n46830 ;
  assign y14307 = ~n46831 ;
  assign y14308 = n46832 ;
  assign y14309 = ~n46835 ;
  assign y14310 = n46840 ;
  assign y14311 = n46841 ;
  assign y14312 = n46842 ;
  assign y14313 = n46845 ;
  assign y14314 = n46848 ;
  assign y14315 = n46849 ;
  assign y14316 = ~n46851 ;
  assign y14317 = n46853 ;
  assign y14318 = ~n46855 ;
  assign y14319 = ~n46857 ;
  assign y14320 = ~n46861 ;
  assign y14321 = n46863 ;
  assign y14322 = n46866 ;
  assign y14323 = n46869 ;
  assign y14324 = ~n46875 ;
  assign y14325 = ~n46876 ;
  assign y14326 = ~n46881 ;
  assign y14327 = ~1'b0 ;
  assign y14328 = ~n46884 ;
  assign y14329 = ~1'b0 ;
  assign y14330 = ~n46889 ;
  assign y14331 = n46891 ;
  assign y14332 = ~n46892 ;
  assign y14333 = n46893 ;
  assign y14334 = ~n46896 ;
  assign y14335 = ~n46897 ;
  assign y14336 = n46900 ;
  assign y14337 = n46905 ;
  assign y14338 = ~1'b0 ;
  assign y14339 = ~n46908 ;
  assign y14340 = ~n46913 ;
  assign y14341 = ~n46914 ;
  assign y14342 = ~n46915 ;
  assign y14343 = ~n46918 ;
  assign y14344 = ~n46921 ;
  assign y14345 = ~n46922 ;
  assign y14346 = n46923 ;
  assign y14347 = n46924 ;
  assign y14348 = n46926 ;
  assign y14349 = ~n46927 ;
  assign y14350 = n46928 ;
  assign y14351 = ~n46929 ;
  assign y14352 = ~n46931 ;
  assign y14353 = ~n33579 ;
  assign y14354 = ~n46933 ;
  assign y14355 = ~1'b0 ;
  assign y14356 = ~1'b0 ;
  assign y14357 = ~n46937 ;
  assign y14358 = n46938 ;
  assign y14359 = n46942 ;
  assign y14360 = n46943 ;
  assign y14361 = ~n46945 ;
  assign y14362 = ~n46950 ;
  assign y14363 = ~n46955 ;
  assign y14364 = n46960 ;
  assign y14365 = ~n46961 ;
  assign y14366 = n46962 ;
  assign y14367 = ~n46964 ;
  assign y14368 = n46965 ;
  assign y14369 = n46969 ;
  assign y14370 = n46976 ;
  assign y14371 = ~n46977 ;
  assign y14372 = ~n46978 ;
  assign y14373 = n46981 ;
  assign y14374 = n46983 ;
  assign y14375 = ~n46984 ;
  assign y14376 = ~n46987 ;
  assign y14377 = n46988 ;
  assign y14378 = n46990 ;
  assign y14379 = n46996 ;
  assign y14380 = n46998 ;
  assign y14381 = n47001 ;
  assign y14382 = n47004 ;
  assign y14383 = ~1'b0 ;
  assign y14384 = ~1'b0 ;
  assign y14385 = n47005 ;
  assign y14386 = ~n47006 ;
  assign y14387 = n47010 ;
  assign y14388 = ~n47013 ;
  assign y14389 = n47020 ;
  assign y14390 = ~n47022 ;
  assign y14391 = ~1'b0 ;
  assign y14392 = ~n47024 ;
  assign y14393 = ~n47026 ;
  assign y14394 = ~n47028 ;
  assign y14395 = n22446 ;
  assign y14396 = n47031 ;
  assign y14397 = ~n47032 ;
  assign y14398 = n47037 ;
  assign y14399 = n47041 ;
  assign y14400 = ~n47044 ;
  assign y14401 = 1'b0 ;
  assign y14402 = n47047 ;
  assign y14403 = n47051 ;
  assign y14404 = n47053 ;
  assign y14405 = ~n47055 ;
  assign y14406 = n47056 ;
  assign y14407 = ~n47059 ;
  assign y14408 = ~n47060 ;
  assign y14409 = ~n47061 ;
  assign y14410 = ~1'b0 ;
  assign y14411 = n47068 ;
  assign y14412 = ~1'b0 ;
  assign y14413 = ~n47069 ;
  assign y14414 = n47071 ;
  assign y14415 = n47075 ;
  assign y14416 = n47076 ;
  assign y14417 = ~n47077 ;
  assign y14418 = ~n47080 ;
  assign y14419 = ~1'b0 ;
  assign y14420 = ~n47087 ;
  assign y14421 = ~n47092 ;
  assign y14422 = ~n47096 ;
  assign y14423 = n47099 ;
  assign y14424 = n47101 ;
  assign y14425 = n47103 ;
  assign y14426 = ~1'b0 ;
  assign y14427 = ~1'b0 ;
  assign y14428 = ~n47104 ;
  assign y14429 = ~n47106 ;
  assign y14430 = ~n47107 ;
  assign y14431 = ~n47110 ;
  assign y14432 = ~n47111 ;
  assign y14433 = ~n47116 ;
  assign y14434 = ~n47120 ;
  assign y14435 = n47122 ;
  assign y14436 = ~n47123 ;
  assign y14437 = ~n47124 ;
  assign y14438 = ~n47125 ;
  assign y14439 = n47126 ;
  assign y14440 = n47127 ;
  assign y14441 = ~n47128 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = ~1'b0 ;
  assign y14444 = ~1'b0 ;
  assign y14445 = ~n47134 ;
  assign y14446 = ~n47135 ;
  assign y14447 = ~n47136 ;
  assign y14448 = n47137 ;
  assign y14449 = ~n47139 ;
  assign y14450 = n47140 ;
  assign y14451 = ~n47148 ;
  assign y14452 = ~n47153 ;
  assign y14453 = ~n47155 ;
  assign y14454 = ~n47158 ;
  assign y14455 = n47159 ;
  assign y14456 = n47162 ;
  assign y14457 = n47163 ;
  assign y14458 = ~n47165 ;
  assign y14459 = ~n47167 ;
  assign y14460 = ~n47175 ;
  assign y14461 = n47179 ;
  assign y14462 = ~1'b0 ;
  assign y14463 = n47181 ;
  assign y14464 = ~1'b0 ;
  assign y14465 = n47183 ;
  assign y14466 = ~n47184 ;
  assign y14467 = ~n47185 ;
  assign y14468 = ~n47186 ;
  assign y14469 = ~n47190 ;
  assign y14470 = ~n47200 ;
  assign y14471 = n47201 ;
  assign y14472 = n47208 ;
  assign y14473 = ~1'b0 ;
  assign y14474 = ~n47216 ;
  assign y14475 = n47221 ;
  assign y14476 = ~n47223 ;
  assign y14477 = n47225 ;
  assign y14478 = n47226 ;
  assign y14479 = ~n47228 ;
  assign y14480 = ~n47232 ;
  assign y14481 = ~n47235 ;
  assign y14482 = n47240 ;
  assign y14483 = ~n47242 ;
  assign y14484 = n47243 ;
  assign y14485 = ~n47247 ;
  assign y14486 = n47248 ;
  assign y14487 = ~1'b0 ;
  assign y14488 = ~n47252 ;
  assign y14489 = ~n47256 ;
  assign y14490 = n47260 ;
  assign y14491 = n47262 ;
  assign y14492 = ~n47263 ;
  assign y14493 = ~n47264 ;
  assign y14494 = n47265 ;
  assign y14495 = n47267 ;
  assign y14496 = n47269 ;
  assign y14497 = ~n47270 ;
  assign y14498 = n47277 ;
  assign y14499 = ~n47278 ;
  assign y14500 = ~n47281 ;
  assign y14501 = n47283 ;
  assign y14502 = n47287 ;
  assign y14503 = n47290 ;
  assign y14504 = ~n47292 ;
  assign y14505 = ~n47293 ;
  assign y14506 = ~n47296 ;
  assign y14507 = ~n47298 ;
  assign y14508 = ~n47301 ;
  assign y14509 = ~1'b0 ;
  assign y14510 = n47306 ;
  assign y14511 = n47307 ;
  assign y14512 = n47309 ;
  assign y14513 = ~n47313 ;
  assign y14514 = ~n47314 ;
  assign y14515 = ~n47317 ;
  assign y14516 = n47318 ;
  assign y14517 = ~1'b0 ;
  assign y14518 = ~n47320 ;
  assign y14519 = n47322 ;
  assign y14520 = ~1'b0 ;
  assign y14521 = n47326 ;
  assign y14522 = ~n47329 ;
  assign y14523 = ~n47331 ;
  assign y14524 = n47334 ;
  assign y14525 = n47337 ;
  assign y14526 = n47342 ;
  assign y14527 = ~n47345 ;
  assign y14528 = ~n47347 ;
  assign y14529 = ~1'b0 ;
  assign y14530 = n47350 ;
  assign y14531 = ~n47352 ;
  assign y14532 = ~n47354 ;
  assign y14533 = n47358 ;
  assign y14534 = ~n47359 ;
  assign y14535 = n47360 ;
  assign y14536 = ~n47362 ;
  assign y14537 = n47364 ;
  assign y14538 = n47370 ;
  assign y14539 = n47371 ;
  assign y14540 = n47374 ;
  assign y14541 = n47375 ;
  assign y14542 = ~n47376 ;
  assign y14543 = ~n47379 ;
  assign y14544 = n47381 ;
  assign y14545 = ~n47383 ;
  assign y14546 = ~1'b0 ;
  assign y14547 = n47385 ;
  assign y14548 = ~n47388 ;
  assign y14549 = ~n47391 ;
  assign y14550 = n47392 ;
  assign y14551 = ~n47396 ;
  assign y14552 = ~n47398 ;
  assign y14553 = n47400 ;
  assign y14554 = n47401 ;
  assign y14555 = ~n47407 ;
  assign y14556 = ~n47409 ;
  assign y14557 = ~1'b0 ;
  assign y14558 = n47412 ;
  assign y14559 = ~n47416 ;
  assign y14560 = n47425 ;
  assign y14561 = n36661 ;
  assign y14562 = ~n47428 ;
  assign y14563 = n47429 ;
  assign y14564 = n47431 ;
  assign y14565 = ~n11913 ;
  assign y14566 = n47433 ;
  assign y14567 = ~n47435 ;
  assign y14568 = n47436 ;
  assign y14569 = n47437 ;
  assign y14570 = n47444 ;
  assign y14571 = n47449 ;
  assign y14572 = n47452 ;
  assign y14573 = n47453 ;
  assign y14574 = n47456 ;
  assign y14575 = ~1'b0 ;
  assign y14576 = n47457 ;
  assign y14577 = ~n47459 ;
  assign y14578 = n47462 ;
  assign y14579 = ~n47465 ;
  assign y14580 = n47467 ;
  assign y14581 = ~n47470 ;
  assign y14582 = n47474 ;
  assign y14583 = ~1'b0 ;
  assign y14584 = ~1'b0 ;
  assign y14585 = ~1'b0 ;
  assign y14586 = n47475 ;
  assign y14587 = ~n47478 ;
  assign y14588 = ~n47479 ;
  assign y14589 = n47481 ;
  assign y14590 = n47484 ;
  assign y14591 = ~n47486 ;
  assign y14592 = ~1'b0 ;
  assign y14593 = ~1'b0 ;
  assign y14594 = ~n47487 ;
  assign y14595 = ~n47488 ;
  assign y14596 = ~n47489 ;
  assign y14597 = ~n47491 ;
  assign y14598 = ~n47495 ;
  assign y14599 = ~n47496 ;
  assign y14600 = ~1'b0 ;
  assign y14601 = ~n47499 ;
  assign y14602 = n47503 ;
  assign y14603 = ~n47508 ;
  assign y14604 = ~n47509 ;
  assign y14605 = ~n47511 ;
  assign y14606 = ~1'b0 ;
  assign y14607 = ~n47513 ;
  assign y14608 = n47514 ;
  assign y14609 = ~n47518 ;
  assign y14610 = n47522 ;
  assign y14611 = ~1'b0 ;
  assign y14612 = ~n47523 ;
  assign y14613 = n47524 ;
  assign y14614 = n47525 ;
  assign y14615 = n47528 ;
  assign y14616 = n47531 ;
  assign y14617 = ~n47536 ;
  assign y14618 = ~1'b0 ;
  assign y14619 = n47539 ;
  assign y14620 = ~n47540 ;
  assign y14621 = ~n47544 ;
  assign y14622 = ~n47546 ;
  assign y14623 = ~n47548 ;
  assign y14624 = ~n47549 ;
  assign y14625 = ~n47551 ;
  assign y14626 = ~n47560 ;
  assign y14627 = ~n47562 ;
  assign y14628 = n47564 ;
  assign y14629 = ~1'b0 ;
  assign y14630 = n47568 ;
  assign y14631 = ~n47573 ;
  assign y14632 = n47574 ;
  assign y14633 = ~n47577 ;
  assign y14634 = ~n47579 ;
  assign y14635 = ~n47587 ;
  assign y14636 = ~n47588 ;
  assign y14637 = ~n47590 ;
  assign y14638 = ~1'b0 ;
  assign y14639 = ~1'b0 ;
  assign y14640 = ~1'b0 ;
  assign y14641 = n47592 ;
  assign y14642 = ~n47594 ;
  assign y14643 = ~n47595 ;
  assign y14644 = n47600 ;
  assign y14645 = n47603 ;
  assign y14646 = n47606 ;
  assign y14647 = ~1'b0 ;
  assign y14648 = n47611 ;
  assign y14649 = n47613 ;
  assign y14650 = ~n47617 ;
  assign y14651 = n47618 ;
  assign y14652 = n47619 ;
  assign y14653 = ~n47625 ;
  assign y14654 = ~n47627 ;
  assign y14655 = ~n47630 ;
  assign y14656 = n47638 ;
  assign y14657 = n47642 ;
  assign y14658 = n47643 ;
  assign y14659 = ~n47644 ;
  assign y14660 = n47646 ;
  assign y14661 = n47647 ;
  assign y14662 = n47648 ;
  assign y14663 = n47650 ;
  assign y14664 = ~n47652 ;
  assign y14665 = n47654 ;
  assign y14666 = ~n47657 ;
  assign y14667 = ~n47658 ;
  assign y14668 = n47663 ;
  assign y14669 = ~n47670 ;
  assign y14670 = n47671 ;
  assign y14671 = ~n47672 ;
  assign y14672 = n47673 ;
  assign y14673 = ~n47675 ;
  assign y14674 = ~1'b0 ;
  assign y14675 = ~n47676 ;
  assign y14676 = ~n47678 ;
  assign y14677 = n47679 ;
  assign y14678 = n47682 ;
  assign y14679 = n47684 ;
  assign y14680 = ~n47690 ;
  assign y14681 = n47693 ;
  assign y14682 = n47696 ;
  assign y14683 = ~n47698 ;
  assign y14684 = ~1'b0 ;
  assign y14685 = ~n47704 ;
  assign y14686 = ~n47707 ;
  assign y14687 = n47708 ;
  assign y14688 = ~n47711 ;
  assign y14689 = ~n47712 ;
  assign y14690 = n47714 ;
  assign y14691 = n47715 ;
  assign y14692 = n47718 ;
  assign y14693 = ~1'b0 ;
  assign y14694 = ~n47720 ;
  assign y14695 = ~n47721 ;
  assign y14696 = n47722 ;
  assign y14697 = ~n47723 ;
  assign y14698 = ~n47725 ;
  assign y14699 = ~n47728 ;
  assign y14700 = ~n47729 ;
  assign y14701 = ~1'b0 ;
  assign y14702 = ~n47731 ;
  assign y14703 = n47733 ;
  assign y14704 = ~1'b0 ;
  assign y14705 = n47734 ;
  assign y14706 = ~n47736 ;
  assign y14707 = ~n47737 ;
  assign y14708 = ~n47741 ;
  assign y14709 = n47744 ;
  assign y14710 = ~n47745 ;
  assign y14711 = ~n47747 ;
  assign y14712 = n47750 ;
  assign y14713 = ~n47753 ;
  assign y14714 = ~1'b0 ;
  assign y14715 = ~n47754 ;
  assign y14716 = ~n47756 ;
  assign y14717 = ~n47761 ;
  assign y14718 = ~n47762 ;
  assign y14719 = n47763 ;
  assign y14720 = ~n47764 ;
  assign y14721 = ~n47770 ;
  assign y14722 = ~n47771 ;
  assign y14723 = ~n47775 ;
  assign y14724 = n47776 ;
  assign y14725 = ~n47777 ;
  assign y14726 = ~n47778 ;
  assign y14727 = ~n47779 ;
  assign y14728 = n47780 ;
  assign y14729 = ~n47781 ;
  assign y14730 = n47782 ;
  assign y14731 = ~n47785 ;
  assign y14732 = n47789 ;
  assign y14733 = ~n47793 ;
  assign y14734 = n47796 ;
  assign y14735 = n47801 ;
  assign y14736 = n47803 ;
  assign y14737 = n47805 ;
  assign y14738 = n47810 ;
  assign y14739 = n47818 ;
  assign y14740 = ~n47819 ;
  assign y14741 = ~n47821 ;
  assign y14742 = n47827 ;
  assign y14743 = ~n47830 ;
  assign y14744 = ~n47831 ;
  assign y14745 = n47832 ;
  assign y14746 = ~n47837 ;
  assign y14747 = ~n47839 ;
  assign y14748 = ~n47840 ;
  assign y14749 = ~n47845 ;
  assign y14750 = ~n47847 ;
  assign y14751 = n47851 ;
  assign y14752 = ~n47854 ;
  assign y14753 = ~n47857 ;
  assign y14754 = ~n47858 ;
  assign y14755 = ~n47859 ;
  assign y14756 = ~n47860 ;
  assign y14757 = ~n47861 ;
  assign y14758 = n47862 ;
  assign y14759 = n47867 ;
  assign y14760 = n47869 ;
  assign y14761 = ~1'b0 ;
  assign y14762 = ~n47871 ;
  assign y14763 = n47872 ;
  assign y14764 = n47873 ;
  assign y14765 = ~n47874 ;
  assign y14766 = n47877 ;
  assign y14767 = ~n47885 ;
  assign y14768 = n47886 ;
  assign y14769 = ~n47888 ;
  assign y14770 = ~n47891 ;
  assign y14771 = ~n47892 ;
  assign y14772 = ~n47893 ;
  assign y14773 = ~n47896 ;
  assign y14774 = ~n47898 ;
  assign y14775 = ~n47899 ;
  assign y14776 = n47904 ;
  assign y14777 = ~n47907 ;
  assign y14778 = ~1'b0 ;
  assign y14779 = n47910 ;
  assign y14780 = ~n47912 ;
  assign y14781 = n47913 ;
  assign y14782 = ~n47914 ;
  assign y14783 = ~n47915 ;
  assign y14784 = n47920 ;
  assign y14785 = n47922 ;
  assign y14786 = n47923 ;
  assign y14787 = n47926 ;
  assign y14788 = n47930 ;
  assign y14789 = n47931 ;
  assign y14790 = ~n47935 ;
  assign y14791 = ~n47936 ;
  assign y14792 = ~n47937 ;
  assign y14793 = n27044 ;
  assign y14794 = ~n47942 ;
  assign y14795 = ~n47944 ;
  assign y14796 = ~1'b0 ;
  assign y14797 = n47947 ;
  assign y14798 = ~n47949 ;
  assign y14799 = n47950 ;
  assign y14800 = n47952 ;
  assign y14801 = ~n47954 ;
  assign y14802 = ~n47956 ;
  assign y14803 = n47959 ;
  assign y14804 = ~n47961 ;
  assign y14805 = n38112 ;
  assign y14806 = ~n47964 ;
  assign y14807 = n47968 ;
  assign y14808 = n47969 ;
  assign y14809 = ~n47971 ;
  assign y14810 = ~1'b0 ;
  assign y14811 = ~1'b0 ;
  assign y14812 = n47975 ;
  assign y14813 = ~n47976 ;
  assign y14814 = n47979 ;
  assign y14815 = n47981 ;
  assign y14816 = ~n47983 ;
  assign y14817 = ~n47984 ;
  assign y14818 = ~n47994 ;
  assign y14819 = n47996 ;
  assign y14820 = ~n47998 ;
  assign y14821 = n48001 ;
  assign y14822 = ~n48003 ;
  assign y14823 = n48004 ;
  assign y14824 = n48008 ;
  assign y14825 = n48009 ;
  assign y14826 = ~n48012 ;
  assign y14827 = ~n48013 ;
  assign y14828 = ~1'b0 ;
  assign y14829 = ~n48016 ;
  assign y14830 = n48018 ;
  assign y14831 = n48019 ;
  assign y14832 = n48022 ;
  assign y14833 = ~n48023 ;
  assign y14834 = ~n48024 ;
  assign y14835 = n48027 ;
  assign y14836 = ~n48028 ;
  assign y14837 = ~n48030 ;
  assign y14838 = ~1'b0 ;
  assign y14839 = n48034 ;
  assign y14840 = ~n48035 ;
  assign y14841 = ~n48041 ;
  assign y14842 = n48042 ;
  assign y14843 = ~n48044 ;
  assign y14844 = n48046 ;
  assign y14845 = ~n48053 ;
  assign y14846 = n48057 ;
  assign y14847 = ~n48062 ;
  assign y14848 = n48063 ;
  assign y14849 = n48064 ;
  assign y14850 = ~1'b0 ;
  assign y14851 = ~1'b0 ;
  assign y14852 = n48069 ;
  assign y14853 = ~n48073 ;
  assign y14854 = n48075 ;
  assign y14855 = ~n48076 ;
  assign y14856 = ~n48080 ;
  assign y14857 = ~n48081 ;
  assign y14858 = ~1'b0 ;
  assign y14859 = ~n48085 ;
  assign y14860 = ~n48087 ;
  assign y14861 = n48089 ;
  assign y14862 = n48091 ;
  assign y14863 = ~n48092 ;
  assign y14864 = ~n48093 ;
  assign y14865 = n48096 ;
  assign y14866 = ~n22882 ;
  assign y14867 = n48100 ;
  assign y14868 = ~n48102 ;
  assign y14869 = ~n48103 ;
  assign y14870 = ~n48106 ;
  assign y14871 = n48107 ;
  assign y14872 = ~n48112 ;
  assign y14873 = n48113 ;
  assign y14874 = ~n48115 ;
  assign y14875 = ~n48116 ;
  assign y14876 = n48119 ;
  assign y14877 = ~n48121 ;
  assign y14878 = ~1'b0 ;
  assign y14879 = n48122 ;
  assign y14880 = n48124 ;
  assign y14881 = ~n48129 ;
  assign y14882 = ~n48132 ;
  assign y14883 = ~n48133 ;
  assign y14884 = ~n39418 ;
  assign y14885 = n48137 ;
  assign y14886 = ~n48140 ;
  assign y14887 = ~n48142 ;
  assign y14888 = ~1'b0 ;
  assign y14889 = n48145 ;
  assign y14890 = n48148 ;
  assign y14891 = n48150 ;
  assign y14892 = ~n48153 ;
  assign y14893 = n48155 ;
  assign y14894 = ~n48158 ;
  assign y14895 = n48161 ;
  assign y14896 = ~n48162 ;
  assign y14897 = n48164 ;
  assign y14898 = ~1'b0 ;
  assign y14899 = n48166 ;
  assign y14900 = ~n48171 ;
  assign y14901 = ~n48173 ;
  assign y14902 = ~n48174 ;
  assign y14903 = n48177 ;
  assign y14904 = ~n48179 ;
  assign y14905 = ~1'b0 ;
  assign y14906 = ~1'b0 ;
  assign y14907 = n48182 ;
  assign y14908 = ~n48184 ;
  assign y14909 = ~n48192 ;
  assign y14910 = n18665 ;
  assign y14911 = ~n48193 ;
  assign y14912 = ~n48196 ;
  assign y14913 = ~n48200 ;
  assign y14914 = ~1'b0 ;
  assign y14915 = ~n48209 ;
  assign y14916 = ~n48211 ;
  assign y14917 = ~n48212 ;
  assign y14918 = ~n48213 ;
  assign y14919 = ~n48214 ;
  assign y14920 = ~n48218 ;
  assign y14921 = ~n48225 ;
  assign y14922 = ~n48226 ;
  assign y14923 = ~n48230 ;
  assign y14924 = ~n48233 ;
  assign y14925 = ~n48235 ;
  assign y14926 = ~n48239 ;
  assign y14927 = n48240 ;
  assign y14928 = ~n48245 ;
  assign y14929 = ~n48247 ;
  assign y14930 = ~n48248 ;
  assign y14931 = ~n48249 ;
  assign y14932 = n10727 ;
  assign y14933 = ~n48250 ;
  assign y14934 = ~n48252 ;
  assign y14935 = n48254 ;
  assign y14936 = ~n48255 ;
  assign y14937 = n48256 ;
  assign y14938 = ~n48261 ;
  assign y14939 = ~n48262 ;
  assign y14940 = ~1'b0 ;
  assign y14941 = n48265 ;
  assign y14942 = ~1'b0 ;
  assign y14943 = ~n48267 ;
  assign y14944 = n48268 ;
  assign y14945 = n48278 ;
  assign y14946 = n48279 ;
  assign y14947 = n48285 ;
  assign y14948 = n48286 ;
  assign y14949 = ~n48288 ;
  assign y14950 = ~n48294 ;
  assign y14951 = ~n48299 ;
  assign y14952 = ~n48301 ;
  assign y14953 = ~n48302 ;
  assign y14954 = n48303 ;
  assign y14955 = ~n32769 ;
  assign y14956 = ~n48304 ;
  assign y14957 = ~n48308 ;
  assign y14958 = ~n48309 ;
  assign y14959 = ~1'b0 ;
  assign y14960 = ~1'b0 ;
  assign y14961 = ~n48315 ;
  assign y14962 = n48316 ;
  assign y14963 = ~n48318 ;
  assign y14964 = n48321 ;
  assign y14965 = n48324 ;
  assign y14966 = n48325 ;
  assign y14967 = n48326 ;
  assign y14968 = ~n48329 ;
  assign y14969 = ~1'b0 ;
  assign y14970 = ~n48334 ;
  assign y14971 = n48338 ;
  assign y14972 = n48339 ;
  assign y14973 = ~n48342 ;
  assign y14974 = ~n48344 ;
  assign y14975 = ~n48346 ;
  assign y14976 = n18000 ;
  assign y14977 = n48349 ;
  assign y14978 = n48351 ;
  assign y14979 = n48354 ;
  assign y14980 = ~n48356 ;
  assign y14981 = ~n48357 ;
  assign y14982 = ~n48360 ;
  assign y14983 = ~n48362 ;
  assign y14984 = ~n48363 ;
  assign y14985 = n48367 ;
  assign y14986 = n48368 ;
  assign y14987 = ~n48370 ;
  assign y14988 = ~1'b0 ;
  assign y14989 = n48372 ;
  assign y14990 = ~n48373 ;
  assign y14991 = n48375 ;
  assign y14992 = n48376 ;
  assign y14993 = ~n48382 ;
  assign y14994 = n48383 ;
  assign y14995 = ~n48394 ;
  assign y14996 = ~n48396 ;
  assign y14997 = n48398 ;
  assign y14998 = ~n48399 ;
  assign y14999 = ~1'b0 ;
  assign y15000 = n48400 ;
  assign y15001 = ~n48401 ;
  assign y15002 = ~n48402 ;
  assign y15003 = ~n48405 ;
  assign y15004 = ~n48406 ;
  assign y15005 = ~n48407 ;
  assign y15006 = n48409 ;
  assign y15007 = ~1'b0 ;
  assign y15008 = ~n48411 ;
  assign y15009 = n48412 ;
  assign y15010 = n2661 ;
  assign y15011 = n48414 ;
  assign y15012 = ~n25050 ;
  assign y15013 = n48415 ;
  assign y15014 = ~n48420 ;
  assign y15015 = ~n48427 ;
  assign y15016 = ~n48428 ;
  assign y15017 = ~n48429 ;
  assign y15018 = ~n48431 ;
  assign y15019 = n48432 ;
  assign y15020 = ~n48433 ;
  assign y15021 = n48434 ;
  assign y15022 = ~n48437 ;
  assign y15023 = ~1'b0 ;
  assign y15024 = ~n48438 ;
  assign y15025 = n48440 ;
  assign y15026 = ~n48447 ;
  assign y15027 = n48452 ;
  assign y15028 = n48454 ;
  assign y15029 = n48457 ;
  assign y15030 = 1'b0 ;
  assign y15031 = n48460 ;
  assign y15032 = ~1'b0 ;
  assign y15033 = n48461 ;
  assign y15034 = ~n48467 ;
  assign y15035 = n48468 ;
  assign y15036 = ~n48469 ;
  assign y15037 = n48471 ;
  assign y15038 = ~n48473 ;
  assign y15039 = n48474 ;
  assign y15040 = n48476 ;
  assign y15041 = ~1'b0 ;
  assign y15042 = n48479 ;
  assign y15043 = n48482 ;
  assign y15044 = ~n48483 ;
  assign y15045 = ~n48485 ;
  assign y15046 = ~n48487 ;
  assign y15047 = n48490 ;
  assign y15048 = n48492 ;
  assign y15049 = ~1'b0 ;
  assign y15050 = ~n48496 ;
  assign y15051 = n48498 ;
  assign y15052 = ~n48502 ;
  assign y15053 = n48503 ;
  assign y15054 = n48505 ;
  assign y15055 = ~n48506 ;
  assign y15056 = ~n48508 ;
  assign y15057 = n48511 ;
  assign y15058 = n48512 ;
  assign y15059 = ~n48514 ;
  assign y15060 = ~n48516 ;
  assign y15061 = n48519 ;
  assign y15062 = ~n48520 ;
  assign y15063 = n48523 ;
  assign y15064 = n48527 ;
  assign y15065 = n48529 ;
  assign y15066 = ~1'b0 ;
  assign y15067 = n48531 ;
  assign y15068 = ~n48534 ;
  assign y15069 = n48536 ;
  assign y15070 = n48537 ;
  assign y15071 = ~n48538 ;
  assign y15072 = n48539 ;
  assign y15073 = ~n48540 ;
  assign y15074 = ~n48541 ;
  assign y15075 = n48543 ;
  assign y15076 = ~n48550 ;
  assign y15077 = n46875 ;
  assign y15078 = ~n48555 ;
  assign y15079 = ~n48558 ;
  assign y15080 = ~n48560 ;
  assign y15081 = n48561 ;
  assign y15082 = ~n48565 ;
  assign y15083 = ~1'b0 ;
  assign y15084 = ~1'b0 ;
  assign y15085 = ~1'b0 ;
  assign y15086 = ~n48567 ;
  assign y15087 = n48568 ;
  assign y15088 = n48569 ;
  assign y15089 = ~n17378 ;
  assign y15090 = n48571 ;
  assign y15091 = n25877 ;
  assign y15092 = n48574 ;
  assign y15093 = ~n48579 ;
  assign y15094 = ~1'b0 ;
  assign y15095 = ~1'b0 ;
  assign y15096 = ~n48580 ;
  assign y15097 = n48581 ;
  assign y15098 = ~n48582 ;
  assign y15099 = n48583 ;
  assign y15100 = n48585 ;
  assign y15101 = ~1'b0 ;
  assign y15102 = n48586 ;
  assign y15103 = ~n48588 ;
  assign y15104 = ~n48590 ;
  assign y15105 = n48594 ;
  assign y15106 = ~n48595 ;
  assign y15107 = ~1'b0 ;
  assign y15108 = n48597 ;
  assign y15109 = n48599 ;
  assign y15110 = n48602 ;
  assign y15111 = n48604 ;
  assign y15112 = ~n48605 ;
  assign y15113 = ~n48607 ;
  assign y15114 = ~n6749 ;
  assign y15115 = ~n48608 ;
  assign y15116 = n48611 ;
  assign y15117 = ~n48614 ;
  assign y15118 = n48616 ;
  assign y15119 = ~1'b0 ;
  assign y15120 = 1'b0 ;
  assign y15121 = n48621 ;
  assign y15122 = ~n48623 ;
  assign y15123 = ~n48625 ;
  assign y15124 = n48626 ;
  assign y15125 = ~n48628 ;
  assign y15126 = n48631 ;
  assign y15127 = ~1'b0 ;
  assign y15128 = ~n48636 ;
  assign y15129 = ~n48638 ;
  assign y15130 = ~n48641 ;
  assign y15131 = ~n48648 ;
  assign y15132 = n48653 ;
  assign y15133 = n48654 ;
  assign y15134 = ~n48655 ;
  assign y15135 = n48661 ;
  assign y15136 = ~n48662 ;
  assign y15137 = n48667 ;
  assign y15138 = ~1'b0 ;
  assign y15139 = n35511 ;
  assign y15140 = ~n48669 ;
  assign y15141 = ~n48670 ;
  assign y15142 = ~n48672 ;
  assign y15143 = ~n48677 ;
  assign y15144 = n48684 ;
  assign y15145 = ~n48685 ;
  assign y15146 = ~n48687 ;
  assign y15147 = ~1'b0 ;
  assign y15148 = n48691 ;
  assign y15149 = n48694 ;
  assign y15150 = ~n48700 ;
  assign y15151 = n48705 ;
  assign y15152 = ~n48708 ;
  assign y15153 = ~n48712 ;
  assign y15154 = n48715 ;
  assign y15155 = ~n48718 ;
  assign y15156 = n48720 ;
  assign y15157 = ~n48721 ;
  assign y15158 = ~1'b0 ;
  assign y15159 = ~n48723 ;
  assign y15160 = n48724 ;
  assign y15161 = n48728 ;
  assign y15162 = n48729 ;
  assign y15163 = ~n48730 ;
  assign y15164 = n48734 ;
  assign y15165 = ~n48735 ;
  assign y15166 = ~1'b0 ;
  assign y15167 = ~1'b0 ;
  assign y15168 = n48736 ;
  assign y15169 = ~n48740 ;
  assign y15170 = ~n48741 ;
  assign y15171 = ~n48746 ;
  assign y15172 = ~n48749 ;
  assign y15173 = n48752 ;
  assign y15174 = ~n48754 ;
  assign y15175 = ~1'b0 ;
  assign y15176 = n48759 ;
  assign y15177 = n48760 ;
  assign y15178 = ~n48766 ;
  assign y15179 = ~n48767 ;
  assign y15180 = ~n48768 ;
  assign y15181 = ~n48778 ;
  assign y15182 = ~n48779 ;
  assign y15183 = ~n48780 ;
  assign y15184 = ~n48783 ;
  assign y15185 = n23614 ;
  assign y15186 = ~n48785 ;
  assign y15187 = ~1'b0 ;
  assign y15188 = n48787 ;
  assign y15189 = n48790 ;
  assign y15190 = n48792 ;
  assign y15191 = n48796 ;
  assign y15192 = n48797 ;
  assign y15193 = n48800 ;
  assign y15194 = n48802 ;
  assign y15195 = n48806 ;
  assign y15196 = ~1'b0 ;
  assign y15197 = n48807 ;
  assign y15198 = ~n48811 ;
  assign y15199 = n48812 ;
  assign y15200 = ~n48813 ;
  assign y15201 = ~n48814 ;
  assign y15202 = n48817 ;
  assign y15203 = ~n48820 ;
  assign y15204 = n48826 ;
  assign y15205 = ~n48827 ;
  assign y15206 = ~1'b0 ;
  assign y15207 = n48829 ;
  assign y15208 = n48830 ;
  assign y15209 = n48832 ;
  assign y15210 = n48839 ;
  assign y15211 = n48840 ;
  assign y15212 = ~n48841 ;
  assign y15213 = ~n48842 ;
  assign y15214 = ~n48844 ;
  assign y15215 = ~1'b0 ;
  assign y15216 = ~1'b0 ;
  assign y15217 = ~n48847 ;
  assign y15218 = n48848 ;
  assign y15219 = ~n48850 ;
  assign y15220 = n48852 ;
  assign y15221 = n48853 ;
  assign y15222 = n48857 ;
  assign y15223 = ~n48863 ;
  assign y15224 = ~1'b0 ;
  assign y15225 = ~1'b0 ;
  assign y15226 = n48865 ;
  assign y15227 = ~n48869 ;
  assign y15228 = n48872 ;
  assign y15229 = n48876 ;
  assign y15230 = ~n48877 ;
  assign y15231 = n48880 ;
  assign y15232 = n48884 ;
  assign y15233 = ~n48885 ;
  assign y15234 = n48886 ;
  assign y15235 = ~1'b0 ;
  assign y15236 = n48888 ;
  assign y15237 = n48891 ;
  assign y15238 = ~n48892 ;
  assign y15239 = ~n48894 ;
  assign y15240 = n48899 ;
  assign y15241 = ~n48903 ;
  assign y15242 = n48904 ;
  assign y15243 = n48906 ;
  assign y15244 = n48910 ;
  assign y15245 = ~n48911 ;
  assign y15246 = ~n48912 ;
  assign y15247 = n48917 ;
  assign y15248 = n48918 ;
  assign y15249 = ~n48920 ;
  assign y15250 = n48921 ;
  assign y15251 = ~1'b0 ;
  assign y15252 = ~n48923 ;
  assign y15253 = n48925 ;
  assign y15254 = ~n28665 ;
  assign y15255 = ~n38658 ;
  assign y15256 = ~n48926 ;
  assign y15257 = n48927 ;
  assign y15258 = n48930 ;
  assign y15259 = ~n48931 ;
  assign y15260 = n48934 ;
  assign y15261 = n48936 ;
  assign y15262 = ~n48939 ;
  assign y15263 = n48940 ;
  assign y15264 = ~n48943 ;
  assign y15265 = ~n48944 ;
  assign y15266 = n48946 ;
  assign y15267 = n48947 ;
  assign y15268 = ~n48949 ;
  assign y15269 = ~n48951 ;
  assign y15270 = ~n20745 ;
  assign y15271 = ~n48953 ;
  assign y15272 = ~n48955 ;
  assign y15273 = n48957 ;
  assign y15274 = ~n48963 ;
  assign y15275 = ~n48967 ;
  assign y15276 = n48968 ;
  assign y15277 = ~n48970 ;
  assign y15278 = n48971 ;
  assign y15279 = n48973 ;
  assign y15280 = ~n48975 ;
  assign y15281 = ~n48977 ;
  assign y15282 = ~n48979 ;
  assign y15283 = ~n48980 ;
  assign y15284 = ~n48983 ;
  assign y15285 = n48986 ;
  assign y15286 = n48987 ;
  assign y15287 = ~n48988 ;
  assign y15288 = ~1'b0 ;
  assign y15289 = ~1'b0 ;
  assign y15290 = ~1'b0 ;
  assign y15291 = ~1'b0 ;
  assign y15292 = ~n48991 ;
  assign y15293 = ~n48993 ;
  assign y15294 = n48994 ;
  assign y15295 = n49003 ;
  assign y15296 = n49004 ;
  assign y15297 = ~n49011 ;
  assign y15298 = n49013 ;
  assign y15299 = n49017 ;
  assign y15300 = ~1'b0 ;
  assign y15301 = ~n49020 ;
  assign y15302 = ~1'b0 ;
  assign y15303 = ~n49021 ;
  assign y15304 = n49022 ;
  assign y15305 = ~n49023 ;
  assign y15306 = ~n49026 ;
  assign y15307 = ~n49027 ;
  assign y15308 = n49028 ;
  assign y15309 = n49029 ;
  assign y15310 = ~n49031 ;
  assign y15311 = ~n49033 ;
  assign y15312 = ~n49036 ;
  assign y15313 = ~n49039 ;
  assign y15314 = n49040 ;
  assign y15315 = n49046 ;
  assign y15316 = ~n49047 ;
  assign y15317 = n49048 ;
  assign y15318 = n49049 ;
  assign y15319 = ~n49050 ;
  assign y15320 = n49056 ;
  assign y15321 = ~1'b0 ;
  assign y15322 = ~1'b0 ;
  assign y15323 = n49057 ;
  assign y15324 = n38408 ;
  assign y15325 = n49058 ;
  assign y15326 = n49060 ;
  assign y15327 = n49063 ;
  assign y15328 = ~n49068 ;
  assign y15329 = ~n49073 ;
  assign y15330 = ~n49076 ;
  assign y15331 = ~1'b0 ;
  assign y15332 = n49078 ;
  assign y15333 = n49081 ;
  assign y15334 = ~n49082 ;
  assign y15335 = ~n49083 ;
  assign y15336 = n49088 ;
  assign y15337 = n49089 ;
  assign y15338 = ~n49092 ;
  assign y15339 = n49096 ;
  assign y15340 = n49098 ;
  assign y15341 = n49099 ;
  assign y15342 = ~n49101 ;
  assign y15343 = ~n49102 ;
  assign y15344 = n49103 ;
  assign y15345 = ~n49105 ;
  assign y15346 = n49108 ;
  assign y15347 = ~n49109 ;
  assign y15348 = n49111 ;
  assign y15349 = ~n49115 ;
  assign y15350 = n49119 ;
  assign y15351 = ~n49123 ;
  assign y15352 = ~1'b0 ;
  assign y15353 = n49125 ;
  assign y15354 = ~n49128 ;
  assign y15355 = n49129 ;
  assign y15356 = ~n49130 ;
  assign y15357 = ~n49133 ;
  assign y15358 = ~n49137 ;
  assign y15359 = ~n49139 ;
  assign y15360 = ~n49143 ;
  assign y15361 = ~1'b0 ;
  assign y15362 = ~n49148 ;
  assign y15363 = ~n49150 ;
  assign y15364 = ~n49152 ;
  assign y15365 = ~n49154 ;
  assign y15366 = ~n49156 ;
  assign y15367 = ~n49158 ;
  assign y15368 = n49159 ;
  assign y15369 = ~n49160 ;
  assign y15370 = ~n49162 ;
  assign y15371 = n49164 ;
  assign y15372 = ~1'b0 ;
  assign y15373 = n49165 ;
  assign y15374 = ~n49171 ;
  assign y15375 = ~n49174 ;
  assign y15376 = ~n49177 ;
  assign y15377 = n49178 ;
  assign y15378 = ~n49179 ;
  assign y15379 = n49180 ;
  assign y15380 = n49182 ;
  assign y15381 = ~n49185 ;
  assign y15382 = ~n49187 ;
  assign y15383 = ~n49188 ;
  assign y15384 = ~n49189 ;
  assign y15385 = ~n49190 ;
  assign y15386 = n49191 ;
  assign y15387 = n49193 ;
  assign y15388 = ~n49196 ;
  assign y15389 = ~1'b0 ;
  assign y15390 = ~n49205 ;
  assign y15391 = n49207 ;
  assign y15392 = ~n49209 ;
  assign y15393 = ~n49212 ;
  assign y15394 = ~n49213 ;
  assign y15395 = n49215 ;
  assign y15396 = ~n49216 ;
  assign y15397 = n49217 ;
  assign y15398 = ~n49218 ;
  assign y15399 = n49220 ;
  assign y15400 = ~n49222 ;
  assign y15401 = n49226 ;
  assign y15402 = ~n49229 ;
  assign y15403 = n49231 ;
  assign y15404 = n49232 ;
  assign y15405 = n49233 ;
  assign y15406 = n49234 ;
  assign y15407 = ~n49236 ;
  assign y15408 = ~n49238 ;
  assign y15409 = n49241 ;
  assign y15410 = n49242 ;
  assign y15411 = ~1'b0 ;
  assign y15412 = n49243 ;
  assign y15413 = ~n49245 ;
  assign y15414 = n49249 ;
  assign y15415 = ~n49250 ;
  assign y15416 = n49251 ;
  assign y15417 = n49254 ;
  assign y15418 = n49256 ;
  assign y15419 = n49259 ;
  assign y15420 = n49261 ;
  assign y15421 = ~n49270 ;
  assign y15422 = ~n49272 ;
  assign y15423 = ~n49273 ;
  assign y15424 = ~n49278 ;
  assign y15425 = n49281 ;
  assign y15426 = ~1'b0 ;
  assign y15427 = ~n49283 ;
  assign y15428 = ~n49286 ;
  assign y15429 = n49289 ;
  assign y15430 = n49290 ;
  assign y15431 = n49291 ;
  assign y15432 = n49295 ;
  assign y15433 = ~n49298 ;
  assign y15434 = ~1'b0 ;
  assign y15435 = ~n49301 ;
  assign y15436 = ~1'b0 ;
  assign y15437 = ~n49303 ;
  assign y15438 = n49308 ;
  assign y15439 = ~n49309 ;
  assign y15440 = ~n49311 ;
  assign y15441 = n49317 ;
  assign y15442 = ~n49322 ;
  assign y15443 = ~n49323 ;
  assign y15444 = ~n49325 ;
  assign y15445 = ~1'b0 ;
  assign y15446 = ~n49327 ;
  assign y15447 = n49328 ;
  assign y15448 = n49331 ;
  assign y15449 = n49337 ;
  assign y15450 = n49339 ;
  assign y15451 = ~n49341 ;
  assign y15452 = n49344 ;
  assign y15453 = n49346 ;
  assign y15454 = ~1'b0 ;
  assign y15455 = ~1'b0 ;
  assign y15456 = ~1'b0 ;
  assign y15457 = n49350 ;
  assign y15458 = n49352 ;
  assign y15459 = ~n49357 ;
  assign y15460 = n49360 ;
  assign y15461 = n49361 ;
  assign y15462 = ~n49365 ;
  assign y15463 = ~1'b0 ;
  assign y15464 = ~n49367 ;
  assign y15465 = ~n49370 ;
  assign y15466 = ~n49377 ;
  assign y15467 = ~n49378 ;
  assign y15468 = ~n49381 ;
  assign y15469 = ~n49383 ;
  assign y15470 = ~n49385 ;
  assign y15471 = n49391 ;
  assign y15472 = ~1'b0 ;
  assign y15473 = n49394 ;
  assign y15474 = ~n49396 ;
  assign y15475 = ~n49399 ;
  assign y15476 = n49402 ;
  assign y15477 = ~n49406 ;
  assign y15478 = ~n49407 ;
  assign y15479 = n49413 ;
  assign y15480 = ~n49414 ;
  assign y15481 = n49421 ;
  assign y15482 = ~1'b0 ;
  assign y15483 = n49422 ;
  assign y15484 = ~1'b0 ;
  assign y15485 = ~1'b0 ;
  assign y15486 = ~n49423 ;
  assign y15487 = ~n49425 ;
  assign y15488 = n49428 ;
  assign y15489 = ~n49429 ;
  assign y15490 = ~n49437 ;
  assign y15491 = n49438 ;
  assign y15492 = n49441 ;
  assign y15493 = n49443 ;
  assign y15494 = ~n49446 ;
  assign y15495 = ~1'b0 ;
  assign y15496 = n49453 ;
  assign y15497 = ~n49454 ;
  assign y15498 = ~n49455 ;
  assign y15499 = n49457 ;
  assign y15500 = n49464 ;
  assign y15501 = ~n49466 ;
  assign y15502 = n49470 ;
  assign y15503 = ~n49473 ;
  assign y15504 = n49475 ;
  assign y15505 = ~n49477 ;
  assign y15506 = ~n49482 ;
  assign y15507 = ~n49486 ;
  assign y15508 = n49490 ;
  assign y15509 = ~n49495 ;
  assign y15510 = ~n49497 ;
  assign y15511 = ~n49498 ;
  assign y15512 = ~n49501 ;
  assign y15513 = ~n49502 ;
  assign y15514 = ~n49504 ;
  assign y15515 = 1'b0 ;
  assign y15516 = n49511 ;
  assign y15517 = n49514 ;
  assign y15518 = ~n49516 ;
  assign y15519 = n49518 ;
  assign y15520 = n49523 ;
  assign y15521 = n49524 ;
  assign y15522 = ~n49527 ;
  assign y15523 = n49529 ;
  assign y15524 = ~1'b0 ;
  assign y15525 = ~1'b0 ;
  assign y15526 = ~n49530 ;
  assign y15527 = ~n7199 ;
  assign y15528 = ~n49532 ;
  assign y15529 = ~n49533 ;
  assign y15530 = ~n49534 ;
  assign y15531 = ~n49535 ;
  assign y15532 = n49538 ;
  assign y15533 = ~n49540 ;
  assign y15534 = n49542 ;
  assign y15535 = ~1'b0 ;
  assign y15536 = n49544 ;
  assign y15537 = ~n49545 ;
  assign y15538 = n49547 ;
  assign y15539 = n49550 ;
  assign y15540 = ~n49553 ;
  assign y15541 = n49556 ;
  assign y15542 = n49558 ;
  assign y15543 = ~n49560 ;
  assign y15544 = ~n49563 ;
  assign y15545 = ~1'b0 ;
  assign y15546 = ~n49569 ;
  assign y15547 = n49570 ;
  assign y15548 = ~n49573 ;
  assign y15549 = ~n49579 ;
  assign y15550 = ~n49581 ;
  assign y15551 = ~n49583 ;
  assign y15552 = ~n49591 ;
  assign y15553 = ~n49593 ;
  assign y15554 = ~n49595 ;
  assign y15555 = ~n49603 ;
  assign y15556 = ~1'b0 ;
  assign y15557 = ~n4836 ;
  assign y15558 = ~n49604 ;
  assign y15559 = ~n49609 ;
  assign y15560 = n49612 ;
  assign y15561 = n49614 ;
  assign y15562 = n49615 ;
  assign y15563 = n49616 ;
  assign y15564 = n49619 ;
  assign y15565 = ~n49620 ;
  assign y15566 = ~1'b0 ;
  assign y15567 = ~n49621 ;
  assign y15568 = n49622 ;
  assign y15569 = ~n49623 ;
  assign y15570 = ~n49625 ;
  assign y15571 = ~n49626 ;
  assign y15572 = ~n49629 ;
  assign y15573 = ~n49630 ;
  assign y15574 = ~n49631 ;
  assign y15575 = ~1'b0 ;
  assign y15576 = ~n49635 ;
  assign y15577 = ~n49639 ;
  assign y15578 = ~n49641 ;
  assign y15579 = ~n49642 ;
  assign y15580 = n49643 ;
  assign y15581 = ~n49645 ;
  assign y15582 = n49647 ;
  assign y15583 = ~n49648 ;
  assign y15584 = ~1'b0 ;
  assign y15585 = ~1'b0 ;
  assign y15586 = ~n49651 ;
  assign y15587 = ~1'b0 ;
  assign y15588 = n49654 ;
  assign y15589 = n49656 ;
  assign y15590 = n49660 ;
  assign y15591 = ~n49663 ;
  assign y15592 = n49666 ;
  assign y15593 = n49671 ;
  assign y15594 = n49673 ;
  assign y15595 = n49675 ;
  assign y15596 = n49679 ;
  assign y15597 = ~1'b0 ;
  assign y15598 = n49682 ;
  assign y15599 = n11785 ;
  assign y15600 = n49693 ;
  assign y15601 = ~n49694 ;
  assign y15602 = ~n49695 ;
  assign y15603 = n49701 ;
  assign y15604 = n49705 ;
  assign y15605 = n49706 ;
  assign y15606 = n49709 ;
  assign y15607 = n49716 ;
  assign y15608 = ~n49718 ;
  assign y15609 = ~n49721 ;
  assign y15610 = n49724 ;
  assign y15611 = n49725 ;
  assign y15612 = ~n49728 ;
  assign y15613 = n49729 ;
  assign y15614 = ~n49731 ;
  assign y15615 = ~1'b0 ;
  assign y15616 = n49736 ;
  assign y15617 = n49737 ;
  assign y15618 = n49738 ;
  assign y15619 = ~n49739 ;
  assign y15620 = ~n49740 ;
  assign y15621 = ~n49743 ;
  assign y15622 = ~n49744 ;
  assign y15623 = n49749 ;
  assign y15624 = ~n49752 ;
  assign y15625 = ~n49755 ;
  assign y15626 = ~1'b0 ;
  assign y15627 = n49757 ;
  assign y15628 = ~n49758 ;
  assign y15629 = ~n49759 ;
  assign y15630 = n24680 ;
  assign y15631 = n49761 ;
  assign y15632 = ~n49766 ;
  assign y15633 = n49771 ;
  assign y15634 = ~n49776 ;
  assign y15635 = n49780 ;
  assign y15636 = ~1'b0 ;
  assign y15637 = n49784 ;
  assign y15638 = ~n49786 ;
  assign y15639 = ~n49787 ;
  assign y15640 = n49788 ;
  assign y15641 = ~n49790 ;
  assign y15642 = n49792 ;
  assign y15643 = ~n49796 ;
  assign y15644 = ~1'b0 ;
  assign y15645 = ~n49797 ;
  assign y15646 = ~1'b0 ;
  assign y15647 = ~1'b0 ;
  assign y15648 = ~n49798 ;
  assign y15649 = n49801 ;
  assign y15650 = n49802 ;
  assign y15651 = n49803 ;
  assign y15652 = n49806 ;
  assign y15653 = n49807 ;
  assign y15654 = ~n49808 ;
  assign y15655 = ~n49810 ;
  assign y15656 = ~n49813 ;
  assign y15657 = ~n49817 ;
  assign y15658 = n49818 ;
  assign y15659 = ~n49824 ;
  assign y15660 = n49827 ;
  assign y15661 = n49828 ;
  assign y15662 = n49831 ;
  assign y15663 = ~n49832 ;
  assign y15664 = ~1'b0 ;
  assign y15665 = ~n49835 ;
  assign y15666 = n49841 ;
  assign y15667 = ~1'b0 ;
  assign y15668 = ~n49842 ;
  assign y15669 = ~n49846 ;
  assign y15670 = ~n49849 ;
  assign y15671 = n49852 ;
  assign y15672 = ~n49853 ;
  assign y15673 = ~n49854 ;
  assign y15674 = ~n49855 ;
  assign y15675 = n49857 ;
  assign y15676 = ~n49862 ;
  assign y15677 = ~n49865 ;
  assign y15678 = ~n49867 ;
  assign y15679 = ~n49872 ;
  assign y15680 = ~n49875 ;
  assign y15681 = ~n49878 ;
  assign y15682 = ~n49882 ;
  assign y15683 = ~n49885 ;
  assign y15684 = ~n49887 ;
  assign y15685 = ~1'b0 ;
  assign y15686 = ~n49889 ;
  assign y15687 = ~n49890 ;
  assign y15688 = ~n49893 ;
  assign y15689 = ~n49896 ;
  assign y15690 = n49898 ;
  assign y15691 = n49900 ;
  assign y15692 = n49903 ;
  assign y15693 = ~n49905 ;
  assign y15694 = n49907 ;
  assign y15695 = ~1'b0 ;
  assign y15696 = ~n49910 ;
  assign y15697 = n49916 ;
  assign y15698 = n49922 ;
  assign y15699 = n49923 ;
  assign y15700 = n49928 ;
  assign y15701 = ~n49931 ;
  assign y15702 = n49932 ;
  assign y15703 = ~n49933 ;
  assign y15704 = ~n49935 ;
  assign y15705 = n49936 ;
  assign y15706 = ~1'b0 ;
  assign y15707 = ~n49937 ;
  assign y15708 = ~n49939 ;
  assign y15709 = n49941 ;
  assign y15710 = ~n49946 ;
  assign y15711 = n49947 ;
  assign y15712 = ~1'b0 ;
  assign y15713 = ~n49956 ;
  assign y15714 = n49961 ;
  assign y15715 = ~n49968 ;
  assign y15716 = n5986 ;
  assign y15717 = n49969 ;
  assign y15718 = ~n49970 ;
  assign y15719 = ~n49971 ;
  assign y15720 = n49974 ;
  assign y15721 = n49975 ;
  assign y15722 = n49976 ;
  assign y15723 = ~1'b0 ;
  assign y15724 = ~n49979 ;
  assign y15725 = n49980 ;
  assign y15726 = n49982 ;
  assign y15727 = ~n49983 ;
  assign y15728 = n49984 ;
  assign y15729 = ~n49985 ;
  assign y15730 = n49986 ;
  assign y15731 = ~n49989 ;
  assign y15732 = ~n49990 ;
  assign y15733 = ~n49994 ;
  assign y15734 = n49999 ;
  assign y15735 = ~n50004 ;
  assign y15736 = ~n50008 ;
  assign y15737 = n50009 ;
  assign y15738 = n50011 ;
  assign y15739 = ~n50015 ;
  assign y15740 = ~n49104 ;
  assign y15741 = n50020 ;
  assign y15742 = ~n50021 ;
  assign y15743 = ~n50023 ;
  assign y15744 = ~1'b0 ;
  assign y15745 = ~n50025 ;
  assign y15746 = n50027 ;
  assign y15747 = n50028 ;
  assign y15748 = n50030 ;
  assign y15749 = n50035 ;
  assign y15750 = n50036 ;
  assign y15751 = n50037 ;
  assign y15752 = n50044 ;
  assign y15753 = ~1'b0 ;
  assign y15754 = n50051 ;
  assign y15755 = n50052 ;
  assign y15756 = n50056 ;
  assign y15757 = ~n50059 ;
  assign y15758 = n50062 ;
  assign y15759 = n50065 ;
  assign y15760 = ~n50066 ;
  assign y15761 = ~n50069 ;
  assign y15762 = ~n50070 ;
  assign y15763 = ~1'b0 ;
  assign y15764 = n50072 ;
  assign y15765 = n50073 ;
  assign y15766 = n50075 ;
  assign y15767 = n50080 ;
  assign y15768 = n50081 ;
  assign y15769 = n50087 ;
  assign y15770 = ~n50090 ;
  assign y15771 = ~n50091 ;
  assign y15772 = n50092 ;
  assign y15773 = ~n50094 ;
  assign y15774 = n50097 ;
  assign y15775 = ~1'b0 ;
  assign y15776 = n50100 ;
  assign y15777 = n17840 ;
  assign y15778 = ~n50101 ;
  assign y15779 = ~n50104 ;
  assign y15780 = n50108 ;
  assign y15781 = ~n50109 ;
  assign y15782 = ~n50110 ;
  assign y15783 = ~n50111 ;
  assign y15784 = n18423 ;
  assign y15785 = n50118 ;
  assign y15786 = ~1'b0 ;
  assign y15787 = ~n50119 ;
  assign y15788 = n50121 ;
  assign y15789 = n50122 ;
  assign y15790 = n50126 ;
  assign y15791 = ~n50128 ;
  assign y15792 = ~n50131 ;
  assign y15793 = ~1'b0 ;
  assign y15794 = ~1'b0 ;
  assign y15795 = ~1'b0 ;
  assign y15796 = ~n50132 ;
  assign y15797 = n50133 ;
  assign y15798 = n50141 ;
  assign y15799 = ~n50142 ;
  assign y15800 = n50144 ;
  assign y15801 = ~n50146 ;
  assign y15802 = ~1'b0 ;
  assign y15803 = n50148 ;
  assign y15804 = n50154 ;
  assign y15805 = ~n50155 ;
  assign y15806 = ~n50156 ;
  assign y15807 = n50157 ;
  assign y15808 = n50158 ;
  assign y15809 = ~n50159 ;
  assign y15810 = ~1'b0 ;
  assign y15811 = 1'b0 ;
  assign y15812 = n50162 ;
  assign y15813 = ~n50164 ;
  assign y15814 = ~n50165 ;
  assign y15815 = ~n50166 ;
  assign y15816 = n50176 ;
  assign y15817 = n50178 ;
  assign y15818 = n50184 ;
  assign y15819 = n50185 ;
  assign y15820 = ~n50188 ;
  assign y15821 = n50194 ;
  assign y15822 = n50195 ;
  assign y15823 = ~1'b0 ;
  assign y15824 = n50196 ;
  assign y15825 = ~n50201 ;
  assign y15826 = ~n958 ;
  assign y15827 = n50203 ;
  assign y15828 = ~n50205 ;
  assign y15829 = ~n50207 ;
  assign y15830 = ~n50209 ;
  assign y15831 = n50211 ;
  assign y15832 = n50215 ;
  assign y15833 = ~1'b0 ;
  assign y15834 = n50220 ;
  assign y15835 = n50226 ;
  assign y15836 = ~n50227 ;
  assign y15837 = ~n50229 ;
  assign y15838 = n50232 ;
  assign y15839 = n50235 ;
  assign y15840 = n50237 ;
  assign y15841 = ~1'b0 ;
  assign y15842 = ~n50238 ;
  assign y15843 = n50242 ;
  assign y15844 = n50244 ;
  assign y15845 = ~n50245 ;
  assign y15846 = n50246 ;
  assign y15847 = ~n50247 ;
  assign y15848 = ~n50248 ;
  assign y15849 = ~n50251 ;
  assign y15850 = n50253 ;
  assign y15851 = ~1'b0 ;
  assign y15852 = ~1'b0 ;
  assign y15853 = ~1'b0 ;
  assign y15854 = ~n50258 ;
  assign y15855 = ~n50259 ;
  assign y15856 = n50261 ;
  assign y15857 = n50263 ;
  assign y15858 = ~n50265 ;
  assign y15859 = ~n50266 ;
  assign y15860 = ~n50269 ;
  assign y15861 = n50271 ;
  assign y15862 = n50275 ;
  assign y15863 = ~1'b0 ;
  assign y15864 = ~n50284 ;
  assign y15865 = n50285 ;
  assign y15866 = ~n50286 ;
  assign y15867 = n50288 ;
  assign y15868 = n50289 ;
  assign y15869 = n50296 ;
  assign y15870 = ~n50298 ;
  assign y15871 = n50303 ;
  assign y15872 = n50307 ;
  assign y15873 = n50309 ;
  assign y15874 = n50312 ;
  assign y15875 = n50315 ;
  assign y15876 = n50318 ;
  assign y15877 = ~n50319 ;
  assign y15878 = ~n50320 ;
  assign y15879 = ~1'b0 ;
  assign y15880 = ~n50322 ;
  assign y15881 = ~n50336 ;
  assign y15882 = n50337 ;
  assign y15883 = ~n50339 ;
  assign y15884 = n50340 ;
  assign y15885 = ~n50342 ;
  assign y15886 = ~n50346 ;
  assign y15887 = n50348 ;
  assign y15888 = ~1'b0 ;
  assign y15889 = ~n50349 ;
  assign y15890 = n50351 ;
  assign y15891 = n50352 ;
  assign y15892 = ~n50353 ;
  assign y15893 = n50355 ;
  assign y15894 = n50357 ;
  assign y15895 = ~n50358 ;
  assign y15896 = ~n50359 ;
  assign y15897 = ~n50360 ;
  assign y15898 = ~n50363 ;
  assign y15899 = ~n50365 ;
  assign y15900 = ~n50367 ;
  assign y15901 = n50369 ;
  assign y15902 = ~n50371 ;
  assign y15903 = n50372 ;
  assign y15904 = ~n50373 ;
  assign y15905 = n50378 ;
  assign y15906 = ~n50379 ;
  assign y15907 = ~1'b0 ;
  assign y15908 = n50382 ;
  assign y15909 = ~n50385 ;
  assign y15910 = ~n50387 ;
  assign y15911 = ~n50388 ;
  assign y15912 = n50390 ;
  assign y15913 = n50394 ;
  assign y15914 = ~n50398 ;
  assign y15915 = ~n50402 ;
  assign y15916 = n50403 ;
  assign y15917 = n50404 ;
  assign y15918 = ~n50406 ;
  assign y15919 = ~n50407 ;
  assign y15920 = ~n50412 ;
  assign y15921 = ~n50414 ;
  assign y15922 = n50417 ;
  assign y15923 = ~n50419 ;
  assign y15924 = n50420 ;
  assign y15925 = n50424 ;
  assign y15926 = ~n50427 ;
  assign y15927 = n50428 ;
  assign y15928 = n50432 ;
  assign y15929 = ~1'b0 ;
  assign y15930 = n50433 ;
  assign y15931 = ~n50435 ;
  assign y15932 = n50440 ;
  assign y15933 = n50443 ;
  assign y15934 = ~1'b0 ;
  assign y15935 = ~n50446 ;
  assign y15936 = ~n50447 ;
  assign y15937 = n50448 ;
  assign y15938 = ~n50449 ;
  assign y15939 = ~n50454 ;
  assign y15940 = ~1'b0 ;
  assign y15941 = ~1'b0 ;
  assign y15942 = n50456 ;
  assign y15943 = n50459 ;
  assign y15944 = n50463 ;
  assign y15945 = n50467 ;
  assign y15946 = ~n50473 ;
  assign y15947 = ~n50474 ;
  assign y15948 = ~n50476 ;
  assign y15949 = ~n50477 ;
  assign y15950 = ~n50478 ;
  assign y15951 = ~1'b0 ;
  assign y15952 = n50481 ;
  assign y15953 = n50482 ;
  assign y15954 = ~n50485 ;
  assign y15955 = ~n50490 ;
  assign y15956 = ~n50499 ;
  assign y15957 = n50500 ;
  assign y15958 = ~n50501 ;
  assign y15959 = ~n50506 ;
  assign y15960 = n50507 ;
  assign y15961 = ~1'b0 ;
  assign y15962 = n50509 ;
  assign y15963 = ~n50510 ;
  assign y15964 = n50511 ;
  assign y15965 = n50513 ;
  assign y15966 = ~n50514 ;
  assign y15967 = ~n50515 ;
  assign y15968 = ~n50519 ;
  assign y15969 = n50520 ;
  assign y15970 = ~n50524 ;
  assign y15971 = n50528 ;
  assign y15972 = n50529 ;
  assign y15973 = ~n50531 ;
  assign y15974 = n50533 ;
  assign y15975 = ~n50534 ;
  assign y15976 = n11323 ;
  assign y15977 = ~n50536 ;
  assign y15978 = ~n50538 ;
  assign y15979 = ~n50539 ;
  assign y15980 = ~1'b0 ;
  assign y15981 = n50541 ;
  assign y15982 = n50542 ;
  assign y15983 = ~n50543 ;
  assign y15984 = n50544 ;
  assign y15985 = ~n50545 ;
  assign y15986 = n50546 ;
  assign y15987 = n50548 ;
  assign y15988 = ~n50554 ;
  assign y15989 = ~n50555 ;
  assign y15990 = 1'b0 ;
  assign y15991 = n50556 ;
  assign y15992 = ~n50559 ;
  assign y15993 = ~n50561 ;
  assign y15994 = n50562 ;
  assign y15995 = n50565 ;
  assign y15996 = n50566 ;
  assign y15997 = ~n50572 ;
  assign y15998 = ~n50576 ;
  assign y15999 = ~n50578 ;
  assign y16000 = ~1'b0 ;
  assign y16001 = n50579 ;
  assign y16002 = n50580 ;
  assign y16003 = ~n50582 ;
  assign y16004 = ~n50585 ;
  assign y16005 = n50588 ;
  assign y16006 = ~n50591 ;
  assign y16007 = n50592 ;
  assign y16008 = ~n50595 ;
  assign y16009 = ~1'b0 ;
  assign y16010 = n50597 ;
  assign y16011 = ~1'b0 ;
  assign y16012 = ~n50599 ;
  assign y16013 = n50600 ;
  assign y16014 = n50602 ;
  assign y16015 = ~n50603 ;
  assign y16016 = n50605 ;
  assign y16017 = ~n50606 ;
  assign y16018 = n50607 ;
  assign y16019 = n50611 ;
  assign y16020 = ~n50615 ;
  assign y16021 = ~n50617 ;
  assign y16022 = n50620 ;
  assign y16023 = ~1'b0 ;
  assign y16024 = n50624 ;
  assign y16025 = n50625 ;
  assign y16026 = ~n50629 ;
  assign y16027 = n50630 ;
  assign y16028 = n50634 ;
  assign y16029 = n50638 ;
  assign y16030 = n50642 ;
  assign y16031 = ~n50644 ;
  assign y16032 = ~n50645 ;
  assign y16033 = ~n50647 ;
  assign y16034 = n50648 ;
  assign y16035 = ~n50649 ;
  assign y16036 = ~n50653 ;
  assign y16037 = ~1'b0 ;
  assign y16038 = ~1'b0 ;
  assign y16039 = n50655 ;
  assign y16040 = ~n50656 ;
  assign y16041 = n50660 ;
  assign y16042 = ~n50666 ;
  assign y16043 = n50668 ;
  assign y16044 = ~n50670 ;
  assign y16045 = n50672 ;
  assign y16046 = ~n50675 ;
  assign y16047 = ~n50676 ;
  assign y16048 = ~n50678 ;
  assign y16049 = n50685 ;
  assign y16050 = ~1'b0 ;
  assign y16051 = n50686 ;
  assign y16052 = ~n50691 ;
  assign y16053 = n50694 ;
  assign y16054 = n50695 ;
  assign y16055 = ~n50697 ;
  assign y16056 = ~n50700 ;
  assign y16057 = ~n50703 ;
  assign y16058 = ~1'b0 ;
  assign y16059 = n50706 ;
  assign y16060 = ~n50710 ;
  assign y16061 = ~1'b0 ;
  assign y16062 = n50713 ;
  assign y16063 = n50716 ;
  assign y16064 = n50720 ;
  assign y16065 = n50721 ;
  assign y16066 = ~n50723 ;
  assign y16067 = n50726 ;
  assign y16068 = n50729 ;
  assign y16069 = ~1'b0 ;
  assign y16070 = ~n50734 ;
  assign y16071 = n50738 ;
  assign y16072 = ~n50739 ;
  assign y16073 = ~n50740 ;
  assign y16074 = n50743 ;
  assign y16075 = n50744 ;
  assign y16076 = n50745 ;
  assign y16077 = n50747 ;
  assign y16078 = ~n50749 ;
  assign y16079 = n50750 ;
  assign y16080 = ~n50752 ;
  assign y16081 = n50753 ;
  assign y16082 = ~n50755 ;
  assign y16083 = ~n50757 ;
  assign y16084 = n50758 ;
  assign y16085 = n50761 ;
  assign y16086 = ~n50766 ;
  assign y16087 = n50768 ;
  assign y16088 = n50771 ;
  assign y16089 = ~n50772 ;
  assign y16090 = n50773 ;
  assign y16091 = ~n50775 ;
  assign y16092 = ~1'b0 ;
  assign y16093 = n50777 ;
  assign y16094 = ~n50778 ;
  assign y16095 = ~n50779 ;
  assign y16096 = ~n50780 ;
  assign y16097 = ~n50786 ;
  assign y16098 = n50787 ;
  assign y16099 = n50789 ;
  assign y16100 = ~1'b0 ;
  assign y16101 = n50794 ;
  assign y16102 = ~n50796 ;
  assign y16103 = n50798 ;
  assign y16104 = n50799 ;
  assign y16105 = n50802 ;
  assign y16106 = n50805 ;
  assign y16107 = n50808 ;
  assign y16108 = n50811 ;
  assign y16109 = n50816 ;
  assign y16110 = ~1'b0 ;
  assign y16111 = ~1'b0 ;
  assign y16112 = ~n50820 ;
  assign y16113 = n50822 ;
  assign y16114 = n50823 ;
  assign y16115 = ~n50824 ;
  assign y16116 = ~n50826 ;
  assign y16117 = n50827 ;
  assign y16118 = ~n50829 ;
  assign y16119 = ~n50832 ;
  assign y16120 = ~1'b0 ;
  assign y16121 = n50834 ;
  assign y16122 = ~1'b0 ;
  assign y16123 = ~n50836 ;
  assign y16124 = ~1'b0 ;
  assign y16125 = ~n50840 ;
  assign y16126 = ~n50841 ;
  assign y16127 = n50844 ;
  assign y16128 = n50846 ;
  assign y16129 = ~n50849 ;
  assign y16130 = ~n50851 ;
  assign y16131 = ~n2958 ;
  assign y16132 = ~1'b0 ;
  assign y16133 = ~1'b0 ;
  assign y16134 = ~1'b0 ;
  assign y16135 = ~1'b0 ;
  assign y16136 = n50853 ;
  assign y16137 = n50855 ;
  assign y16138 = n50856 ;
  assign y16139 = ~n50857 ;
  assign y16140 = ~n50860 ;
  assign y16141 = ~n50865 ;
  assign y16142 = ~n50867 ;
  assign y16143 = n50869 ;
  assign y16144 = n50873 ;
  assign y16145 = ~n50879 ;
  assign y16146 = n50882 ;
  assign y16147 = n50884 ;
  assign y16148 = n50885 ;
  assign y16149 = n50892 ;
  assign y16150 = n50894 ;
  assign y16151 = n50895 ;
  assign y16152 = ~n50896 ;
  assign y16153 = ~n50898 ;
  assign y16154 = ~1'b0 ;
  assign y16155 = ~n50902 ;
  assign y16156 = ~n50903 ;
  assign y16157 = n50905 ;
  assign y16158 = ~n50906 ;
  assign y16159 = ~n50908 ;
  assign y16160 = n50909 ;
  assign y16161 = n50913 ;
  assign y16162 = n50916 ;
  assign y16163 = n50917 ;
  assign y16164 = ~n50923 ;
  assign y16165 = n50924 ;
  assign y16166 = n50926 ;
  assign y16167 = ~n50927 ;
  assign y16168 = n50928 ;
  assign y16169 = n50929 ;
  assign y16170 = n50934 ;
  assign y16171 = n50943 ;
  assign y16172 = ~n50945 ;
  assign y16173 = ~n50948 ;
  assign y16174 = ~n50950 ;
  assign y16175 = ~n50953 ;
  assign y16176 = ~n50954 ;
  assign y16177 = ~n50956 ;
  assign y16178 = n50958 ;
  assign y16179 = ~n50960 ;
  assign y16180 = ~n50961 ;
  assign y16181 = ~n50962 ;
  assign y16182 = n50963 ;
  assign y16183 = ~n50970 ;
  assign y16184 = n50972 ;
  assign y16185 = ~1'b0 ;
  assign y16186 = ~n50977 ;
  assign y16187 = ~1'b0 ;
  assign y16188 = ~n50982 ;
  assign y16189 = ~n50985 ;
  assign y16190 = n50987 ;
  assign y16191 = n50990 ;
  assign y16192 = ~n50994 ;
  assign y16193 = n50996 ;
  assign y16194 = n50999 ;
  assign y16195 = ~1'b0 ;
  assign y16196 = ~n51002 ;
  assign y16197 = ~n51004 ;
  assign y16198 = n51008 ;
  assign y16199 = ~n51010 ;
  assign y16200 = n51012 ;
  assign y16201 = ~n51013 ;
  assign y16202 = ~n51016 ;
  assign y16203 = n51018 ;
  assign y16204 = n51020 ;
  assign y16205 = n51025 ;
  assign y16206 = ~1'b0 ;
  assign y16207 = n51029 ;
  assign y16208 = n51031 ;
  assign y16209 = n51032 ;
  assign y16210 = ~n51033 ;
  assign y16211 = ~n51037 ;
  assign y16212 = n51038 ;
  assign y16213 = ~1'b0 ;
  assign y16214 = ~1'b0 ;
  assign y16215 = ~n51047 ;
  assign y16216 = ~1'b0 ;
  assign y16217 = ~n51048 ;
  assign y16218 = n51050 ;
  assign y16219 = ~n51055 ;
  assign y16220 = ~n51056 ;
  assign y16221 = ~n51057 ;
  assign y16222 = ~n51059 ;
  assign y16223 = ~1'b0 ;
  assign y16224 = ~n51061 ;
  assign y16225 = ~n51062 ;
  assign y16226 = n51063 ;
  assign y16227 = ~n51068 ;
  assign y16228 = n6405 ;
  assign y16229 = n51071 ;
  assign y16230 = ~n51075 ;
  assign y16231 = n51079 ;
  assign y16232 = ~n51082 ;
  assign y16233 = n51084 ;
  assign y16234 = ~n51085 ;
  assign y16235 = n51087 ;
  assign y16236 = ~n51088 ;
  assign y16237 = n51092 ;
  assign y16238 = n7298 ;
  assign y16239 = n51095 ;
  assign y16240 = ~n51097 ;
  assign y16241 = n51098 ;
  assign y16242 = n51100 ;
  assign y16243 = n51104 ;
  assign y16244 = n51114 ;
  assign y16245 = n51115 ;
  assign y16246 = n51116 ;
  assign y16247 = ~n51117 ;
  assign y16248 = n51121 ;
  assign y16249 = ~n51122 ;
  assign y16250 = n51123 ;
  assign y16251 = ~n51124 ;
  assign y16252 = ~n51125 ;
  assign y16253 = ~n51131 ;
  assign y16254 = ~n51134 ;
  assign y16255 = ~n51148 ;
  assign y16256 = ~n51149 ;
  assign y16257 = n51150 ;
  assign y16258 = n51156 ;
  assign y16259 = ~n51161 ;
  assign y16260 = ~n51162 ;
  assign y16261 = n51165 ;
  assign y16262 = n51166 ;
  assign y16263 = n51167 ;
  assign y16264 = n51169 ;
  assign y16265 = ~n51170 ;
  assign y16266 = n51171 ;
  assign y16267 = ~n51173 ;
  assign y16268 = n51175 ;
  assign y16269 = n51177 ;
  assign y16270 = ~n51178 ;
  assign y16271 = ~n51181 ;
  assign y16272 = n51182 ;
  assign y16273 = ~n51184 ;
  assign y16274 = ~n51186 ;
  assign y16275 = ~1'b0 ;
  assign y16276 = ~1'b0 ;
  assign y16277 = ~n51188 ;
  assign y16278 = n51189 ;
  assign y16279 = n51190 ;
  assign y16280 = n51191 ;
  assign y16281 = n51194 ;
  assign y16282 = ~n51195 ;
  assign y16283 = ~n51199 ;
  assign y16284 = ~n51202 ;
  assign y16285 = ~n51204 ;
  assign y16286 = ~n51207 ;
  assign y16287 = ~n51208 ;
  assign y16288 = ~1'b0 ;
  assign y16289 = ~n51210 ;
  assign y16290 = ~n51212 ;
  assign y16291 = ~n51216 ;
  assign y16292 = n51219 ;
  assign y16293 = ~n51225 ;
  assign y16294 = n51226 ;
  assign y16295 = n51228 ;
  assign y16296 = n51230 ;
  assign y16297 = n51232 ;
  assign y16298 = ~1'b0 ;
  assign y16299 = ~1'b0 ;
  assign y16300 = ~n51234 ;
  assign y16301 = ~n51235 ;
  assign y16302 = ~n51236 ;
  assign y16303 = ~n51237 ;
  assign y16304 = n51238 ;
  assign y16305 = n51239 ;
  assign y16306 = ~n51242 ;
  assign y16307 = n51244 ;
  assign y16308 = n51246 ;
  assign y16309 = ~n51249 ;
  assign y16310 = ~n51259 ;
  assign y16311 = ~n51261 ;
  assign y16312 = n51262 ;
  assign y16313 = ~n51266 ;
  assign y16314 = n51268 ;
  assign y16315 = ~n51269 ;
  assign y16316 = ~n51271 ;
  assign y16317 = ~1'b0 ;
  assign y16318 = ~1'b0 ;
  assign y16319 = ~n51273 ;
  assign y16320 = n51275 ;
  assign y16321 = ~n51277 ;
  assign y16322 = ~n51278 ;
  assign y16323 = n51283 ;
  assign y16324 = ~n51285 ;
  assign y16325 = ~n51287 ;
  assign y16326 = ~n51290 ;
  assign y16327 = n51292 ;
  assign y16328 = n51294 ;
  assign y16329 = n51297 ;
  assign y16330 = ~n51299 ;
  assign y16331 = ~1'b0 ;
  assign y16332 = ~n51304 ;
  assign y16333 = ~n51307 ;
  assign y16334 = ~n51310 ;
  assign y16335 = n3678 ;
  assign y16336 = n51313 ;
  assign y16337 = ~n11912 ;
  assign y16338 = n51315 ;
  assign y16339 = ~1'b0 ;
  assign y16340 = ~n51319 ;
  assign y16341 = ~n51320 ;
  assign y16342 = ~n51321 ;
  assign y16343 = ~n51324 ;
  assign y16344 = n51327 ;
  assign y16345 = n51330 ;
  assign y16346 = n51335 ;
  assign y16347 = n51337 ;
  assign y16348 = ~1'b0 ;
  assign y16349 = ~n51340 ;
  assign y16350 = ~n51347 ;
  assign y16351 = n51348 ;
  assign y16352 = n51351 ;
  assign y16353 = ~n51352 ;
  assign y16354 = n51353 ;
  assign y16355 = n51357 ;
  assign y16356 = ~n51361 ;
  assign y16357 = ~n12661 ;
  assign y16358 = ~1'b0 ;
  assign y16359 = n51363 ;
  assign y16360 = ~n51364 ;
  assign y16361 = ~n51367 ;
  assign y16362 = ~n51370 ;
  assign y16363 = n51372 ;
  assign y16364 = ~n51376 ;
  assign y16365 = ~n51381 ;
  assign y16366 = n51382 ;
  assign y16367 = n51383 ;
  assign y16368 = ~n51384 ;
  assign y16369 = n51385 ;
  assign y16370 = n51386 ;
  assign y16371 = ~n51389 ;
  assign y16372 = ~n51391 ;
  assign y16373 = n51392 ;
  assign y16374 = n51394 ;
  assign y16375 = ~n51395 ;
  assign y16376 = n51397 ;
  assign y16377 = n51400 ;
  assign y16378 = ~n51407 ;
  assign y16379 = ~n51411 ;
  assign y16380 = ~n51414 ;
  assign y16381 = ~n51418 ;
  assign y16382 = ~n51420 ;
  assign y16383 = n51423 ;
  assign y16384 = n51426 ;
  assign y16385 = ~n51428 ;
  assign y16386 = ~n51432 ;
  assign y16387 = ~n51433 ;
  assign y16388 = n51436 ;
  assign y16389 = ~n51438 ;
  assign y16390 = ~n51441 ;
  assign y16391 = n51442 ;
  assign y16392 = ~n51443 ;
  assign y16393 = ~n51446 ;
  assign y16394 = n51451 ;
  assign y16395 = ~n51454 ;
  assign y16396 = ~n51457 ;
  assign y16397 = n51459 ;
  assign y16398 = ~1'b0 ;
  assign y16399 = n51462 ;
  assign y16400 = ~n51463 ;
  assign y16401 = n51466 ;
  assign y16402 = ~n51467 ;
  assign y16403 = ~n51468 ;
  assign y16404 = ~n51473 ;
  assign y16405 = ~n51474 ;
  assign y16406 = ~n51476 ;
  assign y16407 = n51479 ;
  assign y16408 = n51485 ;
  assign y16409 = ~n51490 ;
  assign y16410 = ~n51491 ;
  assign y16411 = n51494 ;
  assign y16412 = n51495 ;
  assign y16413 = n51497 ;
  assign y16414 = ~n51501 ;
  assign y16415 = n51502 ;
  assign y16416 = ~n51504 ;
  assign y16417 = ~n51506 ;
  assign y16418 = n51508 ;
  assign y16419 = n51512 ;
  assign y16420 = ~n51513 ;
  assign y16421 = n51515 ;
  assign y16422 = ~n51518 ;
  assign y16423 = ~n51519 ;
  assign y16424 = ~n51520 ;
  assign y16425 = ~n51521 ;
  assign y16426 = ~n48383 ;
  assign y16427 = ~1'b0 ;
  assign y16428 = n51523 ;
  assign y16429 = n51525 ;
  assign y16430 = n51528 ;
  assign y16431 = ~n51530 ;
  assign y16432 = ~n51533 ;
  assign y16433 = n51536 ;
  assign y16434 = n51537 ;
  assign y16435 = ~n51538 ;
  assign y16436 = n51540 ;
  assign y16437 = n51541 ;
  assign y16438 = n51544 ;
  assign y16439 = ~n51548 ;
  assign y16440 = n51550 ;
  assign y16441 = n51555 ;
  assign y16442 = ~n51559 ;
  assign y16443 = ~n51560 ;
  assign y16444 = n51562 ;
  assign y16445 = n51563 ;
  assign y16446 = n51564 ;
  assign y16447 = n51566 ;
  assign y16448 = ~n51570 ;
  assign y16449 = ~n51571 ;
  assign y16450 = n51576 ;
  assign y16451 = n51577 ;
  assign y16452 = n51578 ;
  assign y16453 = ~n51579 ;
  assign y16454 = n51580 ;
  assign y16455 = n51581 ;
  assign y16456 = ~n51584 ;
  assign y16457 = n51586 ;
  assign y16458 = n51593 ;
  assign y16459 = ~n51595 ;
  assign y16460 = ~n51598 ;
  assign y16461 = ~1'b0 ;
  assign y16462 = ~n51599 ;
  assign y16463 = ~n51600 ;
  assign y16464 = n51605 ;
  assign y16465 = ~n51606 ;
  assign y16466 = n51613 ;
  assign y16467 = ~n51621 ;
  assign y16468 = ~1'b0 ;
  assign y16469 = ~1'b0 ;
  assign y16470 = n51622 ;
  assign y16471 = ~n51625 ;
  assign y16472 = ~n51626 ;
  assign y16473 = n51632 ;
  assign y16474 = ~n51633 ;
  assign y16475 = ~n51638 ;
  assign y16476 = ~n51639 ;
  assign y16477 = n51640 ;
  assign y16478 = n5691 ;
  assign y16479 = ~n51643 ;
  assign y16480 = ~n51644 ;
  assign y16481 = ~1'b0 ;
  assign y16482 = ~n51645 ;
  assign y16483 = ~n51647 ;
  assign y16484 = n51648 ;
  assign y16485 = n51650 ;
  assign y16486 = ~n51652 ;
  assign y16487 = ~n51656 ;
  assign y16488 = ~n51659 ;
  assign y16489 = n51666 ;
  assign y16490 = n51668 ;
  assign y16491 = ~1'b0 ;
  assign y16492 = ~n51672 ;
  assign y16493 = n51674 ;
  assign y16494 = ~n51675 ;
  assign y16495 = ~n51676 ;
  assign y16496 = n51677 ;
  assign y16497 = n51680 ;
  assign y16498 = ~n51683 ;
  assign y16499 = ~n51688 ;
  assign y16500 = ~1'b0 ;
  assign y16501 = 1'b0 ;
  assign y16502 = ~1'b0 ;
  assign y16503 = n51689 ;
  assign y16504 = ~n51691 ;
  assign y16505 = ~n51694 ;
  assign y16506 = ~n51699 ;
  assign y16507 = ~n51703 ;
  assign y16508 = ~1'b0 ;
  assign y16509 = ~1'b0 ;
  assign y16510 = n24415 ;
  assign y16511 = ~n51704 ;
  assign y16512 = n51707 ;
  assign y16513 = n51709 ;
  assign y16514 = ~n51711 ;
  assign y16515 = n51714 ;
  assign y16516 = ~n51716 ;
  assign y16517 = ~n51718 ;
  assign y16518 = ~n51721 ;
  assign y16519 = ~n51723 ;
  assign y16520 = n51725 ;
  assign y16521 = n51726 ;
  assign y16522 = n51727 ;
  assign y16523 = ~n51730 ;
  assign y16524 = ~n51732 ;
  assign y16525 = n51733 ;
  assign y16526 = ~n51734 ;
  assign y16527 = n51740 ;
  assign y16528 = ~n51743 ;
  assign y16529 = ~1'b0 ;
  assign y16530 = ~n51746 ;
  assign y16531 = ~n51747 ;
  assign y16532 = ~n51748 ;
  assign y16533 = n51749 ;
  assign y16534 = n51750 ;
  assign y16535 = n51753 ;
  assign y16536 = ~n51757 ;
  assign y16537 = ~n51758 ;
  assign y16538 = ~n51765 ;
  assign y16539 = ~1'b0 ;
  assign y16540 = ~1'b0 ;
  assign y16541 = ~1'b0 ;
  assign y16542 = ~n51766 ;
  assign y16543 = ~1'b0 ;
  assign y16544 = ~n51767 ;
  assign y16545 = n51768 ;
  assign y16546 = ~n51770 ;
  assign y16547 = n51771 ;
  assign y16548 = ~n51772 ;
  assign y16549 = ~n51773 ;
  assign y16550 = ~n51776 ;
  assign y16551 = ~n51777 ;
  assign y16552 = n51780 ;
  assign y16553 = n51781 ;
  assign y16554 = ~n51788 ;
  assign y16555 = ~n51789 ;
  assign y16556 = ~n51792 ;
  assign y16557 = n51796 ;
  assign y16558 = n51803 ;
  assign y16559 = ~1'b0 ;
  assign y16560 = n51806 ;
  assign y16561 = n51807 ;
  assign y16562 = n51808 ;
  assign y16563 = n51812 ;
  assign y16564 = n51813 ;
  assign y16565 = n51814 ;
  assign y16566 = ~n51817 ;
  assign y16567 = ~n51822 ;
  assign y16568 = ~1'b0 ;
  assign y16569 = n51824 ;
  assign y16570 = ~1'b0 ;
  assign y16571 = ~n51831 ;
  assign y16572 = n51832 ;
  assign y16573 = n51833 ;
  assign y16574 = ~n51835 ;
  assign y16575 = ~n51836 ;
  assign y16576 = n51838 ;
  assign y16577 = n51840 ;
  assign y16578 = ~n51842 ;
  assign y16579 = ~1'b0 ;
  assign y16580 = n51844 ;
  assign y16581 = n51846 ;
  assign y16582 = ~n51848 ;
  assign y16583 = n51850 ;
  assign y16584 = n51851 ;
  assign y16585 = ~n51852 ;
  assign y16586 = n51853 ;
  assign y16587 = ~n51854 ;
  assign y16588 = n51860 ;
  assign y16589 = ~n51861 ;
  assign y16590 = ~1'b0 ;
  assign y16591 = n51864 ;
  assign y16592 = ~n51865 ;
  assign y16593 = n51869 ;
  assign y16594 = ~n51874 ;
  assign y16595 = ~n51881 ;
  assign y16596 = ~n51882 ;
  assign y16597 = ~n51884 ;
  assign y16598 = ~1'b0 ;
  assign y16599 = ~1'b0 ;
  assign y16600 = ~n51888 ;
  assign y16601 = ~n51894 ;
  assign y16602 = n51896 ;
  assign y16603 = ~1'b0 ;
  assign y16604 = n51900 ;
  assign y16605 = n51903 ;
  assign y16606 = ~n51904 ;
  assign y16607 = n51908 ;
  assign y16608 = ~n51912 ;
  assign y16609 = ~1'b0 ;
  assign y16610 = n51918 ;
  assign y16611 = n51921 ;
  assign y16612 = n51927 ;
  assign y16613 = ~n51932 ;
  assign y16614 = n51937 ;
  assign y16615 = n51938 ;
  assign y16616 = n51939 ;
  assign y16617 = n51944 ;
  assign y16618 = ~1'b0 ;
  assign y16619 = ~n51946 ;
  assign y16620 = ~n51948 ;
  assign y16621 = ~1'b0 ;
  assign y16622 = n51950 ;
  assign y16623 = n51952 ;
  assign y16624 = ~n51953 ;
  assign y16625 = ~n51956 ;
  assign y16626 = ~n51958 ;
  assign y16627 = ~n51966 ;
  assign y16628 = n51969 ;
  assign y16629 = ~1'b0 ;
  assign y16630 = ~n51971 ;
  assign y16631 = n51975 ;
  assign y16632 = ~1'b0 ;
  assign y16633 = ~n51976 ;
  assign y16634 = ~n51979 ;
  assign y16635 = n51980 ;
  assign y16636 = n51982 ;
  assign y16637 = ~n51983 ;
  assign y16638 = n51985 ;
  assign y16639 = ~n51987 ;
  assign y16640 = ~1'b0 ;
  assign y16641 = ~1'b0 ;
  assign y16642 = ~1'b0 ;
  assign y16643 = ~n51988 ;
  assign y16644 = n51989 ;
  assign y16645 = ~n51991 ;
  assign y16646 = n44812 ;
  assign y16647 = n51993 ;
  assign y16648 = n51996 ;
  assign y16649 = ~1'b0 ;
  assign y16650 = n52001 ;
  assign y16651 = n52002 ;
  assign y16652 = n52003 ;
  assign y16653 = n52005 ;
  assign y16654 = ~n52006 ;
  assign y16655 = n52008 ;
  assign y16656 = n52009 ;
  assign y16657 = ~n52010 ;
  assign y16658 = n52015 ;
  assign y16659 = ~1'b0 ;
  assign y16660 = ~1'b0 ;
  assign y16661 = ~n52016 ;
  assign y16662 = ~1'b0 ;
  assign y16663 = n52017 ;
  assign y16664 = n52020 ;
  assign y16665 = ~n52021 ;
  assign y16666 = ~n52023 ;
  assign y16667 = n52028 ;
  assign y16668 = n52032 ;
  assign y16669 = ~n52033 ;
  assign y16670 = n52040 ;
  assign y16671 = ~n52042 ;
  assign y16672 = ~1'b0 ;
  assign y16673 = n52043 ;
  assign y16674 = ~n52046 ;
  assign y16675 = n52047 ;
  assign y16676 = ~n52050 ;
  assign y16677 = n52051 ;
  assign y16678 = n52052 ;
  assign y16679 = n52053 ;
  assign y16680 = n52055 ;
  assign y16681 = n52058 ;
  assign y16682 = ~n52059 ;
  assign y16683 = ~n52061 ;
  assign y16684 = n52062 ;
  assign y16685 = ~n52064 ;
  assign y16686 = ~1'b0 ;
  assign y16687 = n52067 ;
  assign y16688 = n2989 ;
  assign y16689 = n52068 ;
  assign y16690 = n52070 ;
  assign y16691 = ~n52072 ;
  assign y16692 = ~n52074 ;
  assign y16693 = n25942 ;
  assign y16694 = ~n11893 ;
  assign y16695 = ~n52075 ;
  assign y16696 = n52077 ;
  assign y16697 = n52078 ;
  assign y16698 = ~n52080 ;
  assign y16699 = ~n52083 ;
  assign y16700 = n52086 ;
  assign y16701 = ~n52088 ;
  assign y16702 = ~n52095 ;
  assign y16703 = ~n52099 ;
  assign y16704 = ~1'b0 ;
  assign y16705 = ~n36870 ;
  assign y16706 = ~n52105 ;
  assign y16707 = n52106 ;
  assign y16708 = ~n52107 ;
  assign y16709 = n52111 ;
  assign y16710 = n52113 ;
  assign y16711 = ~1'b0 ;
  assign y16712 = ~n52116 ;
  assign y16713 = ~1'b0 ;
  assign y16714 = ~n52118 ;
  assign y16715 = n52119 ;
  assign y16716 = n52120 ;
  assign y16717 = ~n52121 ;
  assign y16718 = n52125 ;
  assign y16719 = n52126 ;
  assign y16720 = ~n52129 ;
  assign y16721 = n52133 ;
  assign y16722 = n52136 ;
  assign y16723 = n52138 ;
  assign y16724 = n52142 ;
  assign y16725 = n52146 ;
  assign y16726 = ~n52149 ;
  assign y16727 = n52151 ;
  assign y16728 = n52156 ;
  assign y16729 = ~n52157 ;
  assign y16730 = ~n52160 ;
  assign y16731 = n52163 ;
  assign y16732 = n52172 ;
  assign y16733 = ~n52173 ;
  assign y16734 = ~n52174 ;
  assign y16735 = n52176 ;
  assign y16736 = n22484 ;
  assign y16737 = ~n52177 ;
  assign y16738 = ~n52179 ;
  assign y16739 = ~n52183 ;
  assign y16740 = n52184 ;
  assign y16741 = ~n52191 ;
  assign y16742 = ~n52194 ;
  assign y16743 = n52195 ;
  assign y16744 = n52201 ;
  assign y16745 = ~1'b0 ;
  assign y16746 = ~n52205 ;
  assign y16747 = n52206 ;
  assign y16748 = n52207 ;
  assign y16749 = ~n52211 ;
  assign y16750 = n52214 ;
  assign y16751 = n52216 ;
  assign y16752 = n52220 ;
  assign y16753 = n52221 ;
  assign y16754 = ~1'b0 ;
  assign y16755 = n52223 ;
  assign y16756 = n52226 ;
  assign y16757 = ~n52230 ;
  assign y16758 = ~n52231 ;
  assign y16759 = ~n52236 ;
  assign y16760 = ~n52237 ;
  assign y16761 = n52248 ;
  assign y16762 = n52249 ;
  assign y16763 = n52251 ;
  assign y16764 = n52252 ;
  assign y16765 = ~n52253 ;
  assign y16766 = n52257 ;
  assign y16767 = ~n52259 ;
  assign y16768 = ~1'b0 ;
  assign y16769 = ~n52260 ;
  assign y16770 = ~n52261 ;
  assign y16771 = ~n52263 ;
  assign y16772 = ~n52267 ;
  assign y16773 = ~n52272 ;
  assign y16774 = ~n52274 ;
  assign y16775 = ~n52276 ;
  assign y16776 = ~1'b0 ;
  assign y16777 = n52279 ;
  assign y16778 = ~1'b0 ;
  assign y16779 = ~n52281 ;
  assign y16780 = ~n52283 ;
  assign y16781 = ~n52290 ;
  assign y16782 = ~n52292 ;
  assign y16783 = n52294 ;
  assign y16784 = n52295 ;
  assign y16785 = ~n52296 ;
  assign y16786 = ~n52298 ;
  assign y16787 = ~n52307 ;
  assign y16788 = n52309 ;
  assign y16789 = ~n52311 ;
  assign y16790 = n52313 ;
  assign y16791 = ~n52316 ;
  assign y16792 = n52321 ;
  assign y16793 = n52322 ;
  assign y16794 = n52326 ;
  assign y16795 = ~n52328 ;
  assign y16796 = n52329 ;
  assign y16797 = n52331 ;
  assign y16798 = n52333 ;
  assign y16799 = ~n52335 ;
  assign y16800 = n52337 ;
  assign y16801 = n52341 ;
  assign y16802 = n52343 ;
  assign y16803 = n52344 ;
  assign y16804 = ~n52347 ;
  assign y16805 = ~n52348 ;
  assign y16806 = ~n52350 ;
  assign y16807 = ~1'b0 ;
  assign y16808 = n52351 ;
  assign y16809 = ~1'b0 ;
  assign y16810 = ~n52353 ;
  assign y16811 = 1'b0 ;
  assign y16812 = ~n52354 ;
  assign y16813 = n52360 ;
  assign y16814 = n52363 ;
  assign y16815 = n52365 ;
  assign y16816 = ~n52368 ;
  assign y16817 = n52375 ;
  assign y16818 = n52377 ;
  assign y16819 = ~1'b0 ;
  assign y16820 = n52381 ;
  assign y16821 = n52384 ;
  assign y16822 = n52385 ;
  assign y16823 = ~n52390 ;
  assign y16824 = n52396 ;
  assign y16825 = ~n52397 ;
  assign y16826 = ~n52400 ;
  assign y16827 = n52404 ;
  assign y16828 = ~n52406 ;
  assign y16829 = ~n52407 ;
  assign y16830 = ~1'b0 ;
  assign y16831 = ~n52409 ;
  assign y16832 = n52411 ;
  assign y16833 = n52415 ;
  assign y16834 = ~n52416 ;
  assign y16835 = n52419 ;
  assign y16836 = ~n52420 ;
  assign y16837 = ~n52423 ;
  assign y16838 = ~n52425 ;
  assign y16839 = ~1'b0 ;
  assign y16840 = n52427 ;
  assign y16841 = ~n52429 ;
  assign y16842 = ~n52435 ;
  assign y16843 = n52438 ;
  assign y16844 = ~n52440 ;
  assign y16845 = ~n52441 ;
  assign y16846 = ~n52446 ;
  assign y16847 = n52447 ;
  assign y16848 = ~1'b0 ;
  assign y16849 = ~1'b0 ;
  assign y16850 = ~n52450 ;
  assign y16851 = n52453 ;
  assign y16852 = n52457 ;
  assign y16853 = n52459 ;
  assign y16854 = n52460 ;
  assign y16855 = ~n52461 ;
  assign y16856 = ~n52462 ;
  assign y16857 = ~n52465 ;
  assign y16858 = n52467 ;
  assign y16859 = n52469 ;
  assign y16860 = ~1'b0 ;
  assign y16861 = n52475 ;
  assign y16862 = n52477 ;
  assign y16863 = ~n52478 ;
  assign y16864 = n52479 ;
  assign y16865 = n52481 ;
  assign y16866 = n52483 ;
  assign y16867 = n52486 ;
  assign y16868 = n52490 ;
  assign y16869 = ~n52493 ;
  assign y16870 = ~n52495 ;
  assign y16871 = ~n52496 ;
  assign y16872 = ~n20162 ;
  assign y16873 = n52498 ;
  assign y16874 = n52500 ;
  assign y16875 = ~n52503 ;
  assign y16876 = ~n52504 ;
  assign y16877 = ~1'b0 ;
  assign y16878 = ~1'b0 ;
  assign y16879 = ~n52506 ;
  assign y16880 = ~n52507 ;
  assign y16881 = ~n52508 ;
  assign y16882 = ~n52513 ;
  assign y16883 = ~n52515 ;
  assign y16884 = n52518 ;
  assign y16885 = ~n52521 ;
  assign y16886 = n52524 ;
  assign y16887 = ~n52525 ;
  assign y16888 = ~1'b0 ;
  assign y16889 = n52526 ;
  assign y16890 = ~1'b0 ;
  assign y16891 = n52530 ;
  assign y16892 = ~n52532 ;
  assign y16893 = ~n52537 ;
  assign y16894 = n52539 ;
  assign y16895 = n52541 ;
  assign y16896 = ~n52542 ;
  assign y16897 = n52547 ;
  assign y16898 = n52549 ;
  assign y16899 = n52552 ;
  assign y16900 = ~n52554 ;
  assign y16901 = ~n52557 ;
  assign y16902 = ~n52561 ;
  assign y16903 = ~n52564 ;
  assign y16904 = ~n52565 ;
  assign y16905 = ~n52573 ;
  assign y16906 = n52576 ;
  assign y16907 = n52578 ;
  assign y16908 = ~n52581 ;
  assign y16909 = ~n52585 ;
  assign y16910 = ~n52587 ;
  assign y16911 = ~1'b0 ;
  assign y16912 = ~n52589 ;
  assign y16913 = n52591 ;
  assign y16914 = ~n52597 ;
  assign y16915 = ~n52601 ;
  assign y16916 = n52603 ;
  assign y16917 = n52604 ;
  assign y16918 = ~n52606 ;
  assign y16919 = n52607 ;
  assign y16920 = ~1'b0 ;
  assign y16921 = n52608 ;
  assign y16922 = ~n52612 ;
  assign y16923 = ~n52613 ;
  assign y16924 = n52615 ;
  assign y16925 = n52618 ;
  assign y16926 = n52621 ;
  assign y16927 = n52624 ;
  assign y16928 = n52625 ;
  assign y16929 = ~n52628 ;
  assign y16930 = ~n52630 ;
  assign y16931 = ~n52633 ;
  assign y16932 = ~n14875 ;
  assign y16933 = ~n52635 ;
  assign y16934 = ~n52638 ;
  assign y16935 = n52639 ;
  assign y16936 = n52642 ;
  assign y16937 = ~n52645 ;
  assign y16938 = ~n52647 ;
  assign y16939 = ~n52649 ;
  assign y16940 = ~1'b0 ;
  assign y16941 = ~1'b0 ;
  assign y16942 = ~n52651 ;
  assign y16943 = n52652 ;
  assign y16944 = ~n52653 ;
  assign y16945 = ~n52654 ;
  assign y16946 = ~n50839 ;
  assign y16947 = n27684 ;
  assign y16948 = n52658 ;
  assign y16949 = ~1'b0 ;
  assign y16950 = n52662 ;
  assign y16951 = n52664 ;
  assign y16952 = n52666 ;
  assign y16953 = ~n52667 ;
  assign y16954 = ~n52670 ;
  assign y16955 = n52673 ;
  assign y16956 = ~n52675 ;
  assign y16957 = n52678 ;
  assign y16958 = ~n52682 ;
  assign y16959 = ~n52685 ;
  assign y16960 = ~1'b0 ;
  assign y16961 = ~n52688 ;
  assign y16962 = ~n52691 ;
  assign y16963 = n52693 ;
  assign y16964 = ~n52696 ;
  assign y16965 = ~n52698 ;
  assign y16966 = n52699 ;
  assign y16967 = n52701 ;
  assign y16968 = ~n52702 ;
  assign y16969 = n52704 ;
  assign y16970 = ~1'b0 ;
  assign y16971 = n52705 ;
  assign y16972 = n52715 ;
  assign y16973 = n52717 ;
  assign y16974 = ~n52718 ;
  assign y16975 = n52719 ;
  assign y16976 = ~n52720 ;
  assign y16977 = ~n52725 ;
  assign y16978 = ~n13245 ;
  assign y16979 = n52726 ;
  assign y16980 = ~n52728 ;
  assign y16981 = ~n52730 ;
  assign y16982 = n52732 ;
  assign y16983 = ~n52734 ;
  assign y16984 = ~n52737 ;
  assign y16985 = n52741 ;
  assign y16986 = ~n52743 ;
  assign y16987 = n52744 ;
  assign y16988 = ~n52746 ;
  assign y16989 = ~n52748 ;
  assign y16990 = n52752 ;
  assign y16991 = n52754 ;
  assign y16992 = ~n52759 ;
  assign y16993 = ~n52761 ;
  assign y16994 = ~1'b0 ;
  assign y16995 = n52763 ;
  assign y16996 = n52764 ;
  assign y16997 = n52766 ;
  assign y16998 = ~n52767 ;
  assign y16999 = ~1'b0 ;
  assign y17000 = ~n52773 ;
  assign y17001 = ~n52777 ;
  assign y17002 = ~n52778 ;
  assign y17003 = ~n52781 ;
  assign y17004 = n52782 ;
  assign y17005 = ~n52783 ;
  assign y17006 = ~n52788 ;
  assign y17007 = ~n52789 ;
  assign y17008 = ~n52790 ;
  assign y17009 = n52796 ;
  assign y17010 = ~n52800 ;
  assign y17011 = ~n52801 ;
  assign y17012 = ~n52806 ;
  assign y17013 = ~n52813 ;
  assign y17014 = n52818 ;
  assign y17015 = ~n52821 ;
  assign y17016 = ~1'b0 ;
  assign y17017 = n52825 ;
  assign y17018 = ~n52829 ;
  assign y17019 = n52830 ;
  assign y17020 = ~n52835 ;
  assign y17021 = ~n52840 ;
  assign y17022 = n52844 ;
  assign y17023 = n52848 ;
  assign y17024 = n52850 ;
  assign y17025 = n52851 ;
  assign y17026 = n52856 ;
  assign y17027 = n52857 ;
  assign y17028 = ~n52859 ;
  assign y17029 = ~n52860 ;
  assign y17030 = ~n52863 ;
  assign y17031 = ~n52865 ;
  assign y17032 = ~n52870 ;
  assign y17033 = ~n52877 ;
  assign y17034 = ~n52879 ;
  assign y17035 = n52881 ;
  assign y17036 = n52883 ;
  assign y17037 = ~n52885 ;
  assign y17038 = ~n52886 ;
  assign y17039 = n52889 ;
  assign y17040 = n21622 ;
  assign y17041 = ~n52890 ;
  assign y17042 = ~n52891 ;
  assign y17043 = n52895 ;
  assign y17044 = ~n52897 ;
  assign y17045 = ~n52898 ;
  assign y17046 = ~1'b0 ;
  assign y17047 = ~1'b0 ;
  assign y17048 = ~n52901 ;
  assign y17049 = n52903 ;
  assign y17050 = ~n52909 ;
  assign y17051 = ~n52910 ;
  assign y17052 = ~n52913 ;
  assign y17053 = n52914 ;
  assign y17054 = ~n52915 ;
  assign y17055 = ~1'b0 ;
  assign y17056 = n52918 ;
  assign y17057 = ~n52919 ;
  assign y17058 = ~1'b0 ;
  assign y17059 = n52920 ;
  assign y17060 = n52925 ;
  assign y17061 = n52926 ;
  assign y17062 = ~n52927 ;
  assign y17063 = ~n52928 ;
  assign y17064 = n52931 ;
  assign y17065 = ~n52934 ;
  assign y17066 = n52936 ;
  assign y17067 = n52942 ;
  assign y17068 = n52946 ;
  assign y17069 = n52950 ;
  assign y17070 = ~n52952 ;
  assign y17071 = ~n52955 ;
  assign y17072 = n52958 ;
  assign y17073 = ~n52959 ;
  assign y17074 = ~n52961 ;
  assign y17075 = ~1'b0 ;
  assign y17076 = ~n52963 ;
  assign y17077 = n52968 ;
  assign y17078 = n52969 ;
  assign y17079 = n52970 ;
  assign y17080 = n52971 ;
  assign y17081 = n52973 ;
  assign y17082 = ~n52975 ;
  assign y17083 = ~n52976 ;
  assign y17084 = n52979 ;
  assign y17085 = ~n52980 ;
  assign y17086 = ~1'b0 ;
  assign y17087 = n52982 ;
  assign y17088 = n52983 ;
  assign y17089 = ~n52984 ;
  assign y17090 = ~n52985 ;
  assign y17091 = ~n52986 ;
  assign y17092 = ~n52990 ;
  assign y17093 = ~n52991 ;
  assign y17094 = ~n52992 ;
  assign y17095 = ~n52996 ;
  assign y17096 = n52999 ;
  assign y17097 = ~1'b0 ;
  assign y17098 = ~n53001 ;
  assign y17099 = n53002 ;
  assign y17100 = ~n53004 ;
  assign y17101 = ~n53005 ;
  assign y17102 = ~n53007 ;
  assign y17103 = ~n53013 ;
  assign y17104 = ~n53016 ;
  assign y17105 = ~1'b0 ;
  assign y17106 = ~1'b0 ;
  assign y17107 = n53018 ;
  assign y17108 = ~1'b0 ;
  assign y17109 = ~n53024 ;
  assign y17110 = n53026 ;
  assign y17111 = ~n53031 ;
  assign y17112 = n53032 ;
  assign y17113 = ~n53033 ;
  assign y17114 = ~n53036 ;
  assign y17115 = ~n53038 ;
  assign y17116 = ~n49871 ;
  assign y17117 = ~1'b0 ;
  assign y17118 = ~n53040 ;
  assign y17119 = ~n53042 ;
  assign y17120 = ~n53047 ;
  assign y17121 = n53053 ;
  assign y17122 = ~n53054 ;
  assign y17123 = n53058 ;
  assign y17124 = n53062 ;
  assign y17125 = ~n53063 ;
  assign y17126 = ~n53066 ;
  assign y17127 = ~1'b0 ;
  assign y17128 = n53068 ;
  assign y17129 = ~n53070 ;
  assign y17130 = n53071 ;
  assign y17131 = n35651 ;
  assign y17132 = ~n53072 ;
  assign y17133 = n53074 ;
  assign y17134 = ~n53076 ;
  assign y17135 = n53077 ;
  assign y17136 = n53079 ;
  assign y17137 = ~n53081 ;
  assign y17138 = ~n53083 ;
  assign y17139 = n53087 ;
  assign y17140 = n53089 ;
  assign y17141 = ~n53090 ;
  assign y17142 = n53092 ;
  assign y17143 = n53095 ;
  assign y17144 = n53099 ;
  assign y17145 = ~n53100 ;
  assign y17146 = n53102 ;
  assign y17147 = n22795 ;
  assign y17148 = ~n53103 ;
  assign y17149 = ~n53106 ;
  assign y17150 = ~1'b0 ;
  assign y17151 = ~n53109 ;
  assign y17152 = ~n53110 ;
  assign y17153 = ~n53113 ;
  assign y17154 = n53117 ;
  assign y17155 = ~n53118 ;
  assign y17156 = ~n53121 ;
  assign y17157 = ~n53125 ;
  assign y17158 = n53126 ;
  assign y17159 = ~1'b0 ;
  assign y17160 = n53128 ;
  assign y17161 = ~1'b0 ;
  assign y17162 = ~n53130 ;
  assign y17163 = n53131 ;
  assign y17164 = ~n53132 ;
  assign y17165 = n53133 ;
  assign y17166 = ~n53134 ;
  assign y17167 = ~n19048 ;
  assign y17168 = ~n53137 ;
  assign y17169 = n53139 ;
  assign y17170 = ~n53144 ;
  assign y17171 = n53147 ;
  assign y17172 = n53149 ;
  assign y17173 = n53151 ;
  assign y17174 = n53152 ;
  assign y17175 = ~n53153 ;
  assign y17176 = n53154 ;
  assign y17177 = n18399 ;
  assign y17178 = n53158 ;
  assign y17179 = ~n53160 ;
  assign y17180 = n53168 ;
  assign y17181 = ~1'b0 ;
  assign y17182 = ~n53171 ;
  assign y17183 = ~1'b0 ;
  assign y17184 = ~n53172 ;
  assign y17185 = ~n53173 ;
  assign y17186 = n53175 ;
  assign y17187 = n53186 ;
  assign y17188 = n53190 ;
  assign y17189 = ~n53193 ;
  assign y17190 = n53199 ;
  assign y17191 = n53200 ;
  assign y17192 = ~1'b0 ;
  assign y17193 = ~n53205 ;
  assign y17194 = ~1'b0 ;
  assign y17195 = n53207 ;
  assign y17196 = n53210 ;
  assign y17197 = ~n53214 ;
  assign y17198 = ~n53215 ;
  assign y17199 = n53218 ;
  assign y17200 = ~n53221 ;
  assign y17201 = ~n53224 ;
  assign y17202 = n53226 ;
  assign y17203 = n53228 ;
  assign y17204 = ~1'b0 ;
  assign y17205 = ~1'b0 ;
  assign y17206 = ~n53233 ;
  assign y17207 = ~n53237 ;
  assign y17208 = ~n53238 ;
  assign y17209 = n53245 ;
  assign y17210 = n53252 ;
  assign y17211 = n53258 ;
  assign y17212 = n53261 ;
  assign y17213 = ~1'b0 ;
  assign y17214 = ~1'b0 ;
  assign y17215 = ~n53263 ;
  assign y17216 = ~1'b0 ;
  assign y17217 = n53264 ;
  assign y17218 = ~n53272 ;
  assign y17219 = n53274 ;
  assign y17220 = ~n53275 ;
  assign y17221 = n53276 ;
  assign y17222 = n53277 ;
  assign y17223 = ~n53278 ;
  assign y17224 = n53281 ;
  assign y17225 = ~1'b0 ;
  assign y17226 = ~n53283 ;
  assign y17227 = ~1'b0 ;
  assign y17228 = n53284 ;
  assign y17229 = ~n53288 ;
  assign y17230 = n53289 ;
  assign y17231 = n53291 ;
  assign y17232 = ~n53294 ;
  assign y17233 = ~n53297 ;
  assign y17234 = n53299 ;
  assign y17235 = ~1'b0 ;
  assign y17236 = ~n53301 ;
  assign y17237 = ~1'b0 ;
  assign y17238 = ~1'b0 ;
  assign y17239 = ~n53306 ;
  assign y17240 = ~n53307 ;
  assign y17241 = n53310 ;
  assign y17242 = n53316 ;
  assign y17243 = n53319 ;
  assign y17244 = ~n53320 ;
  assign y17245 = n53322 ;
  assign y17246 = ~n53324 ;
  assign y17247 = ~1'b0 ;
  assign y17248 = n53326 ;
  assign y17249 = n53331 ;
  assign y17250 = n53333 ;
  assign y17251 = n53335 ;
  assign y17252 = n53336 ;
  assign y17253 = n53338 ;
  assign y17254 = ~n53339 ;
  assign y17255 = ~n53340 ;
  assign y17256 = ~1'b0 ;
  assign y17257 = n53346 ;
  assign y17258 = ~1'b0 ;
  assign y17259 = n53349 ;
  assign y17260 = n53353 ;
  assign y17261 = n53358 ;
  assign y17262 = ~n53359 ;
  assign y17263 = n53362 ;
  assign y17264 = n53363 ;
  assign y17265 = ~n53364 ;
  assign y17266 = n53369 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~n53371 ;
  assign y17269 = n53373 ;
  assign y17270 = ~n53377 ;
  assign y17271 = n53382 ;
  assign y17272 = n53383 ;
  assign y17273 = n53385 ;
  assign y17274 = n53386 ;
  assign y17275 = ~n53387 ;
  assign y17276 = n53391 ;
  assign y17277 = n53393 ;
  assign y17278 = ~1'b0 ;
  assign y17279 = ~n53394 ;
  assign y17280 = ~n53397 ;
  assign y17281 = n53398 ;
  assign y17282 = ~n14222 ;
  assign y17283 = n53399 ;
  assign y17284 = n53401 ;
  assign y17285 = n53402 ;
  assign y17286 = ~n53407 ;
  assign y17287 = ~n53408 ;
  assign y17288 = ~1'b0 ;
  assign y17289 = n53410 ;
  assign y17290 = n53414 ;
  assign y17291 = n53415 ;
  assign y17292 = ~n53416 ;
  assign y17293 = n53418 ;
  assign y17294 = n53419 ;
  assign y17295 = n53421 ;
  assign y17296 = n53433 ;
  assign y17297 = n53434 ;
  assign y17298 = ~n53437 ;
  assign y17299 = n53438 ;
  assign y17300 = n53440 ;
  assign y17301 = n53442 ;
  assign y17302 = ~n53445 ;
  assign y17303 = ~n53448 ;
  assign y17304 = ~n53449 ;
  assign y17305 = n53454 ;
  assign y17306 = ~n53455 ;
  assign y17307 = n53457 ;
  assign y17308 = ~n53458 ;
  assign y17309 = ~n53459 ;
  assign y17310 = n53463 ;
  assign y17311 = ~n53464 ;
  assign y17312 = ~n53466 ;
  assign y17313 = n53468 ;
  assign y17314 = ~n53470 ;
  assign y17315 = ~n53474 ;
  assign y17316 = n53475 ;
  assign y17317 = n43213 ;
  assign y17318 = ~n53476 ;
  assign y17319 = ~n53479 ;
  assign y17320 = n53481 ;
  assign y17321 = ~n53482 ;
  assign y17322 = ~n53490 ;
  assign y17323 = n53495 ;
  assign y17324 = n53499 ;
  assign y17325 = ~n53500 ;
  assign y17326 = ~n53501 ;
  assign y17327 = n53503 ;
  assign y17328 = n53504 ;
  assign y17329 = ~n53506 ;
  assign y17330 = n53507 ;
  assign y17331 = n53508 ;
  assign y17332 = ~1'b0 ;
  assign y17333 = ~n53510 ;
  assign y17334 = ~1'b0 ;
  assign y17335 = ~n53515 ;
  assign y17336 = n53518 ;
  assign y17337 = ~n53520 ;
  assign y17338 = n53521 ;
  assign y17339 = ~n53522 ;
  assign y17340 = ~n53524 ;
  assign y17341 = n53525 ;
  assign y17342 = n53529 ;
  assign y17343 = ~n53534 ;
  assign y17344 = n53539 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = n53542 ;
  assign y17347 = ~n53543 ;
  assign y17348 = n53546 ;
  assign y17349 = n53548 ;
  assign y17350 = ~n53554 ;
  assign y17351 = ~n53555 ;
  assign y17352 = ~n53556 ;
  assign y17353 = ~1'b0 ;
  assign y17354 = ~n53558 ;
  assign y17355 = ~n53560 ;
  assign y17356 = ~n53562 ;
  assign y17357 = n53564 ;
  assign y17358 = n53565 ;
  assign y17359 = ~n53568 ;
  assign y17360 = ~n53571 ;
  assign y17361 = ~n53572 ;
  assign y17362 = n53577 ;
  assign y17363 = ~n53578 ;
  assign y17364 = ~n53579 ;
  assign y17365 = ~n53581 ;
  assign y17366 = ~1'b0 ;
  assign y17367 = n53583 ;
  assign y17368 = n53584 ;
  assign y17369 = n53585 ;
  assign y17370 = ~n53586 ;
  assign y17371 = n53587 ;
  assign y17372 = n53588 ;
  assign y17373 = n53591 ;
  assign y17374 = n53594 ;
  assign y17375 = ~n53596 ;
  assign y17376 = n53598 ;
  assign y17377 = ~1'b0 ;
  assign y17378 = n53601 ;
  assign y17379 = n53602 ;
  assign y17380 = n53603 ;
  assign y17381 = ~n53608 ;
  assign y17382 = ~n53614 ;
  assign y17383 = ~n53615 ;
  assign y17384 = ~n53616 ;
  assign y17385 = ~n53621 ;
  assign y17386 = ~n53624 ;
  assign y17387 = ~n53625 ;
  assign y17388 = ~n53627 ;
  assign y17389 = ~n53628 ;
  assign y17390 = n53630 ;
  assign y17391 = n53633 ;
  assign y17392 = n53638 ;
  assign y17393 = n53640 ;
  assign y17394 = n53642 ;
  assign y17395 = n53646 ;
  assign y17396 = ~n53650 ;
  assign y17397 = n53652 ;
  assign y17398 = n53654 ;
  assign y17399 = ~n53655 ;
  assign y17400 = n53657 ;
  assign y17401 = ~n53658 ;
  assign y17402 = ~n53659 ;
  assign y17403 = ~n53662 ;
  assign y17404 = ~n53663 ;
  assign y17405 = ~n53666 ;
  assign y17406 = n53668 ;
  assign y17407 = ~n53670 ;
  assign y17408 = ~n53673 ;
  assign y17409 = ~n53674 ;
  assign y17410 = n53675 ;
  assign y17411 = ~n53676 ;
  assign y17412 = n53679 ;
  assign y17413 = ~n53680 ;
  assign y17414 = n53686 ;
  assign y17415 = n53689 ;
  assign y17416 = ~n53691 ;
  assign y17417 = ~n53693 ;
  assign y17418 = n53696 ;
  assign y17419 = ~n53699 ;
  assign y17420 = ~1'b0 ;
  assign y17421 = n53702 ;
  assign y17422 = n53704 ;
  assign y17423 = n53705 ;
  assign y17424 = n53706 ;
  assign y17425 = ~n53707 ;
  assign y17426 = n53708 ;
  assign y17427 = n53709 ;
  assign y17428 = n53711 ;
  assign y17429 = ~n53713 ;
  assign y17430 = n53715 ;
  assign y17431 = ~n53718 ;
  assign y17432 = n53719 ;
  assign y17433 = n53720 ;
  assign y17434 = n53721 ;
  assign y17435 = n53724 ;
  assign y17436 = ~n53725 ;
  assign y17437 = n53730 ;
  assign y17438 = ~1'b0 ;
  assign y17439 = ~1'b0 ;
  assign y17440 = n53732 ;
  assign y17441 = ~n53741 ;
  assign y17442 = n53742 ;
  assign y17443 = ~n53743 ;
  assign y17444 = ~n53746 ;
  assign y17445 = ~n53747 ;
  assign y17446 = n53748 ;
  assign y17447 = ~n53749 ;
  assign y17448 = ~n53757 ;
  assign y17449 = n53761 ;
  assign y17450 = ~1'b0 ;
  assign y17451 = n53762 ;
  assign y17452 = ~1'b0 ;
  assign y17453 = n53765 ;
  assign y17454 = n53766 ;
  assign y17455 = n53770 ;
  assign y17456 = ~n53771 ;
  assign y17457 = n53772 ;
  assign y17458 = n53773 ;
  assign y17459 = ~n53775 ;
  assign y17460 = ~n53777 ;
  assign y17461 = n53779 ;
  assign y17462 = ~1'b0 ;
  assign y17463 = ~n53780 ;
  assign y17464 = n53785 ;
  assign y17465 = ~n53789 ;
  assign y17466 = n53792 ;
  assign y17467 = ~n53793 ;
  assign y17468 = n53795 ;
  assign y17469 = n53798 ;
  assign y17470 = ~n53799 ;
  assign y17471 = n53801 ;
  assign y17472 = n53803 ;
  assign y17473 = ~n53807 ;
  assign y17474 = ~1'b0 ;
  assign y17475 = n53808 ;
  assign y17476 = ~1'b0 ;
  assign y17477 = n53813 ;
  assign y17478 = n53815 ;
  assign y17479 = n53817 ;
  assign y17480 = ~n53822 ;
  assign y17481 = n53824 ;
  assign y17482 = ~n53834 ;
  assign y17483 = n53837 ;
  assign y17484 = ~n53839 ;
  assign y17485 = ~n14318 ;
  assign y17486 = ~n53844 ;
  assign y17487 = ~n53847 ;
  assign y17488 = n53848 ;
  assign y17489 = ~n53852 ;
  assign y17490 = ~n53854 ;
  assign y17491 = ~n53856 ;
  assign y17492 = ~n53857 ;
  assign y17493 = ~n53858 ;
  assign y17494 = ~1'b0 ;
  assign y17495 = ~n53861 ;
  assign y17496 = ~n31832 ;
  assign y17497 = ~n53864 ;
  assign y17498 = n53867 ;
  assign y17499 = ~n53879 ;
  assign y17500 = n53881 ;
  assign y17501 = ~n53885 ;
  assign y17502 = ~n53886 ;
  assign y17503 = n53887 ;
  assign y17504 = ~n53890 ;
  assign y17505 = ~n53892 ;
  assign y17506 = ~1'b0 ;
  assign y17507 = ~1'b0 ;
  assign y17508 = ~n53893 ;
  assign y17509 = n53897 ;
  assign y17510 = n53902 ;
  assign y17511 = ~n53904 ;
  assign y17512 = ~n53905 ;
  assign y17513 = ~n53909 ;
  assign y17514 = ~n53913 ;
  assign y17515 = n53916 ;
  assign y17516 = n53918 ;
  assign y17517 = ~n53920 ;
  assign y17518 = ~1'b0 ;
  assign y17519 = n53921 ;
  assign y17520 = ~n53929 ;
  assign y17521 = ~n24053 ;
  assign y17522 = n53930 ;
  assign y17523 = n53931 ;
  assign y17524 = ~n53933 ;
  assign y17525 = ~n53937 ;
  assign y17526 = ~1'b0 ;
  assign y17527 = ~1'b0 ;
  assign y17528 = ~1'b0 ;
  assign y17529 = ~n53938 ;
  assign y17530 = ~n53939 ;
  assign y17531 = n53945 ;
  assign y17532 = ~n53946 ;
  assign y17533 = n53947 ;
  assign y17534 = ~n53950 ;
  assign y17535 = n16094 ;
  assign y17536 = n53953 ;
  assign y17537 = ~1'b0 ;
  assign y17538 = ~1'b0 ;
  assign y17539 = ~n53955 ;
  assign y17540 = n53957 ;
  assign y17541 = n53960 ;
  assign y17542 = n53962 ;
  assign y17543 = n53963 ;
  assign y17544 = n53967 ;
  assign y17545 = ~n53970 ;
  assign y17546 = n53972 ;
  assign y17547 = ~1'b0 ;
  assign y17548 = ~1'b0 ;
  assign y17549 = ~n53974 ;
  assign y17550 = ~1'b0 ;
  assign y17551 = ~n53980 ;
  assign y17552 = ~n53985 ;
  assign y17553 = ~n53986 ;
  assign y17554 = n53990 ;
  assign y17555 = n53992 ;
  assign y17556 = ~n53993 ;
  assign y17557 = ~n53995 ;
  assign y17558 = ~n53997 ;
  assign y17559 = ~1'b0 ;
  assign y17560 = ~n53998 ;
  assign y17561 = ~n5319 ;
  assign y17562 = ~n54000 ;
  assign y17563 = n54005 ;
  assign y17564 = ~n54006 ;
  assign y17565 = ~n54011 ;
  assign y17566 = n54013 ;
  assign y17567 = ~n54020 ;
  assign y17568 = ~n54023 ;
  assign y17569 = ~n54025 ;
  assign y17570 = n54028 ;
  assign y17571 = ~1'b0 ;
  assign y17572 = ~n54029 ;
  assign y17573 = n54030 ;
  assign y17574 = n40353 ;
  assign y17575 = n54033 ;
  assign y17576 = ~n54035 ;
  assign y17577 = n54039 ;
  assign y17578 = n54045 ;
  assign y17579 = ~n54047 ;
  assign y17580 = ~1'b0 ;
  assign y17581 = ~1'b0 ;
  assign y17582 = ~1'b0 ;
  assign y17583 = n54048 ;
  assign y17584 = n54050 ;
  assign y17585 = ~n54051 ;
  assign y17586 = ~n54061 ;
  assign y17587 = ~n54062 ;
  assign y17588 = ~n54064 ;
  assign y17589 = n54065 ;
  assign y17590 = n54067 ;
  assign y17591 = n54073 ;
  assign y17592 = n54074 ;
  assign y17593 = ~n54076 ;
  assign y17594 = n54078 ;
  assign y17595 = ~n54079 ;
  assign y17596 = n54081 ;
  assign y17597 = n54083 ;
  assign y17598 = n54084 ;
  assign y17599 = ~n54087 ;
  assign y17600 = ~n54089 ;
  assign y17601 = ~n54091 ;
  assign y17602 = n54094 ;
  assign y17603 = ~1'b0 ;
  assign y17604 = ~1'b0 ;
  assign y17605 = ~n54100 ;
  assign y17606 = ~n54101 ;
  assign y17607 = ~n54103 ;
  assign y17608 = ~n54105 ;
  assign y17609 = ~n54111 ;
  assign y17610 = n54113 ;
  assign y17611 = ~n54115 ;
  assign y17612 = n54122 ;
  assign y17613 = n54127 ;
  assign y17614 = n54129 ;
  assign y17615 = ~n54135 ;
  assign y17616 = n54139 ;
  assign y17617 = ~n54140 ;
  assign y17618 = n54144 ;
  assign y17619 = ~n54145 ;
  assign y17620 = ~n54147 ;
  assign y17621 = n54151 ;
  assign y17622 = n54152 ;
  assign y17623 = n54153 ;
  assign y17624 = ~1'b0 ;
  assign y17625 = ~n9062 ;
  assign y17626 = n54157 ;
  assign y17627 = ~n54159 ;
  assign y17628 = ~n54160 ;
  assign y17629 = ~n54162 ;
  assign y17630 = ~n54167 ;
  assign y17631 = ~n54176 ;
  assign y17632 = n54179 ;
  assign y17633 = n54182 ;
  assign y17634 = n54186 ;
  assign y17635 = ~n54188 ;
  assign y17636 = n54189 ;
  assign y17637 = ~n54191 ;
  assign y17638 = n54192 ;
  assign y17639 = n54193 ;
  assign y17640 = ~n54198 ;
  assign y17641 = ~n54200 ;
  assign y17642 = n54204 ;
  assign y17643 = n54206 ;
  assign y17644 = ~1'b0 ;
  assign y17645 = ~n54208 ;
  assign y17646 = ~1'b0 ;
  assign y17647 = n54213 ;
  assign y17648 = n54214 ;
  assign y17649 = ~n54218 ;
  assign y17650 = n54219 ;
  assign y17651 = n54220 ;
  assign y17652 = ~n54222 ;
  assign y17653 = ~n54224 ;
  assign y17654 = ~n54227 ;
  assign y17655 = ~n54229 ;
  assign y17656 = n54231 ;
  assign y17657 = ~n54233 ;
  assign y17658 = n54234 ;
  assign y17659 = n54235 ;
  assign y17660 = n54242 ;
  assign y17661 = ~n54243 ;
  assign y17662 = ~n54248 ;
  assign y17663 = ~n54253 ;
  assign y17664 = n54258 ;
  assign y17665 = ~n54259 ;
  assign y17666 = ~n54261 ;
  assign y17667 = ~1'b0 ;
  assign y17668 = ~n54264 ;
  assign y17669 = ~n54266 ;
  assign y17670 = n54267 ;
  assign y17671 = n54268 ;
  assign y17672 = n54269 ;
  assign y17673 = n54270 ;
  assign y17674 = n54276 ;
  assign y17675 = ~n54278 ;
  assign y17676 = ~n54281 ;
  assign y17677 = ~n54283 ;
  assign y17678 = ~n54287 ;
  assign y17679 = ~n54291 ;
  assign y17680 = ~n54297 ;
  assign y17681 = ~n54298 ;
  assign y17682 = n54299 ;
  assign y17683 = ~n54300 ;
  assign y17684 = n54302 ;
  assign y17685 = ~n54304 ;
  assign y17686 = ~n54311 ;
  assign y17687 = n54313 ;
  assign y17688 = n54315 ;
  assign y17689 = ~1'b0 ;
  assign y17690 = ~n54317 ;
  assign y17691 = ~n54319 ;
  assign y17692 = n54323 ;
  assign y17693 = ~n54326 ;
  assign y17694 = ~n54330 ;
  assign y17695 = n54331 ;
  assign y17696 = n54337 ;
  assign y17697 = n54339 ;
  assign y17698 = n54340 ;
  assign y17699 = ~1'b0 ;
  assign y17700 = ~1'b0 ;
  assign y17701 = n54341 ;
  assign y17702 = n54343 ;
  assign y17703 = ~n54344 ;
  assign y17704 = n54347 ;
  assign y17705 = n54348 ;
  assign y17706 = n54349 ;
  assign y17707 = n54355 ;
  assign y17708 = n54356 ;
  assign y17709 = n54361 ;
  assign y17710 = n54363 ;
  assign y17711 = n54367 ;
  assign y17712 = ~n54369 ;
  assign y17713 = ~n54373 ;
  assign y17714 = n54375 ;
  assign y17715 = n54378 ;
  assign y17716 = ~n54380 ;
  assign y17717 = n54385 ;
  assign y17718 = n54386 ;
  assign y17719 = ~n54387 ;
  assign y17720 = n43363 ;
  assign y17721 = n54391 ;
  assign y17722 = n54394 ;
  assign y17723 = n54396 ;
  assign y17724 = n54397 ;
  assign y17725 = n54399 ;
  assign y17726 = n54400 ;
  assign y17727 = n54401 ;
  assign y17728 = ~n54406 ;
  assign y17729 = ~n4729 ;
  assign y17730 = ~n54409 ;
  assign y17731 = n54412 ;
  assign y17732 = ~1'b0 ;
  assign y17733 = n54414 ;
  assign y17734 = n54416 ;
  assign y17735 = ~1'b0 ;
  assign y17736 = n54417 ;
  assign y17737 = n54419 ;
  assign y17738 = ~n54422 ;
  assign y17739 = ~n54423 ;
  assign y17740 = ~n54424 ;
  assign y17741 = n54425 ;
  assign y17742 = ~n54429 ;
  assign y17743 = ~1'b0 ;
  assign y17744 = ~1'b0 ;
  assign y17745 = ~n54433 ;
  assign y17746 = ~n54434 ;
  assign y17747 = n54437 ;
  assign y17748 = ~n54439 ;
  assign y17749 = ~n54448 ;
  assign y17750 = ~n54449 ;
  assign y17751 = ~n54450 ;
  assign y17752 = ~1'b0 ;
  assign y17753 = ~n54452 ;
  assign y17754 = ~1'b0 ;
  assign y17755 = n54453 ;
  assign y17756 = n54455 ;
  assign y17757 = n54456 ;
  assign y17758 = n54457 ;
  assign y17759 = n54464 ;
  assign y17760 = ~n54465 ;
  assign y17761 = n54466 ;
  assign y17762 = ~n54469 ;
  assign y17763 = ~n54471 ;
  assign y17764 = ~1'b0 ;
  assign y17765 = ~1'b0 ;
  assign y17766 = n54475 ;
  assign y17767 = n54476 ;
  assign y17768 = ~n54477 ;
  assign y17769 = ~n54480 ;
  assign y17770 = ~n54481 ;
  assign y17771 = ~n54487 ;
  assign y17772 = ~n54488 ;
  assign y17773 = n54492 ;
  assign y17774 = n54494 ;
  assign y17775 = ~1'b0 ;
  assign y17776 = ~n54497 ;
  assign y17777 = ~1'b0 ;
  assign y17778 = ~n24374 ;
  assign y17779 = ~n54499 ;
  assign y17780 = ~n54500 ;
  assign y17781 = ~n54501 ;
  assign y17782 = ~n54504 ;
  assign y17783 = n54505 ;
  assign y17784 = ~n54508 ;
  assign y17785 = n54511 ;
  assign y17786 = n54515 ;
  assign y17787 = n54516 ;
  assign y17788 = ~1'b0 ;
  assign y17789 = n54520 ;
  assign y17790 = ~n54521 ;
  assign y17791 = ~n54523 ;
  assign y17792 = ~n54528 ;
  assign y17793 = ~n54529 ;
  assign y17794 = n54532 ;
  assign y17795 = ~n54533 ;
  assign y17796 = ~n54535 ;
  assign y17797 = ~n54537 ;
  assign y17798 = n54538 ;
  assign y17799 = n54539 ;
  assign y17800 = ~n54540 ;
  assign y17801 = ~n54544 ;
  assign y17802 = ~n54548 ;
  assign y17803 = n54549 ;
  assign y17804 = n54553 ;
  assign y17805 = ~n54558 ;
  assign y17806 = ~n54561 ;
  assign y17807 = ~1'b0 ;
  assign y17808 = ~n54563 ;
  assign y17809 = n54565 ;
  assign y17810 = ~1'b0 ;
  assign y17811 = ~n54566 ;
  assign y17812 = n54567 ;
  assign y17813 = n54570 ;
  assign y17814 = ~n54573 ;
  assign y17815 = ~n54574 ;
  assign y17816 = n54575 ;
  assign y17817 = n54576 ;
  assign y17818 = n54578 ;
  assign y17819 = ~n54580 ;
  assign y17820 = ~1'b0 ;
  assign y17821 = n54582 ;
  assign y17822 = ~n54586 ;
  assign y17823 = ~n54590 ;
  assign y17824 = ~n54592 ;
  assign y17825 = n54596 ;
  assign y17826 = ~n54597 ;
  assign y17827 = ~n54599 ;
  assign y17828 = n54601 ;
  assign y17829 = ~n54604 ;
  assign y17830 = ~n54606 ;
  assign y17831 = ~1'b0 ;
  assign y17832 = n54609 ;
  assign y17833 = ~n54614 ;
  assign y17834 = ~1'b0 ;
  assign y17835 = ~n54615 ;
  assign y17836 = n54616 ;
  assign y17837 = ~n54618 ;
  assign y17838 = ~n54619 ;
  assign y17839 = n54620 ;
  assign y17840 = n54623 ;
  assign y17841 = n54625 ;
  assign y17842 = ~n54627 ;
  assign y17843 = n54628 ;
  assign y17844 = ~n54629 ;
  assign y17845 = ~n54630 ;
  assign y17846 = ~n54631 ;
  assign y17847 = n54634 ;
  assign y17848 = n54635 ;
  assign y17849 = n54636 ;
  assign y17850 = ~n54638 ;
  assign y17851 = n54640 ;
  assign y17852 = ~1'b0 ;
  assign y17853 = ~1'b0 ;
  assign y17854 = ~1'b0 ;
  assign y17855 = n54641 ;
  assign y17856 = n54643 ;
  assign y17857 = ~n54645 ;
  assign y17858 = ~n54648 ;
  assign y17859 = n54649 ;
  assign y17860 = ~n54650 ;
  assign y17861 = n54651 ;
  assign y17862 = ~1'b0 ;
  assign y17863 = n54653 ;
  assign y17864 = ~1'b0 ;
  assign y17865 = ~n54659 ;
  assign y17866 = ~n54663 ;
  assign y17867 = ~n54664 ;
  assign y17868 = n54666 ;
  assign y17869 = n54667 ;
  assign y17870 = ~n54670 ;
  assign y17871 = ~n54675 ;
  assign y17872 = ~n54676 ;
  assign y17873 = n54680 ;
  assign y17874 = ~1'b0 ;
  assign y17875 = ~1'b0 ;
  assign y17876 = ~n54682 ;
  assign y17877 = n54684 ;
  assign y17878 = n54685 ;
  assign y17879 = ~n54687 ;
  assign y17880 = n54688 ;
  assign y17881 = n54690 ;
  assign y17882 = ~n54691 ;
  assign y17883 = ~n54692 ;
  assign y17884 = ~n54696 ;
  assign y17885 = n54697 ;
  assign y17886 = n54699 ;
  assign y17887 = ~1'b0 ;
  assign y17888 = n54700 ;
  assign y17889 = ~n54704 ;
  assign y17890 = ~n54705 ;
  assign y17891 = n54711 ;
  assign y17892 = ~n54712 ;
  assign y17893 = n54714 ;
  assign y17894 = ~n54717 ;
  assign y17895 = ~n54722 ;
  assign y17896 = ~n54726 ;
  assign y17897 = ~1'b0 ;
  assign y17898 = n54729 ;
  assign y17899 = ~n54732 ;
  assign y17900 = ~n54734 ;
  assign y17901 = ~n54735 ;
  assign y17902 = ~n54737 ;
  assign y17903 = ~n54739 ;
  assign y17904 = ~n54741 ;
  assign y17905 = n54742 ;
  assign y17906 = ~n54744 ;
  assign y17907 = n54746 ;
  assign y17908 = ~n54748 ;
  assign y17909 = ~n54749 ;
  assign y17910 = ~n54754 ;
  assign y17911 = ~n54756 ;
  assign y17912 = ~n54758 ;
  assign y17913 = n54759 ;
  assign y17914 = ~n54763 ;
  assign y17915 = n28764 ;
  assign y17916 = ~n54770 ;
  assign y17917 = ~n54772 ;
  assign y17918 = ~n54779 ;
  assign y17919 = n54782 ;
  assign y17920 = n54786 ;
  assign y17921 = ~n54787 ;
  assign y17922 = ~n54789 ;
  assign y17923 = ~n54797 ;
  assign y17924 = n54800 ;
  assign y17925 = ~n54801 ;
  assign y17926 = ~n54804 ;
  assign y17927 = n54806 ;
  assign y17928 = ~n54807 ;
  assign y17929 = ~n54808 ;
  assign y17930 = ~1'b0 ;
  assign y17931 = n54810 ;
  assign y17932 = n54811 ;
  assign y17933 = n54814 ;
  assign y17934 = n54816 ;
  assign y17935 = n54817 ;
  assign y17936 = ~n54820 ;
  assign y17937 = n54821 ;
  assign y17938 = n54822 ;
  assign y17939 = ~1'b0 ;
  assign y17940 = ~n54824 ;
  assign y17941 = n54825 ;
  assign y17942 = ~n54826 ;
  assign y17943 = ~n54828 ;
  assign y17944 = ~n54832 ;
  assign y17945 = ~n54834 ;
  assign y17946 = n54835 ;
  assign y17947 = n54837 ;
  assign y17948 = ~n54839 ;
  assign y17949 = ~n54843 ;
  assign y17950 = ~n54849 ;
  assign y17951 = ~n54854 ;
  assign y17952 = n54858 ;
  assign y17953 = n54862 ;
  assign y17954 = n54863 ;
  assign y17955 = ~n54864 ;
  assign y17956 = ~n54868 ;
  assign y17957 = ~n54869 ;
  assign y17958 = ~n54871 ;
  assign y17959 = n54875 ;
  assign y17960 = ~n54877 ;
  assign y17961 = ~1'b0 ;
  assign y17962 = ~n54879 ;
  assign y17963 = ~1'b0 ;
  assign y17964 = ~n54881 ;
  assign y17965 = n54882 ;
  assign y17966 = ~n54885 ;
  assign y17967 = n54886 ;
  assign y17968 = ~n54887 ;
  assign y17969 = ~n54888 ;
  assign y17970 = n54890 ;
  assign y17971 = ~1'b0 ;
  assign y17972 = n54892 ;
  assign y17973 = n54894 ;
  assign y17974 = ~1'b0 ;
  assign y17975 = n54895 ;
  assign y17976 = n54897 ;
  assign y17977 = ~n54898 ;
  assign y17978 = n54899 ;
  assign y17979 = n54900 ;
  assign y17980 = n54904 ;
  assign y17981 = ~n54909 ;
  assign y17982 = ~n54915 ;
  assign y17983 = ~n54917 ;
  assign y17984 = ~n54919 ;
  assign y17985 = ~1'b0 ;
  assign y17986 = ~n54923 ;
  assign y17987 = ~n54929 ;
  assign y17988 = n54930 ;
  assign y17989 = ~n54934 ;
  assign y17990 = ~n54937 ;
  assign y17991 = n54939 ;
  assign y17992 = ~n54945 ;
  assign y17993 = n54946 ;
  assign y17994 = n54949 ;
  assign y17995 = ~n54951 ;
  assign y17996 = ~1'b0 ;
  assign y17997 = n9983 ;
  assign y17998 = n54952 ;
  assign y17999 = n54953 ;
  assign y18000 = n54956 ;
  assign y18001 = n54961 ;
  assign y18002 = n54968 ;
  assign y18003 = n54972 ;
  assign y18004 = ~n54977 ;
  assign y18005 = ~1'b0 ;
  assign y18006 = ~1'b0 ;
  assign y18007 = n54979 ;
  assign y18008 = ~n54985 ;
  assign y18009 = n54987 ;
  assign y18010 = ~n54988 ;
  assign y18011 = n39547 ;
  assign y18012 = ~n54990 ;
  assign y18013 = n54992 ;
  assign y18014 = n54995 ;
  assign y18015 = ~n54999 ;
  assign y18016 = n55003 ;
  assign y18017 = ~n55006 ;
  assign y18018 = ~n55008 ;
  assign y18019 = ~n55011 ;
  assign y18020 = ~n55013 ;
  assign y18021 = ~n55015 ;
  assign y18022 = n55016 ;
  assign y18023 = n55017 ;
  assign y18024 = n55018 ;
  assign y18025 = ~n55019 ;
  assign y18026 = ~n55021 ;
  assign y18027 = ~n55023 ;
  assign y18028 = ~n55028 ;
  assign y18029 = ~n55029 ;
  assign y18030 = ~n55030 ;
  assign y18031 = n55032 ;
  assign y18032 = ~n55033 ;
  assign y18033 = ~n55035 ;
  assign y18034 = ~n55036 ;
  assign y18035 = ~n55038 ;
  assign y18036 = n55039 ;
  assign y18037 = ~n55041 ;
endmodule
