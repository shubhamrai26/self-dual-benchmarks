module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 ;
  assign n129 = ( x5 & x113 ) | ( x5 & ~x120 ) | ( x113 & ~x120 ) ;
  assign n130 = n129 ^ x83 ^ x71 ;
  assign n131 = n130 ^ x95 ^ x73 ;
  assign n132 = x82 ^ x21 ^ x10 ;
  assign n133 = x117 ^ x101 ^ x25 ;
  assign n134 = ( x53 & ~x104 ) | ( x53 & n133 ) | ( ~x104 & n133 ) ;
  assign n135 = ( x83 & ~x97 ) | ( x83 & n134 ) | ( ~x97 & n134 ) ;
  assign n136 = ( x53 & n132 ) | ( x53 & ~n135 ) | ( n132 & ~n135 ) ;
  assign n144 = x75 ^ x50 ^ x47 ;
  assign n145 = ( x62 & ~x105 ) | ( x62 & n144 ) | ( ~x105 & n144 ) ;
  assign n150 = n145 ^ x74 ^ x19 ;
  assign n151 = n150 ^ x28 ^ x9 ;
  assign n149 = ( x9 & ~x18 ) | ( x9 & x125 ) | ( ~x18 & x125 ) ;
  assign n147 = x51 ^ x16 ^ x12 ;
  assign n146 = n145 ^ x69 ^ x9 ;
  assign n137 = ( x1 & ~x39 ) | ( x1 & x126 ) | ( ~x39 & x126 ) ;
  assign n138 = x51 ^ x40 ^ x19 ;
  assign n139 = ( x56 & ~x99 ) | ( x56 & n138 ) | ( ~x99 & n138 ) ;
  assign n140 = ( ~x18 & x44 ) | ( ~x18 & x96 ) | ( x44 & x96 ) ;
  assign n141 = ( x27 & x96 ) | ( x27 & ~n140 ) | ( x96 & ~n140 ) ;
  assign n142 = ( x33 & x47 ) | ( x33 & ~n141 ) | ( x47 & ~n141 ) ;
  assign n143 = ( n137 & n139 ) | ( n137 & n142 ) | ( n139 & n142 ) ;
  assign n148 = n147 ^ n146 ^ n143 ;
  assign n152 = n151 ^ n149 ^ n148 ;
  assign n153 = ( x57 & ~x90 ) | ( x57 & x100 ) | ( ~x90 & x100 ) ;
  assign n154 = n141 ^ x106 ^ x16 ;
  assign n156 = ( x3 & x7 ) | ( x3 & ~x115 ) | ( x7 & ~x115 ) ;
  assign n155 = ( x4 & x35 ) | ( x4 & ~x108 ) | ( x35 & ~x108 ) ;
  assign n157 = n156 ^ n155 ^ x106 ;
  assign n158 = ( x20 & ~x25 ) | ( x20 & x99 ) | ( ~x25 & x99 ) ;
  assign n159 = n158 ^ n137 ^ x77 ;
  assign n160 = ( x46 & x109 ) | ( x46 & ~x125 ) | ( x109 & ~x125 ) ;
  assign n161 = n158 ^ x61 ^ x29 ;
  assign n162 = n161 ^ x116 ^ x30 ;
  assign n163 = ( x87 & n160 ) | ( x87 & ~n162 ) | ( n160 & ~n162 ) ;
  assign n164 = ( ~x40 & n159 ) | ( ~x40 & n163 ) | ( n159 & n163 ) ;
  assign n165 = ( x7 & n157 ) | ( x7 & n164 ) | ( n157 & n164 ) ;
  assign n166 = ( n153 & n154 ) | ( n153 & n165 ) | ( n154 & n165 ) ;
  assign n167 = ( n136 & ~n152 ) | ( n136 & n166 ) | ( ~n152 & n166 ) ;
  assign n184 = n151 ^ x120 ^ x65 ;
  assign n182 = ( x14 & ~x48 ) | ( x14 & x109 ) | ( ~x48 & x109 ) ;
  assign n183 = n182 ^ x126 ^ x6 ;
  assign n178 = x107 ^ x27 ^ x1 ;
  assign n170 = ( ~x93 & x104 ) | ( ~x93 & x117 ) | ( x104 & x117 ) ;
  assign n171 = ( ~x4 & x58 ) | ( ~x4 & n170 ) | ( x58 & n170 ) ;
  assign n179 = n171 ^ n129 ^ x70 ;
  assign n180 = ( x75 & ~n178 ) | ( x75 & n179 ) | ( ~n178 & n179 ) ;
  assign n168 = x126 ^ x97 ^ x34 ;
  assign n169 = ( x27 & ~x89 ) | ( x27 & x104 ) | ( ~x89 & x104 ) ;
  assign n172 = n171 ^ n169 ^ x62 ;
  assign n173 = n172 ^ x74 ^ x73 ;
  assign n174 = x86 ^ x57 ^ x43 ;
  assign n175 = ( ~x17 & x95 ) | ( ~x17 & n174 ) | ( x95 & n174 ) ;
  assign n176 = ( x120 & x122 ) | ( x120 & n175 ) | ( x122 & n175 ) ;
  assign n177 = ( n168 & n173 ) | ( n168 & n176 ) | ( n173 & n176 ) ;
  assign n181 = n180 ^ n177 ^ x26 ;
  assign n185 = n184 ^ n183 ^ n181 ;
  assign n205 = ( x6 & x92 ) | ( x6 & ~x93 ) | ( x92 & ~x93 ) ;
  assign n203 = ( ~x31 & x76 ) | ( ~x31 & x113 ) | ( x76 & x113 ) ;
  assign n204 = n203 ^ x58 ^ x11 ;
  assign n206 = n205 ^ n204 ^ x52 ;
  assign n186 = ( x44 & x108 ) | ( x44 & ~x127 ) | ( x108 & ~x127 ) ;
  assign n201 = n186 ^ n173 ^ x21 ;
  assign n200 = ( x10 & ~x44 ) | ( x10 & x54 ) | ( ~x44 & x54 ) ;
  assign n202 = n201 ^ n200 ^ x11 ;
  assign n187 = ( x99 & x110 ) | ( x99 & ~n186 ) | ( x110 & ~n186 ) ;
  assign n188 = ( ~x106 & x123 ) | ( ~x106 & n178 ) | ( x123 & n178 ) ;
  assign n189 = n188 ^ x115 ^ x54 ;
  assign n192 = n169 ^ n157 ^ x119 ;
  assign n190 = n156 ^ x92 ^ x71 ;
  assign n191 = n190 ^ x78 ^ x34 ;
  assign n193 = n192 ^ n191 ^ x82 ;
  assign n194 = ( x5 & ~x34 ) | ( x5 & x124 ) | ( ~x34 & x124 ) ;
  assign n195 = n194 ^ x114 ^ x37 ;
  assign n196 = ( x21 & ~n153 ) | ( x21 & n195 ) | ( ~n153 & n195 ) ;
  assign n197 = ( ~x37 & x102 ) | ( ~x37 & n196 ) | ( x102 & n196 ) ;
  assign n198 = ( x91 & n193 ) | ( x91 & n197 ) | ( n193 & n197 ) ;
  assign n199 = ( ~n187 & n189 ) | ( ~n187 & n198 ) | ( n189 & n198 ) ;
  assign n207 = n206 ^ n202 ^ n199 ;
  assign n208 = n207 ^ n132 ^ x103 ;
  assign n209 = ( x65 & x82 ) | ( x65 & ~x96 ) | ( x82 & ~x96 ) ;
  assign n210 = n209 ^ n196 ^ x26 ;
  assign n211 = ( n173 & n201 ) | ( n173 & n210 ) | ( n201 & n210 ) ;
  assign n212 = ( n185 & n208 ) | ( n185 & ~n211 ) | ( n208 & ~n211 ) ;
  assign n228 = ( x42 & x94 ) | ( x42 & ~x97 ) | ( x94 & ~x97 ) ;
  assign n229 = n228 ^ x102 ^ x99 ;
  assign n223 = ( x77 & ~x93 ) | ( x77 & x111 ) | ( ~x93 & x111 ) ;
  assign n224 = n223 ^ x94 ^ x15 ;
  assign n225 = x105 ^ x49 ^ x17 ;
  assign n226 = n225 ^ x79 ^ x55 ;
  assign n227 = ( x74 & n224 ) | ( x74 & n226 ) | ( n224 & n226 ) ;
  assign n215 = ( x73 & ~x104 ) | ( x73 & x111 ) | ( ~x104 & x111 ) ;
  assign n219 = ( x96 & ~x103 ) | ( x96 & n205 ) | ( ~x103 & n205 ) ;
  assign n220 = ( ~n137 & n215 ) | ( ~n137 & n219 ) | ( n215 & n219 ) ;
  assign n221 = ( x104 & ~n173 ) | ( x104 & n220 ) | ( ~n173 & n220 ) ;
  assign n213 = x119 ^ x114 ^ x64 ;
  assign n214 = n213 ^ x79 ^ x48 ;
  assign n216 = n215 ^ n159 ^ x19 ;
  assign n217 = ( x4 & n214 ) | ( x4 & ~n216 ) | ( n214 & ~n216 ) ;
  assign n218 = n217 ^ x106 ^ x31 ;
  assign n222 = n221 ^ n218 ^ n172 ;
  assign n230 = n229 ^ n227 ^ n222 ;
  assign n235 = ( ~x62 & x81 ) | ( ~x62 & n200 ) | ( x81 & n200 ) ;
  assign n233 = ( x16 & ~x40 ) | ( x16 & x118 ) | ( ~x40 & x118 ) ;
  assign n234 = n233 ^ x98 ^ x62 ;
  assign n231 = n215 ^ x84 ^ x12 ;
  assign n232 = ( n167 & n180 ) | ( n167 & n231 ) | ( n180 & n231 ) ;
  assign n236 = n235 ^ n234 ^ n232 ;
  assign n239 = ( x41 & x55 ) | ( x41 & ~x115 ) | ( x55 & ~x115 ) ;
  assign n237 = ( x33 & x38 ) | ( x33 & ~x89 ) | ( x38 & ~x89 ) ;
  assign n238 = n237 ^ n187 ^ x3 ;
  assign n240 = n239 ^ n238 ^ x108 ;
  assign n241 = ( x97 & ~n184 ) | ( x97 & n186 ) | ( ~n184 & n186 ) ;
  assign n242 = ( x9 & x13 ) | ( x9 & ~x54 ) | ( x13 & ~x54 ) ;
  assign n243 = ( n240 & n241 ) | ( n240 & ~n242 ) | ( n241 & ~n242 ) ;
  assign n244 = ( n230 & n236 ) | ( n230 & n243 ) | ( n236 & n243 ) ;
  assign n245 = ( n167 & n212 ) | ( n167 & ~n244 ) | ( n212 & ~n244 ) ;
  assign n251 = x116 ^ x113 ^ x91 ;
  assign n252 = ( x65 & x106 ) | ( x65 & n251 ) | ( x106 & n251 ) ;
  assign n253 = n252 ^ n155 ^ x19 ;
  assign n246 = ( ~x64 & x88 ) | ( ~x64 & x97 ) | ( x88 & x97 ) ;
  assign n247 = n246 ^ x54 ^ x48 ;
  assign n248 = ( n161 & n187 ) | ( n161 & n247 ) | ( n187 & n247 ) ;
  assign n249 = x71 ^ x14 ^ x3 ;
  assign n250 = ( n147 & n248 ) | ( n147 & ~n249 ) | ( n248 & ~n249 ) ;
  assign n254 = n253 ^ n250 ^ x56 ;
  assign n318 = x106 ^ x66 ^ x6 ;
  assign n421 = ( x89 & ~x108 ) | ( x89 & n318 ) | ( ~x108 & n318 ) ;
  assign n375 = ( x63 & ~x81 ) | ( x63 & x120 ) | ( ~x81 & x120 ) ;
  assign n422 = ( n157 & ~n178 ) | ( n157 & n375 ) | ( ~n178 & n375 ) ;
  assign n423 = ( x24 & ~x108 ) | ( x24 & n160 ) | ( ~x108 & n160 ) ;
  assign n424 = n423 ^ x66 ^ x30 ;
  assign n425 = x122 ^ x102 ^ x96 ;
  assign n426 = n425 ^ n129 ^ x29 ;
  assign n376 = n375 ^ n203 ^ x21 ;
  assign n377 = n376 ^ x124 ^ x49 ;
  assign n378 = n377 ^ n168 ^ x99 ;
  assign n427 = n426 ^ n378 ^ x72 ;
  assign n428 = ( x27 & n424 ) | ( x27 & ~n427 ) | ( n424 & ~n427 ) ;
  assign n429 = ( n421 & ~n422 ) | ( n421 & n428 ) | ( ~n422 & n428 ) ;
  assign n282 = x121 ^ x30 ^ x23 ;
  assign n283 = n282 ^ x66 ^ x50 ;
  assign n280 = n158 ^ x16 ^ x8 ;
  assign n279 = ( n156 & n173 ) | ( n156 & n174 ) | ( n173 & n174 ) ;
  assign n281 = n280 ^ n279 ^ n215 ;
  assign n284 = n283 ^ n281 ^ x8 ;
  assign n273 = n238 ^ n196 ^ x117 ;
  assign n274 = n273 ^ n194 ^ x71 ;
  assign n285 = ( x53 & x116 ) | ( x53 & n130 ) | ( x116 & n130 ) ;
  assign n286 = x103 ^ x68 ^ x15 ;
  assign n287 = ( x41 & ~x96 ) | ( x41 & n286 ) | ( ~x96 & n286 ) ;
  assign n288 = ( n274 & ~n285 ) | ( n274 & n287 ) | ( ~n285 & n287 ) ;
  assign n289 = ( x124 & ~n284 ) | ( x124 & n288 ) | ( ~n284 & n288 ) ;
  assign n292 = ( ~x54 & x90 ) | ( ~x54 & x91 ) | ( x90 & x91 ) ;
  assign n290 = ( x25 & ~n149 ) | ( x25 & n204 ) | ( ~n149 & n204 ) ;
  assign n259 = x73 ^ x47 ^ x36 ;
  assign n260 = ( x90 & ~n129 ) | ( x90 & n259 ) | ( ~n129 & n259 ) ;
  assign n261 = ( ~x5 & x106 ) | ( ~x5 & n260 ) | ( x106 & n260 ) ;
  assign n291 = n290 ^ n261 ^ x50 ;
  assign n293 = n292 ^ n291 ^ n284 ;
  assign n294 = ( x5 & x118 ) | ( x5 & n195 ) | ( x118 & n195 ) ;
  assign n295 = ( x47 & n161 ) | ( x47 & n294 ) | ( n161 & n294 ) ;
  assign n296 = ( x119 & n238 ) | ( x119 & n295 ) | ( n238 & n295 ) ;
  assign n297 = n296 ^ x62 ^ x12 ;
  assign n298 = ( n156 & ~n198 ) | ( n156 & n297 ) | ( ~n198 & n297 ) ;
  assign n299 = ( x121 & ~n134 ) | ( x121 & n225 ) | ( ~n134 & n225 ) ;
  assign n300 = n280 ^ x98 ^ x86 ;
  assign n301 = ( ~x31 & n210 ) | ( ~x31 & n300 ) | ( n210 & n300 ) ;
  assign n302 = n301 ^ n284 ^ n205 ;
  assign n303 = ( ~x58 & n299 ) | ( ~x58 & n302 ) | ( n299 & n302 ) ;
  assign n304 = ( ~x103 & n228 ) | ( ~x103 & n303 ) | ( n228 & n303 ) ;
  assign n305 = ( n183 & n298 ) | ( n183 & n304 ) | ( n298 & n304 ) ;
  assign n306 = ( ~n289 & n293 ) | ( ~n289 & n305 ) | ( n293 & n305 ) ;
  assign n276 = ( x21 & x59 ) | ( x21 & ~x81 ) | ( x59 & ~x81 ) ;
  assign n277 = n276 ^ x81 ^ x17 ;
  assign n278 = n277 ^ n237 ^ n227 ;
  assign n307 = n306 ^ n285 ^ n278 ;
  assign n270 = ( x50 & n130 ) | ( x50 & ~n158 ) | ( n130 & ~n158 ) ;
  assign n271 = n270 ^ n224 ^ x50 ;
  assign n257 = x118 ^ x112 ^ x90 ;
  assign n256 = x117 ^ x112 ^ x0 ;
  assign n258 = n257 ^ n256 ^ x113 ;
  assign n262 = x107 ^ x100 ^ x56 ;
  assign n263 = ( x74 & ~x88 ) | ( x74 & n262 ) | ( ~x88 & n262 ) ;
  assign n264 = ( x112 & ~n261 ) | ( x112 & n263 ) | ( ~n261 & n263 ) ;
  assign n265 = x106 ^ x59 ^ x44 ;
  assign n266 = ( x39 & ~n187 ) | ( x39 & n265 ) | ( ~n187 & n265 ) ;
  assign n267 = ( x41 & n226 ) | ( x41 & n266 ) | ( n226 & n266 ) ;
  assign n268 = ( n258 & n264 ) | ( n258 & n267 ) | ( n264 & n267 ) ;
  assign n255 = n196 ^ n188 ^ x108 ;
  assign n269 = n268 ^ n255 ^ n169 ;
  assign n272 = n271 ^ n269 ^ x89 ;
  assign n275 = n274 ^ n272 ^ x70 ;
  assign n308 = n307 ^ n299 ^ n275 ;
  assign n416 = ( ~x2 & n135 ) | ( ~x2 & n173 ) | ( n135 & n173 ) ;
  assign n333 = n281 ^ n264 ^ x85 ;
  assign n417 = n416 ^ n333 ^ n144 ;
  assign n409 = n292 ^ x125 ^ x28 ;
  assign n410 = ( ~n168 & n292 ) | ( ~n168 & n409 ) | ( n292 & n409 ) ;
  assign n412 = ( x54 & x99 ) | ( x54 & ~n150 ) | ( x99 & ~n150 ) ;
  assign n327 = n203 ^ n156 ^ n139 ;
  assign n411 = n327 ^ n209 ^ x1 ;
  assign n413 = n412 ^ n411 ^ n180 ;
  assign n340 = n284 ^ x123 ^ x10 ;
  assign n403 = ( n210 & n256 ) | ( n210 & n340 ) | ( n256 & n340 ) ;
  assign n404 = n403 ^ n194 ^ x55 ;
  assign n414 = n404 ^ n233 ^ x107 ;
  assign n415 = ( n410 & n413 ) | ( n410 & ~n414 ) | ( n413 & ~n414 ) ;
  assign n418 = n417 ^ n415 ^ n185 ;
  assign n405 = ( ~x7 & x17 ) | ( ~x7 & x42 ) | ( x17 & x42 ) ;
  assign n406 = ( n146 & n404 ) | ( n146 & ~n405 ) | ( n404 & ~n405 ) ;
  assign n407 = n406 ^ n188 ^ x43 ;
  assign n366 = ( x60 & ~n130 ) | ( x60 & n164 ) | ( ~n130 & n164 ) ;
  assign n402 = ( ~n155 & n170 ) | ( ~n155 & n366 ) | ( n170 & n366 ) ;
  assign n408 = n407 ^ n405 ^ n402 ;
  assign n393 = x61 ^ x11 ^ x5 ;
  assign n394 = ( ~x3 & x71 ) | ( ~x3 & n393 ) | ( x71 & n393 ) ;
  assign n395 = n394 ^ n294 ^ x121 ;
  assign n396 = ( n260 & ~n273 ) | ( n260 & n395 ) | ( ~n273 & n395 ) ;
  assign n397 = n396 ^ n263 ^ n258 ;
  assign n348 = ( x40 & ~x109 ) | ( x40 & n301 ) | ( ~x109 & n301 ) ;
  assign n398 = ( ~x11 & n348 ) | ( ~x11 & n396 ) | ( n348 & n396 ) ;
  assign n399 = n398 ^ n179 ^ x75 ;
  assign n400 = ( n282 & n397 ) | ( n282 & n399 ) | ( n397 & n399 ) ;
  assign n383 = n206 ^ n156 ^ n149 ;
  assign n391 = n383 ^ n215 ^ x113 ;
  assign n357 = x67 ^ x41 ^ x22 ;
  assign n363 = n357 ^ n296 ^ x66 ;
  assign n390 = n363 ^ n293 ^ x1 ;
  assign n330 = n262 ^ x125 ^ x12 ;
  assign n341 = n170 ^ x108 ^ x88 ;
  assign n342 = ( x28 & n330 ) | ( x28 & n341 ) | ( n330 & n341 ) ;
  assign n343 = ( ~n276 & n340 ) | ( ~n276 & n342 ) | ( n340 & n342 ) ;
  assign n344 = n343 ^ x61 ^ x34 ;
  assign n345 = ( n143 & ~n182 ) | ( n143 & n344 ) | ( ~n182 & n344 ) ;
  assign n384 = n239 ^ x35 ^ x33 ;
  assign n385 = ( n246 & ~n251 ) | ( n246 & n384 ) | ( ~n251 & n384 ) ;
  assign n386 = ( ~n251 & n383 ) | ( ~n251 & n385 ) | ( n383 & n385 ) ;
  assign n387 = n260 ^ x111 ^ x79 ;
  assign n388 = ( n345 & n386 ) | ( n345 & ~n387 ) | ( n386 & ~n387 ) ;
  assign n370 = n270 ^ n266 ^ n170 ;
  assign n371 = x117 ^ x90 ^ x14 ;
  assign n372 = n371 ^ n165 ^ n131 ;
  assign n373 = ( ~x115 & x127 ) | ( ~x115 & n175 ) | ( x127 & n175 ) ;
  assign n374 = ( x23 & n270 ) | ( x23 & n373 ) | ( n270 & n373 ) ;
  assign n379 = ( x69 & ~x81 ) | ( x69 & n140 ) | ( ~x81 & n140 ) ;
  assign n380 = ( n177 & n378 ) | ( n177 & ~n379 ) | ( n378 & ~n379 ) ;
  assign n381 = ( n372 & n374 ) | ( n372 & n380 ) | ( n374 & n380 ) ;
  assign n382 = ( x10 & ~n370 ) | ( x10 & n381 ) | ( ~n370 & n381 ) ;
  assign n389 = n388 ^ n382 ^ n373 ;
  assign n392 = n391 ^ n390 ^ n389 ;
  assign n368 = n345 ^ x75 ^ x18 ;
  assign n337 = n219 ^ x107 ^ x14 ;
  assign n338 = n337 ^ x61 ^ x9 ;
  assign n364 = n363 ^ x121 ^ x24 ;
  assign n365 = ( x33 & n338 ) | ( x33 & n364 ) | ( n338 & n364 ) ;
  assign n326 = x80 ^ x55 ^ x40 ;
  assign n328 = n327 ^ n168 ^ n147 ;
  assign n329 = n328 ^ x126 ^ x15 ;
  assign n331 = ( x101 & ~x113 ) | ( x101 & n168 ) | ( ~x113 & n168 ) ;
  assign n332 = ( x91 & ~n330 ) | ( x91 & n331 ) | ( ~n330 & n331 ) ;
  assign n334 = n333 ^ n168 ^ x35 ;
  assign n319 = n318 ^ x82 ^ x49 ;
  assign n335 = n334 ^ n319 ^ x1 ;
  assign n336 = ( ~n149 & n318 ) | ( ~n149 & n335 ) | ( n318 & n335 ) ;
  assign n349 = ( ~x59 & n219 ) | ( ~x59 & n291 ) | ( n219 & n291 ) ;
  assign n350 = ( x58 & ~n171 ) | ( x58 & n349 ) | ( ~n171 & n349 ) ;
  assign n351 = ( x115 & n348 ) | ( x115 & n350 ) | ( n348 & n350 ) ;
  assign n339 = ( x25 & ~x118 ) | ( x25 & n215 ) | ( ~x118 & n215 ) ;
  assign n315 = ( x38 & ~n214 ) | ( x38 & n219 ) | ( ~n214 & n219 ) ;
  assign n316 = ( n195 & n264 ) | ( n195 & ~n315 ) | ( n264 & ~n315 ) ;
  assign n346 = n345 ^ n339 ^ n316 ;
  assign n347 = ( n143 & n274 ) | ( n143 & n346 ) | ( n274 & n346 ) ;
  assign n352 = n351 ^ n347 ^ n152 ;
  assign n353 = ( x65 & n285 ) | ( x65 & n352 ) | ( n285 & n352 ) ;
  assign n354 = ( n203 & n338 ) | ( n203 & ~n353 ) | ( n338 & ~n353 ) ;
  assign n355 = ( ~x67 & x126 ) | ( ~x67 & x127 ) | ( x126 & x127 ) ;
  assign n356 = ( ~x64 & n285 ) | ( ~x64 & n355 ) | ( n285 & n355 ) ;
  assign n358 = n357 ^ n356 ^ n170 ;
  assign n359 = ( x86 & n256 ) | ( x86 & ~n358 ) | ( n256 & ~n358 ) ;
  assign n360 = ( ~n266 & n354 ) | ( ~n266 & n359 ) | ( n354 & n359 ) ;
  assign n361 = ( ~n332 & n336 ) | ( ~n332 & n360 ) | ( n336 & n360 ) ;
  assign n362 = ( n326 & n329 ) | ( n326 & n361 ) | ( n329 & n361 ) ;
  assign n367 = n366 ^ n365 ^ n362 ;
  assign n324 = ( ~x29 & x113 ) | ( ~x29 & n158 ) | ( x113 & n158 ) ;
  assign n309 = n285 ^ n267 ^ x95 ;
  assign n312 = ( x28 & x42 ) | ( x28 & ~n137 ) | ( x42 & ~n137 ) ;
  assign n310 = ( ~x50 & x119 ) | ( ~x50 & n267 ) | ( x119 & n267 ) ;
  assign n311 = ( x89 & n156 ) | ( x89 & ~n310 ) | ( n156 & ~n310 ) ;
  assign n313 = n312 ^ n311 ^ n180 ;
  assign n314 = n313 ^ n288 ^ n247 ;
  assign n317 = n316 ^ n170 ^ x58 ;
  assign n320 = ( x51 & n260 ) | ( x51 & n265 ) | ( n260 & n265 ) ;
  assign n321 = ( ~x0 & n319 ) | ( ~x0 & n320 ) | ( n319 & n320 ) ;
  assign n322 = ( n314 & ~n317 ) | ( n314 & n321 ) | ( ~n317 & n321 ) ;
  assign n323 = ( x102 & ~n309 ) | ( x102 & n322 ) | ( ~n309 & n322 ) ;
  assign n325 = n324 ^ n323 ^ n235 ;
  assign n369 = n368 ^ n367 ^ n325 ;
  assign n401 = n400 ^ n392 ^ n369 ;
  assign n419 = n418 ^ n408 ^ n401 ;
  assign n420 = ( ~x20 & n308 ) | ( ~x20 & n419 ) | ( n308 & n419 ) ;
  assign n430 = n429 ^ n420 ^ n168 ;
  assign n431 = ( n199 & ~n254 ) | ( n199 & n430 ) | ( ~n254 & n430 ) ;
  assign n432 = ( n131 & n245 ) | ( n131 & n431 ) | ( n245 & n431 ) ;
  assign n433 = n327 ^ n320 ^ n311 ;
  assign n434 = n433 ^ n165 ^ x113 ;
  assign n440 = n366 ^ n280 ^ n201 ;
  assign n441 = ( x26 & x38 ) | ( x26 & ~x52 ) | ( x38 & ~x52 ) ;
  assign n442 = ( x6 & n440 ) | ( x6 & n441 ) | ( n440 & n441 ) ;
  assign n436 = ( x65 & n169 ) | ( x65 & n393 ) | ( n169 & n393 ) ;
  assign n437 = ( x127 & n424 ) | ( x127 & n436 ) | ( n424 & n436 ) ;
  assign n438 = ( x69 & n260 ) | ( x69 & ~n437 ) | ( n260 & ~n437 ) ;
  assign n439 = ( ~x102 & n327 ) | ( ~x102 & n438 ) | ( n327 & n438 ) ;
  assign n435 = n380 ^ n183 ^ x36 ;
  assign n443 = n442 ^ n439 ^ n435 ;
  assign n444 = ( x25 & n322 ) | ( x25 & ~n443 ) | ( n322 & ~n443 ) ;
  assign n464 = ( x89 & ~x99 ) | ( x89 & n129 ) | ( ~x99 & n129 ) ;
  assign n460 = ( x6 & n199 ) | ( x6 & n345 ) | ( n199 & n345 ) ;
  assign n461 = n460 ^ n187 ^ x77 ;
  assign n462 = n461 ^ n279 ^ x96 ;
  assign n459 = n161 ^ x97 ^ x65 ;
  assign n456 = ( x56 & x82 ) | ( x56 & n188 ) | ( x82 & n188 ) ;
  assign n454 = ( x3 & n170 ) | ( x3 & ~n171 ) | ( n170 & ~n171 ) ;
  assign n452 = n229 ^ n219 ^ n200 ;
  assign n453 = ( n225 & ~n320 ) | ( n225 & n452 ) | ( ~n320 & n452 ) ;
  assign n455 = n454 ^ n453 ^ n239 ;
  assign n457 = n456 ^ n455 ^ n279 ;
  assign n449 = ( x40 & n319 ) | ( x40 & ~n342 ) | ( n319 & ~n342 ) ;
  assign n445 = ( ~x42 & x93 ) | ( ~x42 & n133 ) | ( x93 & n133 ) ;
  assign n446 = n445 ^ x94 ^ x19 ;
  assign n447 = n446 ^ n139 ^ x101 ;
  assign n448 = ( ~n227 & n345 ) | ( ~n227 & n447 ) | ( n345 & n447 ) ;
  assign n450 = n449 ^ n448 ^ n133 ;
  assign n451 = ( n184 & ~n330 ) | ( n184 & n450 ) | ( ~n330 & n450 ) ;
  assign n458 = n457 ^ n451 ^ n314 ;
  assign n463 = n462 ^ n459 ^ n458 ;
  assign n465 = n464 ^ n463 ^ n273 ;
  assign n466 = ( ~n369 & n444 ) | ( ~n369 & n465 ) | ( n444 & n465 ) ;
  assign n467 = ( ~x127 & n434 ) | ( ~x127 & n466 ) | ( n434 & n466 ) ;
  assign n468 = ( x24 & n250 ) | ( x24 & ~n332 ) | ( n250 & ~n332 ) ;
  assign n469 = ( ~x52 & x111 ) | ( ~x52 & n377 ) | ( x111 & n377 ) ;
  assign n484 = ( x50 & ~x119 ) | ( x50 & n169 ) | ( ~x119 & n169 ) ;
  assign n493 = n484 ^ n162 ^ x56 ;
  assign n494 = ( ~n178 & n192 ) | ( ~n178 & n493 ) | ( n192 & n493 ) ;
  assign n477 = n156 ^ x72 ^ x22 ;
  assign n474 = ( x21 & x57 ) | ( x21 & ~n219 ) | ( x57 & ~n219 ) ;
  assign n475 = n474 ^ n349 ^ x100 ;
  assign n476 = ( n297 & ~n370 ) | ( n297 & n475 ) | ( ~n370 & n475 ) ;
  assign n478 = n477 ^ n476 ^ n186 ;
  assign n485 = n375 ^ n330 ^ n160 ;
  assign n486 = ( n262 & n484 ) | ( n262 & n485 ) | ( n484 & n485 ) ;
  assign n487 = n486 ^ n449 ^ x87 ;
  assign n488 = ( ~n148 & n227 ) | ( ~n148 & n487 ) | ( n227 & n487 ) ;
  assign n489 = ( ~x124 & n255 ) | ( ~x124 & n488 ) | ( n255 & n488 ) ;
  assign n482 = ( x6 & n251 ) | ( x6 & ~n300 ) | ( n251 & ~n300 ) ;
  assign n479 = x68 ^ x29 ^ x23 ;
  assign n480 = n479 ^ x90 ^ x84 ;
  assign n481 = ( n130 & n223 ) | ( n130 & n480 ) | ( n223 & n480 ) ;
  assign n483 = n482 ^ n481 ^ n375 ;
  assign n472 = ( ~x108 & n136 ) | ( ~x108 & n203 ) | ( n136 & n203 ) ;
  assign n490 = n489 ^ n483 ^ n472 ;
  assign n491 = ( x5 & ~n478 ) | ( x5 & n490 ) | ( ~n478 & n490 ) ;
  assign n492 = ( ~x120 & n159 ) | ( ~x120 & n491 ) | ( n159 & n491 ) ;
  assign n470 = n370 ^ x115 ^ x89 ;
  assign n471 = ( ~x109 & n291 ) | ( ~x109 & n470 ) | ( n291 & n470 ) ;
  assign n473 = n472 ^ n471 ^ n324 ;
  assign n495 = n494 ^ n492 ^ n473 ;
  assign n496 = ( x46 & ~n468 ) | ( x46 & n495 ) | ( ~n468 & n495 ) ;
  assign n497 = ( n468 & ~n469 ) | ( n468 & n496 ) | ( ~n469 & n496 ) ;
  assign n498 = ( ~x111 & n467 ) | ( ~x111 & n497 ) | ( n467 & n497 ) ;
  assign n539 = n237 ^ n170 ^ x5 ;
  assign n550 = ( ~n394 & n426 ) | ( ~n394 & n539 ) | ( n426 & n539 ) ;
  assign n565 = n258 ^ x110 ^ x41 ;
  assign n566 = ( ~n358 & n411 ) | ( ~n358 & n565 ) | ( n411 & n565 ) ;
  assign n567 = ( n405 & ~n550 ) | ( n405 & n566 ) | ( ~n550 & n566 ) ;
  assign n576 = n567 ^ n174 ^ x102 ;
  assign n577 = ( n224 & n438 ) | ( n224 & ~n576 ) | ( n438 & ~n576 ) ;
  assign n578 = n577 ^ n454 ^ x30 ;
  assign n588 = ( x65 & ~n162 ) | ( x65 & n184 ) | ( ~n162 & n184 ) ;
  assign n537 = ( n137 & n393 ) | ( n137 & ~n403 ) | ( n393 & ~n403 ) ;
  assign n587 = n537 ^ n206 ^ x101 ;
  assign n557 = x111 ^ x110 ^ x24 ;
  assign n558 = ( ~x22 & x54 ) | ( ~x22 & n258 ) | ( x54 & n258 ) ;
  assign n559 = n558 ^ n486 ^ x40 ;
  assign n560 = ( x68 & ~n178 ) | ( x68 & n559 ) | ( ~n178 & n559 ) ;
  assign n561 = ( x83 & x109 ) | ( x83 & n222 ) | ( x109 & n222 ) ;
  assign n562 = ( n557 & ~n560 ) | ( n557 & n561 ) | ( ~n560 & n561 ) ;
  assign n589 = n588 ^ n587 ^ n562 ;
  assign n590 = ( n224 & ~n423 ) | ( n224 & n589 ) | ( ~n423 & n589 ) ;
  assign n582 = n406 ^ n318 ^ x32 ;
  assign n583 = n582 ^ n154 ^ x43 ;
  assign n580 = n375 ^ x77 ^ x69 ;
  assign n538 = ( x3 & n195 ) | ( x3 & ~n201 ) | ( n195 & ~n201 ) ;
  assign n540 = n539 ^ n538 ^ n240 ;
  assign n579 = ( n141 & n273 ) | ( n141 & n540 ) | ( n273 & n540 ) ;
  assign n581 = n580 ^ n579 ^ n281 ;
  assign n584 = n583 ^ n581 ^ n316 ;
  assign n585 = ( x44 & n142 ) | ( x44 & ~n311 ) | ( n142 & ~n311 ) ;
  assign n586 = ( ~n478 & n584 ) | ( ~n478 & n585 ) | ( n584 & n585 ) ;
  assign n591 = n590 ^ n586 ^ n414 ;
  assign n507 = n360 ^ n260 ^ x42 ;
  assign n508 = ( n219 & n386 ) | ( n219 & ~n507 ) | ( n386 & ~n507 ) ;
  assign n598 = n203 ^ x15 ^ x8 ;
  assign n599 = n598 ^ n538 ^ n159 ;
  assign n596 = ( ~n160 & n169 ) | ( ~n160 & n214 ) | ( n169 & n214 ) ;
  assign n597 = n596 ^ n208 ^ x41 ;
  assign n594 = ( ~x108 & x120 ) | ( ~x108 & n394 ) | ( x120 & n394 ) ;
  assign n593 = ( n138 & ~n187 ) | ( n138 & n343 ) | ( ~n187 & n343 ) ;
  assign n592 = ( x83 & ~n135 ) | ( x83 & n566 ) | ( ~n135 & n566 ) ;
  assign n595 = n594 ^ n593 ^ n592 ;
  assign n600 = n599 ^ n597 ^ n595 ;
  assign n512 = ( n174 & n240 ) | ( n174 & ~n486 ) | ( n240 & ~n486 ) ;
  assign n499 = ( x84 & ~x122 ) | ( x84 & n199 ) | ( ~x122 & n199 ) ;
  assign n601 = n512 ^ n499 ^ x85 ;
  assign n602 = ( n345 & n479 ) | ( n345 & n601 ) | ( n479 & n601 ) ;
  assign n603 = ( ~n508 & n600 ) | ( ~n508 & n602 ) | ( n600 & n602 ) ;
  assign n517 = n474 ^ n256 ^ n158 ;
  assign n518 = ( x79 & n251 ) | ( x79 & ~n517 ) | ( n251 & ~n517 ) ;
  assign n519 = n518 ^ x50 ^ x11 ;
  assign n604 = n603 ^ n519 ^ n341 ;
  assign n605 = ( n578 & n591 ) | ( n578 & n604 ) | ( n591 & n604 ) ;
  assign n529 = ( x2 & ~x104 ) | ( x2 & n184 ) | ( ~x104 & n184 ) ;
  assign n530 = ( x5 & ~n239 ) | ( x5 & n529 ) | ( ~n239 & n529 ) ;
  assign n526 = ( x17 & ~x35 ) | ( x17 & n517 ) | ( ~x35 & n517 ) ;
  assign n521 = n378 ^ n258 ^ x45 ;
  assign n522 = n521 ^ n482 ^ n330 ;
  assign n523 = n522 ^ n411 ^ x19 ;
  assign n516 = ( n256 & n454 ) | ( n256 & ~n485 ) | ( n454 & ~n485 ) ;
  assign n515 = n250 ^ x123 ^ x57 ;
  assign n520 = n519 ^ n516 ^ n515 ;
  assign n524 = n523 ^ n520 ^ n228 ;
  assign n525 = n524 ^ n421 ^ n257 ;
  assign n527 = n526 ^ n525 ^ x60 ;
  assign n513 = n512 ^ n178 ^ x11 ;
  assign n514 = n513 ^ n390 ^ n374 ;
  assign n528 = n527 ^ n514 ^ n230 ;
  assign n505 = ( x31 & ~x112 ) | ( x31 & n493 ) | ( ~x112 & n493 ) ;
  assign n506 = ( n300 & n364 ) | ( n300 & ~n505 ) | ( n364 & ~n505 ) ;
  assign n509 = n508 ^ n506 ^ n428 ;
  assign n510 = n509 ^ n346 ^ n266 ;
  assign n500 = ( x118 & ~n273 ) | ( x118 & n499 ) | ( ~n273 & n499 ) ;
  assign n501 = ( ~x32 & x103 ) | ( ~x32 & n261 ) | ( x103 & n261 ) ;
  assign n502 = ( n289 & n399 ) | ( n289 & n501 ) | ( n399 & n501 ) ;
  assign n503 = ( n220 & n436 ) | ( n220 & ~n502 ) | ( n436 & ~n502 ) ;
  assign n504 = ( ~x0 & n500 ) | ( ~x0 & n503 ) | ( n500 & n503 ) ;
  assign n511 = n510 ^ n504 ^ n264 ;
  assign n531 = n530 ^ n528 ^ n511 ;
  assign n532 = n320 ^ x34 ^ x7 ;
  assign n533 = n532 ^ n350 ^ n176 ;
  assign n534 = ( x19 & ~x117 ) | ( x19 & n263 ) | ( ~x117 & n263 ) ;
  assign n535 = ( n153 & ~n297 ) | ( n153 & n534 ) | ( ~n297 & n534 ) ;
  assign n536 = n535 ^ x104 ^ x65 ;
  assign n541 = n540 ^ n250 ^ n211 ;
  assign n542 = ( ~n391 & n537 ) | ( ~n391 & n541 ) | ( n537 & n541 ) ;
  assign n543 = n542 ^ n377 ^ n206 ;
  assign n544 = ( ~x98 & n202 ) | ( ~x98 & n543 ) | ( n202 & n543 ) ;
  assign n556 = n329 ^ n209 ^ x12 ;
  assign n563 = n562 ^ n556 ^ n294 ;
  assign n568 = ( n288 & n327 ) | ( n288 & n567 ) | ( n327 & n567 ) ;
  assign n564 = ( ~x16 & n362 ) | ( ~x16 & n415 ) | ( n362 & n415 ) ;
  assign n569 = n568 ^ n564 ^ n155 ;
  assign n570 = n569 ^ n299 ^ n289 ;
  assign n571 = ( n399 & ~n563 ) | ( n399 & n570 ) | ( ~n563 & n570 ) ;
  assign n572 = n571 ^ n220 ^ x52 ;
  assign n552 = n246 ^ x27 ^ x2 ;
  assign n549 = n404 ^ n318 ^ n257 ;
  assign n551 = n550 ^ n549 ^ n445 ;
  assign n548 = n517 ^ n264 ^ n166 ;
  assign n553 = n552 ^ n551 ^ n548 ;
  assign n545 = ( ~x40 & n162 ) | ( ~x40 & n298 ) | ( n162 & n298 ) ;
  assign n546 = ( x72 & n213 ) | ( x72 & ~n545 ) | ( n213 & ~n545 ) ;
  assign n547 = ( ~n257 & n440 ) | ( ~n257 & n546 ) | ( n440 & n546 ) ;
  assign n554 = n553 ^ n547 ^ x100 ;
  assign n555 = ( ~n147 & n275 ) | ( ~n147 & n554 ) | ( n275 & n554 ) ;
  assign n573 = n572 ^ n555 ^ n200 ;
  assign n574 = ( n536 & ~n544 ) | ( n536 & n573 ) | ( ~n544 & n573 ) ;
  assign n575 = ( ~n531 & n533 ) | ( ~n531 & n574 ) | ( n533 & n574 ) ;
  assign n606 = n605 ^ n575 ^ n143 ;
  assign n658 = ( n185 & n344 ) | ( n185 & n535 ) | ( n344 & n535 ) ;
  assign n647 = ( x7 & ~n133 ) | ( x7 & n409 ) | ( ~n133 & n409 ) ;
  assign n648 = n647 ^ n477 ^ x35 ;
  assign n649 = n648 ^ n483 ^ n266 ;
  assign n650 = n371 ^ x127 ^ x106 ;
  assign n651 = ( ~x81 & n192 ) | ( ~x81 & n650 ) | ( n192 & n650 ) ;
  assign n652 = ( x39 & x49 ) | ( x39 & ~n651 ) | ( x49 & ~n651 ) ;
  assign n610 = ( ~x99 & n177 ) | ( ~x99 & n338 ) | ( n177 & n338 ) ;
  assign n611 = ( n172 & ~n330 ) | ( n172 & n610 ) | ( ~n330 & n610 ) ;
  assign n612 = n611 ^ n331 ^ x98 ;
  assign n653 = n612 ^ n271 ^ x44 ;
  assign n654 = ( n414 & n652 ) | ( n414 & n653 ) | ( n652 & n653 ) ;
  assign n655 = n654 ^ n324 ^ n139 ;
  assign n656 = n371 ^ n258 ^ n232 ;
  assign n657 = ( n649 & ~n655 ) | ( n649 & n656 ) | ( ~n655 & n656 ) ;
  assign n607 = n132 ^ n130 ^ x63 ;
  assign n608 = ( x49 & ~n222 ) | ( x49 & n607 ) | ( ~n222 & n607 ) ;
  assign n616 = n257 ^ x111 ^ x97 ;
  assign n617 = n616 ^ n177 ^ x125 ;
  assign n618 = n617 ^ n520 ^ x29 ;
  assign n619 = n618 ^ n370 ^ n153 ;
  assign n615 = ( n324 & ~n526 ) | ( n324 & n597 ) | ( ~n526 & n597 ) ;
  assign n620 = n619 ^ n615 ^ n270 ;
  assign n609 = n295 ^ n151 ^ x52 ;
  assign n613 = ( ~n198 & n335 ) | ( ~n198 & n612 ) | ( n335 & n612 ) ;
  assign n614 = ( n330 & ~n609 ) | ( n330 & n613 ) | ( ~n609 & n613 ) ;
  assign n621 = n620 ^ n614 ^ n440 ;
  assign n622 = ( ~n240 & n344 ) | ( ~n240 & n621 ) | ( n344 & n621 ) ;
  assign n623 = ( n441 & n608 ) | ( n441 & n622 ) | ( n608 & n622 ) ;
  assign n624 = ( x20 & n259 ) | ( x20 & ~n371 ) | ( n259 & ~n371 ) ;
  assign n625 = n624 ^ n373 ^ x120 ;
  assign n626 = ( ~x45 & n348 ) | ( ~x45 & n625 ) | ( n348 & n625 ) ;
  assign n627 = n626 ^ n507 ^ n364 ;
  assign n628 = ( n133 & n608 ) | ( n133 & n627 ) | ( n608 & n627 ) ;
  assign n644 = n197 ^ n149 ^ x108 ;
  assign n642 = ( ~n182 & n256 ) | ( ~n182 & n355 ) | ( n256 & n355 ) ;
  assign n643 = n642 ^ x126 ^ x62 ;
  assign n629 = n449 ^ n326 ^ n166 ;
  assign n630 = n629 ^ n204 ^ x4 ;
  assign n631 = n214 ^ x21 ^ x5 ;
  assign n632 = ( x54 & n277 ) | ( x54 & n471 ) | ( n277 & n471 ) ;
  assign n633 = ( x113 & n346 ) | ( x113 & n632 ) | ( n346 & n632 ) ;
  assign n635 = ( ~n247 & n341 ) | ( ~n247 & n440 ) | ( n341 & n440 ) ;
  assign n636 = n635 ^ n251 ^ x95 ;
  assign n634 = n624 ^ n222 ^ x70 ;
  assign n637 = n636 ^ n634 ^ n323 ;
  assign n638 = ( n465 & ~n513 ) | ( n465 & n637 ) | ( ~n513 & n637 ) ;
  assign n639 = ( ~n241 & n633 ) | ( ~n241 & n638 ) | ( n633 & n638 ) ;
  assign n640 = ( n630 & n631 ) | ( n630 & ~n639 ) | ( n631 & ~n639 ) ;
  assign n641 = n640 ^ n495 ^ n330 ;
  assign n645 = n644 ^ n643 ^ n641 ;
  assign n646 = ( n623 & ~n628 ) | ( n623 & n645 ) | ( ~n628 & n645 ) ;
  assign n659 = n658 ^ n657 ^ n646 ;
  assign n660 = ( x103 & n248 ) | ( x103 & ~n253 ) | ( n248 & ~n253 ) ;
  assign n661 = n154 ^ x18 ^ x9 ;
  assign n662 = n661 ^ n438 ^ n260 ;
  assign n680 = ( x82 & x124 ) | ( x82 & n557 ) | ( x124 & n557 ) ;
  assign n681 = ( x65 & x110 ) | ( x65 & ~n680 ) | ( x110 & ~n680 ) ;
  assign n669 = ( n137 & n332 ) | ( n137 & ~n517 ) | ( n332 & ~n517 ) ;
  assign n679 = ( x28 & ~n211 ) | ( x28 & n669 ) | ( ~n211 & n669 ) ;
  assign n675 = n157 ^ x109 ^ x87 ;
  assign n676 = ( ~n276 & n334 ) | ( ~n276 & n675 ) | ( n334 & n675 ) ;
  assign n670 = ( n271 & n480 ) | ( n271 & n669 ) | ( n480 & n669 ) ;
  assign n671 = ( n165 & ~n250 ) | ( n165 & n670 ) | ( ~n250 & n670 ) ;
  assign n667 = ( ~x52 & x53 ) | ( ~x52 & n216 ) | ( x53 & n216 ) ;
  assign n666 = ( ~x25 & x50 ) | ( ~x25 & n261 ) | ( x50 & n261 ) ;
  assign n668 = n667 ^ n666 ^ x25 ;
  assign n672 = n671 ^ n668 ^ n144 ;
  assign n673 = n672 ^ n631 ^ n459 ;
  assign n665 = n595 ^ n457 ^ n292 ;
  assign n663 = n371 ^ n343 ^ n147 ;
  assign n664 = n663 ^ x102 ^ x9 ;
  assign n674 = n673 ^ n665 ^ n664 ;
  assign n677 = n676 ^ n674 ^ x77 ;
  assign n678 = ( ~x92 & n146 ) | ( ~x92 & n677 ) | ( n146 & n677 ) ;
  assign n682 = n681 ^ n679 ^ n678 ;
  assign n683 = ( x115 & n572 ) | ( x115 & ~n682 ) | ( n572 & ~n682 ) ;
  assign n684 = ( ~x97 & n176 ) | ( ~x97 & n185 ) | ( n176 & n185 ) ;
  assign n685 = n684 ^ n643 ^ n487 ;
  assign n686 = ( x118 & n370 ) | ( x118 & n685 ) | ( n370 & n685 ) ;
  assign n687 = ( x5 & n433 ) | ( x5 & ~n686 ) | ( n433 & ~n686 ) ;
  assign n688 = ( ~n662 & n683 ) | ( ~n662 & n687 ) | ( n683 & n687 ) ;
  assign n689 = ( ~n443 & n660 ) | ( ~n443 & n688 ) | ( n660 & n688 ) ;
  assign n841 = ( ~x109 & n274 ) | ( ~x109 & n488 ) | ( n274 & n488 ) ;
  assign n842 = n841 ^ n414 ^ n312 ;
  assign n827 = ( x68 & x110 ) | ( x68 & ~n315 ) | ( x110 & ~n315 ) ;
  assign n828 = ( ~n281 & n319 ) | ( ~n281 & n827 ) | ( n319 & n827 ) ;
  assign n838 = n234 ^ n152 ^ x30 ;
  assign n806 = n485 ^ n374 ^ x92 ;
  assign n759 = n624 ^ n484 ^ n226 ;
  assign n829 = n806 ^ n759 ^ x77 ;
  assign n830 = ( ~x51 & n469 ) | ( ~x51 & n829 ) | ( n469 & n829 ) ;
  assign n831 = ( x108 & n205 ) | ( x108 & n213 ) | ( n205 & n213 ) ;
  assign n701 = ( ~x35 & n276 ) | ( ~x35 & n474 ) | ( n276 & n474 ) ;
  assign n702 = n701 ^ n130 ^ x95 ;
  assign n832 = n831 ^ n702 ^ x7 ;
  assign n833 = ( n304 & n610 ) | ( n304 & n832 ) | ( n610 & n832 ) ;
  assign n834 = n211 ^ n146 ^ x97 ;
  assign n835 = n834 ^ n329 ^ n190 ;
  assign n713 = ( ~x30 & x88 ) | ( ~x30 & n198 ) | ( x88 & n198 ) ;
  assign n714 = ( ~x88 & n294 ) | ( ~x88 & n713 ) | ( n294 & n713 ) ;
  assign n836 = n835 ^ n714 ^ x105 ;
  assign n837 = ( ~n830 & n833 ) | ( ~n830 & n836 ) | ( n833 & n836 ) ;
  assign n839 = n838 ^ n837 ^ n650 ;
  assign n840 = ( n188 & n828 ) | ( n188 & n839 ) | ( n828 & n839 ) ;
  assign n703 = n702 ^ n333 ^ n154 ;
  assign n704 = n703 ^ n207 ^ x4 ;
  assign n705 = n704 ^ n242 ^ x124 ;
  assign n706 = n705 ^ n537 ^ n490 ;
  assign n698 = ( x113 & n161 ) | ( x113 & n600 ) | ( n161 & n600 ) ;
  assign n696 = ( n165 & n296 ) | ( n165 & ~n562 ) | ( n296 & ~n562 ) ;
  assign n697 = n696 ^ n335 ^ x20 ;
  assign n699 = n698 ^ n697 ^ n598 ;
  assign n690 = ( x20 & ~x125 ) | ( x20 & n374 ) | ( ~x125 & n374 ) ;
  assign n691 = ( ~n252 & n379 ) | ( ~n252 & n690 ) | ( n379 & n690 ) ;
  assign n692 = n691 ^ n526 ^ x80 ;
  assign n693 = n317 ^ n175 ^ x33 ;
  assign n694 = ( n414 & n439 ) | ( n414 & n693 ) | ( n439 & n693 ) ;
  assign n695 = ( n393 & n692 ) | ( n393 & n694 ) | ( n692 & n694 ) ;
  assign n700 = n699 ^ n695 ^ x111 ;
  assign n707 = n706 ^ n700 ^ n351 ;
  assign n744 = ( x99 & n333 ) | ( x99 & n636 ) | ( n333 & n636 ) ;
  assign n745 = n192 ^ n178 ^ x121 ;
  assign n746 = ( n213 & ~n561 ) | ( n213 & n745 ) | ( ~n561 & n745 ) ;
  assign n747 = ( n224 & n653 ) | ( n224 & ~n746 ) | ( n653 & ~n746 ) ;
  assign n748 = ( n514 & ~n744 ) | ( n514 & n747 ) | ( ~n744 & n747 ) ;
  assign n719 = ( x71 & n147 ) | ( x71 & ~n442 ) | ( n147 & ~n442 ) ;
  assign n715 = ( x59 & ~x62 ) | ( x59 & x97 ) | ( ~x62 & x97 ) ;
  assign n716 = ( n337 & ~n460 ) | ( n337 & n715 ) | ( ~n460 & n715 ) ;
  assign n717 = ( n650 & n714 ) | ( n650 & ~n716 ) | ( n714 & ~n716 ) ;
  assign n711 = ( n134 & n168 ) | ( n134 & n494 ) | ( n168 & n494 ) ;
  assign n708 = ( x56 & n256 ) | ( x56 & ~n296 ) | ( n256 & ~n296 ) ;
  assign n709 = ( n335 & ~n437 ) | ( n335 & n558 ) | ( ~n437 & n558 ) ;
  assign n710 = ( x9 & n708 ) | ( x9 & ~n709 ) | ( n708 & ~n709 ) ;
  assign n712 = n711 ^ n710 ^ n239 ;
  assign n718 = n717 ^ n712 ^ n440 ;
  assign n720 = n719 ^ n718 ^ x31 ;
  assign n726 = n557 ^ n187 ^ n156 ;
  assign n727 = ( x95 & n377 ) | ( x95 & ~n726 ) | ( n377 & ~n726 ) ;
  assign n723 = ( x42 & x64 ) | ( x42 & n133 ) | ( x64 & n133 ) ;
  assign n721 = n680 ^ n371 ^ n310 ;
  assign n722 = ( n383 & n433 ) | ( n383 & ~n721 ) | ( n433 & ~n721 ) ;
  assign n724 = n723 ^ n722 ^ n288 ;
  assign n725 = ( x9 & ~x107 ) | ( x9 & n724 ) | ( ~x107 & n724 ) ;
  assign n728 = n727 ^ n725 ^ x4 ;
  assign n729 = ( n317 & n630 ) | ( n317 & n728 ) | ( n630 & n728 ) ;
  assign n730 = ( ~x69 & n720 ) | ( ~x69 & n729 ) | ( n720 & n729 ) ;
  assign n741 = ( n363 & n478 ) | ( n363 & ~n549 ) | ( n478 & ~n549 ) ;
  assign n731 = ( ~n139 & n214 ) | ( ~n139 & n518 ) | ( n214 & n518 ) ;
  assign n732 = n201 ^ x83 ^ x36 ;
  assign n733 = n357 ^ x67 ^ x56 ;
  assign n734 = ( n400 & ~n506 ) | ( n400 & n733 ) | ( ~n506 & n733 ) ;
  assign n735 = n266 ^ n213 ^ x7 ;
  assign n736 = n735 ^ n437 ^ n348 ;
  assign n737 = ( ~n732 & n734 ) | ( ~n732 & n736 ) | ( n734 & n736 ) ;
  assign n738 = ( n399 & n663 ) | ( n399 & ~n737 ) | ( n663 & ~n737 ) ;
  assign n739 = ( n394 & ~n731 ) | ( n394 & n738 ) | ( ~n731 & n738 ) ;
  assign n740 = n739 ^ n558 ^ x13 ;
  assign n742 = n741 ^ n740 ^ n160 ;
  assign n743 = ( ~n616 & n730 ) | ( ~n616 & n742 ) | ( n730 & n742 ) ;
  assign n749 = n748 ^ n743 ^ n158 ;
  assign n751 = ( x72 & ~x114 ) | ( x72 & n264 ) | ( ~x114 & n264 ) ;
  assign n750 = n537 ^ n331 ^ n251 ;
  assign n752 = n751 ^ n750 ^ n307 ;
  assign n753 = ( x69 & ~n384 ) | ( x69 & n594 ) | ( ~n384 & n594 ) ;
  assign n754 = n753 ^ x114 ^ x63 ;
  assign n755 = n754 ^ n691 ^ x117 ;
  assign n756 = n576 ^ n225 ^ n146 ;
  assign n757 = n756 ^ n717 ^ x126 ;
  assign n758 = ( x60 & n755 ) | ( x60 & ~n757 ) | ( n755 & ~n757 ) ;
  assign n760 = n171 ^ n145 ^ x49 ;
  assign n761 = ( ~n501 & n759 ) | ( ~n501 & n760 ) | ( n759 & n760 ) ;
  assign n766 = ( ~x29 & x108 ) | ( ~x29 & n220 ) | ( x108 & n220 ) ;
  assign n767 = n766 ^ n175 ^ n137 ;
  assign n768 = ( n182 & n257 ) | ( n182 & ~n767 ) | ( n257 & ~n767 ) ;
  assign n769 = ( n265 & n286 ) | ( n265 & n732 ) | ( n286 & n732 ) ;
  assign n770 = ( n290 & n768 ) | ( n290 & ~n769 ) | ( n768 & ~n769 ) ;
  assign n762 = n558 ^ n147 ^ x37 ;
  assign n763 = ( ~n148 & n186 ) | ( ~n148 & n762 ) | ( n186 & n762 ) ;
  assign n764 = n763 ^ n634 ^ n336 ;
  assign n765 = ( n156 & ~n167 ) | ( n156 & n764 ) | ( ~n167 & n764 ) ;
  assign n771 = n770 ^ n765 ^ n449 ;
  assign n772 = ( n732 & ~n761 ) | ( n732 & n771 ) | ( ~n761 & n771 ) ;
  assign n773 = ( n752 & ~n758 ) | ( n752 & n772 ) | ( ~n758 & n772 ) ;
  assign n777 = n302 ^ n281 ^ x77 ;
  assign n774 = ( ~x41 & x105 ) | ( ~x41 & n146 ) | ( x105 & n146 ) ;
  assign n775 = ( n360 & ~n698 ) | ( n360 & n774 ) | ( ~n698 & n774 ) ;
  assign n776 = n775 ^ n421 ^ n305 ;
  assign n778 = n777 ^ n776 ^ n315 ;
  assign n779 = ( x55 & n370 ) | ( x55 & n778 ) | ( n370 & n778 ) ;
  assign n802 = ( x22 & n352 ) | ( x22 & ~n409 ) | ( n352 & ~n409 ) ;
  assign n800 = n517 ^ n433 ^ n138 ;
  assign n795 = ( ~x49 & x50 ) | ( ~x49 & n474 ) | ( x50 & n474 ) ;
  assign n796 = ( ~n210 & n211 ) | ( ~n210 & n795 ) | ( n211 & n795 ) ;
  assign n797 = n493 ^ n273 ^ x84 ;
  assign n798 = ( n158 & n327 ) | ( n158 & n797 ) | ( n327 & n797 ) ;
  assign n799 = ( n624 & n796 ) | ( n624 & ~n798 ) | ( n796 & ~n798 ) ;
  assign n801 = n800 ^ n799 ^ n247 ;
  assign n780 = n196 ^ x78 ^ x38 ;
  assign n781 = n780 ^ n759 ^ x121 ;
  assign n782 = n440 ^ n144 ^ x55 ;
  assign n783 = ( ~x80 & n335 ) | ( ~x80 & n782 ) | ( n335 & n782 ) ;
  assign n784 = n783 ^ n471 ^ x37 ;
  assign n785 = n281 ^ x99 ^ x25 ;
  assign n786 = n452 ^ n393 ^ x21 ;
  assign n787 = n786 ^ n539 ^ n403 ;
  assign n788 = ( ~n294 & n785 ) | ( ~n294 & n787 ) | ( n785 & n787 ) ;
  assign n790 = n413 ^ n162 ^ x97 ;
  assign n789 = ( x105 & ~n594 ) | ( x105 & n602 ) | ( ~n594 & n602 ) ;
  assign n791 = n790 ^ n789 ^ n179 ;
  assign n792 = n791 ^ n412 ^ n353 ;
  assign n793 = ( n784 & n788 ) | ( n784 & n792 ) | ( n788 & n792 ) ;
  assign n794 = ( ~n243 & n781 ) | ( ~n243 & n793 ) | ( n781 & n793 ) ;
  assign n803 = n802 ^ n801 ^ n794 ;
  assign n820 = n680 ^ n441 ^ x45 ;
  assign n821 = ( x56 & n766 ) | ( x56 & n820 ) | ( n766 & n820 ) ;
  assign n819 = ( x126 & n132 ) | ( x126 & ~n341 ) | ( n132 & ~n341 ) ;
  assign n822 = n821 ^ n819 ^ n651 ;
  assign n816 = x91 ^ x35 ^ x22 ;
  assign n817 = ( x21 & n414 ) | ( x21 & n816 ) | ( n414 & n816 ) ;
  assign n818 = n817 ^ n698 ^ n538 ;
  assign n804 = ( ~x50 & n298 ) | ( ~x50 & n378 ) | ( n298 & n378 ) ;
  assign n805 = ( x120 & n460 ) | ( x120 & n804 ) | ( n460 & n804 ) ;
  assign n809 = ( n251 & ~n350 ) | ( n251 & n379 ) | ( ~n350 & n379 ) ;
  assign n807 = n806 ^ n350 ^ n199 ;
  assign n808 = n807 ^ n703 ^ n133 ;
  assign n810 = n809 ^ n808 ^ n713 ;
  assign n811 = n321 ^ n225 ^ x50 ;
  assign n812 = n703 ^ n158 ^ x45 ;
  assign n813 = n812 ^ n206 ^ x39 ;
  assign n814 = ( ~n810 & n811 ) | ( ~n810 & n813 ) | ( n811 & n813 ) ;
  assign n815 = ( n592 & n805 ) | ( n592 & n814 ) | ( n805 & n814 ) ;
  assign n823 = n822 ^ n818 ^ n815 ;
  assign n824 = ( n489 & n803 ) | ( n489 & ~n823 ) | ( n803 & ~n823 ) ;
  assign n825 = ( n773 & ~n779 ) | ( n773 & n824 ) | ( ~n779 & n824 ) ;
  assign n826 = ( n707 & n749 ) | ( n707 & n825 ) | ( n749 & n825 ) ;
  assign n843 = n842 ^ n840 ^ n826 ;
  assign n905 = n499 ^ x58 ^ x38 ;
  assign n899 = n650 ^ x34 ^ x20 ;
  assign n900 = ( ~n425 & n690 ) | ( ~n425 & n899 ) | ( n690 & n899 ) ;
  assign n901 = ( n143 & n405 ) | ( n143 & n900 ) | ( n405 & n900 ) ;
  assign n902 = n901 ^ n194 ^ x8 ;
  assign n903 = n902 ^ n617 ^ n153 ;
  assign n879 = ( n264 & ~n270 ) | ( n264 & n273 ) | ( ~n270 & n273 ) ;
  assign n848 = ( ~x28 & x95 ) | ( ~x28 & n237 ) | ( x95 & n237 ) ;
  assign n880 = n879 ^ n848 ^ x26 ;
  assign n881 = ( x55 & x100 ) | ( x55 & n880 ) | ( x100 & n880 ) ;
  assign n875 = ( ~x118 & n268 ) | ( ~x118 & n344 ) | ( n268 & n344 ) ;
  assign n876 = n875 ^ n478 ^ n289 ;
  assign n877 = n876 ^ n398 ^ x24 ;
  assign n878 = n877 ^ n759 ^ n365 ;
  assign n882 = n881 ^ n878 ^ n425 ;
  assign n886 = n345 ^ n213 ^ x96 ;
  assign n887 = ( n382 & ~n732 ) | ( n382 & n886 ) | ( ~n732 & n886 ) ;
  assign n888 = n887 ^ n426 ^ n309 ;
  assign n883 = ( ~x20 & n223 ) | ( ~x20 & n493 ) | ( n223 & n493 ) ;
  assign n884 = ( ~n469 & n483 ) | ( ~n469 & n883 ) | ( n483 & n883 ) ;
  assign n844 = n345 ^ n231 ^ x65 ;
  assign n845 = n844 ^ n643 ^ n454 ;
  assign n846 = n845 ^ n620 ^ x14 ;
  assign n847 = ( n233 & n235 ) | ( n233 & n846 ) | ( n235 & n846 ) ;
  assign n885 = n884 ^ n883 ^ n847 ;
  assign n889 = n888 ^ n885 ^ n833 ;
  assign n890 = n889 ^ n531 ^ n491 ;
  assign n891 = n289 ^ n268 ^ x70 ;
  assign n892 = ( ~n331 & n620 ) | ( ~n331 & n891 ) | ( n620 & n891 ) ;
  assign n893 = ( n261 & n454 ) | ( n261 & n892 ) | ( n454 & n892 ) ;
  assign n894 = n546 ^ n384 ^ x101 ;
  assign n895 = n894 ^ n512 ^ n424 ;
  assign n896 = n895 ^ n668 ^ n617 ;
  assign n897 = ( n181 & n893 ) | ( n181 & ~n896 ) | ( n893 & ~n896 ) ;
  assign n898 = ( n882 & ~n890 ) | ( n882 & n897 ) | ( ~n890 & n897 ) ;
  assign n863 = ( n410 & n672 ) | ( n410 & n727 ) | ( n672 & n727 ) ;
  assign n859 = n831 ^ x82 ^ x37 ;
  assign n860 = n611 ^ n265 ^ n148 ;
  assign n861 = n860 ^ n637 ^ n257 ;
  assign n862 = ( n213 & n859 ) | ( n213 & ~n861 ) | ( n859 & ~n861 ) ;
  assign n856 = n426 ^ n395 ^ x44 ;
  assign n857 = ( n208 & n595 ) | ( n208 & ~n856 ) | ( n595 & ~n856 ) ;
  assign n854 = ( n326 & ~n516 ) | ( n326 & n766 ) | ( ~n516 & n766 ) ;
  assign n855 = n854 ^ n828 ^ n277 ;
  assign n858 = n857 ^ n855 ^ n136 ;
  assign n864 = n863 ^ n862 ^ n858 ;
  assign n865 = ( n391 & n734 ) | ( n391 & n864 ) | ( n734 & n864 ) ;
  assign n866 = n623 ^ n318 ^ n285 ;
  assign n867 = ( ~x118 & n353 ) | ( ~x118 & n629 ) | ( n353 & n629 ) ;
  assign n868 = ( ~n351 & n638 ) | ( ~n351 & n867 ) | ( n638 & n867 ) ;
  assign n869 = n562 ^ n427 ^ n197 ;
  assign n870 = ( x60 & ~x65 ) | ( x60 & n522 ) | ( ~x65 & n522 ) ;
  assign n871 = n870 ^ n725 ^ n268 ;
  assign n872 = ( n176 & ~n869 ) | ( n176 & n871 ) | ( ~n869 & n871 ) ;
  assign n873 = ( n866 & n868 ) | ( n866 & ~n872 ) | ( n868 & ~n872 ) ;
  assign n874 = ( n156 & n865 ) | ( n156 & n873 ) | ( n865 & n873 ) ;
  assign n904 = n903 ^ n898 ^ n874 ;
  assign n849 = n848 ^ n506 ^ n205 ;
  assign n850 = ( n217 & n237 ) | ( n217 & ~n398 ) | ( n237 & ~n398 ) ;
  assign n851 = n850 ^ x88 ^ x2 ;
  assign n852 = n851 ^ n559 ^ n512 ;
  assign n853 = ( n847 & n849 ) | ( n847 & ~n852 ) | ( n849 & ~n852 ) ;
  assign n906 = n905 ^ n904 ^ n853 ;
  assign n907 = ( n219 & n348 ) | ( n219 & ~n532 ) | ( n348 & ~n532 ) ;
  assign n908 = ( x111 & n800 ) | ( x111 & ~n907 ) | ( n800 & ~n907 ) ;
  assign n909 = ( n577 & n796 ) | ( n577 & ~n908 ) | ( n796 & ~n908 ) ;
  assign n910 = ( x88 & n577 ) | ( x88 & n909 ) | ( n577 & n909 ) ;
  assign n928 = ( x93 & ~x125 ) | ( x93 & n253 ) | ( ~x125 & n253 ) ;
  assign n926 = ( x15 & n197 ) | ( x15 & ~n241 ) | ( n197 & ~n241 ) ;
  assign n920 = ( ~x13 & x92 ) | ( ~x13 & n582 ) | ( x92 & n582 ) ;
  assign n921 = ( x32 & n326 ) | ( x32 & ~n812 ) | ( n326 & ~n812 ) ;
  assign n922 = ( x97 & n875 ) | ( x97 & ~n921 ) | ( n875 & ~n921 ) ;
  assign n923 = ( n745 & n920 ) | ( n745 & ~n922 ) | ( n920 & ~n922 ) ;
  assign n924 = ( n252 & n670 ) | ( n252 & ~n923 ) | ( n670 & ~n923 ) ;
  assign n925 = ( n188 & ~n450 ) | ( n188 & n924 ) | ( ~n450 & n924 ) ;
  assign n927 = n926 ^ n925 ^ n635 ;
  assign n911 = ( n176 & n259 ) | ( n176 & ~n519 ) | ( n259 & ~n519 ) ;
  assign n912 = n222 ^ n220 ^ x65 ;
  assign n913 = n847 ^ n505 ^ x80 ;
  assign n914 = ( ~x25 & n912 ) | ( ~x25 & n913 ) | ( n912 & n913 ) ;
  assign n915 = ( x11 & ~n137 ) | ( x11 & n151 ) | ( ~n137 & n151 ) ;
  assign n916 = n915 ^ n521 ^ n312 ;
  assign n917 = ( n437 & ~n540 ) | ( n437 & n916 ) | ( ~n540 & n916 ) ;
  assign n918 = n917 ^ n886 ^ n466 ;
  assign n919 = ( n911 & n914 ) | ( n911 & n918 ) | ( n914 & n918 ) ;
  assign n929 = n928 ^ n927 ^ n919 ;
  assign n930 = ( n906 & n910 ) | ( n906 & ~n929 ) | ( n910 & ~n929 ) ;
  assign n1037 = ( x58 & x65 ) | ( x58 & ~n410 ) | ( x65 & ~n410 ) ;
  assign n958 = ( x22 & n138 ) | ( x22 & n675 ) | ( n138 & n675 ) ;
  assign n979 = n958 ^ n374 ^ x37 ;
  assign n980 = n979 ^ n730 ^ n221 ;
  assign n986 = n690 ^ n494 ^ x111 ;
  assign n987 = n986 ^ n263 ^ x41 ;
  assign n988 = ( x58 & n405 ) | ( x58 & n598 ) | ( n405 & n598 ) ;
  assign n989 = n988 ^ n726 ^ n134 ;
  assign n990 = n989 ^ n768 ^ n260 ;
  assign n991 = n881 ^ n508 ^ x113 ;
  assign n992 = ( n987 & n990 ) | ( n987 & n991 ) | ( n990 & n991 ) ;
  assign n950 = n273 ^ n187 ^ x122 ;
  assign n981 = ( n264 & ~n475 ) | ( n264 & n950 ) | ( ~n475 & n950 ) ;
  assign n982 = n471 ^ n357 ^ n253 ;
  assign n983 = ( x21 & x35 ) | ( x21 & ~n982 ) | ( x35 & ~n982 ) ;
  assign n984 = ( x81 & x126 ) | ( x81 & ~n983 ) | ( x126 & ~n983 ) ;
  assign n985 = ( ~n641 & n981 ) | ( ~n641 & n984 ) | ( n981 & n984 ) ;
  assign n993 = n992 ^ n985 ^ n786 ;
  assign n994 = ( n395 & ~n881 ) | ( n395 & n907 ) | ( ~n881 & n907 ) ;
  assign n995 = n543 ^ n426 ^ n273 ;
  assign n996 = ( n459 & ~n994 ) | ( n459 & n995 ) | ( ~n994 & n995 ) ;
  assign n997 = ( ~n368 & n563 ) | ( ~n368 & n996 ) | ( n563 & n996 ) ;
  assign n1006 = n691 ^ n469 ^ n375 ;
  assign n1007 = n1006 ^ n386 ^ n173 ;
  assign n1008 = n1007 ^ n487 ^ x81 ;
  assign n1002 = ( x11 & x26 ) | ( x11 & n768 ) | ( x26 & n768 ) ;
  assign n941 = ( n279 & ~n335 ) | ( n279 & n538 ) | ( ~n335 & n538 ) ;
  assign n998 = ( x11 & ~n480 ) | ( x11 & n941 ) | ( ~n480 & n941 ) ;
  assign n999 = ( ~x103 & n340 ) | ( ~x103 & n411 ) | ( n340 & n411 ) ;
  assign n1000 = ( n242 & n998 ) | ( n242 & n999 ) | ( n998 & n999 ) ;
  assign n1001 = n1000 ^ n861 ^ n317 ;
  assign n1003 = n1002 ^ n1001 ^ n521 ;
  assign n1004 = ( n468 & ~n503 ) | ( n468 & n758 ) | ( ~n503 & n758 ) ;
  assign n1005 = ( n802 & n1003 ) | ( n802 & n1004 ) | ( n1003 & n1004 ) ;
  assign n1009 = n1008 ^ n1005 ^ n543 ;
  assign n1028 = ( x48 & x55 ) | ( x48 & n290 ) | ( x55 & n290 ) ;
  assign n1026 = n723 ^ n424 ^ n143 ;
  assign n1027 = ( x47 & n337 ) | ( x47 & n1026 ) | ( n337 & n1026 ) ;
  assign n1024 = ( ~x125 & n395 ) | ( ~x125 & n702 ) | ( n395 & n702 ) ;
  assign n1020 = n532 ^ n396 ^ n345 ;
  assign n1021 = n1020 ^ n737 ^ n541 ;
  assign n1022 = ( ~x115 & n296 ) | ( ~x115 & n1021 ) | ( n296 & n1021 ) ;
  assign n1023 = ( ~n389 & n427 ) | ( ~n389 & n1022 ) | ( n427 & n1022 ) ;
  assign n1025 = n1024 ^ n1023 ^ n411 ;
  assign n1029 = n1028 ^ n1027 ^ n1025 ;
  assign n951 = ( x54 & n136 ) | ( x54 & n594 ) | ( n136 & n594 ) ;
  assign n952 = ( x99 & n609 ) | ( x99 & ~n951 ) | ( n609 & ~n951 ) ;
  assign n953 = n409 ^ n196 ^ x12 ;
  assign n954 = ( n409 & n952 ) | ( n409 & ~n953 ) | ( n952 & ~n953 ) ;
  assign n1010 = ( x24 & x76 ) | ( x24 & ~n954 ) | ( x76 & ~n954 ) ;
  assign n1011 = n1010 ^ n459 ^ n175 ;
  assign n931 = n921 ^ n524 ^ n226 ;
  assign n1017 = n931 ^ n510 ^ n283 ;
  assign n1013 = ( ~n144 & n301 ) | ( ~n144 & n539 ) | ( n301 & n539 ) ;
  assign n1014 = ( n176 & n350 ) | ( n176 & n1013 ) | ( n350 & n1013 ) ;
  assign n1015 = ( ~n483 & n951 ) | ( ~n483 & n1014 ) | ( n951 & n1014 ) ;
  assign n1012 = n621 ^ n305 ^ x103 ;
  assign n1016 = n1015 ^ n1012 ^ x11 ;
  assign n1018 = n1017 ^ n1016 ^ n767 ;
  assign n1019 = ( x119 & ~n1011 ) | ( x119 & n1018 ) | ( ~n1011 & n1018 ) ;
  assign n1030 = n1029 ^ n1019 ^ x54 ;
  assign n1031 = ( x52 & n157 ) | ( x52 & n412 ) | ( n157 & n412 ) ;
  assign n1032 = n1012 ^ n720 ^ n339 ;
  assign n1033 = ( n673 & n1031 ) | ( n673 & n1032 ) | ( n1031 & n1032 ) ;
  assign n1034 = ( n950 & n1030 ) | ( n950 & n1033 ) | ( n1030 & n1033 ) ;
  assign n1035 = ( n997 & n1009 ) | ( n997 & n1034 ) | ( n1009 & n1034 ) ;
  assign n1036 = ( ~n980 & n993 ) | ( ~n980 & n1035 ) | ( n993 & n1035 ) ;
  assign n932 = n931 ^ n720 ^ n590 ;
  assign n933 = ( ~n347 & n553 ) | ( ~n347 & n932 ) | ( n553 & n932 ) ;
  assign n936 = n252 ^ n247 ^ n160 ;
  assign n934 = n487 ^ n455 ^ x78 ;
  assign n935 = n934 ^ n631 ^ n491 ;
  assign n937 = n936 ^ n935 ^ n787 ;
  assign n938 = n607 ^ n313 ^ x89 ;
  assign n939 = n592 ^ n507 ^ n286 ;
  assign n940 = n939 ^ n589 ^ n405 ;
  assign n943 = ( n224 & ~n350 ) | ( n224 & n543 ) | ( ~n350 & n543 ) ;
  assign n942 = n252 ^ n228 ^ x21 ;
  assign n944 = n943 ^ n942 ^ n370 ;
  assign n945 = ( ~x80 & n170 ) | ( ~x80 & n944 ) | ( n170 & n944 ) ;
  assign n946 = ( n338 & n725 ) | ( n338 & n920 ) | ( n725 & n920 ) ;
  assign n947 = ( n941 & n945 ) | ( n941 & n946 ) | ( n945 & n946 ) ;
  assign n948 = ( ~n938 & n940 ) | ( ~n938 & n947 ) | ( n940 & n947 ) ;
  assign n949 = ( n837 & ~n937 ) | ( n837 & n948 ) | ( ~n937 & n948 ) ;
  assign n975 = n733 ^ x97 ^ x59 ;
  assign n976 = ( n205 & ~n848 ) | ( n205 & n975 ) | ( ~n848 & n975 ) ;
  assign n973 = n396 ^ n131 ^ x103 ;
  assign n971 = ( n298 & ~n428 ) | ( n298 & n517 ) | ( ~n428 & n517 ) ;
  assign n972 = n971 ^ n774 ^ n132 ;
  assign n967 = ( x42 & n188 ) | ( x42 & n252 ) | ( n188 & n252 ) ;
  assign n968 = n967 ^ n642 ^ n394 ;
  assign n969 = ( n171 & ~n509 ) | ( n171 & n968 ) | ( ~n509 & n968 ) ;
  assign n970 = ( x87 & n541 ) | ( x87 & ~n969 ) | ( n541 & ~n969 ) ;
  assign n974 = n973 ^ n972 ^ n970 ;
  assign n955 = n954 ^ n635 ^ x32 ;
  assign n956 = ( n635 & n950 ) | ( n635 & n955 ) | ( n950 & n955 ) ;
  assign n957 = ( n184 & n286 ) | ( n184 & n296 ) | ( n286 & n296 ) ;
  assign n959 = n958 ^ n957 ^ n386 ;
  assign n960 = ( x87 & ~n210 ) | ( x87 & n647 ) | ( ~n210 & n647 ) ;
  assign n961 = ( x11 & x66 ) | ( x11 & n725 ) | ( x66 & n725 ) ;
  assign n962 = ( x115 & n326 ) | ( x115 & n961 ) | ( n326 & n961 ) ;
  assign n963 = ( n425 & n960 ) | ( n425 & n962 ) | ( n960 & n962 ) ;
  assign n964 = ( n609 & n756 ) | ( n609 & n963 ) | ( n756 & n963 ) ;
  assign n965 = ( n729 & n959 ) | ( n729 & n964 ) | ( n959 & n964 ) ;
  assign n966 = ( n533 & ~n956 ) | ( n533 & n965 ) | ( ~n956 & n965 ) ;
  assign n977 = n976 ^ n974 ^ n966 ;
  assign n978 = ( n933 & n949 ) | ( n933 & ~n977 ) | ( n949 & ~n977 ) ;
  assign n1038 = n1037 ^ n1036 ^ n978 ;
  assign n1045 = n454 ^ n141 ^ x48 ;
  assign n1046 = ( x81 & n702 ) | ( x81 & n1045 ) | ( n702 & n1045 ) ;
  assign n1047 = ( x109 & ~n305 ) | ( x109 & n1046 ) | ( ~n305 & n1046 ) ;
  assign n1048 = ( n644 & n870 ) | ( n644 & ~n1047 ) | ( n870 & ~n1047 ) ;
  assign n1042 = ( x9 & n390 ) | ( x9 & ~n914 ) | ( n390 & ~n914 ) ;
  assign n1043 = n1042 ^ n461 ^ x35 ;
  assign n1039 = ( n248 & n442 ) | ( n248 & n746 ) | ( n442 & n746 ) ;
  assign n1040 = ( n206 & n455 ) | ( n206 & n1039 ) | ( n455 & n1039 ) ;
  assign n1041 = ( ~x108 & n533 ) | ( ~x108 & n1040 ) | ( n533 & n1040 ) ;
  assign n1044 = n1043 ^ n1041 ^ x33 ;
  assign n1049 = n1048 ^ n1044 ^ n477 ;
  assign n1072 = ( n353 & n363 ) | ( n353 & ~n601 ) | ( n363 & ~n601 ) ;
  assign n1073 = ( n546 & n922 ) | ( n546 & n1072 ) | ( n922 & n1072 ) ;
  assign n1074 = n1073 ^ n753 ^ n225 ;
  assign n1075 = n1074 ^ n791 ^ n698 ;
  assign n1067 = n944 ^ n259 ^ n193 ;
  assign n1068 = n920 ^ n850 ^ x6 ;
  assign n1069 = ( n360 & ~n473 ) | ( n360 & n1068 ) | ( ~n473 & n1068 ) ;
  assign n1070 = ( ~n272 & n1067 ) | ( ~n272 & n1069 ) | ( n1067 & n1069 ) ;
  assign n1050 = ( ~x76 & n229 ) | ( ~x76 & n385 ) | ( n229 & n385 ) ;
  assign n1051 = n594 ^ x48 ^ x18 ;
  assign n1052 = n1051 ^ x92 ^ x64 ;
  assign n1053 = n812 ^ n175 ^ n138 ;
  assign n1054 = ( ~n174 & n229 ) | ( ~n174 & n253 ) | ( n229 & n253 ) ;
  assign n1055 = n731 ^ n351 ^ n137 ;
  assign n1056 = ( n1053 & ~n1054 ) | ( n1053 & n1055 ) | ( ~n1054 & n1055 ) ;
  assign n1057 = ( n1050 & n1052 ) | ( n1050 & ~n1056 ) | ( n1052 & ~n1056 ) ;
  assign n1058 = ( n278 & ~n296 ) | ( n278 & n397 ) | ( ~n296 & n397 ) ;
  assign n1059 = n1058 ^ n734 ^ n475 ;
  assign n1060 = ( n349 & n946 ) | ( n349 & ~n1059 ) | ( n946 & ~n1059 ) ;
  assign n1061 = ( n261 & ~n1057 ) | ( n261 & n1060 ) | ( ~n1057 & n1060 ) ;
  assign n1064 = ( n227 & n337 ) | ( n227 & n476 ) | ( n337 & n476 ) ;
  assign n1062 = ( ~x39 & n146 ) | ( ~x39 & n355 ) | ( n146 & n355 ) ;
  assign n1063 = n1062 ^ n1057 ^ n323 ;
  assign n1065 = n1064 ^ n1063 ^ n225 ;
  assign n1066 = ( n433 & n1061 ) | ( n433 & ~n1065 ) | ( n1061 & ~n1065 ) ;
  assign n1071 = n1070 ^ n1066 ^ n616 ;
  assign n1076 = n1075 ^ n1071 ^ n184 ;
  assign n1077 = n642 ^ n595 ^ n336 ;
  assign n1078 = ( x5 & x30 ) | ( x5 & ~n1077 ) | ( x30 & ~n1077 ) ;
  assign n1079 = n322 ^ n239 ^ x55 ;
  assign n1080 = ( n293 & n893 ) | ( n293 & n1079 ) | ( n893 & n1079 ) ;
  assign n1081 = n1080 ^ n986 ^ n711 ;
  assign n1082 = ( x82 & ~x106 ) | ( x82 & n223 ) | ( ~x106 & n223 ) ;
  assign n1083 = ( n815 & n877 ) | ( n815 & n1082 ) | ( n877 & n1082 ) ;
  assign n1084 = ( n1078 & n1081 ) | ( n1078 & ~n1083 ) | ( n1081 & ~n1083 ) ;
  assign n1085 = ( ~x13 & x86 ) | ( ~x13 & n1084 ) | ( x86 & n1084 ) ;
  assign n1086 = ( n1049 & ~n1076 ) | ( n1049 & n1085 ) | ( ~n1076 & n1085 ) ;
  assign n1136 = n356 ^ n279 ^ x34 ;
  assign n1137 = n1136 ^ n536 ^ n456 ;
  assign n1138 = n1137 ^ n326 ^ n321 ;
  assign n1139 = ( x113 & ~n476 ) | ( x113 & n613 ) | ( ~n476 & n613 ) ;
  assign n1140 = ( x74 & ~n203 ) | ( x74 & n1139 ) | ( ~n203 & n1139 ) ;
  assign n1103 = n702 ^ n296 ^ x77 ;
  assign n1157 = ( n153 & n387 ) | ( n153 & n1103 ) | ( n387 & n1103 ) ;
  assign n1154 = ( n157 & n422 ) | ( n157 & ~n433 ) | ( n422 & ~n433 ) ;
  assign n1155 = ( x117 & n255 ) | ( x117 & n1154 ) | ( n255 & n1154 ) ;
  assign n1156 = n1155 ^ n363 ^ n332 ;
  assign n1149 = n883 ^ n538 ^ n452 ;
  assign n1150 = n279 ^ n183 ^ x19 ;
  assign n1151 = ( ~x23 & x84 ) | ( ~x23 & n1150 ) | ( x84 & n1150 ) ;
  assign n1152 = ( x118 & n1149 ) | ( x118 & ~n1151 ) | ( n1149 & ~n1151 ) ;
  assign n1146 = n448 ^ n426 ^ x121 ;
  assign n1147 = ( x98 & ~n269 ) | ( x98 & n346 ) | ( ~n269 & n346 ) ;
  assign n1148 = ( ~n812 & n1146 ) | ( ~n812 & n1147 ) | ( n1146 & n1147 ) ;
  assign n1143 = n835 ^ n568 ^ x99 ;
  assign n1144 = n1143 ^ n704 ^ n345 ;
  assign n1141 = n427 ^ n276 ^ n266 ;
  assign n1142 = ( ~x114 & n1002 ) | ( ~x114 & n1141 ) | ( n1002 & n1141 ) ;
  assign n1145 = n1144 ^ n1142 ^ x100 ;
  assign n1153 = n1152 ^ n1148 ^ n1145 ;
  assign n1158 = n1157 ^ n1156 ^ n1153 ;
  assign n1159 = ( ~n1138 & n1140 ) | ( ~n1138 & n1158 ) | ( n1140 & n1158 ) ;
  assign n1132 = n875 ^ n494 ^ n405 ;
  assign n1133 = ( n136 & ~n141 ) | ( n136 & n1132 ) | ( ~n141 & n1132 ) ;
  assign n1134 = ( n698 & ~n893 ) | ( n698 & n1133 ) | ( ~n893 & n1133 ) ;
  assign n1128 = n287 ^ n150 ^ x56 ;
  assign n1129 = n1128 ^ n652 ^ n255 ;
  assign n1127 = ( ~n393 & n623 ) | ( ~n393 & n763 ) | ( n623 & n763 ) ;
  assign n1130 = n1129 ^ n1127 ^ n317 ;
  assign n1131 = n1130 ^ n284 ^ n274 ;
  assign n1135 = n1134 ^ n1131 ^ n872 ;
  assign n1124 = ( n262 & n526 ) | ( n262 & ~n1054 ) | ( n526 & ~n1054 ) ;
  assign n1121 = ( x102 & ~n142 ) | ( x102 & n265 ) | ( ~n142 & n265 ) ;
  assign n1122 = n1121 ^ x99 ^ x25 ;
  assign n1123 = n1122 ^ n744 ^ x28 ;
  assign n1125 = n1124 ^ n1123 ^ n236 ;
  assign n1110 = ( n352 & n357 ) | ( n352 & n510 ) | ( n357 & n510 ) ;
  assign n1114 = ( n292 & ~n375 ) | ( n292 & n652 ) | ( ~n375 & n652 ) ;
  assign n1112 = ( n141 & ~n499 ) | ( n141 & n797 ) | ( ~n499 & n797 ) ;
  assign n1111 = n923 ^ n809 ^ n144 ;
  assign n1113 = n1112 ^ n1111 ^ n365 ;
  assign n1115 = n1114 ^ n1113 ^ x82 ;
  assign n1116 = ( x82 & n407 ) | ( x82 & ~n999 ) | ( n407 & ~n999 ) ;
  assign n1117 = n530 ^ n515 ^ n224 ;
  assign n1118 = n1117 ^ n813 ^ n693 ;
  assign n1119 = ( n986 & n1116 ) | ( n986 & ~n1118 ) | ( n1116 & ~n1118 ) ;
  assign n1120 = ( ~n1110 & n1115 ) | ( ~n1110 & n1119 ) | ( n1115 & n1119 ) ;
  assign n1087 = ( n279 & n732 ) | ( n279 & ~n892 ) | ( n732 & ~n892 ) ;
  assign n1088 = ( n133 & ~n263 ) | ( n133 & n516 ) | ( ~n263 & n516 ) ;
  assign n1089 = ( x80 & n734 ) | ( x80 & ~n1088 ) | ( n734 & ~n1088 ) ;
  assign n1090 = ( x106 & n375 ) | ( x106 & n1089 ) | ( n375 & n1089 ) ;
  assign n1098 = n690 ^ n373 ^ n322 ;
  assign n1097 = n1002 ^ n146 ^ x98 ;
  assign n1091 = n425 ^ n335 ^ x93 ;
  assign n1092 = n1091 ^ n847 ^ x58 ;
  assign n1093 = n616 ^ n208 ^ x46 ;
  assign n1094 = n1093 ^ n757 ^ n224 ;
  assign n1095 = n522 ^ n367 ^ n286 ;
  assign n1096 = ( n1092 & n1094 ) | ( n1092 & ~n1095 ) | ( n1094 & ~n1095 ) ;
  assign n1099 = n1098 ^ n1097 ^ n1096 ;
  assign n1100 = ( ~n532 & n1090 ) | ( ~n532 & n1099 ) | ( n1090 & n1099 ) ;
  assign n1107 = n703 ^ n170 ^ n138 ;
  assign n1104 = ( ~x14 & n283 ) | ( ~x14 & n1103 ) | ( n283 & n1103 ) ;
  assign n1101 = ( x34 & n144 ) | ( x34 & ~n158 ) | ( n144 & ~n158 ) ;
  assign n1102 = n1101 ^ n741 ^ x8 ;
  assign n1105 = n1104 ^ n1102 ^ x80 ;
  assign n1106 = n1105 ^ n475 ^ n444 ;
  assign n1108 = n1107 ^ n1106 ^ n273 ;
  assign n1109 = ( n1087 & ~n1100 ) | ( n1087 & n1108 ) | ( ~n1100 & n1108 ) ;
  assign n1126 = n1125 ^ n1120 ^ n1109 ;
  assign n1160 = n1159 ^ n1135 ^ n1126 ;
  assign n1161 = ( ~n164 & n580 ) | ( ~n164 & n785 ) | ( n580 & n785 ) ;
  assign n1162 = ( ~n151 & n242 ) | ( ~n151 & n257 ) | ( n242 & n257 ) ;
  assign n1163 = ( ~n344 & n621 ) | ( ~n344 & n842 ) | ( n621 & n842 ) ;
  assign n1164 = ( n708 & n1162 ) | ( n708 & ~n1163 ) | ( n1162 & ~n1163 ) ;
  assign n1165 = ( ~n151 & n266 ) | ( ~n151 & n289 ) | ( n266 & n289 ) ;
  assign n1166 = n1165 ^ n819 ^ n306 ;
  assign n1167 = ( n1047 & n1164 ) | ( n1047 & ~n1166 ) | ( n1164 & ~n1166 ) ;
  assign n1168 = ( n278 & n504 ) | ( n278 & ~n950 ) | ( n504 & ~n950 ) ;
  assign n1169 = ( ~n1161 & n1167 ) | ( ~n1161 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = n593 ^ n506 ^ n309 ;
  assign n1171 = n1170 ^ x72 ^ x28 ;
  assign n1172 = n1171 ^ n800 ^ n400 ;
  assign n1173 = ( x119 & n973 ) | ( x119 & ~n1157 ) | ( n973 & ~n1157 ) ;
  assign n1174 = ( ~n167 & n1003 ) | ( ~n167 & n1173 ) | ( n1003 & n1173 ) ;
  assign n1175 = ( ~n1169 & n1172 ) | ( ~n1169 & n1174 ) | ( n1172 & n1174 ) ;
  assign n1177 = ( ~x31 & n152 ) | ( ~x31 & n468 ) | ( n152 & n468 ) ;
  assign n1178 = ( n630 & n711 ) | ( n630 & n1177 ) | ( n711 & n1177 ) ;
  assign n1179 = n848 ^ n291 ^ n187 ;
  assign n1180 = ( ~n545 & n856 ) | ( ~n545 & n1179 ) | ( n856 & n1179 ) ;
  assign n1181 = ( n518 & n1178 ) | ( n518 & ~n1180 ) | ( n1178 & ~n1180 ) ;
  assign n1182 = ( n349 & n765 ) | ( n349 & ~n1181 ) | ( n765 & ~n1181 ) ;
  assign n1176 = n787 ^ n301 ^ n183 ;
  assign n1183 = n1182 ^ n1176 ^ n986 ;
  assign n1190 = n1121 ^ n354 ^ n164 ;
  assign n1191 = ( x79 & n534 ) | ( x79 & ~n1190 ) | ( n534 & ~n1190 ) ;
  assign n1188 = n894 ^ n398 ^ n349 ;
  assign n1189 = ( x65 & n151 ) | ( x65 & ~n1188 ) | ( n151 & ~n1188 ) ;
  assign n1184 = ( ~x100 & n183 ) | ( ~x100 & n301 ) | ( n183 & n301 ) ;
  assign n1185 = n1184 ^ n916 ^ n167 ;
  assign n1186 = n1185 ^ n156 ^ x63 ;
  assign n1187 = ( n504 & n885 ) | ( n504 & ~n1186 ) | ( n885 & ~n1186 ) ;
  assign n1192 = n1191 ^ n1189 ^ n1187 ;
  assign n1193 = ( n965 & n1183 ) | ( n965 & n1192 ) | ( n1183 & n1192 ) ;
  assign n1194 = ( ~n396 & n1175 ) | ( ~n396 & n1193 ) | ( n1175 & n1193 ) ;
  assign n1208 = n215 ^ x111 ^ x26 ;
  assign n1209 = n1208 ^ n471 ^ n335 ;
  assign n1207 = ( n238 & n692 ) | ( n238 & n1146 ) | ( n692 & n1146 ) ;
  assign n1210 = n1209 ^ n1207 ^ n508 ;
  assign n1211 = ( ~x72 & n998 ) | ( ~x72 & n1210 ) | ( n998 & n1210 ) ;
  assign n1212 = ( ~x20 & x49 ) | ( ~x20 & x59 ) | ( x49 & x59 ) ;
  assign n1213 = ( x72 & ~n285 ) | ( x72 & n1212 ) | ( ~n285 & n1212 ) ;
  assign n1214 = n1213 ^ n988 ^ n518 ;
  assign n1215 = ( n732 & n814 ) | ( n732 & n1214 ) | ( n814 & n1214 ) ;
  assign n1216 = ( n706 & n1211 ) | ( n706 & n1215 ) | ( n1211 & n1215 ) ;
  assign n1205 = n1177 ^ n527 ^ n316 ;
  assign n1204 = ( x42 & n350 ) | ( x42 & n599 ) | ( n350 & n599 ) ;
  assign n1201 = ( n248 & n503 ) | ( n248 & ~n1093 ) | ( n503 & ~n1093 ) ;
  assign n1202 = ( x103 & n321 ) | ( x103 & n1201 ) | ( n321 & n1201 ) ;
  assign n1203 = n1202 ^ n1166 ^ n358 ;
  assign n1206 = n1205 ^ n1204 ^ n1203 ;
  assign n1198 = n1015 ^ n599 ^ n341 ;
  assign n1199 = ( n953 & ~n1012 ) | ( n953 & n1198 ) | ( ~n1012 & n1198 ) ;
  assign n1196 = n1107 ^ n321 ^ x62 ;
  assign n1197 = n1196 ^ n355 ^ n224 ;
  assign n1195 = n586 ^ n375 ^ n296 ;
  assign n1200 = n1199 ^ n1197 ^ n1195 ;
  assign n1217 = n1216 ^ n1206 ^ n1200 ;
  assign n1246 = ( x105 & x125 ) | ( x105 & ~n377 ) | ( x125 & ~n377 ) ;
  assign n1244 = n1154 ^ n982 ^ n339 ;
  assign n1245 = n1244 ^ n489 ^ n254 ;
  assign n1247 = n1246 ^ n1245 ^ n535 ;
  assign n1243 = ( x20 & ~x31 ) | ( x20 & n733 ) | ( ~x31 & n733 ) ;
  assign n1241 = n1132 ^ n583 ^ x125 ;
  assign n1238 = ( n207 & n501 ) | ( n207 & n542 ) | ( n501 & n542 ) ;
  assign n1239 = n1238 ^ n1000 ^ n417 ;
  assign n1237 = ( n448 & ~n708 ) | ( n448 & n1180 ) | ( ~n708 & n1180 ) ;
  assign n1240 = n1239 ^ n1237 ^ n339 ;
  assign n1242 = n1241 ^ n1240 ^ x65 ;
  assign n1248 = n1247 ^ n1243 ^ n1242 ;
  assign n1249 = ( ~x110 & x125 ) | ( ~x110 & n1248 ) | ( x125 & n1248 ) ;
  assign n1230 = n986 ^ n599 ^ x61 ;
  assign n1227 = ( n333 & n452 ) | ( n333 & n741 ) | ( n452 & n741 ) ;
  assign n1228 = ( ~n500 & n720 ) | ( ~n500 & n1227 ) | ( n720 & n1227 ) ;
  assign n1229 = n1228 ^ n220 ^ n162 ;
  assign n1224 = ( n352 & ~n637 ) | ( n352 & n957 ) | ( ~n637 & n957 ) ;
  assign n1225 = n1091 ^ x111 ^ x40 ;
  assign n1226 = ( n311 & n1224 ) | ( n311 & n1225 ) | ( n1224 & n1225 ) ;
  assign n1231 = n1230 ^ n1229 ^ n1226 ;
  assign n1233 = n1178 ^ n1146 ^ n713 ;
  assign n1232 = n1095 ^ n891 ^ x96 ;
  assign n1234 = n1233 ^ n1232 ^ n746 ;
  assign n1235 = ( n478 & ~n1231 ) | ( n478 & n1234 ) | ( ~n1231 & n1234 ) ;
  assign n1218 = n685 ^ n624 ^ x16 ;
  assign n1219 = ( n561 & n690 ) | ( n561 & ~n857 ) | ( n690 & ~n857 ) ;
  assign n1220 = ( n446 & ~n999 ) | ( n446 & n1219 ) | ( ~n999 & n1219 ) ;
  assign n1221 = n893 ^ n811 ^ n652 ;
  assign n1222 = n1221 ^ n1149 ^ n462 ;
  assign n1223 = ( n1218 & n1220 ) | ( n1218 & ~n1222 ) | ( n1220 & ~n1222 ) ;
  assign n1236 = n1235 ^ n1223 ^ n333 ;
  assign n1250 = n1249 ^ n1236 ^ n395 ;
  assign n1251 = n295 ^ x50 ^ x22 ;
  assign n1252 = ( n160 & n436 ) | ( n160 & n542 ) | ( n436 & n542 ) ;
  assign n1253 = ( n509 & ~n608 ) | ( n509 & n1252 ) | ( ~n608 & n1252 ) ;
  assign n1254 = ( x43 & ~n1251 ) | ( x43 & n1253 ) | ( ~n1251 & n1253 ) ;
  assign n1255 = ( ~n298 & n637 ) | ( ~n298 & n1254 ) | ( n637 & n1254 ) ;
  assign n1256 = ( n389 & n392 ) | ( n389 & n1002 ) | ( n392 & n1002 ) ;
  assign n1258 = ( ~n266 & n581 ) | ( ~n266 & n635 ) | ( n581 & n635 ) ;
  assign n1257 = n526 ^ n490 ^ n223 ;
  assign n1259 = n1258 ^ n1257 ^ n876 ;
  assign n1276 = n610 ^ n441 ^ n177 ;
  assign n1277 = n540 ^ n332 ^ n272 ;
  assign n1278 = ( ~n411 & n953 ) | ( ~n411 & n1277 ) | ( n953 & n1277 ) ;
  assign n1279 = ( x103 & n1276 ) | ( x103 & ~n1278 ) | ( n1276 & ~n1278 ) ;
  assign n1273 = ( x56 & x82 ) | ( x56 & ~n1133 ) | ( x82 & ~n1133 ) ;
  assign n1270 = n484 ^ n237 ^ n201 ;
  assign n1269 = ( ~x82 & n215 ) | ( ~x82 & n383 ) | ( n215 & n383 ) ;
  assign n1271 = n1270 ^ n1269 ^ x45 ;
  assign n1272 = n1271 ^ n418 ^ x107 ;
  assign n1274 = n1273 ^ n1272 ^ n523 ;
  assign n1275 = n1274 ^ n404 ^ n129 ;
  assign n1267 = ( x20 & x48 ) | ( x20 & n580 ) | ( x48 & n580 ) ;
  assign n1263 = ( n297 & ~n333 ) | ( n297 & n488 ) | ( ~n333 & n488 ) ;
  assign n1264 = ( n595 & n1048 ) | ( n595 & ~n1263 ) | ( n1048 & ~n1263 ) ;
  assign n1265 = n1264 ^ n936 ^ n471 ;
  assign n1266 = ( n421 & n871 ) | ( n421 & ~n1265 ) | ( n871 & ~n1265 ) ;
  assign n1261 = ( n289 & n367 ) | ( n289 & n722 ) | ( n367 & n722 ) ;
  assign n1260 = ( ~n233 & n775 ) | ( ~n233 & n1114 ) | ( n775 & n1114 ) ;
  assign n1262 = n1261 ^ n1260 ^ n1186 ;
  assign n1268 = n1267 ^ n1266 ^ n1262 ;
  assign n1280 = n1279 ^ n1275 ^ n1268 ;
  assign n1281 = ( x83 & n392 ) | ( x83 & n1280 ) | ( n392 & n1280 ) ;
  assign n1282 = ( ~n1256 & n1259 ) | ( ~n1256 & n1281 ) | ( n1259 & n1281 ) ;
  assign n1332 = n538 ^ n349 ^ n347 ;
  assign n1333 = n1332 ^ n197 ^ x1 ;
  assign n1334 = n931 ^ n583 ^ x79 ;
  assign n1335 = n905 ^ n867 ^ n516 ;
  assign n1336 = n1335 ^ n593 ^ n308 ;
  assign n1337 = ( n600 & n1334 ) | ( n600 & ~n1336 ) | ( n1334 & ~n1336 ) ;
  assign n1338 = ( x120 & ~n1333 ) | ( x120 & n1337 ) | ( ~n1333 & n1337 ) ;
  assign n1339 = ( n280 & ~n343 ) | ( n280 & n1338 ) | ( ~n343 & n1338 ) ;
  assign n1326 = n263 ^ n202 ^ x54 ;
  assign n1327 = ( n397 & n684 ) | ( n397 & n1263 ) | ( n684 & n1263 ) ;
  assign n1328 = ( ~n131 & n654 ) | ( ~n131 & n1327 ) | ( n654 & n1327 ) ;
  assign n1329 = ( n268 & n877 ) | ( n268 & ~n1328 ) | ( n877 & ~n1328 ) ;
  assign n1330 = ( ~n412 & n1326 ) | ( ~n412 & n1329 ) | ( n1326 & n1329 ) ;
  assign n1321 = ( n224 & n375 ) | ( n224 & ~n670 ) | ( n375 & ~n670 ) ;
  assign n1322 = n1321 ^ n357 ^ x118 ;
  assign n1323 = ( n790 & n838 ) | ( n790 & ~n1322 ) | ( n838 & ~n1322 ) ;
  assign n1324 = ( ~n740 & n1185 ) | ( ~n740 & n1323 ) | ( n1185 & n1323 ) ;
  assign n1317 = n1117 ^ n774 ^ n540 ;
  assign n1318 = ( n347 & n1050 ) | ( n347 & ~n1317 ) | ( n1050 & ~n1317 ) ;
  assign n1312 = x116 ^ x79 ^ x25 ;
  assign n1313 = n1312 ^ n462 ^ n212 ;
  assign n1314 = ( n410 & ~n809 ) | ( n410 & n1313 ) | ( ~n809 & n1313 ) ;
  assign n1310 = ( n469 & ~n827 ) | ( n469 & n1110 ) | ( ~n827 & n1110 ) ;
  assign n1311 = n1310 ^ n1233 ^ n763 ;
  assign n1315 = n1314 ^ n1311 ^ n179 ;
  assign n1309 = n818 ^ n580 ^ n471 ;
  assign n1316 = n1315 ^ n1309 ^ n654 ;
  assign n1319 = n1318 ^ n1316 ^ x122 ;
  assign n1320 = ( n973 & n989 ) | ( n973 & n1319 ) | ( n989 & n1319 ) ;
  assign n1325 = n1324 ^ n1320 ^ n719 ;
  assign n1331 = n1330 ^ n1325 ^ n997 ;
  assign n1283 = ( x86 & ~n449 ) | ( x86 & n751 ) | ( ~n449 & n751 ) ;
  assign n1284 = n856 ^ n741 ^ n142 ;
  assign n1285 = n701 ^ n204 ^ n144 ;
  assign n1289 = ( n267 & n786 ) | ( n267 & ~n807 ) | ( n786 & ~n807 ) ;
  assign n1290 = ( n488 & ~n515 ) | ( n488 & n1289 ) | ( ~n515 & n1289 ) ;
  assign n1291 = ( ~x80 & n739 ) | ( ~x80 & n1290 ) | ( n739 & n1290 ) ;
  assign n1287 = n817 ^ n259 ^ n157 ;
  assign n1286 = ( n222 & n829 ) | ( n222 & n1028 ) | ( n829 & n1028 ) ;
  assign n1288 = n1287 ^ n1286 ^ x30 ;
  assign n1292 = n1291 ^ n1288 ^ n797 ;
  assign n1293 = ( n690 & ~n1285 ) | ( n690 & n1292 ) | ( ~n1285 & n1292 ) ;
  assign n1294 = ( n1283 & ~n1284 ) | ( n1283 & n1293 ) | ( ~n1284 & n1293 ) ;
  assign n1295 = ( ~n213 & n326 ) | ( ~n213 & n616 ) | ( n326 & n616 ) ;
  assign n1296 = ( n149 & n835 ) | ( n149 & ~n1295 ) | ( n835 & ~n1295 ) ;
  assign n1297 = n253 ^ n187 ^ x57 ;
  assign n1298 = n1297 ^ n900 ^ n224 ;
  assign n1299 = n1298 ^ n642 ^ n293 ;
  assign n1300 = ( n341 & n1296 ) | ( n341 & n1299 ) | ( n1296 & n1299 ) ;
  assign n1301 = n1300 ^ n1294 ^ n263 ;
  assign n1302 = ( n170 & ~n472 ) | ( n170 & n795 ) | ( ~n472 & n795 ) ;
  assign n1303 = n1302 ^ n812 ^ n211 ;
  assign n1304 = ( n135 & ~n675 ) | ( n135 & n775 ) | ( ~n675 & n775 ) ;
  assign n1305 = n611 ^ n163 ^ x39 ;
  assign n1306 = ( ~n303 & n1304 ) | ( ~n303 & n1305 ) | ( n1304 & n1305 ) ;
  assign n1307 = ( n838 & n1303 ) | ( n838 & ~n1306 ) | ( n1303 & ~n1306 ) ;
  assign n1308 = ( n1294 & n1301 ) | ( n1294 & ~n1307 ) | ( n1301 & ~n1307 ) ;
  assign n1340 = n1339 ^ n1331 ^ n1308 ;
  assign n1395 = ( x107 & n888 ) | ( x107 & ~n1026 ) | ( n888 & ~n1026 ) ;
  assign n1396 = n1298 ^ n844 ^ n158 ;
  assign n1397 = ( n1115 & n1395 ) | ( n1115 & ~n1396 ) | ( n1395 & ~n1396 ) ;
  assign n1391 = n550 ^ n540 ^ n374 ;
  assign n1392 = ( n501 & n828 ) | ( n501 & ~n1121 ) | ( n828 & ~n1121 ) ;
  assign n1393 = ( ~n1133 & n1391 ) | ( ~n1133 & n1392 ) | ( n1391 & n1392 ) ;
  assign n1387 = ( n210 & n220 ) | ( n210 & n714 ) | ( n220 & n714 ) ;
  assign n1386 = ( ~x48 & n503 ) | ( ~x48 & n995 ) | ( n503 & n995 ) ;
  assign n1388 = n1387 ^ n1386 ^ n137 ;
  assign n1389 = ( n750 & n1070 ) | ( n750 & n1388 ) | ( n1070 & n1388 ) ;
  assign n1381 = ( ~n205 & n296 ) | ( ~n205 & n516 ) | ( n296 & n516 ) ;
  assign n1382 = n1381 ^ n651 ^ n227 ;
  assign n1383 = n738 ^ n485 ^ n384 ;
  assign n1384 = n1383 ^ n403 ^ n305 ;
  assign n1385 = ( n626 & n1382 ) | ( n626 & ~n1384 ) | ( n1382 & ~n1384 ) ;
  assign n1390 = n1389 ^ n1385 ^ n663 ;
  assign n1378 = n653 ^ n642 ^ n193 ;
  assign n1379 = ( n778 & ~n857 ) | ( n778 & n1378 ) | ( ~n857 & n1378 ) ;
  assign n1375 = ( ~x95 & n204 ) | ( ~x95 & n1047 ) | ( n204 & n1047 ) ;
  assign n1376 = n1375 ^ n598 ^ n314 ;
  assign n1377 = ( n440 & ~n759 ) | ( n440 & n1376 ) | ( ~n759 & n1376 ) ;
  assign n1353 = ( x89 & n1191 ) | ( x89 & ~n1290 ) | ( n1191 & ~n1290 ) ;
  assign n1354 = n1353 ^ n1087 ^ x72 ;
  assign n1355 = n652 ^ n588 ^ n141 ;
  assign n1356 = ( ~x26 & n181 ) | ( ~x26 & n1246 ) | ( n181 & n1246 ) ;
  assign n1357 = ( n317 & ~n1355 ) | ( n317 & n1356 ) | ( ~n1355 & n1356 ) ;
  assign n1358 = ( ~n744 & n1161 ) | ( ~n744 & n1357 ) | ( n1161 & n1357 ) ;
  assign n1359 = ( ~n521 & n1354 ) | ( ~n521 & n1358 ) | ( n1354 & n1358 ) ;
  assign n1360 = ( x42 & ~n616 ) | ( x42 & n1167 ) | ( ~n616 & n1167 ) ;
  assign n1361 = ( x7 & ~n1353 ) | ( x7 & n1360 ) | ( ~n1353 & n1360 ) ;
  assign n1362 = ( n362 & n1359 ) | ( n362 & n1361 ) | ( n1359 & n1361 ) ;
  assign n1369 = ( x54 & n547 ) | ( x54 & n860 ) | ( n547 & n860 ) ;
  assign n1370 = n1369 ^ n237 ^ n234 ;
  assign n1371 = n1370 ^ n845 ^ n712 ;
  assign n1367 = n1238 ^ n789 ^ x112 ;
  assign n1366 = n945 ^ n224 ^ n193 ;
  assign n1363 = ( ~n202 & n300 ) | ( ~n202 & n1046 ) | ( n300 & n1046 ) ;
  assign n1364 = ( n782 & n1070 ) | ( n782 & ~n1363 ) | ( n1070 & ~n1363 ) ;
  assign n1365 = n1364 ^ n1042 ^ n700 ;
  assign n1368 = n1367 ^ n1366 ^ n1365 ;
  assign n1372 = n1371 ^ n1368 ^ n345 ;
  assign n1373 = ( n139 & ~n1264 ) | ( n139 & n1372 ) | ( ~n1264 & n1372 ) ;
  assign n1374 = ( n1180 & ~n1362 ) | ( n1180 & n1373 ) | ( ~n1362 & n1373 ) ;
  assign n1380 = n1379 ^ n1377 ^ n1374 ;
  assign n1394 = n1393 ^ n1390 ^ n1380 ;
  assign n1341 = n216 ^ n168 ^ x21 ;
  assign n1342 = n1017 ^ n1014 ^ x119 ;
  assign n1343 = ( x95 & n523 ) | ( x95 & ~n1342 ) | ( n523 & ~n1342 ) ;
  assign n1348 = n1208 ^ n163 ^ x25 ;
  assign n1349 = ( ~x91 & n411 ) | ( ~x91 & n1348 ) | ( n411 & n1348 ) ;
  assign n1346 = n784 ^ n759 ^ x34 ;
  assign n1347 = n1346 ^ n1207 ^ n952 ;
  assign n1344 = ( ~n599 & n835 ) | ( ~n599 & n920 ) | ( n835 & n920 ) ;
  assign n1345 = ( n649 & n902 ) | ( n649 & ~n1344 ) | ( n902 & ~n1344 ) ;
  assign n1350 = n1349 ^ n1347 ^ n1345 ;
  assign n1351 = ( n1341 & n1343 ) | ( n1341 & ~n1350 ) | ( n1343 & ~n1350 ) ;
  assign n1352 = ( n376 & ~n750 ) | ( n376 & n1351 ) | ( ~n750 & n1351 ) ;
  assign n1398 = n1397 ^ n1394 ^ n1352 ;
  assign n1405 = ( x74 & ~n495 ) | ( x74 & n1012 ) | ( ~n495 & n1012 ) ;
  assign n1407 = ( x76 & x115 ) | ( x76 & n783 ) | ( x115 & n783 ) ;
  assign n1406 = ( ~n162 & n225 ) | ( ~n162 & n831 ) | ( n225 & n831 ) ;
  assign n1408 = n1407 ^ n1406 ^ n844 ;
  assign n1409 = n660 ^ n594 ^ x30 ;
  assign n1410 = ( ~n1314 & n1408 ) | ( ~n1314 & n1409 ) | ( n1408 & n1409 ) ;
  assign n1411 = ( n1121 & n1405 ) | ( n1121 & ~n1410 ) | ( n1405 & ~n1410 ) ;
  assign n1399 = ( x119 & ~n356 ) | ( x119 & n820 ) | ( ~n356 & n820 ) ;
  assign n1401 = ( n327 & ~n503 ) | ( n327 & n920 ) | ( ~n503 & n920 ) ;
  assign n1402 = ( ~n170 & n1031 ) | ( ~n170 & n1401 ) | ( n1031 & n1401 ) ;
  assign n1400 = n352 ^ n258 ^ x5 ;
  assign n1403 = n1402 ^ n1400 ^ n832 ;
  assign n1404 = ( ~n379 & n1399 ) | ( ~n379 & n1403 ) | ( n1399 & n1403 ) ;
  assign n1412 = n1411 ^ n1404 ^ n501 ;
  assign n1481 = ( x88 & n383 ) | ( x88 & n913 ) | ( n383 & n913 ) ;
  assign n1421 = ( n390 & n859 ) | ( n390 & n1150 ) | ( n859 & n1150 ) ;
  assign n1422 = ( n480 & n764 ) | ( n480 & n1421 ) | ( n764 & n1421 ) ;
  assign n1482 = n1481 ^ n1422 ^ x1 ;
  assign n1437 = ( ~x126 & n338 ) | ( ~x126 & n845 ) | ( n338 & n845 ) ;
  assign n1438 = ( n202 & ~n614 ) | ( n202 & n1437 ) | ( ~n614 & n1437 ) ;
  assign n1439 = n1438 ^ n762 ^ x48 ;
  assign n1483 = ( n183 & n422 ) | ( n183 & n1439 ) | ( n422 & n1439 ) ;
  assign n1490 = n596 ^ n441 ^ n152 ;
  assign n1488 = ( ~x35 & n846 ) | ( ~x35 & n1297 ) | ( n846 & n1297 ) ;
  assign n1485 = ( ~x69 & x96 ) | ( ~x69 & n292 ) | ( x96 & n292 ) ;
  assign n1486 = n1485 ^ n513 ^ n434 ;
  assign n1487 = n1486 ^ n675 ^ n227 ;
  assign n1489 = n1488 ^ n1487 ^ x54 ;
  assign n1484 = ( x52 & ~x109 ) | ( x52 & n392 ) | ( ~x109 & n392 ) ;
  assign n1491 = n1490 ^ n1489 ^ n1484 ;
  assign n1492 = ( n1482 & ~n1483 ) | ( n1482 & n1491 ) | ( ~n1483 & n1491 ) ;
  assign n1460 = n150 ^ x98 ^ x75 ;
  assign n1459 = ( x46 & n303 ) | ( x46 & ~n1091 ) | ( n303 & ~n1091 ) ;
  assign n1448 = ( ~x112 & n309 ) | ( ~x112 & n519 ) | ( n309 & n519 ) ;
  assign n1449 = n1448 ^ n1008 ^ n428 ;
  assign n1450 = ( n507 & n1285 ) | ( n507 & n1449 ) | ( n1285 & n1449 ) ;
  assign n1451 = n1450 ^ n856 ^ n336 ;
  assign n1446 = n1137 ^ n1000 ^ n841 ;
  assign n1447 = n1446 ^ n850 ^ n514 ;
  assign n1443 = ( x25 & ~n447 ) | ( x25 & n569 ) | ( ~n447 & n569 ) ;
  assign n1444 = n1443 ^ n1022 ^ n670 ;
  assign n1445 = ( x97 & n975 ) | ( x97 & n1444 ) | ( n975 & n1444 ) ;
  assign n1452 = n1451 ^ n1447 ^ n1445 ;
  assign n1453 = ( x6 & ~x11 ) | ( x6 & n216 ) | ( ~x11 & n216 ) ;
  assign n1454 = ( ~x49 & n272 ) | ( ~x49 & n622 ) | ( n272 & n622 ) ;
  assign n1455 = ( n548 & ~n1453 ) | ( n548 & n1454 ) | ( ~n1453 & n1454 ) ;
  assign n1456 = ( n198 & n1149 ) | ( n198 & n1455 ) | ( n1149 & n1455 ) ;
  assign n1457 = ( n208 & n1276 ) | ( n208 & ~n1456 ) | ( n1276 & ~n1456 ) ;
  assign n1458 = ( ~n160 & n1452 ) | ( ~n160 & n1457 ) | ( n1452 & n1457 ) ;
  assign n1461 = n1460 ^ n1459 ^ n1458 ;
  assign n1462 = n717 ^ n469 ^ x112 ;
  assign n1463 = ( n197 & n285 ) | ( n197 & n570 ) | ( n285 & n570 ) ;
  assign n1464 = n1463 ^ n475 ^ n256 ;
  assign n1475 = n860 ^ n583 ^ n268 ;
  assign n1467 = ( ~n330 & n343 ) | ( ~n330 & n856 ) | ( n343 & n856 ) ;
  assign n1468 = ( x92 & n888 ) | ( x92 & n1467 ) | ( n888 & n1467 ) ;
  assign n1474 = n1468 ^ n1165 ^ n557 ;
  assign n1473 = n1191 ^ n992 ^ n775 ;
  assign n1476 = n1475 ^ n1474 ^ n1473 ;
  assign n1470 = n1111 ^ n380 ^ x20 ;
  assign n1471 = ( n640 & ~n1072 ) | ( n640 & n1470 ) | ( ~n1072 & n1470 ) ;
  assign n1469 = ( ~n712 & n1333 ) | ( ~n712 & n1468 ) | ( n1333 & n1468 ) ;
  assign n1465 = ( n548 & ~n619 ) | ( n548 & n739 ) | ( ~n619 & n739 ) ;
  assign n1466 = n1465 ^ n413 ^ n196 ;
  assign n1472 = n1471 ^ n1469 ^ n1466 ;
  assign n1477 = n1476 ^ n1472 ^ n1132 ;
  assign n1478 = ( ~n144 & n1464 ) | ( ~n144 & n1477 ) | ( n1464 & n1477 ) ;
  assign n1479 = ( n1382 & n1462 ) | ( n1382 & ~n1478 ) | ( n1462 & ~n1478 ) ;
  assign n1480 = ( n629 & n1461 ) | ( n629 & n1479 ) | ( n1461 & n1479 ) ;
  assign n1436 = n1239 ^ n1212 ^ n579 ;
  assign n1440 = n1439 ^ n1436 ^ n543 ;
  assign n1441 = n1440 ^ n648 ^ n272 ;
  assign n1430 = ( n411 & n506 ) | ( n411 & n831 ) | ( n506 & n831 ) ;
  assign n1431 = ( ~n309 & n394 ) | ( ~n309 & n1430 ) | ( n394 & n1430 ) ;
  assign n1432 = ( n385 & n509 ) | ( n385 & ~n1431 ) | ( n509 & ~n1431 ) ;
  assign n1433 = ( ~n388 & n1376 ) | ( ~n388 & n1432 ) | ( n1376 & n1432 ) ;
  assign n1429 = n1357 ^ n1070 ^ x80 ;
  assign n1434 = n1433 ^ n1429 ^ n1007 ;
  assign n1435 = n1434 ^ n1201 ^ n1019 ;
  assign n1424 = ( n162 & n360 ) | ( n162 & n404 ) | ( n360 & n404 ) ;
  assign n1425 = ( ~x94 & n891 ) | ( ~x94 & n1424 ) | ( n891 & n1424 ) ;
  assign n1426 = n1425 ^ n569 ^ x93 ;
  assign n1427 = ( n330 & n1054 ) | ( n330 & n1426 ) | ( n1054 & n1426 ) ;
  assign n1419 = n416 ^ n227 ^ x38 ;
  assign n1420 = n1419 ^ n1002 ^ n230 ;
  assign n1423 = n1422 ^ n1420 ^ n653 ;
  assign n1417 = n1239 ^ n220 ^ n191 ;
  assign n1418 = n1417 ^ n186 ^ x79 ;
  assign n1428 = n1427 ^ n1423 ^ n1418 ;
  assign n1442 = n1441 ^ n1435 ^ n1428 ;
  assign n1493 = n1492 ^ n1480 ^ n1442 ;
  assign n1413 = ( x95 & n135 ) | ( x95 & n820 ) | ( n135 & n820 ) ;
  assign n1414 = ( ~n427 & n468 ) | ( ~n427 & n1413 ) | ( n468 & n1413 ) ;
  assign n1415 = ( n175 & ~n286 ) | ( n175 & n1414 ) | ( ~n286 & n1414 ) ;
  assign n1416 = ( n401 & ~n645 ) | ( n401 & n1415 ) | ( ~n645 & n1415 ) ;
  assign n1494 = n1493 ^ n1416 ^ n1167 ;
  assign n1504 = ( x99 & n727 ) | ( x99 & ~n962 ) | ( n727 & ~n962 ) ;
  assign n1506 = ( n179 & n294 ) | ( n179 & ~n669 ) | ( n294 & ~n669 ) ;
  assign n1507 = n1506 ^ n335 ^ x99 ;
  assign n1505 = n926 ^ n770 ^ n375 ;
  assign n1508 = n1507 ^ n1505 ^ n404 ;
  assign n1509 = n452 ^ n447 ^ n131 ;
  assign n1510 = n1509 ^ n893 ^ n836 ;
  assign n1511 = ( n1045 & n1508 ) | ( n1045 & n1510 ) | ( n1508 & n1510 ) ;
  assign n1513 = n218 ^ x68 ^ x55 ;
  assign n1512 = n1305 ^ n1134 ^ n516 ;
  assign n1514 = n1513 ^ n1512 ^ n932 ;
  assign n1515 = ( n1504 & ~n1511 ) | ( n1504 & n1514 ) | ( ~n1511 & n1514 ) ;
  assign n1495 = ( ~n486 & n737 ) | ( ~n486 & n1332 ) | ( n737 & n1332 ) ;
  assign n1496 = n1188 ^ n363 ^ x62 ;
  assign n1497 = ( n198 & ~n364 ) | ( n198 & n1496 ) | ( ~n364 & n1496 ) ;
  assign n1498 = ( n681 & n1495 ) | ( n681 & ~n1497 ) | ( n1495 & ~n1497 ) ;
  assign n1499 = ( ~n363 & n422 ) | ( ~n363 & n580 ) | ( n422 & n580 ) ;
  assign n1500 = n465 ^ n348 ^ n290 ;
  assign n1501 = ( ~n744 & n1499 ) | ( ~n744 & n1500 ) | ( n1499 & n1500 ) ;
  assign n1502 = n1501 ^ n274 ^ x15 ;
  assign n1503 = ( n1411 & n1498 ) | ( n1411 & ~n1502 ) | ( n1498 & ~n1502 ) ;
  assign n1516 = n1515 ^ n1503 ^ n135 ;
  assign n1517 = ( n666 & n1489 ) | ( n666 & n1516 ) | ( n1489 & n1516 ) ;
  assign n1518 = ( ~n1412 & n1494 ) | ( ~n1412 & n1517 ) | ( n1494 & n1517 ) ;
  assign n1519 = ( n536 & n1359 ) | ( n536 & ~n1364 ) | ( n1359 & ~n1364 ) ;
  assign n1535 = n476 ^ x73 ^ x42 ;
  assign n1534 = n191 ^ n144 ^ x124 ;
  assign n1536 = n1535 ^ n1534 ^ n675 ;
  assign n1537 = ( x99 & n633 ) | ( x99 & n1536 ) | ( n633 & n1536 ) ;
  assign n1520 = ( ~n928 & n1173 ) | ( ~n928 & n1465 ) | ( n1173 & n1465 ) ;
  assign n1521 = ( n616 & n707 ) | ( n616 & ~n1520 ) | ( n707 & ~n1520 ) ;
  assign n1522 = ( n272 & n1422 ) | ( n272 & n1507 ) | ( n1422 & n1507 ) ;
  assign n1523 = ( ~x53 & n963 ) | ( ~x53 & n1522 ) | ( n963 & n1522 ) ;
  assign n1524 = n1523 ^ n1356 ^ n1010 ;
  assign n1526 = ( n386 & n629 ) | ( n386 & n1208 ) | ( n629 & n1208 ) ;
  assign n1525 = ( n590 & n958 ) | ( n590 & n1290 ) | ( n958 & n1290 ) ;
  assign n1527 = n1526 ^ n1525 ^ n634 ;
  assign n1528 = ( n208 & n1410 ) | ( n208 & ~n1482 ) | ( n1410 & ~n1482 ) ;
  assign n1529 = ( x76 & x86 ) | ( x76 & ~n215 ) | ( x86 & ~n215 ) ;
  assign n1530 = n1529 ^ n645 ^ x103 ;
  assign n1531 = ( n1527 & n1528 ) | ( n1527 & ~n1530 ) | ( n1528 & ~n1530 ) ;
  assign n1532 = ( ~n233 & n1524 ) | ( ~n233 & n1531 ) | ( n1524 & n1531 ) ;
  assign n1533 = ( x76 & ~n1521 ) | ( x76 & n1532 ) | ( ~n1521 & n1532 ) ;
  assign n1538 = n1537 ^ n1533 ^ n705 ;
  assign n1542 = n618 ^ n566 ^ n363 ;
  assign n1543 = n1542 ^ n892 ^ x12 ;
  assign n1544 = n1543 ^ n875 ^ n258 ;
  assign n1545 = n850 ^ x62 ^ x23 ;
  assign n1546 = ( n218 & n303 ) | ( n218 & ~n1545 ) | ( n303 & ~n1545 ) ;
  assign n1547 = ( n414 & n1544 ) | ( n414 & ~n1546 ) | ( n1544 & ~n1546 ) ;
  assign n1539 = n964 ^ n520 ^ n385 ;
  assign n1540 = n1539 ^ n762 ^ n394 ;
  assign n1541 = ( n293 & n658 ) | ( n293 & ~n1540 ) | ( n658 & ~n1540 ) ;
  assign n1548 = n1547 ^ n1541 ^ n794 ;
  assign n1557 = ( n172 & ~n876 ) | ( n172 & n901 ) | ( ~n876 & n901 ) ;
  assign n1558 = n1557 ^ n1026 ^ n751 ;
  assign n1559 = n1558 ^ n1229 ^ n387 ;
  assign n1551 = n1481 ^ n1405 ^ n884 ;
  assign n1552 = n1273 ^ n812 ^ x127 ;
  assign n1553 = ( n735 & ~n747 ) | ( n735 & n1552 ) | ( ~n747 & n1552 ) ;
  assign n1554 = ( n1383 & ~n1551 ) | ( n1383 & n1553 ) | ( ~n1551 & n1553 ) ;
  assign n1555 = ( n1004 & ~n1182 ) | ( n1004 & n1554 ) | ( ~n1182 & n1554 ) ;
  assign n1556 = n1555 ^ n138 ^ x29 ;
  assign n1549 = ( ~x19 & n1169 ) | ( ~x19 & n1441 ) | ( n1169 & n1441 ) ;
  assign n1550 = n1549 ^ n285 ^ x83 ;
  assign n1560 = n1559 ^ n1556 ^ n1550 ;
  assign n1570 = ( n412 & n911 ) | ( n412 & ~n1437 ) | ( n911 & ~n1437 ) ;
  assign n1571 = n1570 ^ n388 ^ x19 ;
  assign n1564 = n483 ^ n313 ^ n286 ;
  assign n1565 = n1564 ^ n351 ^ x62 ;
  assign n1566 = ( n751 & n889 ) | ( n751 & n1565 ) | ( n889 & n1565 ) ;
  assign n1567 = ( n152 & n255 ) | ( n152 & ~n747 ) | ( n255 & ~n747 ) ;
  assign n1568 = ( n1232 & ~n1383 ) | ( n1232 & n1567 ) | ( ~n1383 & n1567 ) ;
  assign n1569 = ( ~x103 & n1566 ) | ( ~x103 & n1568 ) | ( n1566 & n1568 ) ;
  assign n1561 = n817 ^ x102 ^ x20 ;
  assign n1562 = ( n630 & n1244 ) | ( n630 & n1561 ) | ( n1244 & n1561 ) ;
  assign n1563 = ( ~n472 & n742 ) | ( ~n472 & n1562 ) | ( n742 & n1562 ) ;
  assign n1572 = n1571 ^ n1569 ^ n1563 ;
  assign n1573 = ( n958 & n1560 ) | ( n958 & ~n1572 ) | ( n1560 & ~n1572 ) ;
  assign n1574 = ( n735 & n792 ) | ( n735 & ~n1573 ) | ( n792 & ~n1573 ) ;
  assign n1575 = ( ~n487 & n536 ) | ( ~n487 & n1470 ) | ( n536 & n1470 ) ;
  assign n1577 = n153 ^ x94 ^ x23 ;
  assign n1576 = n1543 ^ n469 ^ x22 ;
  assign n1578 = n1577 ^ n1576 ^ n670 ;
  assign n1579 = n1578 ^ n1513 ^ n263 ;
  assign n1581 = ( n251 & n1240 ) | ( n251 & n1537 ) | ( n1240 & n1537 ) ;
  assign n1580 = ( ~n348 & n485 ) | ( ~n348 & n731 ) | ( n485 & n731 ) ;
  assign n1582 = n1581 ^ n1580 ^ n915 ;
  assign n1589 = ( x107 & n334 ) | ( x107 & ~n1078 ) | ( n334 & ~n1078 ) ;
  assign n1587 = n1112 ^ x121 ^ x53 ;
  assign n1585 = n309 ^ n229 ^ n135 ;
  assign n1586 = n1585 ^ n1031 ^ n673 ;
  assign n1583 = ( n573 & ~n1075 ) | ( n573 & n1348 ) | ( ~n1075 & n1348 ) ;
  assign n1584 = ( n165 & n551 ) | ( n165 & ~n1583 ) | ( n551 & ~n1583 ) ;
  assign n1588 = n1587 ^ n1586 ^ n1584 ;
  assign n1590 = n1589 ^ n1588 ^ x62 ;
  assign n1591 = n1185 ^ n372 ^ n342 ;
  assign n1592 = ( ~n156 & n182 ) | ( ~n156 & n1591 ) | ( n182 & n1591 ) ;
  assign n1593 = ( n536 & n549 ) | ( n536 & ~n1592 ) | ( n549 & ~n1592 ) ;
  assign n1594 = n1124 ^ n832 ^ n140 ;
  assign n1595 = n716 ^ n386 ^ n164 ;
  assign n1596 = n1595 ^ n712 ^ n633 ;
  assign n1597 = ( n147 & ~n1336 ) | ( n147 & n1596 ) | ( ~n1336 & n1596 ) ;
  assign n1598 = n1597 ^ n571 ^ n322 ;
  assign n1599 = n1598 ^ n1251 ^ n972 ;
  assign n1600 = ( n566 & n1180 ) | ( n566 & ~n1599 ) | ( n1180 & ~n1599 ) ;
  assign n1601 = ( n1593 & n1594 ) | ( n1593 & n1600 ) | ( n1594 & n1600 ) ;
  assign n1602 = ( n394 & ~n652 ) | ( n394 & n1031 ) | ( ~n652 & n1031 ) ;
  assign n1603 = n366 ^ n240 ^ x40 ;
  assign n1604 = n841 ^ n795 ^ n405 ;
  assign n1605 = ( x58 & ~n1603 ) | ( x58 & n1604 ) | ( ~n1603 & n1604 ) ;
  assign n1606 = ( n1050 & n1602 ) | ( n1050 & n1605 ) | ( n1602 & n1605 ) ;
  assign n1607 = ( n475 & n1079 ) | ( n475 & ~n1139 ) | ( n1079 & ~n1139 ) ;
  assign n1608 = n922 ^ n766 ^ n624 ;
  assign n1609 = ( n318 & n1001 ) | ( n318 & ~n1509 ) | ( n1001 & ~n1509 ) ;
  assign n1610 = ( ~n928 & n1608 ) | ( ~n928 & n1609 ) | ( n1608 & n1609 ) ;
  assign n1611 = ( n1042 & n1607 ) | ( n1042 & ~n1610 ) | ( n1607 & ~n1610 ) ;
  assign n1612 = ( ~n235 & n273 ) | ( ~n235 & n1611 ) | ( n273 & n1611 ) ;
  assign n1613 = ( n924 & n1306 ) | ( n924 & ~n1528 ) | ( n1306 & ~n1528 ) ;
  assign n1614 = ( n230 & n240 ) | ( n230 & n1510 ) | ( n240 & n1510 ) ;
  assign n1615 = ( ~n1612 & n1613 ) | ( ~n1612 & n1614 ) | ( n1613 & n1614 ) ;
  assign n1616 = ( n1601 & n1606 ) | ( n1601 & ~n1615 ) | ( n1606 & ~n1615 ) ;
  assign n1617 = ( n1582 & ~n1590 ) | ( n1582 & n1616 ) | ( ~n1590 & n1616 ) ;
  assign n1618 = ( n1575 & n1579 ) | ( n1575 & ~n1617 ) | ( n1579 & ~n1617 ) ;
  assign n1655 = ( n159 & n1177 ) | ( n159 & n1443 ) | ( n1177 & n1443 ) ;
  assign n1656 = n1655 ^ n1578 ^ n551 ;
  assign n1653 = n1238 ^ n469 ^ n328 ;
  assign n1654 = n1653 ^ n1222 ^ n406 ;
  assign n1657 = n1656 ^ n1654 ^ x95 ;
  assign n1619 = ( n312 & n358 ) | ( n312 & ~n564 ) | ( n358 & ~n564 ) ;
  assign n1620 = ( ~n407 & n1190 ) | ( ~n407 & n1619 ) | ( n1190 & n1619 ) ;
  assign n1621 = ( n208 & n222 ) | ( n208 & n277 ) | ( n222 & n277 ) ;
  assign n1622 = ( x36 & ~n298 ) | ( x36 & n653 ) | ( ~n298 & n653 ) ;
  assign n1623 = n1622 ^ n711 ^ n706 ;
  assign n1624 = n650 ^ x120 ^ x24 ;
  assign n1625 = ( ~n1621 & n1623 ) | ( ~n1621 & n1624 ) | ( n1623 & n1624 ) ;
  assign n1626 = ( n347 & n862 ) | ( n347 & n1417 ) | ( n862 & n1417 ) ;
  assign n1649 = ( n510 & n747 ) | ( n510 & ~n979 ) | ( n747 & ~n979 ) ;
  assign n1646 = n331 ^ n268 ^ n162 ;
  assign n1647 = ( n391 & n445 ) | ( n391 & ~n1646 ) | ( n445 & ~n1646 ) ;
  assign n1643 = ( ~x28 & x53 ) | ( ~x28 & n527 ) | ( x53 & n527 ) ;
  assign n1642 = ( x49 & n1052 ) | ( x49 & ~n1525 ) | ( n1052 & ~n1525 ) ;
  assign n1639 = n1302 ^ n429 ^ x34 ;
  assign n1640 = ( n346 & n985 ) | ( n346 & ~n1639 ) | ( n985 & ~n1639 ) ;
  assign n1637 = ( ~n172 & n267 ) | ( ~n172 & n309 ) | ( n267 & n309 ) ;
  assign n1638 = ( n726 & n1265 ) | ( n726 & ~n1637 ) | ( n1265 & ~n1637 ) ;
  assign n1632 = n1050 ^ n561 ^ x13 ;
  assign n1631 = ( n1074 & n1075 ) | ( n1074 & n1413 ) | ( n1075 & n1413 ) ;
  assign n1629 = ( n260 & ~n1184 ) | ( n260 & n1321 ) | ( ~n1184 & n1321 ) ;
  assign n1627 = ( x64 & n671 ) | ( x64 & n999 ) | ( n671 & n999 ) ;
  assign n1628 = n1627 ^ n691 ^ x100 ;
  assign n1630 = n1629 ^ n1628 ^ n353 ;
  assign n1633 = n1632 ^ n1631 ^ n1630 ;
  assign n1634 = ( ~n545 & n1421 ) | ( ~n545 & n1633 ) | ( n1421 & n1633 ) ;
  assign n1635 = n1634 ^ n918 ^ n681 ;
  assign n1636 = n1635 ^ n1488 ^ n560 ;
  assign n1641 = n1640 ^ n1638 ^ n1636 ;
  assign n1644 = n1643 ^ n1642 ^ n1641 ;
  assign n1645 = ( n1011 & n1215 ) | ( n1011 & n1644 ) | ( n1215 & n1644 ) ;
  assign n1648 = n1647 ^ n1645 ^ n1242 ;
  assign n1650 = n1649 ^ n1648 ^ n1638 ;
  assign n1651 = ( ~x97 & n1626 ) | ( ~x97 & n1650 ) | ( n1626 & n1650 ) ;
  assign n1652 = ( n1620 & n1625 ) | ( n1620 & n1651 ) | ( n1625 & n1651 ) ;
  assign n1658 = n1657 ^ n1652 ^ n1114 ;
  assign n1659 = ( ~n504 & n1408 ) | ( ~n504 & n1501 ) | ( n1408 & n1501 ) ;
  assign n1662 = n737 ^ n579 ^ n378 ;
  assign n1660 = n1180 ^ n871 ^ n702 ;
  assign n1661 = ( n628 & n871 ) | ( n628 & ~n1660 ) | ( n871 & ~n1660 ) ;
  assign n1663 = n1662 ^ n1661 ^ n310 ;
  assign n1664 = n1663 ^ n1129 ^ n1125 ;
  assign n1666 = n310 ^ n279 ^ n156 ;
  assign n1667 = n1666 ^ n603 ^ n249 ;
  assign n1668 = n1667 ^ n671 ^ n307 ;
  assign n1665 = n1285 ^ n305 ^ n228 ;
  assign n1669 = n1668 ^ n1665 ^ x112 ;
  assign n1680 = ( n369 & n435 ) | ( n369 & n1526 ) | ( n435 & n1526 ) ;
  assign n1676 = ( x12 & n562 ) | ( x12 & ~n952 ) | ( n562 & ~n952 ) ;
  assign n1677 = ( n672 & ~n938 ) | ( n672 & n1676 ) | ( ~n938 & n1676 ) ;
  assign n1678 = ( n738 & ~n1127 ) | ( n738 & n1179 ) | ( ~n1127 & n1179 ) ;
  assign n1679 = ( n348 & n1677 ) | ( n348 & ~n1678 ) | ( n1677 & ~n1678 ) ;
  assign n1673 = n1567 ^ n724 ^ n157 ;
  assign n1674 = ( x120 & n790 ) | ( x120 & ~n1673 ) | ( n790 & ~n1673 ) ;
  assign n1670 = n1121 ^ n445 ^ n348 ;
  assign n1671 = n1670 ^ n241 ^ n160 ;
  assign n1672 = n1671 ^ n1201 ^ n319 ;
  assign n1675 = n1674 ^ n1672 ^ n511 ;
  assign n1681 = n1680 ^ n1679 ^ n1675 ;
  assign n1682 = n703 ^ n248 ^ x80 ;
  assign n1683 = ( x115 & n537 ) | ( x115 & ~n1424 ) | ( n537 & ~n1424 ) ;
  assign n1684 = n1683 ^ n956 ^ n831 ;
  assign n1685 = ( n231 & ~n1682 ) | ( n231 & n1684 ) | ( ~n1682 & n1684 ) ;
  assign n1686 = ( n1669 & n1681 ) | ( n1669 & ~n1685 ) | ( n1681 & ~n1685 ) ;
  assign n1687 = ( ~n1659 & n1664 ) | ( ~n1659 & n1686 ) | ( n1664 & n1686 ) ;
  assign n1688 = ( ~x124 & n597 ) | ( ~x124 & n954 ) | ( n597 & n954 ) ;
  assign n1689 = n1688 ^ n1012 ^ n981 ;
  assign n1690 = ( n717 & n838 ) | ( n717 & n1571 ) | ( n838 & n1571 ) ;
  assign n1692 = n1002 ^ n786 ^ n403 ;
  assign n1691 = ( x26 & n522 ) | ( x26 & n806 ) | ( n522 & n806 ) ;
  assign n1693 = n1692 ^ n1691 ^ n231 ;
  assign n1694 = n450 ^ n404 ^ n310 ;
  assign n1695 = ( n1268 & ~n1693 ) | ( n1268 & n1694 ) | ( ~n1693 & n1694 ) ;
  assign n1696 = ( n892 & n1690 ) | ( n892 & n1695 ) | ( n1690 & n1695 ) ;
  assign n1706 = x70 ^ x39 ^ x21 ;
  assign n1707 = ( n352 & n845 ) | ( n352 & n1706 ) | ( n845 & n1706 ) ;
  assign n1708 = ( ~x4 & x105 ) | ( ~x4 & n1707 ) | ( x105 & n1707 ) ;
  assign n1697 = ( x103 & n477 ) | ( x103 & n648 ) | ( n477 & n648 ) ;
  assign n1698 = ( ~x105 & n229 ) | ( ~x105 & n1697 ) | ( n229 & n1697 ) ;
  assign n1699 = ( n165 & n311 ) | ( n165 & n1698 ) | ( n311 & n1698 ) ;
  assign n1702 = n709 ^ n304 ^ x3 ;
  assign n1701 = n1536 ^ n613 ^ n144 ;
  assign n1700 = n847 ^ n715 ^ n651 ;
  assign n1703 = n1702 ^ n1701 ^ n1700 ;
  assign n1704 = n1703 ^ n798 ^ x41 ;
  assign n1705 = ( n1059 & ~n1699 ) | ( n1059 & n1704 ) | ( ~n1699 & n1704 ) ;
  assign n1709 = n1708 ^ n1705 ^ n243 ;
  assign n1710 = ( ~n1689 & n1696 ) | ( ~n1689 & n1709 ) | ( n1696 & n1709 ) ;
  assign n1711 = n1710 ^ n846 ^ n211 ;
  assign n1712 = ( n301 & n855 ) | ( n301 & n1238 ) | ( n855 & n1238 ) ;
  assign n1713 = ( ~x112 & n411 ) | ( ~x112 & n827 ) | ( n411 & n827 ) ;
  assign n1714 = ( n859 & ~n1712 ) | ( n859 & n1713 ) | ( ~n1712 & n1713 ) ;
  assign n1715 = n1714 ^ n920 ^ n888 ;
  assign n1716 = n1715 ^ n1104 ^ n531 ;
  assign n1717 = ( n224 & n744 ) | ( n224 & n1716 ) | ( n744 & n1716 ) ;
  assign n1719 = n383 ^ n268 ^ n246 ;
  assign n1718 = ( n538 & n579 ) | ( n538 & ~n802 ) | ( n579 & ~n802 ) ;
  assign n1720 = n1719 ^ n1718 ^ n1400 ;
  assign n1721 = n869 ^ n737 ^ n173 ;
  assign n1722 = n1721 ^ n439 ^ n172 ;
  assign n1723 = n1722 ^ n632 ^ n364 ;
  assign n1724 = n1723 ^ n754 ^ n424 ;
  assign n1725 = ( n444 & n1720 ) | ( n444 & n1724 ) | ( n1720 & n1724 ) ;
  assign n1726 = ( ~n389 & n1717 ) | ( ~n389 & n1725 ) | ( n1717 & n1725 ) ;
  assign n1727 = n1571 ^ n360 ^ x44 ;
  assign n1728 = ( x10 & n812 ) | ( x10 & n903 ) | ( n812 & n903 ) ;
  assign n1729 = ( n478 & n844 ) | ( n478 & ~n1728 ) | ( n844 & ~n1728 ) ;
  assign n1743 = ( n351 & n632 ) | ( n351 & n1082 ) | ( n632 & n1082 ) ;
  assign n1744 = n1743 ^ n1463 ^ n794 ;
  assign n1741 = ( ~n594 & n858 ) | ( ~n594 & n895 ) | ( n858 & n895 ) ;
  assign n1740 = n1695 ^ n1450 ^ n1405 ;
  assign n1733 = n409 ^ x72 ^ x30 ;
  assign n1732 = n777 ^ n676 ^ n222 ;
  assign n1730 = n223 ^ n209 ^ n194 ;
  assign n1731 = n1730 ^ n495 ^ n176 ;
  assign n1734 = n1733 ^ n1732 ^ n1731 ;
  assign n1735 = n1629 ^ n665 ^ n425 ;
  assign n1736 = ( n781 & n1424 ) | ( n781 & ~n1660 ) | ( n1424 & ~n1660 ) ;
  assign n1737 = ( n768 & ~n1223 ) | ( n768 & n1370 ) | ( ~n1223 & n1370 ) ;
  assign n1738 = ( n1735 & ~n1736 ) | ( n1735 & n1737 ) | ( ~n1736 & n1737 ) ;
  assign n1739 = ( n777 & ~n1734 ) | ( n777 & n1738 ) | ( ~n1734 & n1738 ) ;
  assign n1742 = n1741 ^ n1740 ^ n1739 ;
  assign n1745 = n1744 ^ n1742 ^ n1381 ;
  assign n1746 = ( n1727 & n1729 ) | ( n1727 & ~n1745 ) | ( n1729 & ~n1745 ) ;
  assign n1760 = ( x97 & n308 ) | ( x97 & n552 ) | ( n308 & n552 ) ;
  assign n1753 = ( x50 & n921 ) | ( x50 & ~n953 ) | ( n921 & ~n953 ) ;
  assign n1754 = ( n808 & n1375 ) | ( n808 & n1753 ) | ( n1375 & n1753 ) ;
  assign n1755 = ( n1075 & n1476 ) | ( n1075 & ~n1754 ) | ( n1476 & ~n1754 ) ;
  assign n1756 = n1213 ^ n911 ^ n370 ;
  assign n1757 = ( ~x124 & n1470 ) | ( ~x124 & n1756 ) | ( n1470 & n1756 ) ;
  assign n1758 = n1757 ^ n1258 ^ n622 ;
  assign n1759 = ( n1304 & n1755 ) | ( n1304 & n1758 ) | ( n1755 & n1758 ) ;
  assign n1750 = n1443 ^ n920 ^ n150 ;
  assign n1748 = n1101 ^ n770 ^ n546 ;
  assign n1747 = n1529 ^ n392 ^ n174 ;
  assign n1749 = n1748 ^ n1747 ^ x118 ;
  assign n1751 = n1750 ^ n1749 ^ n1579 ;
  assign n1752 = n1751 ^ n1270 ^ n212 ;
  assign n1761 = n1760 ^ n1759 ^ n1752 ;
  assign n1762 = ( n421 & n543 ) | ( n421 & ~n835 ) | ( n543 & ~n835 ) ;
  assign n1763 = ( n425 & n848 ) | ( n425 & ~n1762 ) | ( n848 & ~n1762 ) ;
  assign n1764 = ( n638 & ~n1040 ) | ( n638 & n1763 ) | ( ~n1040 & n1763 ) ;
  assign n1777 = n1647 ^ n450 ^ n259 ;
  assign n1776 = n899 ^ n729 ^ x0 ;
  assign n1768 = ( n176 & n440 ) | ( n176 & ~n1054 ) | ( n440 & ~n1054 ) ;
  assign n1769 = n1768 ^ n279 ^ x109 ;
  assign n1765 = n594 ^ n489 ^ n352 ;
  assign n1766 = n1765 ^ n781 ^ n480 ;
  assign n1767 = n1766 ^ n1290 ^ n755 ;
  assign n1770 = n1769 ^ n1767 ^ n888 ;
  assign n1771 = ( n441 & n1334 ) | ( n441 & ~n1378 ) | ( n1334 & ~n1378 ) ;
  assign n1772 = n1771 ^ n846 ^ n277 ;
  assign n1773 = ( n245 & ~n312 ) | ( n245 & n1384 ) | ( ~n312 & n1384 ) ;
  assign n1774 = n1773 ^ n1058 ^ n435 ;
  assign n1775 = ( n1770 & n1772 ) | ( n1770 & n1774 ) | ( n1772 & n1774 ) ;
  assign n1778 = n1777 ^ n1776 ^ n1775 ;
  assign n1779 = ( n1187 & n1764 ) | ( n1187 & ~n1778 ) | ( n1764 & ~n1778 ) ;
  assign n1780 = n610 ^ n480 ^ x18 ;
  assign n1781 = n1780 ^ n318 ^ n130 ;
  assign n1782 = ( n175 & n1355 ) | ( n175 & n1781 ) | ( n1355 & n1781 ) ;
  assign n1783 = ( n414 & ~n440 ) | ( n414 & n1298 ) | ( ~n440 & n1298 ) ;
  assign n1784 = ( n468 & n1147 ) | ( n468 & ~n1783 ) | ( n1147 & ~n1783 ) ;
  assign n1785 = n1784 ^ n1393 ^ n590 ;
  assign n1789 = ( x117 & n138 ) | ( x117 & ~n256 ) | ( n138 & ~n256 ) ;
  assign n1790 = ( n499 & n639 ) | ( n499 & n1789 ) | ( n639 & n1789 ) ;
  assign n1786 = ( ~n510 & n902 ) | ( ~n510 & n998 ) | ( n902 & n998 ) ;
  assign n1787 = n1786 ^ n1188 ^ n1015 ;
  assign n1788 = n1787 ^ n1748 ^ n1655 ;
  assign n1791 = n1790 ^ n1788 ^ n1090 ;
  assign n1792 = ( n1782 & ~n1785 ) | ( n1782 & n1791 ) | ( ~n1785 & n1791 ) ;
  assign n1793 = n1792 ^ n1607 ^ n557 ;
  assign n1794 = ( n519 & n735 ) | ( n519 & ~n795 ) | ( n735 & ~n795 ) ;
  assign n1795 = n1794 ^ n788 ^ n205 ;
  assign n1796 = ( n221 & n1793 ) | ( n221 & n1795 ) | ( n1793 & n1795 ) ;
  assign n1797 = ( ~n1761 & n1779 ) | ( ~n1761 & n1796 ) | ( n1779 & n1796 ) ;
  assign n1825 = ( ~x75 & n1031 ) | ( ~x75 & n1189 ) | ( n1031 & n1189 ) ;
  assign n1822 = ( x33 & ~n304 ) | ( x33 & n759 ) | ( ~n304 & n759 ) ;
  assign n1823 = n1363 ^ n842 ^ n750 ;
  assign n1824 = ( n600 & n1822 ) | ( n600 & n1823 ) | ( n1822 & n1823 ) ;
  assign n1798 = ( n366 & n788 ) | ( n366 & n1321 ) | ( n788 & n1321 ) ;
  assign n1799 = ( n368 & n1682 ) | ( n368 & n1798 ) | ( n1682 & n1798 ) ;
  assign n1800 = n1799 ^ n1499 ^ n298 ;
  assign n1801 = n354 ^ x98 ^ x65 ;
  assign n1802 = ( ~n615 & n1140 ) | ( ~n615 & n1801 ) | ( n1140 & n1801 ) ;
  assign n1803 = n1802 ^ n1624 ^ n189 ;
  assign n1818 = ( ~n299 & n438 ) | ( ~n299 & n1026 ) | ( n438 & n1026 ) ;
  assign n1817 = ( n193 & n901 ) | ( n193 & n934 ) | ( n901 & n934 ) ;
  assign n1819 = n1818 ^ n1817 ^ n425 ;
  assign n1808 = ( n138 & n538 ) | ( n138 & ~n1237 ) | ( n538 & ~n1237 ) ;
  assign n1809 = n1808 ^ n1654 ^ n1382 ;
  assign n1810 = ( n407 & n581 ) | ( n407 & n1180 ) | ( n581 & n1180 ) ;
  assign n1811 = ( n160 & n177 ) | ( n160 & n1460 ) | ( n177 & n1460 ) ;
  assign n1812 = n1811 ^ x111 ^ x49 ;
  assign n1813 = n1812 ^ n1413 ^ n362 ;
  assign n1814 = ( n592 & n1810 ) | ( n592 & ~n1813 ) | ( n1810 & ~n1813 ) ;
  assign n1815 = ( n443 & ~n528 ) | ( n443 & n1814 ) | ( ~n528 & n1814 ) ;
  assign n1816 = ( ~n348 & n1809 ) | ( ~n348 & n1815 ) | ( n1809 & n1815 ) ;
  assign n1804 = ( ~n315 & n349 ) | ( ~n315 & n982 ) | ( n349 & n982 ) ;
  assign n1805 = ( ~n1210 & n1335 ) | ( ~n1210 & n1804 ) | ( n1335 & n1804 ) ;
  assign n1806 = n1805 ^ n1602 ^ n831 ;
  assign n1807 = ( n469 & n1126 ) | ( n469 & n1806 ) | ( n1126 & n1806 ) ;
  assign n1820 = n1819 ^ n1816 ^ n1807 ;
  assign n1821 = ( n1800 & n1803 ) | ( n1800 & n1820 ) | ( n1803 & n1820 ) ;
  assign n1826 = n1825 ^ n1824 ^ n1821 ;
  assign n1827 = ( ~x68 & n934 ) | ( ~x68 & n1591 ) | ( n934 & n1591 ) ;
  assign n1828 = n1827 ^ n776 ^ n159 ;
  assign n1829 = n142 ^ x127 ^ x40 ;
  assign n1830 = ( n339 & n753 ) | ( n339 & ~n1721 ) | ( n753 & ~n1721 ) ;
  assign n1831 = n1830 ^ n1451 ^ n525 ;
  assign n1835 = n1095 ^ n719 ^ n648 ;
  assign n1832 = ( ~n578 & n1090 ) | ( ~n578 & n1220 ) | ( n1090 & n1220 ) ;
  assign n1833 = ( ~n212 & n394 ) | ( ~n212 & n1832 ) | ( n394 & n1832 ) ;
  assign n1834 = ( ~x90 & n1509 ) | ( ~x90 & n1833 ) | ( n1509 & n1833 ) ;
  assign n1836 = n1835 ^ n1834 ^ n1445 ;
  assign n1837 = ( n1829 & n1831 ) | ( n1829 & ~n1836 ) | ( n1831 & ~n1836 ) ;
  assign n1846 = n417 ^ n300 ^ x118 ;
  assign n1847 = n1846 ^ n1131 ^ n411 ;
  assign n1838 = n505 ^ n136 ^ x50 ;
  assign n1839 = ( x13 & ~n377 ) | ( x13 & n1838 ) | ( ~n377 & n1838 ) ;
  assign n1840 = n1839 ^ n1349 ^ n802 ;
  assign n1841 = ( n178 & n625 ) | ( n178 & ~n850 ) | ( n625 & ~n850 ) ;
  assign n1842 = ( n169 & n266 ) | ( n169 & ~n1543 ) | ( n266 & ~n1543 ) ;
  assign n1843 = ( n1624 & n1841 ) | ( n1624 & ~n1842 ) | ( n1841 & ~n1842 ) ;
  assign n1844 = ( ~n1415 & n1840 ) | ( ~n1415 & n1843 ) | ( n1840 & n1843 ) ;
  assign n1845 = n1844 ^ n1631 ^ n340 ;
  assign n1848 = n1847 ^ n1845 ^ n1296 ;
  assign n1849 = ( n1828 & ~n1837 ) | ( n1828 & n1848 ) | ( ~n1837 & n1848 ) ;
  assign n1852 = ( x44 & ~n350 ) | ( x44 & n1670 ) | ( ~n350 & n1670 ) ;
  assign n1853 = n1852 ^ x111 ^ x44 ;
  assign n1851 = ( ~x2 & x75 ) | ( ~x2 & n859 ) | ( x75 & n859 ) ;
  assign n1854 = n1853 ^ n1851 ^ n337 ;
  assign n1855 = ( n1143 & n1375 ) | ( n1143 & n1854 ) | ( n1375 & n1854 ) ;
  assign n1850 = n1825 ^ n1784 ^ n527 ;
  assign n1856 = n1855 ^ n1850 ^ n1469 ;
  assign n1881 = ( ~n278 & n363 ) | ( ~n278 & n867 ) | ( n363 & n867 ) ;
  assign n1882 = ( x116 & n242 ) | ( x116 & ~n1124 ) | ( n242 & ~n1124 ) ;
  assign n1883 = n293 ^ n242 ^ n205 ;
  assign n1884 = ( n666 & ~n1882 ) | ( n666 & n1883 ) | ( ~n1882 & n1883 ) ;
  assign n1885 = ( x45 & ~n292 ) | ( x45 & n650 ) | ( ~n292 & n650 ) ;
  assign n1886 = ( ~n293 & n1468 ) | ( ~n293 & n1885 ) | ( n1468 & n1885 ) ;
  assign n1887 = ( ~n1570 & n1884 ) | ( ~n1570 & n1886 ) | ( n1884 & n1886 ) ;
  assign n1888 = n1887 ^ n1615 ^ n592 ;
  assign n1889 = ( n1032 & n1881 ) | ( n1032 & n1888 ) | ( n1881 & n1888 ) ;
  assign n1872 = n1512 ^ n727 ^ n565 ;
  assign n1866 = ( n476 & n507 ) | ( n476 & ~n521 ) | ( n507 & ~n521 ) ;
  assign n1867 = ( n478 & n829 ) | ( n478 & n1866 ) | ( n829 & n1866 ) ;
  assign n1868 = ( x5 & n159 ) | ( x5 & ~n251 ) | ( n159 & ~n251 ) ;
  assign n1869 = ( n428 & n608 ) | ( n428 & ~n1868 ) | ( n608 & ~n1868 ) ;
  assign n1870 = ( x39 & ~n1867 ) | ( x39 & n1869 ) | ( ~n1867 & n1869 ) ;
  assign n1871 = ( n230 & n1462 ) | ( n230 & ~n1870 ) | ( n1462 & ~n1870 ) ;
  assign n1873 = n1872 ^ n1871 ^ n1523 ;
  assign n1877 = n168 ^ n161 ^ n159 ;
  assign n1876 = n616 ^ n132 ^ x124 ;
  assign n1878 = n1877 ^ n1876 ^ n215 ;
  assign n1874 = n1010 ^ n511 ^ n258 ;
  assign n1875 = ( x6 & n855 ) | ( x6 & n1874 ) | ( n855 & n1874 ) ;
  assign n1879 = n1878 ^ n1875 ^ n340 ;
  assign n1880 = ( x92 & ~n1873 ) | ( x92 & n1879 ) | ( ~n1873 & n1879 ) ;
  assign n1857 = n1733 ^ n726 ^ n584 ;
  assign n1858 = n1857 ^ n711 ^ n133 ;
  assign n1859 = n1801 ^ n1719 ^ n362 ;
  assign n1860 = n541 ^ n354 ^ n159 ;
  assign n1861 = ( n304 & n331 ) | ( n304 & ~n1860 ) | ( n331 & ~n1860 ) ;
  assign n1862 = ( n134 & n1358 ) | ( n134 & ~n1861 ) | ( n1358 & ~n1861 ) ;
  assign n1863 = ( n1289 & ~n1859 ) | ( n1289 & n1862 ) | ( ~n1859 & n1862 ) ;
  assign n1864 = ( n287 & ~n1668 ) | ( n287 & n1732 ) | ( ~n1668 & n1732 ) ;
  assign n1865 = ( ~n1858 & n1863 ) | ( ~n1858 & n1864 ) | ( n1863 & n1864 ) ;
  assign n1890 = n1889 ^ n1880 ^ n1865 ;
  assign n1916 = ( ~n775 & n1508 ) | ( ~n775 & n1838 ) | ( n1508 & n1838 ) ;
  assign n1914 = n1390 ^ n1052 ^ n339 ;
  assign n1915 = n1914 ^ n1303 ^ x16 ;
  assign n1917 = n1916 ^ n1915 ^ n632 ;
  assign n1911 = n1718 ^ n771 ^ n187 ;
  assign n1912 = ( n219 & ~n1005 ) | ( n219 & n1911 ) | ( ~n1005 & n1911 ) ;
  assign n1895 = ( n353 & n381 ) | ( n353 & ~n1426 ) | ( n381 & ~n1426 ) ;
  assign n1906 = ( n205 & n580 ) | ( n205 & ~n941 ) | ( n580 & ~n941 ) ;
  assign n1907 = ( ~n918 & n1445 ) | ( ~n918 & n1906 ) | ( n1445 & n1906 ) ;
  assign n1905 = ( x91 & n1180 ) | ( x91 & n1365 ) | ( n1180 & n1365 ) ;
  assign n1903 = n1129 ^ n195 ^ n181 ;
  assign n1904 = n1903 ^ n1825 ^ n848 ;
  assign n1908 = n1907 ^ n1905 ^ n1904 ;
  assign n1898 = n1766 ^ n1587 ^ n344 ;
  assign n1896 = n440 ^ x123 ^ x17 ;
  assign n1897 = ( n328 & n761 ) | ( n328 & ~n1896 ) | ( n761 & ~n1896 ) ;
  assign n1899 = n1898 ^ n1897 ^ n815 ;
  assign n1900 = n1487 ^ n1467 ^ n290 ;
  assign n1901 = n1900 ^ n1515 ^ n461 ;
  assign n1902 = ( n1881 & n1899 ) | ( n1881 & n1901 ) | ( n1899 & n1901 ) ;
  assign n1909 = n1908 ^ n1902 ^ n1206 ;
  assign n1910 = ( ~n613 & n1895 ) | ( ~n613 & n1909 ) | ( n1895 & n1909 ) ;
  assign n1891 = n1460 ^ n1155 ^ n999 ;
  assign n1892 = n1891 ^ n1660 ^ n228 ;
  assign n1893 = n1892 ^ n1431 ^ n983 ;
  assign n1894 = ( n899 & n1363 ) | ( n899 & ~n1893 ) | ( n1363 & ~n1893 ) ;
  assign n1913 = n1912 ^ n1910 ^ n1894 ;
  assign n1918 = n1917 ^ n1913 ^ n1328 ;
  assign n1919 = ( n493 & n541 ) | ( n493 & n556 ) | ( n541 & n556 ) ;
  assign n1931 = ( n773 & n1067 ) | ( n773 & n1498 ) | ( n1067 & n1498 ) ;
  assign n1928 = n841 ^ n359 ^ x56 ;
  assign n1929 = n1928 ^ n1535 ^ n1015 ;
  assign n1924 = n999 ^ n797 ^ n161 ;
  assign n1925 = ( ~x105 & n774 ) | ( ~x105 & n1924 ) | ( n774 & n1924 ) ;
  assign n1926 = n1925 ^ n921 ^ n258 ;
  assign n1927 = ( n1424 & n1628 ) | ( n1424 & n1926 ) | ( n1628 & n1926 ) ;
  assign n1930 = n1929 ^ n1927 ^ n1513 ;
  assign n1920 = ( n161 & n774 ) | ( n161 & n1422 ) | ( n774 & n1422 ) ;
  assign n1921 = ( x2 & n562 ) | ( x2 & n1920 ) | ( n562 & n1920 ) ;
  assign n1922 = ( n544 & n1512 ) | ( n544 & ~n1921 ) | ( n1512 & ~n1921 ) ;
  assign n1923 = ( n289 & ~n1433 ) | ( n289 & n1922 ) | ( ~n1433 & n1922 ) ;
  assign n1932 = n1931 ^ n1930 ^ n1923 ;
  assign n1933 = n1932 ^ n1836 ^ n676 ;
  assign n1941 = ( n254 & n536 ) | ( n254 & n585 ) | ( n536 & n585 ) ;
  assign n1942 = n1941 ^ n894 ^ n854 ;
  assign n1934 = ( ~x122 & n276 ) | ( ~x122 & n989 ) | ( n276 & n989 ) ;
  assign n1936 = ( n129 & n984 ) | ( n129 & n1238 ) | ( n984 & n1238 ) ;
  assign n1935 = ( n257 & ~n666 ) | ( n257 & n1928 ) | ( ~n666 & n1928 ) ;
  assign n1937 = n1936 ^ n1935 ^ n156 ;
  assign n1938 = n1937 ^ n1678 ^ n898 ;
  assign n1939 = ( n1176 & ~n1646 ) | ( n1176 & n1938 ) | ( ~n1646 & n1938 ) ;
  assign n1940 = ( n695 & n1934 ) | ( n695 & n1939 ) | ( n1934 & n1939 ) ;
  assign n1943 = n1942 ^ n1940 ^ n1730 ;
  assign n1959 = ( x47 & ~n523 ) | ( x47 & n1151 ) | ( ~n523 & n1151 ) ;
  assign n1958 = ( ~n1293 & n1539 ) | ( ~n1293 & n1765 ) | ( n1539 & n1765 ) ;
  assign n1960 = n1959 ^ n1958 ^ n369 ;
  assign n1944 = ( x116 & n285 ) | ( x116 & n953 ) | ( n285 & n953 ) ;
  assign n1945 = n1015 ^ n881 ^ n235 ;
  assign n1946 = n1765 ^ n397 ^ n331 ;
  assign n1947 = n1706 ^ n1020 ^ n729 ;
  assign n1948 = ( ~n767 & n1536 ) | ( ~n767 & n1947 ) | ( n1536 & n1947 ) ;
  assign n1949 = ( n746 & n1446 ) | ( n746 & ~n1948 ) | ( n1446 & ~n1948 ) ;
  assign n1950 = ( ~n1557 & n1946 ) | ( ~n1557 & n1949 ) | ( n1946 & n1949 ) ;
  assign n1951 = ( n1113 & ~n1945 ) | ( n1113 & n1950 ) | ( ~n1945 & n1950 ) ;
  assign n1955 = ( n546 & ~n723 ) | ( n546 & n1595 ) | ( ~n723 & n1595 ) ;
  assign n1953 = ( ~n226 & n227 ) | ( ~n226 & n1243 ) | ( n227 & n1243 ) ;
  assign n1952 = ( n864 & ~n1583 ) | ( n864 & n1602 ) | ( ~n1583 & n1602 ) ;
  assign n1954 = n1953 ^ n1952 ^ n138 ;
  assign n1956 = n1955 ^ n1954 ^ n1808 ;
  assign n1957 = ( ~n1944 & n1951 ) | ( ~n1944 & n1956 ) | ( n1951 & n1956 ) ;
  assign n1961 = n1960 ^ n1957 ^ n1527 ;
  assign n1962 = ( n1933 & ~n1943 ) | ( n1933 & n1961 ) | ( ~n1943 & n1961 ) ;
  assign n1963 = ( n1772 & n1919 ) | ( n1772 & n1962 ) | ( n1919 & n1962 ) ;
  assign n1964 = ( ~n240 & n441 ) | ( ~n240 & n1166 ) | ( n441 & n1166 ) ;
  assign n1965 = n1964 ^ n777 ^ n694 ;
  assign n1967 = n1321 ^ n567 ^ n537 ;
  assign n1966 = n1290 ^ n1020 ^ n912 ;
  assign n1968 = n1967 ^ n1966 ^ n1214 ;
  assign n1969 = n1017 ^ n178 ^ x66 ;
  assign n1970 = ( n1965 & n1968 ) | ( n1965 & n1969 ) | ( n1968 & n1969 ) ;
  assign n1971 = n383 ^ n190 ^ x120 ;
  assign n1972 = n808 ^ x87 ^ x21 ;
  assign n1973 = ( n337 & n1971 ) | ( n337 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1974 = n1882 ^ n1822 ^ n741 ;
  assign n1975 = ( n1721 & n1973 ) | ( n1721 & n1974 ) | ( n1973 & n1974 ) ;
  assign n1976 = ( n406 & n1016 ) | ( n406 & n1975 ) | ( n1016 & n1975 ) ;
  assign n1977 = n818 ^ n351 ^ x1 ;
  assign n1978 = ( n213 & ~n1393 ) | ( n213 & n1977 ) | ( ~n1393 & n1977 ) ;
  assign n1982 = n527 ^ n448 ^ x76 ;
  assign n1983 = n1982 ^ n1661 ^ n601 ;
  assign n1980 = ( x66 & n502 ) | ( x66 & ~n1124 ) | ( n502 & ~n1124 ) ;
  assign n1979 = ( ~n324 & n1220 ) | ( ~n324 & n1931 ) | ( n1220 & n1931 ) ;
  assign n1981 = n1980 ^ n1979 ^ n1055 ;
  assign n1984 = n1983 ^ n1981 ^ n1833 ;
  assign n2000 = n1736 ^ n1566 ^ n1049 ;
  assign n1998 = n1770 ^ n662 ^ n603 ;
  assign n1999 = ( ~n807 & n1921 ) | ( ~n807 & n1998 ) | ( n1921 & n1998 ) ;
  assign n2001 = n2000 ^ n1999 ^ n1805 ;
  assign n1994 = ( n285 & n377 ) | ( n285 & ~n470 ) | ( n377 & ~n470 ) ;
  assign n1995 = ( n946 & n1162 ) | ( n946 & ~n1994 ) | ( n1162 & ~n1994 ) ;
  assign n1996 = ( n390 & ~n1011 ) | ( n390 & n1995 ) | ( ~n1011 & n1995 ) ;
  assign n1997 = ( n984 & n1750 ) | ( n984 & n1996 ) | ( n1750 & n1996 ) ;
  assign n1988 = n1321 ^ n404 ^ n275 ;
  assign n1990 = ( n375 & n690 ) | ( n375 & ~n1000 ) | ( n690 & ~n1000 ) ;
  assign n1989 = n837 ^ n409 ^ n265 ;
  assign n1991 = n1990 ^ n1989 ^ n207 ;
  assign n1992 = n1919 ^ n1581 ^ n1020 ;
  assign n1993 = ( n1988 & n1991 ) | ( n1988 & n1992 ) | ( n1991 & n1992 ) ;
  assign n2002 = n2001 ^ n1997 ^ n1993 ;
  assign n1985 = n1273 ^ n738 ^ n272 ;
  assign n1986 = n1611 ^ n438 ^ n264 ;
  assign n1987 = ( n163 & n1985 ) | ( n163 & ~n1986 ) | ( n1985 & ~n1986 ) ;
  assign n2003 = n2002 ^ n1987 ^ n358 ;
  assign n2004 = ( n1978 & n1984 ) | ( n1978 & ~n2003 ) | ( n1984 & ~n2003 ) ;
  assign n2029 = ( n196 & ~n230 ) | ( n196 & n1298 ) | ( ~n230 & n1298 ) ;
  assign n2027 = ( ~n708 & n774 ) | ( ~n708 & n1264 ) | ( n774 & n1264 ) ;
  assign n2028 = n2027 ^ n1092 ^ n555 ;
  assign n2030 = n2029 ^ n2028 ^ n736 ;
  assign n2020 = n1213 ^ n1208 ^ x24 ;
  assign n2021 = n1884 ^ n1092 ^ n1053 ;
  assign n2022 = ( n1039 & n1231 ) | ( n1039 & n2021 ) | ( n1231 & n2021 ) ;
  assign n2023 = n1668 ^ n1023 ^ n719 ;
  assign n2024 = ( n813 & n2022 ) | ( n813 & n2023 ) | ( n2022 & n2023 ) ;
  assign n2025 = ( n492 & n2020 ) | ( n492 & ~n2024 ) | ( n2020 & ~n2024 ) ;
  assign n2007 = ( n352 & ~n588 ) | ( n352 & n1860 ) | ( ~n588 & n1860 ) ;
  assign n2006 = n334 ^ x113 ^ x44 ;
  assign n2005 = n1444 ^ n513 ^ x18 ;
  assign n2008 = n2007 ^ n2006 ^ n2005 ;
  assign n2009 = n1633 ^ n723 ^ x90 ;
  assign n2012 = n1936 ^ n1631 ^ n1427 ;
  assign n2010 = ( ~n416 & n1525 ) | ( ~n416 & n1653 ) | ( n1525 & n1653 ) ;
  assign n2011 = ( n148 & n873 ) | ( n148 & n2010 ) | ( n873 & n2010 ) ;
  assign n2013 = n2012 ^ n2011 ^ n1566 ;
  assign n2014 = n686 ^ n529 ^ n443 ;
  assign n2015 = n2014 ^ n891 ^ n732 ;
  assign n2016 = n2015 ^ n1676 ^ n402 ;
  assign n2017 = ( n2009 & n2013 ) | ( n2009 & n2016 ) | ( n2013 & n2016 ) ;
  assign n2018 = ( n1209 & n2008 ) | ( n1209 & n2017 ) | ( n2008 & n2017 ) ;
  assign n2019 = n2018 ^ n1722 ^ n1630 ;
  assign n2026 = n2025 ^ n2019 ^ n1034 ;
  assign n2031 = n2030 ^ n2026 ^ n1747 ;
  assign n2032 = ( ~n283 & n1296 ) | ( ~n283 & n1504 ) | ( n1296 & n1504 ) ;
  assign n2041 = n1906 ^ n1133 ^ n666 ;
  assign n2042 = n1178 ^ n850 ^ x2 ;
  assign n2043 = n2042 ^ n1431 ^ n231 ;
  assign n2044 = ( ~x5 & x96 ) | ( ~x5 & n681 ) | ( x96 & n681 ) ;
  assign n2045 = n2044 ^ n269 ^ x120 ;
  assign n2046 = n2045 ^ n1835 ^ n477 ;
  assign n2047 = ( ~n614 & n2043 ) | ( ~n614 & n2046 ) | ( n2043 & n2046 ) ;
  assign n2048 = ( n200 & n2041 ) | ( n200 & ~n2047 ) | ( n2041 & ~n2047 ) ;
  assign n2040 = ( n151 & n1201 ) | ( n151 & n1777 ) | ( n1201 & n1777 ) ;
  assign n2035 = n1252 ^ n1243 ^ n835 ;
  assign n2036 = ( n416 & n1511 ) | ( n416 & n2035 ) | ( n1511 & n2035 ) ;
  assign n2033 = ( n361 & ~n459 ) | ( n361 & n939 ) | ( ~n459 & n939 ) ;
  assign n2034 = n2033 ^ n1777 ^ n1117 ;
  assign n2037 = n2036 ^ n2034 ^ n883 ;
  assign n2038 = n2037 ^ n1899 ^ n1449 ;
  assign n2039 = ( n1258 & n1346 ) | ( n1258 & ~n2038 ) | ( n1346 & ~n2038 ) ;
  assign n2049 = n2048 ^ n2040 ^ n2039 ;
  assign n2059 = ( ~n321 & n381 ) | ( ~n321 & n1267 ) | ( n381 & n1267 ) ;
  assign n2060 = n2059 ^ n813 ^ n564 ;
  assign n2061 = n2060 ^ n539 ^ x50 ;
  assign n2058 = ( n649 & ~n1172 ) | ( n649 & n1644 ) | ( ~n1172 & n1644 ) ;
  assign n2056 = ( ~n1132 & n1332 ) | ( ~n1132 & n1513 ) | ( n1332 & n1513 ) ;
  assign n2050 = n440 ^ n408 ^ x125 ;
  assign n2051 = ( ~n140 & n1026 ) | ( ~n140 & n1628 ) | ( n1026 & n1628 ) ;
  assign n2052 = n2051 ^ n1784 ^ n353 ;
  assign n2053 = ( ~n306 & n944 ) | ( ~n306 & n954 ) | ( n944 & n954 ) ;
  assign n2054 = n2053 ^ n1354 ^ n434 ;
  assign n2055 = ( n2050 & n2052 ) | ( n2050 & ~n2054 ) | ( n2052 & ~n2054 ) ;
  assign n2057 = n2056 ^ n2055 ^ n148 ;
  assign n2062 = n2061 ^ n2058 ^ n2057 ;
  assign n2063 = ( n2032 & ~n2049 ) | ( n2032 & n2062 ) | ( ~n2049 & n2062 ) ;
  assign n2076 = ( n319 & n561 ) | ( n319 & ~n1453 ) | ( n561 & ~n1453 ) ;
  assign n2075 = ( n501 & ~n1050 ) | ( n501 & n1284 ) | ( ~n1050 & n1284 ) ;
  assign n2077 = n2076 ^ n2075 ^ n822 ;
  assign n2065 = ( ~n513 & n812 ) | ( ~n513 & n848 ) | ( n812 & n848 ) ;
  assign n2066 = n2065 ^ n785 ^ n373 ;
  assign n2067 = ( ~x65 & n366 ) | ( ~x65 & n2066 ) | ( n366 & n2066 ) ;
  assign n2068 = ( ~n176 & n800 ) | ( ~n176 & n1149 ) | ( n800 & n1149 ) ;
  assign n2069 = n2068 ^ n744 ^ n307 ;
  assign n2070 = ( n415 & ~n452 ) | ( n415 & n2069 ) | ( ~n452 & n2069 ) ;
  assign n2071 = ( n461 & n770 ) | ( n461 & ~n1990 ) | ( n770 & ~n1990 ) ;
  assign n2072 = n2071 ^ n1771 ^ n517 ;
  assign n2073 = ( ~n1260 & n2070 ) | ( ~n1260 & n2072 ) | ( n2070 & n2072 ) ;
  assign n2074 = ( n893 & n2067 ) | ( n893 & ~n2073 ) | ( n2067 & ~n2073 ) ;
  assign n2064 = ( x104 & n425 ) | ( x104 & ~n1677 ) | ( n425 & ~n1677 ) ;
  assign n2078 = n2077 ^ n2074 ^ n2064 ;
  assign n2082 = ( ~x105 & n1944 ) | ( ~x105 & n1945 ) | ( n1944 & n1945 ) ;
  assign n2083 = ( n590 & n891 ) | ( n590 & ~n2082 ) | ( n891 & ~n2082 ) ;
  assign n2084 = n2083 ^ n1258 ^ n991 ;
  assign n2079 = n1602 ^ n1137 ^ n796 ;
  assign n2080 = ( ~x53 & n319 ) | ( ~x53 & n1113 ) | ( n319 & n1113 ) ;
  assign n2081 = ( ~n804 & n2079 ) | ( ~n804 & n2080 ) | ( n2079 & n2080 ) ;
  assign n2085 = n2084 ^ n2081 ^ n1451 ;
  assign n2086 = n2085 ^ n2018 ^ n1821 ;
  assign n2099 = ( ~n1275 & n1426 ) | ( ~n1275 & n1776 ) | ( n1426 & n1776 ) ;
  assign n2097 = n1765 ^ n1297 ^ n1043 ;
  assign n2094 = n1781 ^ n690 ^ x19 ;
  assign n2095 = ( n460 & n802 ) | ( n460 & n2094 ) | ( n802 & n2094 ) ;
  assign n2096 = n2095 ^ n1625 ^ n1409 ;
  assign n2091 = ( ~n549 & n746 ) | ( ~n549 & n1762 ) | ( n746 & n1762 ) ;
  assign n2090 = n1240 ^ n849 ^ n567 ;
  assign n2089 = n1488 ^ n975 ^ n816 ;
  assign n2092 = n2091 ^ n2090 ^ n2089 ;
  assign n2087 = ( ~n149 & n592 ) | ( ~n149 & n861 ) | ( n592 & n861 ) ;
  assign n2088 = ( x86 & ~n1831 ) | ( x86 & n2087 ) | ( ~n1831 & n2087 ) ;
  assign n2093 = n2092 ^ n2088 ^ n376 ;
  assign n2098 = n2097 ^ n2096 ^ n2093 ;
  assign n2100 = n2099 ^ n2098 ^ n737 ;
  assign n2123 = n1882 ^ n1091 ^ n332 ;
  assign n2132 = ( ~x28 & n1444 ) | ( ~x28 & n1656 ) | ( n1444 & n1656 ) ;
  assign n2128 = n1186 ^ x106 ^ x91 ;
  assign n2129 = n2128 ^ n2027 ^ n1141 ;
  assign n2130 = ( n362 & n672 ) | ( n362 & ~n2129 ) | ( n672 & ~n2129 ) ;
  assign n2131 = ( n496 & n1498 ) | ( n496 & ~n2130 ) | ( n1498 & ~n2130 ) ;
  assign n2124 = ( n465 & n1007 ) | ( n465 & n1388 ) | ( n1007 & n1388 ) ;
  assign n2125 = n898 ^ n747 ^ n680 ;
  assign n2126 = n2125 ^ n1021 ^ n189 ;
  assign n2127 = ( n177 & n2124 ) | ( n177 & n2126 ) | ( n2124 & n2126 ) ;
  assign n2133 = n2132 ^ n2131 ^ n2127 ;
  assign n2134 = ( n787 & ~n2123 ) | ( n787 & n2133 ) | ( ~n2123 & n2133 ) ;
  assign n2119 = ( n313 & n912 ) | ( n313 & ~n1219 ) | ( n912 & ~n1219 ) ;
  assign n2120 = n2119 ^ n1013 ^ n495 ;
  assign n2121 = n2120 ^ n1368 ^ n1019 ;
  assign n2101 = ( x84 & ~x107 ) | ( x84 & n2065 ) | ( ~x107 & n2065 ) ;
  assign n2102 = ( n314 & n1246 ) | ( n314 & ~n2101 ) | ( n1246 & ~n2101 ) ;
  assign n2103 = ( n418 & n449 ) | ( n418 & n932 ) | ( n449 & n932 ) ;
  assign n2104 = n2103 ^ n1522 ^ x64 ;
  assign n2105 = ( x40 & ~n1287 ) | ( x40 & n2104 ) | ( ~n1287 & n2104 ) ;
  assign n2106 = n2105 ^ n1926 ^ n1224 ;
  assign n2107 = ( n1327 & n2102 ) | ( n1327 & n2106 ) | ( n2102 & n2106 ) ;
  assign n2111 = ( n157 & n1001 ) | ( n157 & n1929 ) | ( n1001 & n1929 ) ;
  assign n2112 = ( n143 & n630 ) | ( n143 & ~n2111 ) | ( n630 & ~n2111 ) ;
  assign n2109 = n1766 ^ n1150 ^ n533 ;
  assign n2108 = ( n565 & ~n817 ) | ( n565 & n1166 ) | ( ~n817 & n1166 ) ;
  assign n2110 = n2109 ^ n2108 ^ n679 ;
  assign n2113 = n2112 ^ n2110 ^ n779 ;
  assign n2114 = ( x33 & ~n541 ) | ( x33 & n753 ) | ( ~n541 & n753 ) ;
  assign n2115 = ( n303 & n926 ) | ( n303 & ~n2114 ) | ( n926 & ~n2114 ) ;
  assign n2116 = n2115 ^ n1383 ^ n1345 ;
  assign n2117 = ( n450 & n680 ) | ( n450 & n2116 ) | ( n680 & n2116 ) ;
  assign n2118 = ( ~n2107 & n2113 ) | ( ~n2107 & n2117 ) | ( n2113 & n2117 ) ;
  assign n2122 = n2121 ^ n2118 ^ n1283 ;
  assign n2135 = n2134 ^ n2122 ^ n965 ;
  assign n2139 = ( x106 & n344 ) | ( x106 & n417 ) | ( n344 & n417 ) ;
  assign n2140 = ( n611 & n658 ) | ( n611 & n1972 ) | ( n658 & n1972 ) ;
  assign n2141 = ( n302 & ~n2139 ) | ( n302 & n2140 ) | ( ~n2139 & n2140 ) ;
  assign n2142 = ( n475 & ~n607 ) | ( n475 & n2141 ) | ( ~n607 & n2141 ) ;
  assign n2136 = ( n525 & n625 ) | ( n525 & n1205 ) | ( n625 & n1205 ) ;
  assign n2137 = n1443 ^ n1247 ^ n757 ;
  assign n2138 = ( n1438 & n2136 ) | ( n1438 & ~n2137 ) | ( n2136 & ~n2137 ) ;
  assign n2143 = n2142 ^ n2138 ^ n2121 ;
  assign n2148 = ( n1383 & n1396 ) | ( n1383 & n1947 ) | ( n1396 & n1947 ) ;
  assign n2144 = n1141 ^ n495 ^ n338 ;
  assign n2145 = n2144 ^ x101 ^ x87 ;
  assign n2146 = n2145 ^ n1877 ^ n165 ;
  assign n2147 = n2146 ^ n1456 ^ n1009 ;
  assign n2149 = n2148 ^ n2147 ^ n1306 ;
  assign n2150 = ( n480 & ~n750 ) | ( n480 & n1667 ) | ( ~n750 & n1667 ) ;
  assign n2151 = n1059 ^ n443 ^ x123 ;
  assign n2152 = n2151 ^ n726 ^ n284 ;
  assign n2153 = ( ~x103 & n274 ) | ( ~x103 & n2152 ) | ( n274 & n2152 ) ;
  assign n2168 = ( ~n998 & n1071 ) | ( ~n998 & n1655 ) | ( n1071 & n1655 ) ;
  assign n2166 = n1977 ^ n1112 ^ n355 ;
  assign n2167 = n2166 ^ n1706 ^ n882 ;
  assign n2169 = n2168 ^ n2167 ^ x115 ;
  assign n2154 = ( x44 & n507 ) | ( x44 & n1104 ) | ( n507 & n1104 ) ;
  assign n2155 = ( n427 & n1259 ) | ( n427 & n2154 ) | ( n1259 & n2154 ) ;
  assign n2156 = ( x27 & n175 ) | ( x27 & ~n336 ) | ( n175 & ~n336 ) ;
  assign n2157 = n1101 ^ n947 ^ x84 ;
  assign n2158 = n1564 ^ n1059 ^ n200 ;
  assign n2159 = ( n1012 & n1185 ) | ( n1012 & ~n2158 ) | ( n1185 & ~n2158 ) ;
  assign n2160 = ( n1583 & n2157 ) | ( n1583 & n2159 ) | ( n2157 & n2159 ) ;
  assign n2161 = n2160 ^ n1260 ^ x90 ;
  assign n2162 = ( n499 & n2156 ) | ( n499 & ~n2161 ) | ( n2156 & ~n2161 ) ;
  assign n2163 = ( n534 & n2155 ) | ( n534 & ~n2162 ) | ( n2155 & ~n2162 ) ;
  assign n2164 = n2163 ^ n1418 ^ n635 ;
  assign n2165 = ( n188 & ~n1792 ) | ( n188 & n2164 ) | ( ~n1792 & n2164 ) ;
  assign n2170 = n2169 ^ n2165 ^ x110 ;
  assign n2171 = ( n2150 & n2153 ) | ( n2150 & n2170 ) | ( n2153 & n2170 ) ;
  assign n2172 = ( n2143 & n2149 ) | ( n2143 & n2171 ) | ( n2149 & n2171 ) ;
  assign n2173 = ( n555 & n572 ) | ( n555 & ~n1357 ) | ( n572 & ~n1357 ) ;
  assign n2174 = ( ~n228 & n405 ) | ( ~n228 & n1008 ) | ( n405 & n1008 ) ;
  assign n2175 = n2174 ^ n876 ^ x17 ;
  assign n2176 = n2175 ^ n472 ^ n425 ;
  assign n2177 = ( n298 & n663 ) | ( n298 & ~n2176 ) | ( n663 & ~n2176 ) ;
  assign n2178 = ( ~n726 & n1354 ) | ( ~n726 & n2177 ) | ( n1354 & n2177 ) ;
  assign n2179 = n2178 ^ n1181 ^ x4 ;
  assign n2180 = n1509 ^ n1328 ^ x39 ;
  assign n2181 = n2103 ^ n1912 ^ n622 ;
  assign n2183 = n530 ^ n384 ^ n238 ;
  assign n2182 = ( n350 & ~n1104 ) | ( n350 & n1107 ) | ( ~n1104 & n1107 ) ;
  assign n2184 = n2183 ^ n2182 ^ n741 ;
  assign n2185 = n741 ^ n347 ^ x15 ;
  assign n2186 = ( n1173 & ~n1230 ) | ( n1173 & n1290 ) | ( ~n1230 & n1290 ) ;
  assign n2187 = n2186 ^ n237 ^ x110 ;
  assign n2188 = ( n1447 & n2185 ) | ( n1447 & n2187 ) | ( n2185 & n2187 ) ;
  assign n2189 = ( ~n658 & n2184 ) | ( ~n658 & n2188 ) | ( n2184 & n2188 ) ;
  assign n2190 = ( n1173 & ~n1696 ) | ( n1173 & n2189 ) | ( ~n1696 & n2189 ) ;
  assign n2191 = ( n2180 & ~n2181 ) | ( n2180 & n2190 ) | ( ~n2181 & n2190 ) ;
  assign n2192 = ( n2173 & n2179 ) | ( n2173 & ~n2191 ) | ( n2179 & ~n2191 ) ;
  assign n2250 = ( n673 & ~n1040 ) | ( n673 & n1078 ) | ( ~n1040 & n1078 ) ;
  assign n2240 = n1092 ^ n934 ^ n397 ;
  assign n2241 = n2240 ^ n871 ^ n244 ;
  assign n2242 = n2241 ^ n1819 ^ n1050 ;
  assign n2243 = n519 ^ n397 ^ n209 ;
  assign n2244 = n2243 ^ n1373 ^ n1098 ;
  assign n2245 = ( n1501 & n1879 ) | ( n1501 & ~n2244 ) | ( n1879 & ~n2244 ) ;
  assign n2247 = ( ~x88 & n148 ) | ( ~x88 & n493 ) | ( n148 & n493 ) ;
  assign n2246 = ( x33 & n1413 ) | ( x33 & n1525 ) | ( n1413 & n1525 ) ;
  assign n2248 = n2247 ^ n2246 ^ n989 ;
  assign n2249 = ( n2242 & n2245 ) | ( n2242 & ~n2248 ) | ( n2245 & ~n2248 ) ;
  assign n2193 = n667 ^ n419 ^ n158 ;
  assign n2194 = ( n1053 & ~n1196 ) | ( n1053 & n2193 ) | ( ~n1196 & n2193 ) ;
  assign n2198 = ( ~n518 & n1090 ) | ( ~n518 & n1238 ) | ( n1090 & n1238 ) ;
  assign n2197 = n1317 ^ n1031 ^ n628 ;
  assign n2199 = n2198 ^ n2197 ^ n480 ;
  assign n2195 = n2174 ^ n1626 ^ n1063 ;
  assign n2196 = ( ~n701 & n1303 ) | ( ~n701 & n2195 ) | ( n1303 & n2195 ) ;
  assign n2200 = n2199 ^ n2196 ^ n1991 ;
  assign n2214 = n1426 ^ n1104 ^ x6 ;
  assign n2211 = n804 ^ n524 ^ n281 ;
  assign n2212 = ( x122 & n1512 ) | ( x122 & ~n2211 ) | ( n1512 & ~n2211 ) ;
  assign n2208 = ( x107 & n529 ) | ( x107 & ~n675 ) | ( n529 & ~n675 ) ;
  assign n2209 = ( x89 & ~n219 ) | ( x89 & n2208 ) | ( ~n219 & n2208 ) ;
  assign n2207 = n1971 ^ n191 ^ x72 ;
  assign n2206 = ( n1552 & n1942 ) | ( n1552 & ~n2186 ) | ( n1942 & ~n2186 ) ;
  assign n2210 = n2209 ^ n2207 ^ n2206 ;
  assign n2213 = n2212 ^ n2210 ^ n1929 ;
  assign n2215 = n2214 ^ n2213 ^ n1543 ;
  assign n2204 = ( n275 & n397 ) | ( n275 & n1022 ) | ( n397 & n1022 ) ;
  assign n2201 = n907 ^ n406 ^ x52 ;
  assign n2202 = ( n623 & ~n1133 ) | ( n623 & n2201 ) | ( ~n1133 & n2201 ) ;
  assign n2203 = ( n1439 & n1642 ) | ( n1439 & n2202 ) | ( n1642 & n2202 ) ;
  assign n2205 = n2204 ^ n2203 ^ x126 ;
  assign n2216 = n2215 ^ n2205 ^ n1638 ;
  assign n2217 = ( n424 & n2200 ) | ( n424 & ~n2216 ) | ( n2200 & ~n2216 ) ;
  assign n2218 = ( ~n367 & n634 ) | ( ~n367 & n1328 ) | ( n634 & n1328 ) ;
  assign n2219 = ( n412 & n1089 ) | ( n412 & ~n2218 ) | ( n1089 & ~n2218 ) ;
  assign n2220 = ( n171 & n889 ) | ( n171 & n2059 ) | ( n889 & n2059 ) ;
  assign n2221 = ( n554 & ~n1202 ) | ( n554 & n2220 ) | ( ~n1202 & n2220 ) ;
  assign n2226 = n1425 ^ n1146 ^ n559 ;
  assign n2222 = n1535 ^ n1462 ^ x119 ;
  assign n2223 = ( ~n524 & n854 ) | ( ~n524 & n2222 ) | ( n854 & n2222 ) ;
  assign n2224 = ( ~n1053 & n1291 ) | ( ~n1053 & n2223 ) | ( n1291 & n2223 ) ;
  assign n2225 = ( n379 & n1780 ) | ( n379 & ~n2224 ) | ( n1780 & ~n2224 ) ;
  assign n2227 = n2226 ^ n2225 ^ n1774 ;
  assign n2233 = ( n187 & ~n627 ) | ( n187 & n1794 ) | ( ~n627 & n1794 ) ;
  assign n2234 = ( ~n759 & n1539 ) | ( ~n759 & n2233 ) | ( n1539 & n2233 ) ;
  assign n2235 = ( ~n1671 & n2033 ) | ( ~n1671 & n2234 ) | ( n2033 & n2234 ) ;
  assign n2228 = ( x91 & n685 ) | ( x91 & n744 ) | ( n685 & n744 ) ;
  assign n2229 = n2228 ^ n1552 ^ n1054 ;
  assign n2230 = ( n202 & n1169 ) | ( n202 & n1272 ) | ( n1169 & n1272 ) ;
  assign n2231 = ( n728 & n2229 ) | ( n728 & n2230 ) | ( n2229 & n2230 ) ;
  assign n2232 = ( n130 & n792 ) | ( n130 & ~n2231 ) | ( n792 & ~n2231 ) ;
  assign n2236 = n2235 ^ n2232 ^ n2194 ;
  assign n2237 = ( ~n388 & n2227 ) | ( ~n388 & n2236 ) | ( n2227 & n2236 ) ;
  assign n2238 = ( n2219 & n2221 ) | ( n2219 & n2237 ) | ( n2221 & n2237 ) ;
  assign n2239 = ( ~n2194 & n2217 ) | ( ~n2194 & n2238 ) | ( n2217 & n2238 ) ;
  assign n2251 = n2250 ^ n2249 ^ n2239 ;
  assign n2252 = n1104 ^ n713 ^ n453 ;
  assign n2253 = ( n224 & n1000 ) | ( n224 & n2252 ) | ( n1000 & n2252 ) ;
  assign n2254 = n2253 ^ n681 ^ n344 ;
  assign n2255 = n1169 ^ n1056 ^ n162 ;
  assign n2256 = ( n384 & n921 ) | ( n384 & n1150 ) | ( n921 & n1150 ) ;
  assign n2257 = n2256 ^ n855 ^ n552 ;
  assign n2258 = n2257 ^ n818 ^ n235 ;
  assign n2259 = n1830 ^ n1529 ^ n331 ;
  assign n2262 = ( ~n189 & n481 ) | ( ~n189 & n1045 ) | ( n481 & n1045 ) ;
  assign n2260 = ( n519 & n681 ) | ( n519 & ~n924 ) | ( n681 & ~n924 ) ;
  assign n2261 = n2260 ^ n844 ^ n338 ;
  assign n2263 = n2262 ^ n2261 ^ x81 ;
  assign n2264 = ( x117 & n1137 ) | ( x117 & n2263 ) | ( n1137 & n2263 ) ;
  assign n2265 = ( ~n535 & n2259 ) | ( ~n535 & n2264 ) | ( n2259 & n2264 ) ;
  assign n2266 = ( n1263 & n2258 ) | ( n1263 & ~n2265 ) | ( n2258 & ~n2265 ) ;
  assign n2267 = ( n2254 & n2255 ) | ( n2254 & n2266 ) | ( n2255 & n2266 ) ;
  assign n2269 = ( ~x50 & n1258 ) | ( ~x50 & n2178 ) | ( n1258 & n2178 ) ;
  assign n2270 = ( ~n501 & n784 ) | ( ~n501 & n2269 ) | ( n784 & n2269 ) ;
  assign n2271 = ( n549 & n1682 ) | ( n549 & n2270 ) | ( n1682 & n2270 ) ;
  assign n2268 = ( n1129 & n1144 ) | ( n1129 & ~n1495 ) | ( n1144 & ~n1495 ) ;
  assign n2272 = n2271 ^ n2268 ^ n2104 ;
  assign n2303 = n920 ^ n782 ^ n322 ;
  assign n2304 = ( n237 & n875 ) | ( n237 & n2303 ) | ( n875 & n2303 ) ;
  assign n2305 = ( n503 & n1218 ) | ( n503 & ~n1971 ) | ( n1218 & ~n1971 ) ;
  assign n2306 = n2305 ^ n1708 ^ n621 ;
  assign n2307 = ( ~x100 & n1438 ) | ( ~x100 & n2306 ) | ( n1438 & n2306 ) ;
  assign n2308 = n2307 ^ n1805 ^ n692 ;
  assign n2309 = ( n1174 & ~n2304 ) | ( n1174 & n2308 ) | ( ~n2304 & n2308 ) ;
  assign n2310 = n2309 ^ n677 ^ x94 ;
  assign n2294 = n1046 ^ n290 ^ n276 ;
  assign n2295 = n2294 ^ n1437 ^ n919 ;
  assign n2296 = n1766 ^ n500 ^ n454 ;
  assign n2297 = n2296 ^ n350 ^ n241 ;
  assign n2298 = ( ~n997 & n2184 ) | ( ~n997 & n2297 ) | ( n2184 & n2297 ) ;
  assign n2299 = ( n237 & n489 ) | ( n237 & ~n2298 ) | ( n489 & ~n2298 ) ;
  assign n2300 = ( n224 & n543 ) | ( n224 & n925 ) | ( n543 & n925 ) ;
  assign n2301 = n2300 ^ n813 ^ n451 ;
  assign n2302 = ( ~n2295 & n2299 ) | ( ~n2295 & n2301 ) | ( n2299 & n2301 ) ;
  assign n2292 = ( n401 & n833 ) | ( n401 & ~n866 ) | ( n833 & ~n866 ) ;
  assign n2290 = ( x81 & n1155 ) | ( x81 & n2150 ) | ( n1155 & n2150 ) ;
  assign n2291 = ( ~n247 & n547 ) | ( ~n247 & n2290 ) | ( n547 & n2290 ) ;
  assign n2293 = n2292 ^ n2291 ^ n679 ;
  assign n2311 = n2310 ^ n2302 ^ n2293 ;
  assign n2288 = n2075 ^ n1872 ^ n1750 ;
  assign n2277 = n987 ^ n781 ^ n393 ;
  assign n2278 = n2277 ^ n1163 ^ n407 ;
  assign n2279 = ( n443 & n924 ) | ( n443 & n1121 ) | ( n924 & n1121 ) ;
  assign n2280 = ( n266 & ~n2278 ) | ( n266 & n2279 ) | ( ~n2278 & n2279 ) ;
  assign n2281 = ( x95 & n524 ) | ( x95 & n836 ) | ( n524 & n836 ) ;
  assign n2282 = ( n185 & n1381 ) | ( n185 & n2281 ) | ( n1381 & n2281 ) ;
  assign n2283 = n2282 ^ n1251 ^ n976 ;
  assign n2284 = ( x36 & n1621 ) | ( x36 & n2070 ) | ( n1621 & n2070 ) ;
  assign n2285 = ( ~n448 & n2283 ) | ( ~n448 & n2284 ) | ( n2283 & n2284 ) ;
  assign n2286 = ( n1205 & n2280 ) | ( n1205 & n2285 ) | ( n2280 & n2285 ) ;
  assign n2287 = ( ~n949 & n2115 ) | ( ~n949 & n2286 ) | ( n2115 & n2286 ) ;
  assign n2273 = ( n666 & n855 ) | ( n666 & n913 ) | ( n855 & n913 ) ;
  assign n2274 = n1205 ^ n656 ^ n292 ;
  assign n2275 = ( n1575 & ~n2273 ) | ( n1575 & n2274 ) | ( ~n2273 & n2274 ) ;
  assign n2276 = ( ~n1440 & n1958 ) | ( ~n1440 & n2275 ) | ( n1958 & n2275 ) ;
  assign n2289 = n2288 ^ n2287 ^ n2276 ;
  assign n2312 = n2311 ^ n2289 ^ n2185 ;
  assign n2314 = ( ~x58 & n195 ) | ( ~x58 & n264 ) | ( n195 & n264 ) ;
  assign n2313 = n820 ^ n658 ^ n275 ;
  assign n2315 = n2314 ^ n2313 ^ n334 ;
  assign n2316 = n2315 ^ n1491 ^ n935 ;
  assign n2317 = n1419 ^ n1237 ^ n434 ;
  assign n2318 = ( n314 & n1173 ) | ( n314 & ~n2317 ) | ( n1173 & ~n2317 ) ;
  assign n2319 = n2318 ^ n1279 ^ x11 ;
  assign n2320 = ( ~n847 & n980 ) | ( ~n847 & n2319 ) | ( n980 & n2319 ) ;
  assign n2321 = ( n294 & ~n2316 ) | ( n294 & n2320 ) | ( ~n2316 & n2320 ) ;
  assign n2323 = ( n143 & n318 ) | ( n143 & n810 ) | ( n318 & n810 ) ;
  assign n2322 = ( n367 & ~n1298 ) | ( n367 & n1388 ) | ( ~n1298 & n1388 ) ;
  assign n2324 = n2323 ^ n2322 ^ n1343 ;
  assign n2325 = ( n616 & ~n2321 ) | ( n616 & n2324 ) | ( ~n2321 & n2324 ) ;
  assign n2326 = ( n168 & n1412 ) | ( n168 & ~n2325 ) | ( n1412 & ~n2325 ) ;
  assign n2335 = ( n811 & n1335 ) | ( n811 & ~n1635 ) | ( n1335 & ~n1635 ) ;
  assign n2336 = n2335 ^ n2183 ^ n919 ;
  assign n2337 = n2336 ^ n1672 ^ n516 ;
  assign n2327 = ( ~n348 & n711 ) | ( ~n348 & n1177 ) | ( n711 & n1177 ) ;
  assign n2328 = n2327 ^ n855 ^ x7 ;
  assign n2329 = n2328 ^ n1768 ^ n585 ;
  assign n2330 = ( n628 & n653 ) | ( n628 & ~n2329 ) | ( n653 & ~n2329 ) ;
  assign n2331 = ( ~x117 & n320 ) | ( ~x117 & n848 ) | ( n320 & n848 ) ;
  assign n2332 = ( n951 & ~n1508 ) | ( n951 & n2331 ) | ( ~n1508 & n2331 ) ;
  assign n2333 = ( n1024 & ~n2330 ) | ( n1024 & n2332 ) | ( ~n2330 & n2332 ) ;
  assign n2334 = n2333 ^ n1413 ^ n1261 ;
  assign n2338 = n2337 ^ n2334 ^ n335 ;
  assign n2346 = ( n134 & n647 ) | ( n134 & n964 ) | ( n647 & n964 ) ;
  assign n2345 = n1830 ^ n1704 ^ n1178 ;
  assign n2347 = n2346 ^ n2345 ^ n527 ;
  assign n2343 = n802 ^ x117 ^ x94 ;
  assign n2339 = n2014 ^ n391 ^ n357 ;
  assign n2340 = n588 ^ n576 ^ n512 ;
  assign n2341 = n2340 ^ n2254 ^ n963 ;
  assign n2342 = ( n1210 & n2339 ) | ( n1210 & n2341 ) | ( n2339 & n2341 ) ;
  assign n2344 = n2343 ^ n2342 ^ n1390 ;
  assign n2348 = n2347 ^ n2344 ^ n1037 ;
  assign n2349 = ( ~n221 & n1347 ) | ( ~n221 & n2348 ) | ( n1347 & n2348 ) ;
  assign n2350 = ( n2326 & ~n2338 ) | ( n2326 & n2349 ) | ( ~n2338 & n2349 ) ;
  assign n2351 = n1903 ^ n1469 ^ n676 ;
  assign n2374 = ( x125 & n703 ) | ( x125 & n1166 ) | ( n703 & n1166 ) ;
  assign n2373 = n2059 ^ n1056 ^ n532 ;
  assign n2375 = n2374 ^ n2373 ^ n1472 ;
  assign n2376 = n726 ^ n476 ^ n439 ;
  assign n2377 = ( ~x57 & n1406 ) | ( ~x57 & n2376 ) | ( n1406 & n2376 ) ;
  assign n2378 = n2377 ^ n2184 ^ n792 ;
  assign n2379 = n2378 ^ n466 ^ n300 ;
  assign n2380 = ( n369 & n2375 ) | ( n369 & ~n2379 ) | ( n2375 & ~n2379 ) ;
  assign n2364 = n1586 ^ n713 ^ n301 ;
  assign n2368 = ( ~n307 & n485 ) | ( ~n307 & n1267 ) | ( n485 & n1267 ) ;
  assign n2369 = n2368 ^ n1062 ^ n426 ;
  assign n2370 = ( n300 & n572 ) | ( n300 & n2369 ) | ( n572 & n2369 ) ;
  assign n2365 = n2243 ^ n1789 ^ n384 ;
  assign n2366 = ( ~n225 & n311 ) | ( ~n225 & n1304 ) | ( n311 & n1304 ) ;
  assign n2367 = ( n416 & n2365 ) | ( n416 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2371 = n2370 ^ n2367 ^ n1551 ;
  assign n2372 = ( n1805 & n2364 ) | ( n1805 & ~n2371 ) | ( n2364 & ~n2371 ) ;
  assign n2352 = ( n288 & ~n644 ) | ( n288 & n2156 ) | ( ~n644 & n2156 ) ;
  assign n2353 = n2352 ^ n1699 ^ n1111 ;
  assign n2354 = n2175 ^ n720 ^ n544 ;
  assign n2355 = ( n1025 & ~n1643 ) | ( n1025 & n2354 ) | ( ~n1643 & n2354 ) ;
  assign n2357 = ( x88 & n266 ) | ( x88 & n273 ) | ( n266 & n273 ) ;
  assign n2356 = ( n549 & n994 ) | ( n549 & ~n2228 ) | ( n994 & ~n2228 ) ;
  assign n2358 = n2357 ^ n2356 ^ n463 ;
  assign n2359 = ( n1701 & n2355 ) | ( n1701 & n2358 ) | ( n2355 & n2358 ) ;
  assign n2360 = n2359 ^ n2180 ^ n423 ;
  assign n2361 = n2300 ^ n1661 ^ n1047 ;
  assign n2362 = ( n627 & ~n2226 ) | ( n627 & n2361 ) | ( ~n2226 & n2361 ) ;
  assign n2363 = ( n2353 & n2360 ) | ( n2353 & ~n2362 ) | ( n2360 & ~n2362 ) ;
  assign n2381 = n2380 ^ n2372 ^ n2363 ;
  assign n2382 = ( ~n1888 & n2351 ) | ( ~n1888 & n2381 ) | ( n2351 & n2381 ) ;
  assign n2385 = ( x16 & ~n307 ) | ( x16 & n1853 ) | ( ~n307 & n1853 ) ;
  assign n2386 = ( n261 & n590 ) | ( n261 & ~n947 ) | ( n590 & ~n947 ) ;
  assign n2388 = n1769 ^ n1400 ^ x88 ;
  assign n2387 = n1396 ^ n1027 ^ n536 ;
  assign n2389 = n2388 ^ n2387 ^ n988 ;
  assign n2390 = ( n2385 & ~n2386 ) | ( n2385 & n2389 ) | ( ~n2386 & n2389 ) ;
  assign n2391 = n2390 ^ n2221 ^ n1388 ;
  assign n2383 = n1488 ^ n744 ^ n374 ;
  assign n2384 = ( n1127 & ~n1168 ) | ( n1127 & n2383 ) | ( ~n1168 & n2383 ) ;
  assign n2392 = n2391 ^ n2384 ^ n275 ;
  assign n2393 = ( n591 & n728 ) | ( n591 & ~n1198 ) | ( n728 & ~n1198 ) ;
  assign n2394 = ( n389 & n1409 ) | ( n389 & ~n2393 ) | ( n1409 & ~n2393 ) ;
  assign n2423 = n1453 ^ n835 ^ n152 ;
  assign n2420 = ( x116 & n775 ) | ( x116 & ~n1213 ) | ( n775 & ~n1213 ) ;
  assign n2416 = n551 ^ n417 ^ x100 ;
  assign n2417 = ( x118 & n170 ) | ( x118 & ~n1117 ) | ( n170 & ~n1117 ) ;
  assign n2418 = ( x36 & n2416 ) | ( x36 & ~n2417 ) | ( n2416 & ~n2417 ) ;
  assign n2419 = ( n600 & n1024 ) | ( n600 & n2418 ) | ( n1024 & n2418 ) ;
  assign n2421 = n2420 ^ n2419 ^ n239 ;
  assign n2414 = n2207 ^ n1069 ^ n900 ;
  assign n2413 = n1737 ^ n292 ^ n195 ;
  assign n2415 = n2414 ^ n2413 ^ n488 ;
  assign n2408 = ( x43 & n242 ) | ( x43 & ~n437 ) | ( n242 & ~n437 ) ;
  assign n2409 = ( n802 & n1431 ) | ( n802 & ~n2408 ) | ( n1431 & ~n2408 ) ;
  assign n2410 = ( ~n360 & n1735 ) | ( ~n360 & n2409 ) | ( n1735 & n2409 ) ;
  assign n2403 = ( n288 & n385 ) | ( n288 & n1007 ) | ( n385 & n1007 ) ;
  assign n2404 = ( n585 & ~n2151 ) | ( n585 & n2403 ) | ( ~n2151 & n2403 ) ;
  assign n2405 = n2369 ^ n956 ^ n914 ;
  assign n2406 = n2405 ^ n1886 ^ n447 ;
  assign n2407 = ( ~n224 & n2404 ) | ( ~n224 & n2406 ) | ( n2404 & n2406 ) ;
  assign n2411 = n2410 ^ n2407 ^ n1431 ;
  assign n2412 = ( n2035 & n2077 ) | ( n2035 & n2411 ) | ( n2077 & n2411 ) ;
  assign n2422 = n2421 ^ n2415 ^ n2412 ;
  assign n2424 = n2423 ^ n2422 ^ n1863 ;
  assign n2400 = n1215 ^ n685 ^ x61 ;
  assign n2401 = n2400 ^ n762 ^ n212 ;
  assign n2397 = ( n298 & n1545 ) | ( n298 & ~n2068 ) | ( n1545 & ~n2068 ) ;
  assign n2398 = ( n209 & n309 ) | ( n209 & n721 ) | ( n309 & n721 ) ;
  assign n2399 = ( n1172 & n2397 ) | ( n1172 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2395 = n2209 ^ n896 ^ n692 ;
  assign n2396 = n2395 ^ n1475 ^ n1098 ;
  assign n2402 = n2401 ^ n2399 ^ n2396 ;
  assign n2425 = n2424 ^ n2402 ^ n576 ;
  assign n2426 = ( n1464 & n2394 ) | ( n1464 & n2425 ) | ( n2394 & n2425 ) ;
  assign n2427 = n1378 ^ n337 ^ x58 ;
  assign n2430 = ( n287 & n784 ) | ( n287 & ~n851 ) | ( n784 & ~n851 ) ;
  assign n2428 = ( ~n744 & n808 ) | ( ~n744 & n1509 ) | ( n808 & n1509 ) ;
  assign n2429 = n2428 ^ n580 ^ n395 ;
  assign n2431 = n2430 ^ n2429 ^ n1702 ;
  assign n2432 = ( n981 & ~n2427 ) | ( n981 & n2431 ) | ( ~n2427 & n2431 ) ;
  assign n2437 = n2275 ^ n1867 ^ n808 ;
  assign n2433 = ( n1091 & n1336 ) | ( n1091 & ~n1422 ) | ( n1336 & ~n1422 ) ;
  assign n2434 = n2433 ^ n730 ^ n311 ;
  assign n2435 = ( n1382 & ~n2198 ) | ( n1382 & n2434 ) | ( ~n2198 & n2434 ) ;
  assign n2436 = n2435 ^ n1152 ^ n891 ;
  assign n2438 = n2437 ^ n2436 ^ n455 ;
  assign n2439 = ( n1409 & n1551 ) | ( n1409 & n1892 ) | ( n1551 & n1892 ) ;
  assign n2440 = ( ~n1036 & n1177 ) | ( ~n1036 & n2439 ) | ( n1177 & n2439 ) ;
  assign n2441 = ( n306 & n2438 ) | ( n306 & n2440 ) | ( n2438 & n2440 ) ;
  assign n2442 = ( n2322 & ~n2432 ) | ( n2322 & n2441 ) | ( ~n2432 & n2441 ) ;
  assign n2443 = ( n895 & ~n1857 ) | ( n895 & n2442 ) | ( ~n1857 & n2442 ) ;
  assign n2468 = n1768 ^ n879 ^ n489 ;
  assign n2469 = ( ~n1431 & n2197 ) | ( ~n1431 & n2468 ) | ( n2197 & n2468 ) ;
  assign n2461 = ( x99 & ~n796 ) | ( x99 & n2182 ) | ( ~n796 & n2182 ) ;
  assign n2459 = n2420 ^ n1859 ^ n1163 ;
  assign n2457 = ( n755 & ~n961 ) | ( n755 & n1157 ) | ( ~n961 & n1157 ) ;
  assign n2458 = ( n327 & n564 ) | ( n327 & n2457 ) | ( n564 & n2457 ) ;
  assign n2460 = n2459 ^ n2458 ^ n1891 ;
  assign n2462 = n2461 ^ n2460 ^ n604 ;
  assign n2463 = ( ~x32 & x63 ) | ( ~x32 & n917 ) | ( x63 & n917 ) ;
  assign n2464 = n2463 ^ n1349 ^ n312 ;
  assign n2465 = ( n464 & n1000 ) | ( n464 & ~n2464 ) | ( n1000 & ~n2464 ) ;
  assign n2466 = ( n719 & n795 ) | ( n719 & n2465 ) | ( n795 & n2465 ) ;
  assign n2467 = ( n2043 & n2462 ) | ( n2043 & n2466 ) | ( n2462 & n2466 ) ;
  assign n2470 = n2469 ^ n2467 ^ n1597 ;
  assign n2454 = ( ~n743 & n1147 ) | ( ~n743 & n1483 ) | ( n1147 & n1483 ) ;
  assign n2455 = ( n568 & ~n1156 ) | ( n568 & n2454 ) | ( ~n1156 & n2454 ) ;
  assign n2452 = n1026 ^ n279 ^ n192 ;
  assign n2453 = n2452 ^ n2009 ^ n1715 ;
  assign n2449 = n1391 ^ n750 ^ n426 ;
  assign n2446 = ( n134 & n1670 ) | ( n134 & n2259 ) | ( n1670 & n2259 ) ;
  assign n2447 = n2446 ^ n2352 ^ n234 ;
  assign n2448 = ( n485 & n957 ) | ( n485 & ~n2447 ) | ( n957 & ~n2447 ) ;
  assign n2450 = n2449 ^ n2448 ^ n351 ;
  assign n2444 = ( x82 & n887 ) | ( x82 & n917 ) | ( n887 & n917 ) ;
  assign n2445 = ( n1078 & ~n1869 ) | ( n1078 & n2444 ) | ( ~n1869 & n2444 ) ;
  assign n2451 = n2450 ^ n2445 ^ n1805 ;
  assign n2456 = n2455 ^ n2453 ^ n2451 ;
  assign n2471 = n2470 ^ n2456 ^ x60 ;
  assign n2499 = n1124 ^ n456 ^ n372 ;
  assign n2495 = n2449 ^ n1051 ^ n189 ;
  assign n2496 = n2495 ^ n1813 ^ n649 ;
  assign n2497 = ( x46 & n594 ) | ( x46 & n2496 ) | ( n594 & n2496 ) ;
  assign n2498 = ( n621 & ~n2088 ) | ( n621 & n2497 ) | ( ~n2088 & n2497 ) ;
  assign n2489 = ( ~n1060 & n1133 ) | ( ~n1060 & n2045 ) | ( n1133 & n2045 ) ;
  assign n2490 = ( n405 & n485 ) | ( n405 & n2489 ) | ( n485 & n2489 ) ;
  assign n2487 = n529 ^ n300 ^ n186 ;
  assign n2488 = n2487 ^ n1495 ^ x48 ;
  assign n2486 = n2388 ^ n698 ^ x50 ;
  assign n2491 = n2490 ^ n2488 ^ n2486 ;
  assign n2492 = ( n1110 & n1602 ) | ( n1110 & ~n1758 ) | ( n1602 & ~n1758 ) ;
  assign n2493 = ( ~n725 & n2491 ) | ( ~n725 & n2492 ) | ( n2491 & n2492 ) ;
  assign n2484 = n1145 ^ n320 ^ n274 ;
  assign n2482 = ( x117 & ~n701 ) | ( x117 & n2050 ) | ( ~n701 & n2050 ) ;
  assign n2483 = ( n306 & n1954 ) | ( n306 & n2482 ) | ( n1954 & n2482 ) ;
  assign n2480 = n2253 ^ n1198 ^ n601 ;
  assign n2479 = n660 ^ n589 ^ n168 ;
  assign n2481 = n2480 ^ n2479 ^ n786 ;
  assign n2485 = n2484 ^ n2483 ^ n2481 ;
  assign n2472 = n1437 ^ n493 ^ n240 ;
  assign n2475 = n914 ^ n795 ^ n767 ;
  assign n2473 = ( ~x118 & n543 ) | ( ~x118 & n1239 ) | ( n543 & n1239 ) ;
  assign n2474 = ( n249 & n1487 ) | ( n249 & ~n2473 ) | ( n1487 & ~n2473 ) ;
  assign n2476 = n2475 ^ n2474 ^ n1885 ;
  assign n2477 = ( n1043 & n1401 ) | ( n1043 & ~n2476 ) | ( n1401 & ~n2476 ) ;
  assign n2478 = ( ~n1633 & n2472 ) | ( ~n1633 & n2477 ) | ( n2472 & n2477 ) ;
  assign n2494 = n2493 ^ n2485 ^ n2478 ;
  assign n2500 = n2499 ^ n2498 ^ n2494 ;
  assign n2501 = ( ~n198 & n330 ) | ( ~n198 & n896 ) | ( n330 & n896 ) ;
  assign n2502 = n2501 ^ n2331 ^ n631 ;
  assign n2503 = n2202 ^ n495 ^ n321 ;
  assign n2504 = n594 ^ n229 ^ x67 ;
  assign n2505 = ( n192 & n229 ) | ( n192 & n1196 ) | ( n229 & n1196 ) ;
  assign n2506 = n2505 ^ n1370 ^ n380 ;
  assign n2507 = ( n1042 & n2504 ) | ( n1042 & ~n2506 ) | ( n2504 & ~n2506 ) ;
  assign n2508 = ( n1731 & n2503 ) | ( n1731 & ~n2507 ) | ( n2503 & ~n2507 ) ;
  assign n2509 = n2352 ^ n1477 ^ n1209 ;
  assign n2510 = ( n2502 & n2508 ) | ( n2502 & ~n2509 ) | ( n2508 & ~n2509 ) ;
  assign n2541 = ( x58 & n650 ) | ( x58 & n1180 ) | ( n650 & n1180 ) ;
  assign n2542 = ( n744 & ~n1186 ) | ( n744 & n2541 ) | ( ~n1186 & n2541 ) ;
  assign n2535 = ( x92 & n318 ) | ( x92 & n2250 ) | ( n318 & n2250 ) ;
  assign n2536 = ( x113 & n1325 ) | ( x113 & n2535 ) | ( n1325 & n2535 ) ;
  assign n2537 = n1629 ^ n1013 ^ n523 ;
  assign n2538 = n2537 ^ n1662 ^ n310 ;
  assign n2539 = ( x113 & n493 ) | ( x113 & ~n1589 ) | ( n493 & ~n1589 ) ;
  assign n2540 = ( n2536 & n2538 ) | ( n2536 & ~n2539 ) | ( n2538 & ~n2539 ) ;
  assign n2543 = n2542 ^ n2540 ^ n1988 ;
  assign n2511 = ( n141 & ~n725 ) | ( n141 & n902 ) | ( ~n725 & n902 ) ;
  assign n2512 = n540 ^ n233 ^ n185 ;
  assign n2513 = ( n236 & n249 ) | ( n236 & n2512 ) | ( n249 & n2512 ) ;
  assign n2514 = ( n739 & n880 ) | ( n739 & ~n2513 ) | ( n880 & ~n2513 ) ;
  assign n2515 = n2514 ^ n1429 ^ x90 ;
  assign n2516 = ( x21 & n2511 ) | ( x21 & n2515 ) | ( n2511 & n2515 ) ;
  assign n2517 = ( n246 & n1167 ) | ( n246 & ~n2070 ) | ( n1167 & ~n2070 ) ;
  assign n2518 = n1432 ^ n658 ^ n533 ;
  assign n2519 = n2254 ^ n2103 ^ n1444 ;
  assign n2520 = ( x126 & n2518 ) | ( x126 & n2519 ) | ( n2518 & n2519 ) ;
  assign n2521 = ( x82 & ~n453 ) | ( x82 & n2520 ) | ( ~n453 & n2520 ) ;
  assign n2522 = ( n726 & n1464 ) | ( n726 & ~n2521 ) | ( n1464 & ~n2521 ) ;
  assign n2525 = n1486 ^ n1024 ^ x82 ;
  assign n2524 = n1634 ^ n220 ^ n163 ;
  assign n2523 = ( n738 & n894 ) | ( n738 & n1068 ) | ( n894 & n1068 ) ;
  assign n2526 = n2525 ^ n2524 ^ n2523 ;
  assign n2527 = n1230 ^ n622 ^ n438 ;
  assign n2528 = ( n1603 & n2221 ) | ( n1603 & ~n2527 ) | ( n2221 & ~n2527 ) ;
  assign n2529 = ( n1268 & n1854 ) | ( n1268 & n2102 ) | ( n1854 & n2102 ) ;
  assign n2530 = n2125 ^ n856 ^ n178 ;
  assign n2531 = ( x112 & n617 ) | ( x112 & ~n2530 ) | ( n617 & ~n2530 ) ;
  assign n2532 = ( n2528 & ~n2529 ) | ( n2528 & n2531 ) | ( ~n2529 & n2531 ) ;
  assign n2533 = ( n2522 & ~n2526 ) | ( n2522 & n2532 ) | ( ~n2526 & n2532 ) ;
  assign n2534 = ( n2516 & n2517 ) | ( n2516 & n2533 ) | ( n2517 & n2533 ) ;
  assign n2544 = n2543 ^ n2534 ^ n526 ;
  assign n2549 = n1177 ^ n883 ^ n763 ;
  assign n2545 = ( ~n907 & n1088 ) | ( ~n907 & n2007 ) | ( n1088 & n2007 ) ;
  assign n2546 = ( n148 & n788 ) | ( n148 & n2545 ) | ( n788 & n2545 ) ;
  assign n2547 = n2546 ^ n750 ^ n452 ;
  assign n2548 = ( n2273 & n2307 ) | ( n2273 & ~n2547 ) | ( n2307 & ~n2547 ) ;
  assign n2550 = n2549 ^ n2548 ^ n2369 ;
  assign n2551 = n2550 ^ n2464 ^ n1773 ;
  assign n2612 = n1870 ^ n1721 ^ n474 ;
  assign n2607 = ( n681 & ~n1102 ) | ( n681 & n1334 ) | ( ~n1102 & n1334 ) ;
  assign n2608 = ( n422 & n1296 ) | ( n422 & ~n2607 ) | ( n1296 & ~n2607 ) ;
  assign n2606 = n677 ^ n615 ^ n409 ;
  assign n2609 = n2608 ^ n2606 ^ n2250 ;
  assign n2610 = ( ~n1576 & n2479 ) | ( ~n1576 & n2609 ) | ( n2479 & n2609 ) ;
  assign n2603 = ( n134 & n428 ) | ( n134 & ~n1332 ) | ( n428 & ~n1332 ) ;
  assign n2602 = n1841 ^ n1288 ^ x64 ;
  assign n2604 = n2603 ^ n2602 ^ n1096 ;
  assign n2605 = ( n999 & n1848 ) | ( n999 & n2604 ) | ( n1848 & n2604 ) ;
  assign n2611 = n2610 ^ n2605 ^ n579 ;
  assign n2600 = n2010 ^ n1972 ^ x37 ;
  assign n2594 = n1860 ^ n796 ^ n493 ;
  assign n2595 = n2594 ^ n1077 ^ n379 ;
  assign n2596 = ( ~n1411 & n1515 ) | ( ~n1411 & n2595 ) | ( n1515 & n2595 ) ;
  assign n2597 = n287 ^ n240 ^ n170 ;
  assign n2598 = ( n1919 & ~n2331 ) | ( n1919 & n2597 ) | ( ~n2331 & n2597 ) ;
  assign n2599 = ( n2117 & ~n2596 ) | ( n2117 & n2598 ) | ( ~n2596 & n2598 ) ;
  assign n2591 = ( n203 & n373 ) | ( n203 & n489 ) | ( n373 & n489 ) ;
  assign n2592 = ( x99 & n138 ) | ( x99 & n2591 ) | ( n138 & n2591 ) ;
  assign n2578 = n1934 ^ n582 ^ n515 ;
  assign n2579 = n2436 ^ n504 ^ x86 ;
  assign n2583 = ( x125 & ~n491 ) | ( x125 & n634 ) | ( ~n491 & n634 ) ;
  assign n2584 = n2583 ^ n1134 ^ n612 ;
  assign n2585 = n2584 ^ n550 ^ n166 ;
  assign n2580 = ( n202 & ~n1877 ) | ( n202 & n1883 ) | ( ~n1877 & n1883 ) ;
  assign n2581 = ( n377 & n471 ) | ( n377 & n2580 ) | ( n471 & n2580 ) ;
  assign n2582 = ( n2105 & n2446 ) | ( n2105 & n2581 ) | ( n2446 & n2581 ) ;
  assign n2586 = n2585 ^ n2582 ^ n1332 ;
  assign n2587 = ( n2578 & n2579 ) | ( n2578 & n2586 ) | ( n2579 & n2586 ) ;
  assign n2588 = ( n190 & n2052 ) | ( n190 & n2587 ) | ( n2052 & n2587 ) ;
  assign n2589 = n2588 ^ n1102 ^ n228 ;
  assign n2590 = ( n1181 & ~n1198 ) | ( n1181 & n2589 ) | ( ~n1198 & n2589 ) ;
  assign n2574 = ( n666 & ~n1592 ) | ( n666 & n1853 ) | ( ~n1592 & n1853 ) ;
  assign n2575 = n2574 ^ n1356 ^ n695 ;
  assign n2572 = n1274 ^ n776 ^ x115 ;
  assign n2569 = ( n191 & n1098 ) | ( n191 & ~n2265 ) | ( n1098 & ~n2265 ) ;
  assign n2568 = n593 ^ n500 ^ n247 ;
  assign n2570 = n2569 ^ n2568 ^ n579 ;
  assign n2571 = n2570 ^ n682 ^ n636 ;
  assign n2563 = ( n610 & n1002 ) | ( n610 & n1448 ) | ( n1002 & n1448 ) ;
  assign n2564 = n2563 ^ n2256 ^ n1350 ;
  assign n2565 = ( ~x120 & n1001 ) | ( ~x120 & n2564 ) | ( n1001 & n2564 ) ;
  assign n2566 = n2565 ^ n1404 ^ n625 ;
  assign n2552 = n1719 ^ n821 ^ n290 ;
  assign n2556 = n1279 ^ n690 ^ x49 ;
  assign n2553 = ( n214 & n259 ) | ( n214 & n1629 ) | ( n259 & n1629 ) ;
  assign n2554 = n2553 ^ n1534 ^ n278 ;
  assign n2555 = ( n729 & ~n2416 ) | ( n729 & n2554 ) | ( ~n2416 & n2554 ) ;
  assign n2557 = n2556 ^ n2555 ^ n2109 ;
  assign n2558 = n2557 ^ n1594 ^ n177 ;
  assign n2559 = ( ~n991 & n2552 ) | ( ~n991 & n2558 ) | ( n2552 & n2558 ) ;
  assign n2560 = n2559 ^ n638 ^ n237 ;
  assign n2561 = ( n847 & n1167 ) | ( n847 & ~n2560 ) | ( n1167 & ~n2560 ) ;
  assign n2562 = ( n840 & n2194 ) | ( n840 & n2561 ) | ( n2194 & n2561 ) ;
  assign n2567 = n2566 ^ n2562 ^ n405 ;
  assign n2573 = n2572 ^ n2571 ^ n2567 ;
  assign n2576 = n2575 ^ n2573 ^ n338 ;
  assign n2577 = n2576 ^ n236 ^ x55 ;
  assign n2593 = n2592 ^ n2590 ^ n2577 ;
  assign n2601 = n2600 ^ n2599 ^ n2593 ;
  assign n2613 = n2612 ^ n2611 ^ n2601 ;
  assign n2614 = n1267 ^ n375 ^ n130 ;
  assign n2616 = ( ~n700 & n1293 ) | ( ~n700 & n2256 ) | ( n1293 & n2256 ) ;
  assign n2615 = ( n951 & n1300 ) | ( n951 & ~n2104 ) | ( n1300 & ~n2104 ) ;
  assign n2617 = n2616 ^ n2615 ^ n1817 ;
  assign n2618 = ( n2327 & ~n2614 ) | ( n2327 & n2617 ) | ( ~n2614 & n2617 ) ;
  assign n2619 = n938 ^ n192 ^ x90 ;
  assign n2620 = ( n834 & n2022 ) | ( n834 & n2619 ) | ( n2022 & n2619 ) ;
  assign n2621 = n1237 ^ n656 ^ n332 ;
  assign n2622 = n2621 ^ n1313 ^ n400 ;
  assign n2623 = n2622 ^ n871 ^ n625 ;
  assign n2624 = ( n833 & ~n2620 ) | ( n833 & n2623 ) | ( ~n2620 & n2623 ) ;
  assign n2625 = n2624 ^ n2215 ^ n1430 ;
  assign n2639 = ( x60 & n135 ) | ( x60 & ~n1772 ) | ( n135 & ~n1772 ) ;
  assign n2628 = ( x78 & n716 ) | ( x78 & ~n857 ) | ( n716 & ~n857 ) ;
  assign n2627 = n1505 ^ n492 ^ n444 ;
  assign n2626 = n2501 ^ n1218 ^ n873 ;
  assign n2629 = n2628 ^ n2627 ^ n2626 ;
  assign n2630 = ( n527 & n1978 ) | ( n527 & ~n2629 ) | ( n1978 & ~n2629 ) ;
  assign n2631 = ( n1000 & n1069 ) | ( n1000 & ~n1762 ) | ( n1069 & ~n1762 ) ;
  assign n2632 = ( n347 & n2059 ) | ( n347 & ~n2631 ) | ( n2059 & ~n2631 ) ;
  assign n2633 = n2632 ^ n2051 ^ x124 ;
  assign n2634 = ( n178 & n800 ) | ( n178 & n2160 ) | ( n800 & n2160 ) ;
  assign n2635 = ( ~n1297 & n2633 ) | ( ~n1297 & n2634 ) | ( n2633 & n2634 ) ;
  assign n2636 = n2631 ^ n1791 ^ n1341 ;
  assign n2637 = ( n1902 & ~n2635 ) | ( n1902 & n2636 ) | ( ~n2635 & n2636 ) ;
  assign n2638 = ( ~n778 & n2630 ) | ( ~n778 & n2637 ) | ( n2630 & n2637 ) ;
  assign n2640 = n2639 ^ n2638 ^ n2176 ;
  assign n2642 = n1102 ^ n581 ^ n274 ;
  assign n2641 = n729 ^ n633 ^ n563 ;
  assign n2643 = n2642 ^ n2641 ^ n2131 ;
  assign n2644 = n2307 ^ x62 ^ x32 ;
  assign n2645 = ( n199 & n526 ) | ( n199 & n2644 ) | ( n526 & n2644 ) ;
  assign n2646 = ( n738 & n1176 ) | ( n738 & n1280 ) | ( n1176 & n1280 ) ;
  assign n2647 = n2646 ^ n1167 ^ n402 ;
  assign n2648 = ( n998 & n1110 ) | ( n998 & n2647 ) | ( n1110 & n2647 ) ;
  assign n2649 = ( n942 & ~n1782 ) | ( n942 & n2142 ) | ( ~n1782 & n2142 ) ;
  assign n2650 = n2649 ^ n1298 ^ n976 ;
  assign n2651 = ( ~n280 & n363 ) | ( ~n280 & n2650 ) | ( n363 & n2650 ) ;
  assign n2652 = ( n2645 & ~n2648 ) | ( n2645 & n2651 ) | ( ~n2648 & n2651 ) ;
  assign n2653 = ( n1485 & n2643 ) | ( n1485 & ~n2652 ) | ( n2643 & ~n2652 ) ;
  assign n2654 = ( n423 & n1056 ) | ( n423 & n2468 ) | ( n1056 & n2468 ) ;
  assign n2655 = n2654 ^ n1227 ^ n1223 ;
  assign n2697 = ( n475 & n739 ) | ( n475 & n1304 ) | ( n739 & n1304 ) ;
  assign n2698 = ( n544 & n1627 ) | ( n544 & ~n2697 ) | ( n1627 & ~n2697 ) ;
  assign n2699 = ( n1000 & n2314 ) | ( n1000 & ~n2698 ) | ( n2314 & ~n2698 ) ;
  assign n2684 = n878 ^ n593 ^ n198 ;
  assign n2685 = n2684 ^ n1433 ^ n173 ;
  assign n2686 = n2685 ^ n2527 ^ n1700 ;
  assign n2687 = n454 ^ n277 ^ x46 ;
  assign n2688 = ( x105 & ~n1179 ) | ( x105 & n2687 ) | ( ~n1179 & n2687 ) ;
  assign n2689 = n2688 ^ n858 ^ n483 ;
  assign n2692 = ( x59 & ~n182 ) | ( x59 & n505 ) | ( ~n182 & n505 ) ;
  assign n2693 = n998 ^ n387 ^ x51 ;
  assign n2694 = ( n501 & n2692 ) | ( n501 & ~n2693 ) | ( n2692 & ~n2693 ) ;
  assign n2690 = ( n553 & ~n941 ) | ( n553 & n1023 ) | ( ~n941 & n1023 ) ;
  assign n2691 = ( ~n1179 & n1623 ) | ( ~n1179 & n2690 ) | ( n1623 & n2690 ) ;
  assign n2695 = n2694 ^ n2691 ^ n2438 ;
  assign n2696 = ( n2686 & n2689 ) | ( n2686 & n2695 ) | ( n2689 & n2695 ) ;
  assign n2680 = ( n226 & n472 ) | ( n226 & ~n1381 ) | ( n472 & ~n1381 ) ;
  assign n2681 = ( ~n947 & n1361 ) | ( ~n947 & n2680 ) | ( n1361 & n2680 ) ;
  assign n2682 = n2681 ^ n2366 ^ n970 ;
  assign n2659 = n1289 ^ n1140 ^ n599 ;
  assign n2660 = ( ~x38 & n868 ) | ( ~x38 & n1595 ) | ( n868 & n1595 ) ;
  assign n2661 = n1799 ^ n847 ^ n517 ;
  assign n2662 = ( n956 & n1967 ) | ( n956 & n2661 ) | ( n1967 & n2661 ) ;
  assign n2663 = n2662 ^ n1678 ^ n819 ;
  assign n2664 = ( ~n2535 & n2660 ) | ( ~n2535 & n2663 ) | ( n2660 & n2663 ) ;
  assign n2665 = ( ~n507 & n2659 ) | ( ~n507 & n2664 ) | ( n2659 & n2664 ) ;
  assign n2673 = ( ~n229 & n394 ) | ( ~n229 & n830 ) | ( n394 & n830 ) ;
  assign n2674 = n424 ^ n255 ^ x38 ;
  assign n2675 = ( n881 & ~n887 ) | ( n881 & n2674 ) | ( ~n887 & n2674 ) ;
  assign n2676 = ( ~n1147 & n2673 ) | ( ~n1147 & n2675 ) | ( n2673 & n2675 ) ;
  assign n2666 = ( x26 & ~n533 ) | ( x26 & n578 ) | ( ~n533 & n578 ) ;
  assign n2667 = n2666 ^ n784 ^ n546 ;
  assign n2668 = ( n847 & n1561 ) | ( n847 & ~n1634 ) | ( n1561 & ~n1634 ) ;
  assign n2669 = ( n1475 & ~n2327 ) | ( n1475 & n2628 ) | ( ~n2327 & n2628 ) ;
  assign n2670 = n2669 ^ n1150 ^ n301 ;
  assign n2671 = n2670 ^ n2444 ^ n1214 ;
  assign n2672 = ( n2667 & n2668 ) | ( n2667 & n2671 ) | ( n2668 & n2671 ) ;
  assign n2677 = n2676 ^ n2672 ^ n2266 ;
  assign n2678 = ( n1229 & n2665 ) | ( n1229 & n2677 ) | ( n2665 & n2677 ) ;
  assign n2656 = ( ~n131 & n163 ) | ( ~n131 & n469 ) | ( n163 & n469 ) ;
  assign n2657 = ( n591 & ~n2515 ) | ( n591 & n2656 ) | ( ~n2515 & n2656 ) ;
  assign n2658 = n2657 ^ n1690 ^ n1591 ;
  assign n2679 = n2678 ^ n2658 ^ n1811 ;
  assign n2683 = n2682 ^ n2679 ^ n2530 ;
  assign n2700 = n2699 ^ n2696 ^ n2683 ;
  assign n2705 = ( n898 & n2553 ) | ( n898 & n2671 ) | ( n2553 & n2671 ) ;
  assign n2701 = n2554 ^ n1698 ^ n1631 ;
  assign n2702 = n1375 ^ n711 ^ n686 ;
  assign n2703 = ( n254 & ~n1129 ) | ( n254 & n1284 ) | ( ~n1129 & n1284 ) ;
  assign n2704 = ( ~n2701 & n2702 ) | ( ~n2701 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2706 = n2705 ^ n2704 ^ n2528 ;
  assign n2707 = n2453 ^ n2104 ^ n378 ;
  assign n2708 = ( n530 & n2146 ) | ( n530 & n2707 ) | ( n2146 & n2707 ) ;
  assign n2709 = ( n1556 & ~n2706 ) | ( n1556 & n2708 ) | ( ~n2706 & n2708 ) ;
  assign n2715 = ( n840 & n1816 ) | ( n840 & n1823 ) | ( n1816 & n1823 ) ;
  assign n2710 = ( ~x27 & n227 ) | ( ~x27 & n2115 ) | ( n227 & n2115 ) ;
  assign n2711 = ( n1111 & n1670 ) | ( n1111 & ~n2710 ) | ( n1670 & ~n2710 ) ;
  assign n2712 = n1621 ^ n1162 ^ n598 ;
  assign n2713 = n2712 ^ n1965 ^ n481 ;
  assign n2714 = ( ~n534 & n2711 ) | ( ~n534 & n2713 ) | ( n2711 & n2713 ) ;
  assign n2716 = n2715 ^ n2714 ^ n1275 ;
  assign n2717 = n1818 ^ n1595 ^ x126 ;
  assign n2718 = n2717 ^ n1140 ^ x49 ;
  assign n2722 = ( n564 & ~n1322 ) | ( n564 & n2068 ) | ( ~n1322 & n2068 ) ;
  assign n2723 = ( n1276 & ~n1496 ) | ( n1276 & n2722 ) | ( ~n1496 & n2722 ) ;
  assign n2719 = ( x2 & ~n765 ) | ( x2 & n2253 ) | ( ~n765 & n2253 ) ;
  assign n2720 = n2719 ^ n2280 ^ n493 ;
  assign n2721 = ( ~n226 & n833 ) | ( ~n226 & n2720 ) | ( n833 & n2720 ) ;
  assign n2724 = n2723 ^ n2721 ^ n2226 ;
  assign n2725 = ( n979 & n2718 ) | ( n979 & n2724 ) | ( n2718 & n2724 ) ;
  assign n2726 = ( x34 & n1248 ) | ( x34 & n1251 ) | ( n1248 & n1251 ) ;
  assign n2727 = n2726 ^ n1926 ^ n422 ;
  assign n2728 = ( n928 & n2725 ) | ( n928 & n2727 ) | ( n2725 & n2727 ) ;
  assign n2729 = n2728 ^ n2278 ^ n1818 ;
  assign n2730 = n2292 ^ n1290 ^ n944 ;
  assign n2731 = ( n144 & ~n1712 ) | ( n144 & n2730 ) | ( ~n1712 & n2730 ) ;
  assign n2732 = n2095 ^ n1557 ^ n1285 ;
  assign n2737 = ( n962 & n1644 ) | ( n962 & n2056 ) | ( n1644 & n2056 ) ;
  assign n2733 = ( n570 & n2212 ) | ( n570 & ~n2457 ) | ( n2212 & ~n2457 ) ;
  assign n2734 = n2733 ^ n2674 ^ n879 ;
  assign n2735 = n2734 ^ n1836 ^ n1474 ;
  assign n2736 = n2735 ^ n2600 ^ n1197 ;
  assign n2738 = n2737 ^ n2736 ^ n2626 ;
  assign n2739 = ( n1129 & n2732 ) | ( n1129 & ~n2738 ) | ( n2732 & ~n2738 ) ;
  assign n2740 = ( n470 & n2731 ) | ( n470 & n2739 ) | ( n2731 & n2739 ) ;
  assign n2753 = n1838 ^ n1132 ^ n620 ;
  assign n2754 = n2753 ^ n1068 ^ x18 ;
  assign n2755 = n2754 ^ n2140 ^ n604 ;
  assign n2752 = ( ~n494 & n587 ) | ( ~n494 & n2501 ) | ( n587 & n2501 ) ;
  assign n2750 = ( n1269 & ~n2091 ) | ( n1269 & n2434 ) | ( ~n2091 & n2434 ) ;
  assign n2744 = n747 ^ n652 ^ n625 ;
  assign n2745 = n729 ^ n359 ^ n294 ;
  assign n2746 = ( x113 & ~n1078 ) | ( x113 & n2210 ) | ( ~n1078 & n2210 ) ;
  assign n2747 = ( ~n2744 & n2745 ) | ( ~n2744 & n2746 ) | ( n2745 & n2746 ) ;
  assign n2741 = ( ~x53 & n1276 ) | ( ~x53 & n1504 ) | ( n1276 & n1504 ) ;
  assign n2742 = ( n1434 & n2087 ) | ( n1434 & ~n2741 ) | ( n2087 & ~n2741 ) ;
  assign n2743 = n2742 ^ n1171 ^ n662 ;
  assign n2748 = n2747 ^ n2743 ^ n1053 ;
  assign n2749 = ( ~n645 & n2315 ) | ( ~n645 & n2748 ) | ( n2315 & n2748 ) ;
  assign n2751 = n2750 ^ n2749 ^ n2573 ;
  assign n2756 = n2755 ^ n2752 ^ n2751 ;
  assign n2757 = n2691 ^ n2198 ^ n619 ;
  assign n2758 = n2757 ^ n1173 ^ x17 ;
  assign n2759 = ( ~n547 & n700 ) | ( ~n547 & n1272 ) | ( n700 & n1272 ) ;
  assign n2760 = n2759 ^ n668 ^ x45 ;
  assign n2761 = ( ~n804 & n2205 ) | ( ~n804 & n2760 ) | ( n2205 & n2760 ) ;
  assign n2762 = n1073 ^ n1045 ^ n389 ;
  assign n2763 = ( n433 & ~n1604 ) | ( n433 & n2762 ) | ( ~n1604 & n2762 ) ;
  assign n2764 = ( n1434 & ~n1462 ) | ( n1434 & n1577 ) | ( ~n1462 & n1577 ) ;
  assign n2765 = n2764 ^ n1271 ^ n392 ;
  assign n2766 = n2765 ^ n2224 ^ n620 ;
  assign n2767 = ( n2529 & n2763 ) | ( n2529 & ~n2766 ) | ( n2763 & ~n2766 ) ;
  assign n2768 = n2767 ^ n623 ^ x72 ;
  assign n2769 = n2384 ^ n2055 ^ n1594 ;
  assign n2770 = ( ~n2761 & n2768 ) | ( ~n2761 & n2769 ) | ( n2768 & n2769 ) ;
  assign n2771 = ( n259 & n483 ) | ( n259 & n521 ) | ( n483 & n521 ) ;
  assign n2772 = n2771 ^ n698 ^ n306 ;
  assign n2773 = n2772 ^ n1405 ^ n337 ;
  assign n2774 = ( ~n631 & n2608 ) | ( ~n631 & n2773 ) | ( n2608 & n2773 ) ;
  assign n2775 = ( n2758 & ~n2770 ) | ( n2758 & n2774 ) | ( ~n2770 & n2774 ) ;
  assign n2821 = n1839 ^ n1075 ^ n313 ;
  assign n2818 = ( ~n369 & n1237 ) | ( ~n369 & n2343 ) | ( n1237 & n2343 ) ;
  assign n2819 = ( n333 & n1046 ) | ( n333 & ~n2818 ) | ( n1046 & ~n2818 ) ;
  assign n2817 = ( n748 & n1828 ) | ( n748 & n2594 ) | ( n1828 & n2594 ) ;
  assign n2820 = n2819 ^ n2817 ^ n310 ;
  assign n2822 = n2821 ^ n2820 ^ x53 ;
  assign n2815 = n2208 ^ n587 ^ n439 ;
  assign n2794 = ( x115 & n139 ) | ( x115 & n761 ) | ( n139 & n761 ) ;
  assign n2812 = ( n586 & n734 ) | ( n586 & n864 ) | ( n734 & n864 ) ;
  assign n2813 = ( n614 & ~n715 ) | ( n614 & n2644 ) | ( ~n715 & n2644 ) ;
  assign n2814 = ( n2794 & n2812 ) | ( n2794 & ~n2813 ) | ( n2812 & ~n2813 ) ;
  assign n2809 = ( ~x49 & n1099 ) | ( ~x49 & n1871 ) | ( n1099 & n1871 ) ;
  assign n2807 = ( n221 & n1148 ) | ( n221 & n2366 ) | ( n1148 & n2366 ) ;
  assign n2808 = n2807 ^ n2150 ^ n441 ;
  assign n2810 = n2809 ^ n2808 ^ n1174 ;
  assign n2803 = ( n651 & n746 ) | ( n651 & ~n1053 ) | ( n746 & ~n1053 ) ;
  assign n2804 = n2803 ^ n2280 ^ n2023 ;
  assign n2802 = n1012 ^ n694 ^ n257 ;
  assign n2805 = n2804 ^ n2802 ^ n2749 ;
  assign n2806 = n2805 ^ n1834 ^ n1829 ;
  assign n2811 = n2810 ^ n2806 ^ n1074 ;
  assign n2816 = n2815 ^ n2814 ^ n2811 ;
  assign n2776 = ( ~n450 & n1115 ) | ( ~n450 & n1278 ) | ( n1115 & n1278 ) ;
  assign n2795 = n2794 ^ n1674 ^ n816 ;
  assign n2792 = ( ~x21 & n186 ) | ( ~x21 & n1052 ) | ( n186 & n1052 ) ;
  assign n2793 = n2792 ^ n494 ^ n289 ;
  assign n2796 = n2795 ^ n2793 ^ n2051 ;
  assign n2797 = n2223 ^ n1693 ^ n240 ;
  assign n2798 = ( n234 & n1733 ) | ( n234 & n2797 ) | ( n1733 & n2797 ) ;
  assign n2799 = ( n1063 & ~n2796 ) | ( n1063 & n2798 ) | ( ~n2796 & n2798 ) ;
  assign n2790 = n1005 ^ n811 ^ n371 ;
  assign n2791 = ( ~n1314 & n2102 ) | ( ~n1314 & n2790 ) | ( n2102 & n2790 ) ;
  assign n2788 = ( n217 & n511 ) | ( n217 & n845 ) | ( n511 & n845 ) ;
  assign n2783 = ( ~n170 & n311 ) | ( ~n170 & n512 ) | ( n311 & n512 ) ;
  assign n2784 = n1464 ^ n186 ^ x19 ;
  assign n2785 = ( n1867 & ~n2783 ) | ( n1867 & n2784 ) | ( ~n2783 & n2784 ) ;
  assign n2781 = ( ~n953 & n957 ) | ( ~n953 & n2029 ) | ( n957 & n2029 ) ;
  assign n2782 = n2781 ^ n2112 ^ n1418 ;
  assign n2786 = n2785 ^ n2782 ^ n1173 ;
  assign n2787 = n2786 ^ n1781 ^ n1706 ;
  assign n2777 = ( n408 & n533 ) | ( n408 & ~n787 ) | ( n533 & ~n787 ) ;
  assign n2778 = n2777 ^ n396 ^ n297 ;
  assign n2779 = n2778 ^ n1233 ^ n886 ;
  assign n2780 = ( n265 & n2733 ) | ( n265 & n2779 ) | ( n2733 & n2779 ) ;
  assign n2789 = n2788 ^ n2787 ^ n2780 ;
  assign n2800 = n2799 ^ n2791 ^ n2789 ;
  assign n2801 = ( n1146 & n2776 ) | ( n1146 & n2800 ) | ( n2776 & n2800 ) ;
  assign n2823 = n2822 ^ n2816 ^ n2801 ;
  assign n2824 = n2128 ^ n1091 ^ n254 ;
  assign n2825 = ( n300 & ~n2487 ) | ( n300 & n2824 ) | ( ~n2487 & n2824 ) ;
  assign n2830 = ( ~n571 & n1448 ) | ( ~n571 & n1466 ) | ( n1448 & n1466 ) ;
  assign n2831 = ( n1866 & n2730 ) | ( n1866 & ~n2830 ) | ( n2730 & ~n2830 ) ;
  assign n2826 = ( ~n748 & n1551 ) | ( ~n748 & n2499 ) | ( n1551 & n2499 ) ;
  assign n2827 = ( ~n1376 & n2275 ) | ( ~n1376 & n2826 ) | ( n2275 & n2826 ) ;
  assign n2828 = ( ~n872 & n2009 ) | ( ~n872 & n2827 ) | ( n2009 & n2827 ) ;
  assign n2829 = n2828 ^ n647 ^ n591 ;
  assign n2832 = n2831 ^ n2829 ^ n471 ;
  assign n2833 = n2832 ^ n2777 ^ n254 ;
  assign n2844 = ( n148 & n932 ) | ( n148 & n2298 ) | ( n932 & n2298 ) ;
  assign n2845 = ( ~n273 & n2773 ) | ( ~n273 & n2844 ) | ( n2773 & n2844 ) ;
  assign n2846 = ( ~n1393 & n1902 ) | ( ~n1393 & n2845 ) | ( n1902 & n2845 ) ;
  assign n2834 = n2546 ^ n1021 ^ n672 ;
  assign n2835 = n2834 ^ n2329 ^ n1201 ;
  assign n2836 = ( n470 & n979 ) | ( n470 & ~n1929 ) | ( n979 & ~n1929 ) ;
  assign n2837 = n1851 ^ n1814 ^ n288 ;
  assign n2838 = ( ~n1271 & n2742 ) | ( ~n1271 & n2837 ) | ( n2742 & n2837 ) ;
  assign n2840 = n835 ^ n489 ^ n271 ;
  assign n2839 = ( x61 & ~n361 ) | ( x61 & n623 ) | ( ~n361 & n623 ) ;
  assign n2841 = n2840 ^ n2839 ^ n1850 ;
  assign n2842 = ( n2836 & ~n2838 ) | ( n2836 & n2841 ) | ( ~n2838 & n2841 ) ;
  assign n2843 = ( n1304 & n2835 ) | ( n1304 & ~n2842 ) | ( n2835 & ~n2842 ) ;
  assign n2847 = n2846 ^ n2843 ^ n913 ;
  assign n2848 = ( n632 & n950 ) | ( n632 & ~n1877 ) | ( n950 & ~n1877 ) ;
  assign n2849 = n1707 ^ n499 ^ n342 ;
  assign n2850 = ( ~n2339 & n2848 ) | ( ~n2339 & n2849 ) | ( n2848 & n2849 ) ;
  assign n2851 = ( n1529 & ~n1748 ) | ( n1529 & n2850 ) | ( ~n1748 & n2850 ) ;
  assign n2889 = n2262 ^ n1897 ^ x75 ;
  assign n2890 = n2687 ^ n2300 ^ n129 ;
  assign n2891 = n2890 ^ n859 ^ x124 ;
  assign n2892 = n2891 ^ n1170 ^ n329 ;
  assign n2893 = ( ~n1801 & n2889 ) | ( ~n1801 & n2892 ) | ( n2889 & n2892 ) ;
  assign n2894 = n2893 ^ n2759 ^ n778 ;
  assign n2885 = ( n806 & n986 ) | ( n806 & ~n1389 ) | ( n986 & ~n1389 ) ;
  assign n2886 = n2885 ^ n807 ^ n722 ;
  assign n2883 = ( x13 & n1901 ) | ( x13 & n2041 ) | ( n1901 & n2041 ) ;
  assign n2884 = n2883 ^ n1656 ^ x9 ;
  assign n2887 = n2886 ^ n2884 ^ n1143 ;
  assign n2879 = ( ~x30 & x117 ) | ( ~x30 & n787 ) | ( x117 & n787 ) ;
  assign n2880 = n1414 ^ n1080 ^ x59 ;
  assign n2881 = ( n1130 & n2879 ) | ( n1130 & ~n2880 ) | ( n2879 & ~n2880 ) ;
  assign n2882 = ( ~n287 & n978 ) | ( ~n287 & n2881 ) | ( n978 & n2881 ) ;
  assign n2876 = ( ~n299 & n2104 ) | ( ~n299 & n2347 ) | ( n2104 & n2347 ) ;
  assign n2877 = n2876 ^ n935 ^ x121 ;
  assign n2867 = ( n755 & n988 ) | ( n755 & ~n1161 ) | ( n988 & ~n1161 ) ;
  assign n2872 = ( n1083 & n2256 ) | ( n1083 & ~n2418 ) | ( n2256 & ~n2418 ) ;
  assign n2871 = ( n822 & n1355 ) | ( n822 & n2750 ) | ( n1355 & n2750 ) ;
  assign n2868 = ( ~n676 & n1512 ) | ( ~n676 & n2369 ) | ( n1512 & n2369 ) ;
  assign n2869 = n2868 ^ n1682 ^ n1118 ;
  assign n2870 = n2869 ^ n1432 ^ n655 ;
  assign n2873 = n2872 ^ n2871 ^ n2870 ;
  assign n2874 = n2873 ^ n651 ^ n224 ;
  assign n2875 = ( ~n1536 & n2867 ) | ( ~n1536 & n2874 ) | ( n2867 & n2874 ) ;
  assign n2878 = n2877 ^ n2875 ^ n1966 ;
  assign n2888 = n2887 ^ n2882 ^ n2878 ;
  assign n2855 = ( n294 & n624 ) | ( n294 & ~n1189 ) | ( n624 & ~n1189 ) ;
  assign n2854 = n2434 ^ n2274 ^ n2173 ;
  assign n2852 = n811 ^ n444 ^ n322 ;
  assign n2853 = n2852 ^ n2489 ^ n861 ;
  assign n2856 = n2855 ^ n2854 ^ n2853 ;
  assign n2857 = n2856 ^ n1914 ^ n1413 ;
  assign n2859 = ( n339 & n766 ) | ( n339 & ~n1322 ) | ( n766 & ~n1322 ) ;
  assign n2860 = ( n131 & n1513 ) | ( n131 & ~n1668 ) | ( n1513 & ~n1668 ) ;
  assign n2861 = ( n796 & ~n2859 ) | ( n796 & n2860 ) | ( ~n2859 & n2860 ) ;
  assign n2862 = n2861 ^ n2294 ^ x36 ;
  assign n2858 = n2490 ^ n2319 ^ n1013 ;
  assign n2863 = n2862 ^ n2858 ^ n1173 ;
  assign n2864 = ( ~n348 & n855 ) | ( ~n348 & n1437 ) | ( n855 & n1437 ) ;
  assign n2865 = ( n299 & n1396 ) | ( n299 & n2864 ) | ( n1396 & n2864 ) ;
  assign n2866 = ( ~n2857 & n2863 ) | ( ~n2857 & n2865 ) | ( n2863 & n2865 ) ;
  assign n2895 = n2894 ^ n2888 ^ n2866 ;
  assign n2896 = n679 ^ n195 ^ x119 ;
  assign n2897 = n970 ^ n911 ^ n437 ;
  assign n2898 = n1122 ^ x114 ^ x22 ;
  assign n2899 = n2296 ^ n1630 ^ n1118 ;
  assign n2900 = ( ~n1580 & n2898 ) | ( ~n1580 & n2899 ) | ( n2898 & n2899 ) ;
  assign n2901 = ( n252 & n2897 ) | ( n252 & n2900 ) | ( n2897 & n2900 ) ;
  assign n2904 = n809 ^ n191 ^ x118 ;
  assign n2905 = ( n146 & ~n1388 ) | ( n146 & n2904 ) | ( ~n1388 & n2904 ) ;
  assign n2906 = ( n816 & ~n1662 ) | ( n816 & n2905 ) | ( ~n1662 & n2905 ) ;
  assign n2902 = n1400 ^ n959 ^ n461 ;
  assign n2903 = ( n327 & ~n1677 ) | ( n327 & n2902 ) | ( ~n1677 & n2902 ) ;
  assign n2907 = n2906 ^ n2903 ^ n580 ;
  assign n2908 = ( ~n2896 & n2901 ) | ( ~n2896 & n2907 ) | ( n2901 & n2907 ) ;
  assign n2909 = ( ~n985 & n2217 ) | ( ~n985 & n2908 ) | ( n2217 & n2908 ) ;
  assign n2910 = n1363 ^ n725 ^ n710 ;
  assign n2911 = ( n281 & n1602 ) | ( n281 & ~n2910 ) | ( n1602 & ~n2910 ) ;
  assign n2912 = n1575 ^ n1020 ^ n709 ;
  assign n2913 = n2388 ^ n1316 ^ n272 ;
  assign n2916 = ( ~n686 & n1445 ) | ( ~n686 & n1571 ) | ( n1445 & n1571 ) ;
  assign n2914 = n2746 ^ n1145 ^ n1039 ;
  assign n2915 = ( n464 & ~n2750 ) | ( n464 & n2914 ) | ( ~n2750 & n2914 ) ;
  assign n2917 = n2916 ^ n2915 ^ n1071 ;
  assign n2918 = n1527 ^ n500 ^ n321 ;
  assign n2919 = n2918 ^ n994 ^ n964 ;
  assign n2920 = ( ~n1703 & n2917 ) | ( ~n1703 & n2919 ) | ( n2917 & n2919 ) ;
  assign n2921 = ( n458 & n2913 ) | ( n458 & n2920 ) | ( n2913 & n2920 ) ;
  assign n2922 = ( ~n2911 & n2912 ) | ( ~n2911 & n2921 ) | ( n2912 & n2921 ) ;
  assign n2923 = n959 ^ n201 ^ x50 ;
  assign n2924 = n2923 ^ n2051 ^ x69 ;
  assign n2927 = ( x71 & ~n771 ) | ( x71 & n878 ) | ( ~n771 & n878 ) ;
  assign n2928 = n2243 ^ n337 ^ x69 ;
  assign n2929 = ( n190 & ~n451 ) | ( n190 & n1467 ) | ( ~n451 & n1467 ) ;
  assign n2930 = ( n2109 & n2513 ) | ( n2109 & n2929 ) | ( n2513 & n2929 ) ;
  assign n2931 = ( x75 & ~n440 ) | ( x75 & n2930 ) | ( ~n440 & n2930 ) ;
  assign n2932 = ( n2629 & n2928 ) | ( n2629 & ~n2931 ) | ( n2928 & ~n2931 ) ;
  assign n2933 = ( ~n1719 & n2927 ) | ( ~n1719 & n2932 ) | ( n2927 & n2932 ) ;
  assign n2925 = ( ~n171 & n434 ) | ( ~n171 & n1887 ) | ( n434 & n1887 ) ;
  assign n2926 = n2925 ^ n1673 ^ n894 ;
  assign n2934 = n2933 ^ n2926 ^ n417 ;
  assign n2935 = ( n578 & n2924 ) | ( n578 & n2934 ) | ( n2924 & n2934 ) ;
  assign n2936 = n2935 ^ n1876 ^ n221 ;
  assign n2937 = ( n346 & ~n774 ) | ( n346 & n1138 ) | ( ~n774 & n1138 ) ;
  assign n2938 = n2931 ^ n967 ^ n955 ;
  assign n2939 = n2938 ^ n466 ^ n136 ;
  assign n2940 = ( n2028 & n2937 ) | ( n2028 & n2939 ) | ( n2937 & n2939 ) ;
  assign n2962 = ( n691 & ~n782 ) | ( n691 & n920 ) | ( ~n782 & n920 ) ;
  assign n2961 = n2466 ^ n1030 ^ n627 ;
  assign n2941 = n2240 ^ n2194 ^ n444 ;
  assign n2942 = n2941 ^ n198 ^ x8 ;
  assign n2943 = ( n1273 & ~n2691 ) | ( n1273 & n2942 ) | ( ~n2691 & n2942 ) ;
  assign n2958 = ( x29 & n164 ) | ( x29 & ~n167 ) | ( n164 & ~n167 ) ;
  assign n2952 = n516 ^ n377 ^ n145 ;
  assign n2953 = n2952 ^ n1602 ^ n542 ;
  assign n2954 = ( ~n849 & n1769 ) | ( ~n849 & n2953 ) | ( n1769 & n2953 ) ;
  assign n2955 = n2125 ^ n897 ^ n853 ;
  assign n2956 = n2955 ^ n1631 ^ n678 ;
  assign n2957 = ( n2794 & n2954 ) | ( n2794 & ~n2956 ) | ( n2954 & ~n2956 ) ;
  assign n2944 = ( n1253 & n1668 ) | ( n1253 & ~n2527 ) | ( n1668 & ~n2527 ) ;
  assign n2946 = n1052 ^ n481 ^ n157 ;
  assign n2947 = ( n186 & ~n474 ) | ( n186 & n755 ) | ( ~n474 & n755 ) ;
  assign n2948 = ( n822 & n2946 ) | ( n822 & ~n2947 ) | ( n2946 & ~n2947 ) ;
  assign n2945 = n1809 ^ n419 ^ n394 ;
  assign n2949 = n2948 ^ n2945 ^ n1930 ;
  assign n2950 = ( ~n1061 & n2944 ) | ( ~n1061 & n2949 ) | ( n2944 & n2949 ) ;
  assign n2951 = ( ~n599 & n1076 ) | ( ~n599 & n2950 ) | ( n1076 & n2950 ) ;
  assign n2959 = n2958 ^ n2957 ^ n2951 ;
  assign n2960 = ( ~n841 & n2943 ) | ( ~n841 & n2959 ) | ( n2943 & n2959 ) ;
  assign n2963 = n2962 ^ n2961 ^ n2960 ;
  assign n2975 = n1434 ^ n1219 ^ n686 ;
  assign n2976 = ( n912 & n2257 ) | ( n912 & ~n2975 ) | ( n2257 & ~n2975 ) ;
  assign n2977 = n2976 ^ n1370 ^ n349 ;
  assign n2978 = n2977 ^ n1645 ^ n918 ;
  assign n2972 = ( n578 & n1712 ) | ( n578 & n2398 ) | ( n1712 & n2398 ) ;
  assign n2971 = ( ~n199 & n1476 ) | ( ~n199 & n2219 ) | ( n1476 & n2219 ) ;
  assign n2973 = n2972 ^ n2971 ^ n1604 ;
  assign n2969 = ( n491 & ~n1786 ) | ( n491 & n2368 ) | ( ~n1786 & n2368 ) ;
  assign n2968 = n1234 ^ n298 ^ x82 ;
  assign n2970 = n2969 ^ n2968 ^ n1454 ;
  assign n2967 = ( n524 & ~n2045 ) | ( n524 & n2923 ) | ( ~n2045 & n2923 ) ;
  assign n2974 = n2973 ^ n2970 ^ n2967 ;
  assign n2964 = n2876 ^ n2248 ^ n1752 ;
  assign n2965 = n2964 ^ n2193 ^ n1109 ;
  assign n2966 = n2965 ^ n2732 ^ n334 ;
  assign n2979 = n2978 ^ n2974 ^ n2966 ;
  assign n2980 = ( n499 & n529 ) | ( n499 & n1564 ) | ( n529 & n1564 ) ;
  assign n2990 = n2952 ^ n2258 ^ n748 ;
  assign n2981 = ( n1937 & ~n2439 ) | ( n1937 & n2642 ) | ( ~n2439 & n2642 ) ;
  assign n2982 = ( ~n394 & n752 ) | ( ~n394 & n1973 ) | ( n752 & n1973 ) ;
  assign n2983 = ( n421 & n2981 ) | ( n421 & ~n2982 ) | ( n2981 & ~n2982 ) ;
  assign n2986 = ( n230 & ~n234 ) | ( n230 & n1682 ) | ( ~n234 & n1682 ) ;
  assign n2987 = ( n1767 & ~n2090 ) | ( n1767 & n2986 ) | ( ~n2090 & n2986 ) ;
  assign n2984 = n2545 ^ n2370 ^ n443 ;
  assign n2985 = ( n1815 & n2437 ) | ( n1815 & n2984 ) | ( n2437 & n2984 ) ;
  assign n2988 = n2987 ^ n2985 ^ n2162 ;
  assign n2989 = ( n1209 & ~n2983 ) | ( n1209 & n2988 ) | ( ~n2983 & n2988 ) ;
  assign n2991 = n2990 ^ n2989 ^ n1156 ;
  assign n2992 = ( n469 & ~n2317 ) | ( n469 & n2991 ) | ( ~n2317 & n2991 ) ;
  assign n3010 = n2750 ^ n2307 ^ n1833 ;
  assign n3011 = n3010 ^ n1147 ^ n1047 ;
  assign n2993 = ( ~n617 & n1003 ) | ( ~n617 & n1924 ) | ( n1003 & n1924 ) ;
  assign n2994 = n2986 ^ n1396 ^ n143 ;
  assign n2995 = ( ~n628 & n972 ) | ( ~n628 & n2994 ) | ( n972 & n2994 ) ;
  assign n2996 = ( n481 & n2048 ) | ( n481 & n2995 ) | ( n2048 & n2995 ) ;
  assign n2997 = n2996 ^ n1674 ^ n712 ;
  assign n2998 = n2997 ^ n2007 ^ n1396 ;
  assign n3006 = n1662 ^ n1147 ^ n928 ;
  assign n3005 = n1827 ^ n1691 ^ x110 ;
  assign n3007 = n3006 ^ n3005 ^ n1765 ;
  assign n3004 = ( ~n1045 & n1060 ) | ( ~n1045 & n1146 ) | ( n1060 & n1146 ) ;
  assign n2999 = ( x39 & x90 ) | ( x39 & n471 ) | ( x90 & n471 ) ;
  assign n3000 = n999 ^ n959 ^ n595 ;
  assign n3001 = n3000 ^ n2512 ^ n1149 ;
  assign n3002 = ( n181 & n1594 ) | ( n181 & ~n2123 ) | ( n1594 & ~n2123 ) ;
  assign n3003 = ( n2999 & n3001 ) | ( n2999 & n3002 ) | ( n3001 & n3002 ) ;
  assign n3008 = n3007 ^ n3004 ^ n3003 ;
  assign n3009 = ( n2993 & n2998 ) | ( n2993 & n3008 ) | ( n2998 & n3008 ) ;
  assign n3012 = n3011 ^ n3009 ^ n550 ;
  assign n3029 = ( x32 & ~n760 ) | ( x32 & n1860 ) | ( ~n760 & n1860 ) ;
  assign n3030 = n3029 ^ n2536 ^ n980 ;
  assign n3022 = ( n1073 & n1382 ) | ( n1073 & ~n2619 ) | ( n1382 & ~n2619 ) ;
  assign n3021 = n2574 ^ n1568 ^ n876 ;
  assign n3014 = n776 ^ n369 ^ n189 ;
  assign n3015 = ( n374 & ~n1840 ) | ( n374 & n1882 ) | ( ~n1840 & n1882 ) ;
  assign n3016 = n3015 ^ n1043 ^ n1012 ;
  assign n3017 = ( ~n679 & n1487 ) | ( ~n679 & n2898 ) | ( n1487 & n2898 ) ;
  assign n3018 = ( n383 & n3016 ) | ( n383 & ~n3017 ) | ( n3016 & ~n3017 ) ;
  assign n3019 = ( ~n333 & n3014 ) | ( ~n333 & n3018 ) | ( n3014 & n3018 ) ;
  assign n3020 = n3019 ^ n1754 ^ n1296 ;
  assign n3023 = n3022 ^ n3021 ^ n3020 ;
  assign n3024 = ( x40 & n620 ) | ( x40 & ~n1392 ) | ( n620 & ~n1392 ) ;
  assign n3025 = ( ~n388 & n1522 ) | ( ~n388 & n1810 ) | ( n1522 & n1810 ) ;
  assign n3026 = ( ~n131 & n1515 ) | ( ~n131 & n3025 ) | ( n1515 & n3025 ) ;
  assign n3027 = ( ~n2118 & n3024 ) | ( ~n2118 & n3026 ) | ( n3024 & n3026 ) ;
  assign n3028 = ( n2928 & n3023 ) | ( n2928 & ~n3027 ) | ( n3023 & ~n3027 ) ;
  assign n3031 = n3030 ^ n3028 ^ n2586 ;
  assign n3013 = ( n1583 & ~n1738 ) | ( n1583 & n3003 ) | ( ~n1738 & n3003 ) ;
  assign n3032 = n3031 ^ n3013 ^ n2154 ;
  assign n3038 = n1118 ^ n792 ^ n660 ;
  assign n3039 = ( n1561 & n2197 ) | ( n1561 & n3038 ) | ( n2197 & n3038 ) ;
  assign n3033 = ( n260 & ~n710 ) | ( n260 & n1046 ) | ( ~n710 & n1046 ) ;
  assign n3034 = n639 ^ n618 ^ n439 ;
  assign n3035 = ( n674 & n2641 ) | ( n674 & ~n3034 ) | ( n2641 & ~n3034 ) ;
  assign n3036 = n1833 ^ n752 ^ n530 ;
  assign n3037 = ( n3033 & n3035 ) | ( n3033 & n3036 ) | ( n3035 & n3036 ) ;
  assign n3040 = n3039 ^ n3037 ^ n161 ;
  assign n3061 = n3033 ^ n506 ^ x66 ;
  assign n3062 = ( n791 & n1632 ) | ( n791 & ~n3061 ) | ( n1632 & ~n3061 ) ;
  assign n3071 = ( n610 & ~n745 ) | ( n610 & n1317 ) | ( ~n745 & n1317 ) ;
  assign n3069 = n795 ^ n676 ^ x119 ;
  assign n3066 = ( n264 & n1578 ) | ( n264 & ~n1768 ) | ( n1578 & ~n1768 ) ;
  assign n3067 = n3066 ^ n2079 ^ n1094 ;
  assign n3068 = ( n2116 & n2294 ) | ( n2116 & n3067 ) | ( n2294 & n3067 ) ;
  assign n3070 = n3069 ^ n3068 ^ n1062 ;
  assign n3063 = n2313 ^ n1589 ^ n1168 ;
  assign n3064 = n3063 ^ n2299 ^ n2277 ;
  assign n3065 = ( ~n1098 & n2126 ) | ( ~n1098 & n3064 ) | ( n2126 & n3064 ) ;
  assign n3072 = n3071 ^ n3070 ^ n3065 ;
  assign n3073 = ( n623 & n3062 ) | ( n623 & ~n3072 ) | ( n3062 & ~n3072 ) ;
  assign n3074 = n3073 ^ n1528 ^ n1172 ;
  assign n3045 = ( x123 & ~n998 ) | ( x123 & n2772 ) | ( ~n998 & n2772 ) ;
  assign n3043 = ( n817 & n1093 ) | ( n817 & n1575 ) | ( n1093 & n1575 ) ;
  assign n3044 = n3043 ^ n1972 ^ n1598 ;
  assign n3041 = ( ~x27 & n967 ) | ( ~x27 & n2376 ) | ( n967 & n2376 ) ;
  assign n3042 = ( n1824 & n3018 ) | ( n1824 & n3041 ) | ( n3018 & n3041 ) ;
  assign n3046 = n3045 ^ n3044 ^ n3042 ;
  assign n3057 = n2898 ^ n1511 ^ n675 ;
  assign n3058 = ( n2317 & ~n2353 ) | ( n2317 & n3057 ) | ( ~n2353 & n3057 ) ;
  assign n3054 = ( ~n1364 & n1580 ) | ( ~n1364 & n2202 ) | ( n1580 & n2202 ) ;
  assign n3055 = n3054 ^ n2459 ^ n956 ;
  assign n3056 = ( n1674 & n2368 ) | ( n1674 & ~n3055 ) | ( n2368 & ~n3055 ) ;
  assign n3051 = n2692 ^ n1289 ^ n777 ;
  assign n3052 = n3051 ^ n2365 ^ n1769 ;
  assign n3047 = ( n454 & ~n918 ) | ( n454 & n2627 ) | ( ~n918 & n2627 ) ;
  assign n3048 = ( ~n189 & n672 ) | ( ~n189 & n3047 ) | ( n672 & n3047 ) ;
  assign n3049 = n3048 ^ n2819 ^ n2221 ;
  assign n3050 = ( n398 & n2336 ) | ( n398 & ~n3049 ) | ( n2336 & ~n3049 ) ;
  assign n3053 = n3052 ^ n3050 ^ n797 ;
  assign n3059 = n3058 ^ n3056 ^ n3053 ;
  assign n3060 = ( ~n1449 & n3046 ) | ( ~n1449 & n3059 ) | ( n3046 & n3059 ) ;
  assign n3075 = n3074 ^ n3060 ^ n796 ;
  assign n3098 = n1371 ^ n1168 ^ n475 ;
  assign n3090 = ( ~x33 & n1318 ) | ( ~x33 & n2156 ) | ( n1318 & n2156 ) ;
  assign n3094 = n2136 ^ n1505 ^ n131 ;
  assign n3092 = ( ~n162 & n783 ) | ( ~n162 & n1297 ) | ( n783 & n1297 ) ;
  assign n3091 = ( n896 & ~n1157 ) | ( n896 & n2053 ) | ( ~n1157 & n2053 ) ;
  assign n3093 = n3092 ^ n3091 ^ n1583 ;
  assign n3095 = n3094 ^ n3093 ^ n791 ;
  assign n3096 = n3095 ^ n1920 ^ x54 ;
  assign n3097 = ( ~n819 & n3090 ) | ( ~n819 & n3096 ) | ( n3090 & n3096 ) ;
  assign n3085 = n2480 ^ n2201 ^ n608 ;
  assign n3086 = n3085 ^ n2300 ^ n958 ;
  assign n3087 = n1753 ^ n1337 ^ n1286 ;
  assign n3088 = ( n267 & n3086 ) | ( n267 & ~n3087 ) | ( n3086 & ~n3087 ) ;
  assign n3079 = n2475 ^ n2015 ^ n230 ;
  assign n3080 = ( n1882 & n2273 ) | ( n1882 & ~n3079 ) | ( n2273 & ~n3079 ) ;
  assign n3081 = n3080 ^ n2790 ^ n1159 ;
  assign n3077 = ( n242 & ~n1071 ) | ( n242 & n2817 ) | ( ~n1071 & n2817 ) ;
  assign n3078 = ( x94 & ~n1235 ) | ( x94 & n3077 ) | ( ~n1235 & n3077 ) ;
  assign n3082 = n3081 ^ n3078 ^ n200 ;
  assign n3076 = ( n213 & ~n542 ) | ( n213 & n2237 ) | ( ~n542 & n2237 ) ;
  assign n3083 = n3082 ^ n3076 ^ n160 ;
  assign n3084 = n3083 ^ n2869 ^ n1749 ;
  assign n3089 = n3088 ^ n3084 ^ n1170 ;
  assign n3099 = n3098 ^ n3097 ^ n3089 ;
  assign n3100 = n1290 ^ n1154 ^ n766 ;
  assign n3101 = ( ~n170 & n1266 ) | ( ~n170 & n1679 ) | ( n1266 & n1679 ) ;
  assign n3102 = ( n259 & n466 ) | ( n259 & ~n3101 ) | ( n466 & ~n3101 ) ;
  assign n3103 = ( n1247 & n1580 ) | ( n1247 & ~n2128 ) | ( n1580 & ~n2128 ) ;
  assign n3104 = n3103 ^ n2595 ^ n2094 ;
  assign n3105 = ( ~n380 & n1173 ) | ( ~n380 & n1459 ) | ( n1173 & n1459 ) ;
  assign n3106 = n3105 ^ n2029 ^ n1425 ;
  assign n3107 = ( n712 & n1692 ) | ( n712 & n2436 ) | ( n1692 & n2436 ) ;
  assign n3108 = n3107 ^ n1986 ^ n576 ;
  assign n3109 = ( n3085 & ~n3106 ) | ( n3085 & n3108 ) | ( ~n3106 & n3108 ) ;
  assign n3113 = n1052 ^ n1027 ^ n172 ;
  assign n3112 = n1813 ^ n1688 ^ n174 ;
  assign n3110 = ( ~n1399 & n1545 ) | ( ~n1399 & n1636 ) | ( n1545 & n1636 ) ;
  assign n3111 = n3110 ^ n1257 ^ n787 ;
  assign n3114 = n3113 ^ n3112 ^ n3111 ;
  assign n3116 = ( n1101 & n1721 ) | ( n1101 & n2142 ) | ( n1721 & n2142 ) ;
  assign n3115 = ( n817 & n1089 ) | ( n817 & n1235 ) | ( n1089 & n1235 ) ;
  assign n3117 = n3116 ^ n3115 ^ n525 ;
  assign n3118 = n3117 ^ n1293 ^ n488 ;
  assign n3119 = ( ~n3109 & n3114 ) | ( ~n3109 & n3118 ) | ( n3114 & n3118 ) ;
  assign n3120 = ( ~n1275 & n3104 ) | ( ~n1275 & n3119 ) | ( n3104 & n3119 ) ;
  assign n3121 = ( n3100 & ~n3102 ) | ( n3100 & n3120 ) | ( ~n3102 & n3120 ) ;
  assign n3122 = ( n393 & n3069 ) | ( n393 & n3094 ) | ( n3069 & n3094 ) ;
  assign n3123 = n3122 ^ n2187 ^ n651 ;
  assign n3126 = ( n340 & n539 ) | ( n340 & n548 ) | ( n539 & n548 ) ;
  assign n3127 = n3126 ^ n419 ^ n380 ;
  assign n3128 = ( n940 & n1334 ) | ( n940 & n3127 ) | ( n1334 & n3127 ) ;
  assign n3129 = n3128 ^ n1245 ^ x99 ;
  assign n3137 = n1551 ^ n1104 ^ n485 ;
  assign n3138 = ( n900 & n1900 ) | ( n900 & n3137 ) | ( n1900 & n3137 ) ;
  assign n3139 = ( x76 & n1512 ) | ( x76 & ~n3138 ) | ( n1512 & ~n3138 ) ;
  assign n3140 = ( n347 & n722 ) | ( n347 & ~n3139 ) | ( n722 & ~n3139 ) ;
  assign n3141 = ( n413 & ~n1450 ) | ( n413 & n2259 ) | ( ~n1450 & n2259 ) ;
  assign n3142 = ( n3129 & n3140 ) | ( n3129 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3135 = n2197 ^ n1731 ^ n1339 ;
  assign n3136 = ( n603 & ~n1847 ) | ( n603 & n3135 ) | ( ~n1847 & n3135 ) ;
  assign n3143 = n3142 ^ n3136 ^ n2665 ;
  assign n3144 = n3143 ^ n1896 ^ n493 ;
  assign n3124 = ( n229 & n940 ) | ( n229 & ~n2986 ) | ( n940 & ~n2986 ) ;
  assign n3125 = ( ~n2356 & n2633 ) | ( ~n2356 & n3124 ) | ( n2633 & n3124 ) ;
  assign n3130 = n365 ^ n160 ^ x32 ;
  assign n3131 = ( n1074 & n3129 ) | ( n1074 & ~n3130 ) | ( n3129 & ~n3130 ) ;
  assign n3132 = ( n447 & n3125 ) | ( n447 & n3131 ) | ( n3125 & n3131 ) ;
  assign n3133 = n3132 ^ n985 ^ x16 ;
  assign n3134 = ( n1795 & n2050 ) | ( n1795 & n3133 ) | ( n2050 & n3133 ) ;
  assign n3145 = n3144 ^ n3134 ^ n2650 ;
  assign n3146 = ( n676 & n3123 ) | ( n676 & ~n3145 ) | ( n3123 & ~n3145 ) ;
  assign n3156 = ( n784 & n2269 ) | ( n784 & ~n2896 ) | ( n2269 & ~n2896 ) ;
  assign n3157 = ( ~n1154 & n1266 ) | ( ~n1154 & n3156 ) | ( n1266 & n3156 ) ;
  assign n3147 = ( x41 & ~n847 ) | ( x41 & n2306 ) | ( ~n847 & n2306 ) ;
  assign n3148 = ( n951 & n1294 ) | ( n951 & n1394 ) | ( n1294 & n1394 ) ;
  assign n3149 = ( ~n263 & n411 ) | ( ~n263 & n1502 ) | ( n411 & n1502 ) ;
  assign n3150 = n3149 ^ n2491 ^ n1847 ;
  assign n3151 = n3150 ^ n2151 ^ x46 ;
  assign n3152 = ( n1152 & n1388 ) | ( n1152 & n2262 ) | ( n1388 & n2262 ) ;
  assign n3153 = n3152 ^ n1954 ^ n1528 ;
  assign n3154 = ( ~n2079 & n3151 ) | ( ~n2079 & n3153 ) | ( n3151 & n3153 ) ;
  assign n3155 = ( n3147 & n3148 ) | ( n3147 & ~n3154 ) | ( n3148 & ~n3154 ) ;
  assign n3158 = n3157 ^ n3155 ^ n1796 ;
  assign n3167 = ( n1054 & n1136 ) | ( n1054 & n1643 ) | ( n1136 & n1643 ) ;
  assign n3168 = ( n1133 & ~n2228 ) | ( n1133 & n3167 ) | ( ~n2228 & n3167 ) ;
  assign n3169 = ( n920 & ~n1455 ) | ( n920 & n3168 ) | ( ~n1455 & n3168 ) ;
  assign n3165 = ( x0 & ~n187 ) | ( x0 & n1286 ) | ( ~n187 & n1286 ) ;
  assign n3160 = n1734 ^ n571 ^ n425 ;
  assign n3161 = n555 ^ n250 ^ n199 ;
  assign n3162 = ( n2291 & ~n3160 ) | ( n2291 & n3161 ) | ( ~n3160 & n3161 ) ;
  assign n3163 = n3162 ^ n2759 ^ n216 ;
  assign n3164 = ( n1690 & ~n2328 ) | ( n1690 & n3163 ) | ( ~n2328 & n3163 ) ;
  assign n3159 = n2691 ^ n2125 ^ n1727 ;
  assign n3166 = n3165 ^ n3164 ^ n3159 ;
  assign n3170 = n3169 ^ n3166 ^ n586 ;
  assign n3171 = ( n1573 & n1999 ) | ( n1573 & ~n3170 ) | ( n1999 & ~n3170 ) ;
  assign n3172 = n483 ^ n323 ^ n151 ;
  assign n3173 = n3172 ^ n2037 ^ n429 ;
  assign n3174 = n2952 ^ n1334 ^ n376 ;
  assign n3175 = ( n266 & n952 ) | ( n266 & ~n3174 ) | ( n952 & ~n3174 ) ;
  assign n3176 = n3175 ^ n2324 ^ n1012 ;
  assign n3178 = ( n416 & ~n1897 ) | ( n416 & n2759 ) | ( ~n1897 & n2759 ) ;
  assign n3179 = n3178 ^ n2853 ^ n2124 ;
  assign n3177 = ( ~n1346 & n2438 ) | ( ~n1346 & n2995 ) | ( n2438 & n2995 ) ;
  assign n3180 = n3179 ^ n3177 ^ n2624 ;
  assign n3193 = ( n959 & n1313 ) | ( n959 & ~n1684 ) | ( n1313 & ~n1684 ) ;
  assign n3181 = ( ~n685 & n971 ) | ( ~n685 & n1269 ) | ( n971 & n1269 ) ;
  assign n3182 = n874 ^ n803 ^ n595 ;
  assign n3183 = n3182 ^ n3010 ^ n1336 ;
  assign n3184 = ( ~x68 & n2291 ) | ( ~x68 & n3183 ) | ( n2291 & n3183 ) ;
  assign n3187 = ( x11 & n614 ) | ( x11 & ~n620 ) | ( n614 & ~n620 ) ;
  assign n3186 = n1753 ^ n282 ^ n221 ;
  assign n3185 = ( n301 & n932 ) | ( n301 & n2607 ) | ( n932 & n2607 ) ;
  assign n3188 = n3187 ^ n3186 ^ n3185 ;
  assign n3189 = ( ~n547 & n910 ) | ( ~n547 & n2408 ) | ( n910 & n2408 ) ;
  assign n3190 = n1452 ^ n414 ^ n171 ;
  assign n3191 = ( n3188 & n3189 ) | ( n3188 & ~n3190 ) | ( n3189 & ~n3190 ) ;
  assign n3192 = ( n3181 & n3184 ) | ( n3181 & ~n3191 ) | ( n3184 & ~n3191 ) ;
  assign n3194 = n3193 ^ n3192 ^ n1517 ;
  assign n3195 = ( n1096 & n3180 ) | ( n1096 & ~n3194 ) | ( n3180 & ~n3194 ) ;
  assign n3196 = ( n591 & n1597 ) | ( n591 & n1948 ) | ( n1597 & n1948 ) ;
  assign n3197 = ( n532 & n3101 ) | ( n532 & ~n3196 ) | ( n3101 & ~n3196 ) ;
  assign n3198 = n1322 ^ n226 ^ x27 ;
  assign n3199 = n2407 ^ n1057 ^ n230 ;
  assign n3200 = ( ~n1116 & n1593 ) | ( ~n1116 & n3199 ) | ( n1593 & n3199 ) ;
  assign n3201 = n3200 ^ n2732 ^ n2301 ;
  assign n3219 = n1433 ^ n954 ^ n685 ;
  assign n3220 = n3219 ^ n1591 ^ n1576 ;
  assign n3221 = n3220 ^ n1534 ^ n899 ;
  assign n3217 = n832 ^ n469 ^ x73 ;
  assign n3216 = ( n131 & n135 ) | ( n131 & ~n1350 ) | ( n135 & ~n1350 ) ;
  assign n3215 = n3014 ^ n2094 ^ n1764 ;
  assign n3218 = n3217 ^ n3216 ^ n3215 ;
  assign n3202 = n1453 ^ n221 ^ x6 ;
  assign n3203 = ( n154 & n1733 ) | ( n154 & ~n3052 ) | ( n1733 & ~n3052 ) ;
  assign n3210 = ( ~n293 & n816 ) | ( ~n293 & n1485 ) | ( n816 & n1485 ) ;
  assign n3211 = ( n2020 & n2475 ) | ( n2020 & ~n3210 ) | ( n2475 & ~n3210 ) ;
  assign n3212 = n3211 ^ n2126 ^ n1552 ;
  assign n3206 = ( x57 & ~n647 ) | ( x57 & n982 ) | ( ~n647 & n982 ) ;
  assign n3204 = n1621 ^ n381 ^ n257 ;
  assign n3205 = ( n1130 & n3033 ) | ( n1130 & n3204 ) | ( n3033 & n3204 ) ;
  assign n3207 = n3206 ^ n3205 ^ n1887 ;
  assign n3208 = ( ~n573 & n2154 ) | ( ~n573 & n3207 ) | ( n2154 & n3207 ) ;
  assign n3209 = n3208 ^ n2897 ^ x54 ;
  assign n3213 = n3212 ^ n3209 ^ n279 ;
  assign n3214 = ( n3202 & n3203 ) | ( n3202 & n3213 ) | ( n3203 & n3213 ) ;
  assign n3222 = n3221 ^ n3218 ^ n3214 ;
  assign n3223 = ( n3198 & n3201 ) | ( n3198 & n3222 ) | ( n3201 & n3222 ) ;
  assign n3224 = n3223 ^ n1612 ^ n970 ;
  assign n3247 = ( ~x90 & n472 ) | ( ~x90 & n1002 ) | ( n472 & n1002 ) ;
  assign n3248 = ( n330 & n714 ) | ( n330 & n3247 ) | ( n714 & n3247 ) ;
  assign n3249 = n3248 ^ n2367 ^ n1208 ;
  assign n3250 = ( ~x51 & n144 ) | ( ~x51 & n3249 ) | ( n144 & n3249 ) ;
  assign n3245 = n3130 ^ n820 ^ n639 ;
  assign n3237 = n983 ^ n830 ^ n459 ;
  assign n3238 = n3237 ^ n557 ^ n188 ;
  assign n3241 = ( n846 & n865 ) | ( n846 & n2252 ) | ( n865 & n2252 ) ;
  assign n3239 = ( ~x119 & n1227 ) | ( ~x119 & n2490 ) | ( n1227 & n2490 ) ;
  assign n3240 = n3239 ^ n690 ^ n367 ;
  assign n3242 = n3241 ^ n3240 ^ n674 ;
  assign n3243 = ( n2403 & n3238 ) | ( n2403 & ~n3242 ) | ( n3238 & ~n3242 ) ;
  assign n3244 = ( n650 & n2240 ) | ( n650 & ~n3243 ) | ( n2240 & ~n3243 ) ;
  assign n3246 = n3245 ^ n3244 ^ n1503 ;
  assign n3225 = ( ~x6 & n496 ) | ( ~x6 & n1251 ) | ( n496 & n1251 ) ;
  assign n3226 = n3225 ^ n374 ^ n252 ;
  assign n3227 = ( n1020 & n2060 ) | ( n1020 & n3226 ) | ( n2060 & n3226 ) ;
  assign n3233 = n3186 ^ n1846 ^ n306 ;
  assign n3234 = n3233 ^ n1713 ^ x45 ;
  assign n3231 = ( n602 & ~n961 ) | ( n602 & n1860 ) | ( ~n961 & n1860 ) ;
  assign n3230 = ( n1523 & n1665 ) | ( n1523 & n2480 ) | ( n1665 & n2480 ) ;
  assign n3228 = n2942 ^ n1022 ^ n968 ;
  assign n3229 = n3228 ^ n807 ^ x41 ;
  assign n3232 = n3231 ^ n3230 ^ n3229 ;
  assign n3235 = n3234 ^ n3232 ^ n1049 ;
  assign n3236 = ( n1897 & n3227 ) | ( n1897 & ~n3235 ) | ( n3227 & ~n3235 ) ;
  assign n3251 = n3250 ^ n3246 ^ n3236 ;
  assign n3263 = ( n287 & ~n759 ) | ( n287 & n1188 ) | ( ~n759 & n1188 ) ;
  assign n3264 = n3263 ^ n2103 ^ x72 ;
  assign n3259 = n1639 ^ n1428 ^ n1157 ;
  assign n3260 = ( n1241 & ~n1568 ) | ( n1241 & n2981 ) | ( ~n1568 & n2981 ) ;
  assign n3261 = ( x30 & ~n966 ) | ( x30 & n3260 ) | ( ~n966 & n3260 ) ;
  assign n3262 = ( ~n1927 & n3259 ) | ( ~n1927 & n3261 ) | ( n3259 & n3261 ) ;
  assign n3265 = n3264 ^ n3262 ^ n2942 ;
  assign n3256 = n2923 ^ n2352 ^ n1274 ;
  assign n3254 = n2454 ^ n2257 ^ n414 ;
  assign n3255 = n3254 ^ n2094 ^ n1431 ;
  assign n3252 = n3229 ^ n1059 ^ n586 ;
  assign n3253 = n3252 ^ n3091 ^ n1504 ;
  assign n3257 = n3256 ^ n3255 ^ n3253 ;
  assign n3258 = ( n1427 & n3203 ) | ( n1427 & ~n3257 ) | ( n3203 & ~n3257 ) ;
  assign n3266 = n3265 ^ n3258 ^ n343 ;
  assign n3267 = n2465 ^ n1642 ^ n1383 ;
  assign n3268 = n3267 ^ n2821 ^ n765 ;
  assign n3269 = ( ~n1401 & n2274 ) | ( ~n1401 & n3268 ) | ( n2274 & n3268 ) ;
  assign n3273 = n2473 ^ n1507 ^ x64 ;
  assign n3274 = ( n1413 & n2817 ) | ( n1413 & ~n3273 ) | ( n2817 & ~n3273 ) ;
  assign n3275 = ( n1635 & n3188 ) | ( n1635 & ~n3274 ) | ( n3188 & ~n3274 ) ;
  assign n3270 = n1974 ^ n1835 ^ n1395 ;
  assign n3271 = n2563 ^ n2038 ^ n1825 ;
  assign n3272 = ( n1158 & ~n3270 ) | ( n1158 & n3271 ) | ( ~n3270 & n3271 ) ;
  assign n3276 = n3275 ^ n3272 ^ n470 ;
  assign n3277 = n3276 ^ n1831 ^ n557 ;
  assign n3278 = n3277 ^ n1188 ^ n422 ;
  assign n3279 = ( n2045 & ~n3269 ) | ( n2045 & n3278 ) | ( ~n3269 & n3278 ) ;
  assign n3301 = ( ~n487 & n902 ) | ( ~n487 & n1001 ) | ( n902 & n1001 ) ;
  assign n3297 = ( n1020 & n2627 ) | ( n1020 & ~n2763 ) | ( n2627 & ~n2763 ) ;
  assign n3298 = n3297 ^ n1046 ^ n233 ;
  assign n3294 = ( n197 & n474 ) | ( n197 & ~n1357 ) | ( n474 & ~n1357 ) ;
  assign n3292 = n1670 ^ n1170 ^ n807 ;
  assign n3293 = n3292 ^ n3057 ^ n446 ;
  assign n3290 = n2806 ^ n1700 ^ n441 ;
  assign n3280 = ( n620 & n2128 ) | ( n620 & n3047 ) | ( n2128 & n3047 ) ;
  assign n3281 = n3280 ^ n1263 ^ n703 ;
  assign n3282 = ( n1401 & ~n2269 ) | ( n1401 & n2753 ) | ( ~n2269 & n2753 ) ;
  assign n3286 = ( ~n458 & n1131 ) | ( ~n458 & n1529 ) | ( n1131 & n1529 ) ;
  assign n3284 = ( n398 & ~n469 ) | ( n398 & n973 ) | ( ~n469 & n973 ) ;
  assign n3285 = ( ~n582 & n1182 ) | ( ~n582 & n3284 ) | ( n1182 & n3284 ) ;
  assign n3287 = n3286 ^ n3285 ^ n647 ;
  assign n3283 = ( n974 & n1136 ) | ( n974 & ~n2603 ) | ( n1136 & ~n2603 ) ;
  assign n3288 = n3287 ^ n3283 ^ x101 ;
  assign n3289 = ( n3281 & n3282 ) | ( n3281 & ~n3288 ) | ( n3282 & ~n3288 ) ;
  assign n3291 = n3290 ^ n3289 ^ n1383 ;
  assign n3295 = n3294 ^ n3293 ^ n3291 ;
  assign n3296 = n3295 ^ n1772 ^ n1740 ;
  assign n3299 = n3298 ^ n3296 ^ n523 ;
  assign n3300 = n3299 ^ n1805 ^ n769 ;
  assign n3302 = n3301 ^ n3300 ^ n2069 ;
  assign n3318 = n2834 ^ n880 ^ n192 ;
  assign n3319 = n3318 ^ n796 ^ n303 ;
  assign n3320 = ( ~n234 & n599 ) | ( ~n234 & n2065 ) | ( n599 & n2065 ) ;
  assign n3321 = ( n1124 & n3319 ) | ( n1124 & ~n3320 ) | ( n3319 & ~n3320 ) ;
  assign n3322 = n3321 ^ n788 ^ n355 ;
  assign n3314 = ( ~n494 & n541 ) | ( ~n494 & n655 ) | ( n541 & n655 ) ;
  assign n3315 = n3314 ^ n1011 ^ n609 ;
  assign n3316 = ( n207 & ~n766 ) | ( n207 & n1782 ) | ( ~n766 & n1782 ) ;
  assign n3317 = ( n1914 & n3315 ) | ( n1914 & ~n3316 ) | ( n3315 & ~n3316 ) ;
  assign n3310 = ( n1070 & ~n1676 ) | ( n1070 & n2430 ) | ( ~n1676 & n2430 ) ;
  assign n3306 = ( n942 & n1014 ) | ( n942 & ~n1846 ) | ( n1014 & ~n1846 ) ;
  assign n3307 = ( n266 & n1222 ) | ( n266 & n3306 ) | ( n1222 & n3306 ) ;
  assign n3308 = ( ~n1015 & n2719 ) | ( ~n1015 & n3307 ) | ( n2719 & n3307 ) ;
  assign n3303 = ( ~n321 & n595 ) | ( ~n321 & n1124 ) | ( n595 & n1124 ) ;
  assign n3304 = ( n318 & ~n667 ) | ( n318 & n3303 ) | ( ~n667 & n3303 ) ;
  assign n3305 = ( x37 & n2913 ) | ( x37 & n3304 ) | ( n2913 & n3304 ) ;
  assign n3309 = n3308 ^ n3305 ^ n275 ;
  assign n3311 = n3310 ^ n3309 ^ n3018 ;
  assign n3312 = ( n845 & ~n2010 ) | ( n845 & n3311 ) | ( ~n2010 & n3311 ) ;
  assign n3313 = ( ~n314 & n409 ) | ( ~n314 & n3312 ) | ( n409 & n3312 ) ;
  assign n3323 = n3322 ^ n3317 ^ n3313 ;
  assign n3324 = n3323 ^ n2449 ^ n339 ;
  assign n3325 = ( n1413 & n2064 ) | ( n1413 & n3324 ) | ( n2064 & n3324 ) ;
  assign n3326 = n3085 ^ n2269 ^ n2065 ;
  assign n3327 = n3326 ^ n519 ^ n491 ;
  assign n3328 = ( ~n801 & n1535 ) | ( ~n801 & n3061 ) | ( n1535 & n3061 ) ;
  assign n3329 = ( n3004 & n3327 ) | ( n3004 & n3328 ) | ( n3327 & n3328 ) ;
  assign n3330 = ( n2432 & ~n3325 ) | ( n2432 & n3329 ) | ( ~n3325 & n3329 ) ;
  assign n3331 = n1413 ^ n1224 ^ n924 ;
  assign n3332 = n3331 ^ n2449 ^ n330 ;
  assign n3333 = n925 ^ n597 ^ n158 ;
  assign n3334 = ( n563 & n830 ) | ( n563 & n3333 ) | ( n830 & n3333 ) ;
  assign n3335 = ( n1608 & n2837 ) | ( n1608 & ~n3334 ) | ( n2837 & ~n3334 ) ;
  assign n3336 = ( ~n1986 & n2050 ) | ( ~n1986 & n3335 ) | ( n2050 & n3335 ) ;
  assign n3337 = ( n3026 & n3332 ) | ( n3026 & ~n3336 ) | ( n3332 & ~n3336 ) ;
  assign n3338 = ( n135 & n262 ) | ( n135 & n2473 ) | ( n262 & n2473 ) ;
  assign n3339 = n3338 ^ n190 ^ x100 ;
  assign n3340 = n3339 ^ n3033 ^ n1090 ;
  assign n3341 = n1860 ^ n781 ^ n267 ;
  assign n3342 = n1355 ^ n1045 ^ n476 ;
  assign n3343 = ( n2009 & n3341 ) | ( n2009 & ~n3342 ) | ( n3341 & ~n3342 ) ;
  assign n3344 = n3021 ^ n1511 ^ n316 ;
  assign n3348 = ( n1015 & n1483 ) | ( n1015 & ~n2356 ) | ( n1483 & ~n2356 ) ;
  assign n3345 = n2174 ^ n398 ^ n249 ;
  assign n3346 = n3345 ^ n2075 ^ n828 ;
  assign n3347 = ( x91 & n1638 ) | ( x91 & ~n3346 ) | ( n1638 & ~n3346 ) ;
  assign n3349 = n3348 ^ n3347 ^ n1782 ;
  assign n3350 = ( n2115 & ~n3344 ) | ( n2115 & n3349 ) | ( ~n3344 & n3349 ) ;
  assign n3355 = ( ~n415 & n428 ) | ( ~n415 & n875 ) | ( n428 & n875 ) ;
  assign n3356 = n3355 ^ n2050 ^ n1647 ;
  assign n3351 = n2414 ^ n1075 ^ n672 ;
  assign n3352 = ( n330 & n1287 ) | ( n330 & ~n1586 ) | ( n1287 & ~n1586 ) ;
  assign n3353 = n1155 ^ n633 ^ x26 ;
  assign n3354 = ( n3351 & n3352 ) | ( n3351 & ~n3353 ) | ( n3352 & ~n3353 ) ;
  assign n3357 = n3356 ^ n3354 ^ n2457 ;
  assign n3358 = ( n3343 & ~n3350 ) | ( n3343 & n3357 ) | ( ~n3350 & n3357 ) ;
  assign n3379 = ( n1289 & n1357 ) | ( n1289 & ~n1643 ) | ( n1357 & ~n1643 ) ;
  assign n3380 = n1568 ^ n1261 ^ n318 ;
  assign n3381 = n3380 ^ n2938 ^ x127 ;
  assign n3382 = n3381 ^ n1842 ^ n1584 ;
  assign n3383 = ( ~x42 & n189 ) | ( ~x42 & n830 ) | ( n189 & n830 ) ;
  assign n3384 = ( x15 & n590 ) | ( x15 & n3383 ) | ( n590 & n3383 ) ;
  assign n3385 = ( n470 & ~n1111 ) | ( n470 & n3384 ) | ( ~n1111 & n3384 ) ;
  assign n3386 = ( ~n304 & n1291 ) | ( ~n304 & n3385 ) | ( n1291 & n3385 ) ;
  assign n3387 = ( n1306 & n2029 ) | ( n1306 & ~n3386 ) | ( n2029 & ~n3386 ) ;
  assign n3388 = ( n3379 & n3382 ) | ( n3379 & n3387 ) | ( n3382 & n3387 ) ;
  assign n3370 = n715 ^ n551 ^ x29 ;
  assign n3367 = n2826 ^ n1941 ^ n347 ;
  assign n3368 = ( n138 & n2583 ) | ( n138 & ~n3367 ) | ( n2583 & ~n3367 ) ;
  assign n3369 = ( ~n1355 & n1451 ) | ( ~n1355 & n3368 ) | ( n1451 & n3368 ) ;
  assign n3371 = n3370 ^ n3369 ^ n755 ;
  assign n3372 = n1620 ^ n1438 ^ n406 ;
  assign n3373 = ( n865 & ~n920 ) | ( n865 & n1184 ) | ( ~n920 & n1184 ) ;
  assign n3374 = ( x9 & n854 ) | ( x9 & ~n3373 ) | ( n854 & ~n3373 ) ;
  assign n3375 = ( n1567 & n3372 ) | ( n1567 & n3374 ) | ( n3372 & n3374 ) ;
  assign n3376 = n3375 ^ n2648 ^ n2404 ;
  assign n3377 = ( n322 & n1683 ) | ( n322 & n3376 ) | ( n1683 & n3376 ) ;
  assign n3378 = ( n2570 & n3371 ) | ( n2570 & n3377 ) | ( n3371 & n3377 ) ;
  assign n3359 = n2549 ^ n1757 ^ n1230 ;
  assign n3360 = n3359 ^ n2704 ^ n2290 ;
  assign n3361 = n3360 ^ n2918 ^ n2848 ;
  assign n3362 = ( ~n247 & n358 ) | ( ~n247 & n1794 ) | ( n358 & n1794 ) ;
  assign n3363 = ( n693 & ~n3285 ) | ( n693 & n3362 ) | ( ~n3285 & n3362 ) ;
  assign n3364 = ( n1882 & n2075 ) | ( n1882 & ~n3363 ) | ( n2075 & ~n3363 ) ;
  assign n3365 = ( ~n2089 & n2173 ) | ( ~n2089 & n3364 ) | ( n2173 & n3364 ) ;
  assign n3366 = ( n1092 & n3361 ) | ( n1092 & ~n3365 ) | ( n3361 & ~n3365 ) ;
  assign n3389 = n3388 ^ n3378 ^ n3366 ;
  assign n3390 = ( n3340 & ~n3358 ) | ( n3340 & n3389 ) | ( ~n3358 & n3389 ) ;
  assign n3401 = ( n1790 & n2182 ) | ( n1790 & ~n2256 ) | ( n2182 & ~n2256 ) ;
  assign n3391 = n3187 ^ n1075 ^ n799 ;
  assign n3392 = ( ~n651 & n934 ) | ( ~n651 & n1575 ) | ( n934 & n1575 ) ;
  assign n3393 = n1508 ^ n1443 ^ n1153 ;
  assign n3394 = ( n1050 & ~n1731 ) | ( n1050 & n3393 ) | ( ~n1731 & n3393 ) ;
  assign n3395 = ( n2111 & ~n3392 ) | ( n2111 & n3394 ) | ( ~n3392 & n3394 ) ;
  assign n3396 = n2087 ^ n280 ^ n199 ;
  assign n3397 = ( n304 & n1840 ) | ( n304 & ~n1948 ) | ( n1840 & ~n1948 ) ;
  assign n3398 = ( n1240 & ~n3396 ) | ( n1240 & n3397 ) | ( ~n3396 & n3397 ) ;
  assign n3399 = n3398 ^ n2482 ^ n1091 ;
  assign n3400 = ( n3391 & n3395 ) | ( n3391 & ~n3399 ) | ( n3395 & ~n3399 ) ;
  assign n3402 = n3401 ^ n3400 ^ n2409 ;
  assign n3403 = n2199 ^ n763 ^ x79 ;
  assign n3404 = n3403 ^ n2840 ^ n1988 ;
  assign n3405 = ( n1488 & ~n2176 ) | ( n1488 & n2676 ) | ( ~n2176 & n2676 ) ;
  assign n3406 = ( n799 & n1989 ) | ( n799 & n3373 ) | ( n1989 & n3373 ) ;
  assign n3407 = n3406 ^ n3388 ^ n3101 ;
  assign n3408 = ( n2008 & n3405 ) | ( n2008 & n3407 ) | ( n3405 & n3407 ) ;
  assign n3409 = ( ~n2235 & n3404 ) | ( ~n2235 & n3408 ) | ( n3404 & n3408 ) ;
  assign n3410 = n3409 ^ n3382 ^ n643 ;
  assign n3411 = ( n1026 & n1301 ) | ( n1026 & n3398 ) | ( n1301 & n3398 ) ;
  assign n3412 = n669 ^ n525 ^ n146 ;
  assign n3413 = n3412 ^ n1653 ^ n1037 ;
  assign n3414 = ( ~n1991 & n2468 ) | ( ~n1991 & n3413 ) | ( n2468 & n3413 ) ;
  assign n3415 = n3414 ^ n3049 ^ n800 ;
  assign n3463 = ( n1141 & n1799 ) | ( n1141 & n2114 ) | ( n1799 & n2114 ) ;
  assign n3464 = n3463 ^ n2977 ^ n1437 ;
  assign n3462 = ( n1384 & n2296 ) | ( n1384 & ~n3320 ) | ( n2296 & ~n3320 ) ;
  assign n3425 = n3061 ^ n131 ^ x103 ;
  assign n3426 = n3425 ^ n1710 ^ n647 ;
  assign n3429 = n1942 ^ n884 ^ n327 ;
  assign n3430 = ( ~x78 & n1785 ) | ( ~x78 & n3429 ) | ( n1785 & n3429 ) ;
  assign n3431 = ( x97 & ~n805 ) | ( x97 & n3430 ) | ( ~n805 & n3430 ) ;
  assign n3427 = n2519 ^ n2005 ^ n215 ;
  assign n3428 = n3427 ^ n1898 ^ n1410 ;
  assign n3432 = n3431 ^ n3428 ^ x88 ;
  assign n3416 = ( n135 & n170 ) | ( n135 & ~n3362 ) | ( n170 & ~n3362 ) ;
  assign n3417 = n3416 ^ n2154 ^ n1431 ;
  assign n3446 = ( ~n1239 & n2295 ) | ( ~n1239 & n3417 ) | ( n2295 & n3417 ) ;
  assign n3447 = n3446 ^ n3057 ^ n178 ;
  assign n3451 = ( n589 & n791 ) | ( n589 & ~n1167 ) | ( n791 & ~n1167 ) ;
  assign n3448 = ( n179 & n941 ) | ( n179 & ~n2409 ) | ( n941 & ~n2409 ) ;
  assign n3449 = ( n884 & n2398 ) | ( n884 & ~n3086 ) | ( n2398 & ~n3086 ) ;
  assign n3450 = ( n2687 & n3448 ) | ( n2687 & ~n3449 ) | ( n3448 & ~n3449 ) ;
  assign n3452 = n3451 ^ n3450 ^ n665 ;
  assign n3453 = ( n884 & n2260 ) | ( n884 & n3452 ) | ( n2260 & n3452 ) ;
  assign n3456 = n2527 ^ n1733 ^ n1018 ;
  assign n3454 = n1025 ^ n718 ^ n425 ;
  assign n3455 = ( n1018 & n1232 ) | ( n1018 & ~n3454 ) | ( n1232 & ~n3454 ) ;
  assign n3457 = n3456 ^ n3455 ^ n3035 ;
  assign n3458 = ( ~n3447 & n3453 ) | ( ~n3447 & n3457 ) | ( n3453 & n3457 ) ;
  assign n3418 = ( ~n820 & n2256 ) | ( ~n820 & n3167 ) | ( n2256 & n3167 ) ;
  assign n3419 = ( ~n2633 & n3112 ) | ( ~n2633 & n3418 ) | ( n3112 & n3418 ) ;
  assign n3420 = ( x22 & n2335 ) | ( x22 & ~n2634 ) | ( n2335 & ~n2634 ) ;
  assign n3421 = n3420 ^ n3016 ^ n1088 ;
  assign n3422 = ( n2315 & ~n2826 ) | ( n2315 & n3421 ) | ( ~n2826 & n3421 ) ;
  assign n3423 = ( n3368 & n3419 ) | ( n3368 & n3422 ) | ( n3419 & n3422 ) ;
  assign n3436 = n3045 ^ n618 ^ x49 ;
  assign n3437 = n3436 ^ n1413 ^ n1067 ;
  assign n3438 = n3437 ^ n766 ^ x61 ;
  assign n3433 = ( n1244 & ~n1801 ) | ( n1244 & n2091 ) | ( ~n1801 & n2091 ) ;
  assign n3434 = n3206 ^ n1713 ^ n1552 ;
  assign n3435 = ( x105 & n3433 ) | ( x105 & n3434 ) | ( n3433 & n3434 ) ;
  assign n3439 = n3438 ^ n3435 ^ n2279 ;
  assign n3440 = ( n891 & ~n1147 ) | ( n891 & n2046 ) | ( ~n1147 & n2046 ) ;
  assign n3441 = ( ~x7 & n443 ) | ( ~x7 & n945 ) | ( n443 & n945 ) ;
  assign n3442 = n3441 ^ n1225 ^ n754 ;
  assign n3443 = n3442 ^ n1782 ^ n297 ;
  assign n3444 = ( n880 & n3440 ) | ( n880 & n3443 ) | ( n3440 & n3443 ) ;
  assign n3445 = ( n3423 & n3439 ) | ( n3423 & ~n3444 ) | ( n3439 & ~n3444 ) ;
  assign n3459 = n3458 ^ n3445 ^ n602 ;
  assign n3460 = ( n3426 & ~n3432 ) | ( n3426 & n3459 ) | ( ~n3432 & n3459 ) ;
  assign n3424 = ( ~n993 & n3417 ) | ( ~n993 & n3423 ) | ( n3417 & n3423 ) ;
  assign n3461 = n3460 ^ n3424 ^ n1046 ;
  assign n3465 = n3464 ^ n3462 ^ n3461 ;
  assign n3466 = ( n756 & ~n1467 ) | ( n756 & n1621 ) | ( ~n1467 & n1621 ) ;
  assign n3467 = n3466 ^ n670 ^ n444 ;
  assign n3468 = ( x39 & n881 ) | ( x39 & ~n1227 ) | ( n881 & ~n1227 ) ;
  assign n3469 = n1756 ^ n1285 ^ n256 ;
  assign n3470 = n3469 ^ n3106 ^ n840 ;
  assign n3471 = ( n2324 & n3468 ) | ( n2324 & ~n3470 ) | ( n3468 & ~n3470 ) ;
  assign n3472 = n3471 ^ n1899 ^ x17 ;
  assign n3473 = ( n214 & ~n2512 ) | ( n214 & n3472 ) | ( ~n2512 & n3472 ) ;
  assign n3474 = ( n3163 & ~n3467 ) | ( n3163 & n3473 ) | ( ~n3467 & n3473 ) ;
  assign n3498 = n3237 ^ n2483 ^ n1081 ;
  assign n3495 = ( n639 & ~n947 ) | ( n639 & n1313 ) | ( ~n947 & n1313 ) ;
  assign n3493 = ( n392 & ~n2198 ) | ( n392 & n2947 ) | ( ~n2198 & n2947 ) ;
  assign n3494 = ( n473 & n1451 ) | ( n473 & ~n3493 ) | ( n1451 & ~n3493 ) ;
  assign n3496 = n3495 ^ n3494 ^ n3413 ;
  assign n3497 = ( n504 & n599 ) | ( n504 & ~n3496 ) | ( n599 & ~n3496 ) ;
  assign n3499 = n3498 ^ n3497 ^ x101 ;
  assign n3488 = ( n712 & n1785 ) | ( n712 & n2270 ) | ( n1785 & n2270 ) ;
  assign n3489 = n3488 ^ n2479 ^ n1585 ;
  assign n3490 = ( ~n176 & n1872 ) | ( ~n176 & n3489 ) | ( n1872 & n3489 ) ;
  assign n3491 = ( x0 & n1527 ) | ( x0 & ~n3490 ) | ( n1527 & ~n3490 ) ;
  assign n3492 = n3491 ^ n2948 ^ n1630 ;
  assign n3475 = ( n326 & n1225 ) | ( n326 & ~n2368 ) | ( n1225 & ~n2368 ) ;
  assign n3476 = n3475 ^ n1295 ^ n1237 ;
  assign n3477 = ( ~n536 & n859 ) | ( ~n536 & n3476 ) | ( n859 & n3476 ) ;
  assign n3478 = n1296 ^ n1287 ^ n1137 ;
  assign n3479 = ( n3454 & ~n3477 ) | ( n3454 & n3478 ) | ( ~n3477 & n3478 ) ;
  assign n3480 = ( n303 & n461 ) | ( n303 & n1577 ) | ( n461 & n1577 ) ;
  assign n3481 = n3480 ^ n641 ^ n519 ;
  assign n3482 = ( ~n2279 & n2473 ) | ( ~n2279 & n2947 ) | ( n2473 & n2947 ) ;
  assign n3483 = n3482 ^ n3125 ^ n791 ;
  assign n3484 = ( n1145 & ~n3481 ) | ( n1145 & n3483 ) | ( ~n3481 & n3483 ) ;
  assign n3485 = n3484 ^ n1734 ^ n1561 ;
  assign n3486 = n3485 ^ n2377 ^ n662 ;
  assign n3487 = ( n3088 & n3479 ) | ( n3088 & ~n3486 ) | ( n3479 & ~n3486 ) ;
  assign n3500 = n3499 ^ n3492 ^ n3487 ;
  assign n3535 = ( ~n1382 & n2176 ) | ( ~n1382 & n2717 ) | ( n2176 & n2717 ) ;
  assign n3536 = n3535 ^ n1838 ^ n960 ;
  assign n3537 = n3536 ^ n2973 ^ n1949 ;
  assign n3527 = n3463 ^ n2091 ^ n1585 ;
  assign n3525 = ( ~n143 & n1468 ) | ( ~n143 & n1948 ) | ( n1468 & n1948 ) ;
  assign n3526 = ( n971 & ~n3093 ) | ( n971 & n3525 ) | ( ~n3093 & n3525 ) ;
  assign n3528 = n3527 ^ n3526 ^ n992 ;
  assign n3529 = ( n159 & n1111 ) | ( n159 & ~n1376 ) | ( n1111 & ~n1376 ) ;
  assign n3530 = n3529 ^ n2896 ^ n228 ;
  assign n3531 = ( ~x43 & n3528 ) | ( ~x43 & n3530 ) | ( n3528 & n3530 ) ;
  assign n3522 = ( n417 & n1092 ) | ( n417 & ~n1312 ) | ( n1092 & ~n1312 ) ;
  assign n3523 = n3522 ^ n1712 ^ n1335 ;
  assign n3524 = n3523 ^ n2971 ^ n2190 ;
  assign n3519 = n2839 ^ n1199 ^ x67 ;
  assign n3520 = ( ~n1372 & n2644 ) | ( ~n1372 & n3519 ) | ( n2644 & n3519 ) ;
  assign n3516 = ( n880 & n1747 ) | ( n880 & ~n2141 ) | ( n1747 & ~n2141 ) ;
  assign n3517 = ( n1409 & n3227 ) | ( n1409 & ~n3516 ) | ( n3227 & ~n3516 ) ;
  assign n3512 = n2689 ^ n2309 ^ n338 ;
  assign n3511 = n2849 ^ n1355 ^ n1065 ;
  assign n3513 = n3512 ^ n3511 ^ n474 ;
  assign n3514 = n2213 ^ n1197 ^ n494 ;
  assign n3515 = ( n1101 & ~n3513 ) | ( n1101 & n3514 ) | ( ~n3513 & n3514 ) ;
  assign n3518 = n3517 ^ n3515 ^ n3369 ;
  assign n3501 = ( n846 & ~n1647 ) | ( n846 & n1852 ) | ( ~n1647 & n1852 ) ;
  assign n3506 = n1852 ^ n1634 ^ n698 ;
  assign n3507 = n3506 ^ n979 ^ n732 ;
  assign n3502 = n1744 ^ n1668 ^ n1336 ;
  assign n3503 = n3502 ^ n1305 ^ n980 ;
  assign n3504 = n3503 ^ n2208 ^ n156 ;
  assign n3505 = ( n1292 & ~n2130 ) | ( n1292 & n3504 ) | ( ~n2130 & n3504 ) ;
  assign n3508 = n3507 ^ n3505 ^ n2021 ;
  assign n3509 = ( n2836 & n3501 ) | ( n2836 & ~n3508 ) | ( n3501 & ~n3508 ) ;
  assign n3510 = ( n813 & n1028 ) | ( n813 & ~n3509 ) | ( n1028 & ~n3509 ) ;
  assign n3521 = n3520 ^ n3518 ^ n3510 ;
  assign n3532 = n3531 ^ n3524 ^ n3521 ;
  assign n3533 = n3532 ^ n467 ^ n455 ;
  assign n3534 = n3533 ^ n1302 ^ n466 ;
  assign n3538 = n3537 ^ n3534 ^ n198 ;
  assign n3556 = n1211 ^ n458 ^ n298 ;
  assign n3557 = ( n971 & ~n2051 ) | ( n971 & n3556 ) | ( ~n2051 & n3556 ) ;
  assign n3552 = n336 ^ n133 ^ x88 ;
  assign n3551 = ( x95 & n875 ) | ( x95 & n2254 ) | ( n875 & n2254 ) ;
  assign n3553 = n3552 ^ n3551 ^ n2650 ;
  assign n3554 = ( ~n268 & n576 ) | ( ~n268 & n3553 ) | ( n576 & n3553 ) ;
  assign n3555 = n3554 ^ n1586 ^ n1136 ;
  assign n3547 = n3185 ^ n1842 ^ n1228 ;
  assign n3548 = n3547 ^ n881 ^ n442 ;
  assign n3543 = n2397 ^ n1920 ^ n257 ;
  assign n3539 = n490 ^ n215 ^ n187 ;
  assign n3540 = ( x54 & n505 ) | ( x54 & ~n1934 ) | ( n505 & ~n1934 ) ;
  assign n3541 = ( n2211 & ~n3539 ) | ( n2211 & n3540 ) | ( ~n3539 & n3540 ) ;
  assign n3542 = ( x44 & ~n2304 ) | ( x44 & n3541 ) | ( ~n2304 & n3541 ) ;
  assign n3544 = n3543 ^ n3542 ^ n1851 ;
  assign n3545 = n3544 ^ n1527 ^ x42 ;
  assign n3546 = n3545 ^ n1421 ^ n617 ;
  assign n3549 = n3548 ^ n3546 ^ n1899 ;
  assign n3550 = ( n1651 & n2819 ) | ( n1651 & n3549 ) | ( n2819 & n3549 ) ;
  assign n3558 = n3557 ^ n3555 ^ n3550 ;
  assign n3561 = ( ~n642 & n1119 ) | ( ~n642 & n2574 ) | ( n1119 & n2574 ) ;
  assign n3560 = ( n431 & n1339 ) | ( n431 & ~n2199 ) | ( n1339 & ~n2199 ) ;
  assign n3559 = n1869 ^ n574 ^ n420 ;
  assign n3562 = n3561 ^ n3560 ^ n3559 ;
  assign n3563 = n3562 ^ n3468 ^ n925 ;
  assign n3564 = n3563 ^ n1253 ^ n534 ;
  assign n3565 = ( n367 & n575 ) | ( n367 & n2671 ) | ( n575 & n2671 ) ;
  assign n3566 = n1686 ^ n675 ^ n436 ;
  assign n3567 = ( x89 & n975 ) | ( x89 & n1364 ) | ( n975 & n1364 ) ;
  assign n3568 = n3567 ^ n2046 ^ n1221 ;
  assign n3569 = ( ~n1585 & n1965 ) | ( ~n1585 & n3568 ) | ( n1965 & n3568 ) ;
  assign n3570 = ( n362 & n1443 ) | ( n362 & n2602 ) | ( n1443 & n2602 ) ;
  assign n3571 = ( ~n1977 & n3569 ) | ( ~n1977 & n3570 ) | ( n3569 & n3570 ) ;
  assign n3572 = ( n3565 & n3566 ) | ( n3565 & n3571 ) | ( n3566 & n3571 ) ;
  assign n3573 = ( n2296 & ~n3564 ) | ( n2296 & n3572 ) | ( ~n3564 & n3572 ) ;
  assign n3575 = n2732 ^ n823 ^ n657 ;
  assign n3574 = ( n1846 & ~n2112 ) | ( n1846 & n2505 ) | ( ~n2112 & n2505 ) ;
  assign n3576 = n3575 ^ n3574 ^ n1073 ;
  assign n3577 = ( ~n2490 & n2744 ) | ( ~n2490 & n3045 ) | ( n2744 & n3045 ) ;
  assign n3578 = n3577 ^ n3003 ^ n1097 ;
  assign n3579 = ( n2363 & n3576 ) | ( n2363 & n3578 ) | ( n3576 & n3578 ) ;
  assign n3580 = ( n1748 & n3093 ) | ( n1748 & ~n3579 ) | ( n3093 & ~n3579 ) ;
  assign n3581 = n2694 ^ n351 ^ x16 ;
  assign n3582 = ( n1881 & ~n2557 ) | ( n1881 & n2619 ) | ( ~n2557 & n2619 ) ;
  assign n3583 = ( n1926 & n3581 ) | ( n1926 & ~n3582 ) | ( n3581 & ~n3582 ) ;
  assign n3584 = ( n1137 & ~n1138 ) | ( n1137 & n1496 ) | ( ~n1138 & n1496 ) ;
  assign n3585 = n3438 ^ n2785 ^ n2497 ;
  assign n3586 = ( ~n1835 & n3584 ) | ( ~n1835 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3587 = n1174 ^ n1032 ^ n889 ;
  assign n3594 = ( ~n445 & n749 ) | ( ~n445 & n2403 ) | ( n749 & n2403 ) ;
  assign n3591 = ( n401 & n1284 ) | ( n401 & ~n1689 ) | ( n1284 & ~n1689 ) ;
  assign n3588 = ( ~n2218 & n2719 ) | ( ~n2218 & n2733 ) | ( n2719 & n2733 ) ;
  assign n3589 = ( n378 & ~n1231 ) | ( n378 & n3588 ) | ( ~n1231 & n3588 ) ;
  assign n3590 = n3589 ^ n2803 ^ n1026 ;
  assign n3592 = n3591 ^ n3590 ^ n714 ;
  assign n3593 = n3592 ^ n1773 ^ x65 ;
  assign n3595 = n3594 ^ n3593 ^ n1403 ;
  assign n3596 = ( n3011 & n3587 ) | ( n3011 & ~n3595 ) | ( n3587 & ~n3595 ) ;
  assign n3597 = ( x31 & n784 ) | ( x31 & n3551 ) | ( n784 & n3551 ) ;
  assign n3598 = n3597 ^ n2791 ^ n1539 ;
  assign n3599 = ( ~n3586 & n3596 ) | ( ~n3586 & n3598 ) | ( n3596 & n3598 ) ;
  assign n3602 = n609 ^ n476 ^ n456 ;
  assign n3600 = ( n476 & n2699 ) | ( n476 & n2831 ) | ( n2699 & n2831 ) ;
  assign n3601 = n3600 ^ n1077 ^ n1024 ;
  assign n3603 = n3602 ^ n3601 ^ n1300 ;
  assign n3604 = n3603 ^ n604 ^ n566 ;
  assign n3613 = n3433 ^ n3216 ^ n1501 ;
  assign n3614 = n3613 ^ n2358 ^ n300 ;
  assign n3605 = n3162 ^ n768 ^ n719 ;
  assign n3606 = n3605 ^ n3292 ^ n1979 ;
  assign n3610 = n3240 ^ n2314 ^ n272 ;
  assign n3608 = ( n671 & n1181 ) | ( n671 & n2061 ) | ( n1181 & n2061 ) ;
  assign n3607 = ( ~x79 & n366 ) | ( ~x79 & n2060 ) | ( n366 & n2060 ) ;
  assign n3609 = n3608 ^ n3607 ^ n1923 ;
  assign n3611 = n3610 ^ n3609 ^ n1771 ;
  assign n3612 = ( ~n3058 & n3606 ) | ( ~n3058 & n3611 ) | ( n3606 & n3611 ) ;
  assign n3615 = n3614 ^ n3612 ^ n1876 ;
  assign n3616 = n3338 ^ n3221 ^ n1401 ;
  assign n3617 = ( n388 & ~n2364 ) | ( n388 & n3616 ) | ( ~n2364 & n3616 ) ;
  assign n3618 = ( ~n236 & n1321 ) | ( ~n236 & n3617 ) | ( n1321 & n3617 ) ;
  assign n3619 = ( n224 & n387 ) | ( n224 & n808 ) | ( n387 & n808 ) ;
  assign n3620 = ( ~n886 & n3514 ) | ( ~n886 & n3619 ) | ( n3514 & n3619 ) ;
  assign n3621 = ( ~x2 & n2656 ) | ( ~x2 & n3620 ) | ( n2656 & n3620 ) ;
  assign n3622 = n3621 ^ n1966 ^ n1808 ;
  assign n3623 = ( n1641 & ~n3618 ) | ( n1641 & n3622 ) | ( ~n3618 & n3622 ) ;
  assign n3626 = ( n736 & n756 ) | ( n736 & ~n1155 ) | ( n756 & ~n1155 ) ;
  assign n3627 = n3626 ^ n1066 ^ n158 ;
  assign n3624 = ( n1145 & n3014 ) | ( n1145 & ~n3281 ) | ( n3014 & ~n3281 ) ;
  assign n3625 = n3624 ^ n2656 ^ n473 ;
  assign n3628 = n3627 ^ n3625 ^ n2415 ;
  assign n3644 = n2697 ^ n1052 ^ n721 ;
  assign n3643 = n2634 ^ n1706 ^ n1436 ;
  assign n3631 = n2911 ^ n917 ^ n348 ;
  assign n3629 = n1578 ^ n372 ^ n285 ;
  assign n3630 = n3629 ^ n985 ^ n200 ;
  assign n3632 = n3631 ^ n3630 ^ n2899 ;
  assign n3633 = ( ~n2173 & n3488 ) | ( ~n2173 & n3632 ) | ( n3488 & n3632 ) ;
  assign n3634 = ( n311 & ~n1755 ) | ( n311 & n2308 ) | ( ~n1755 & n2308 ) ;
  assign n3639 = n2403 ^ n1409 ^ n434 ;
  assign n3635 = ( n600 & n2547 ) | ( n600 & n2812 ) | ( n2547 & n2812 ) ;
  assign n3636 = ( n1526 & ~n1677 ) | ( n1526 & n3635 ) | ( ~n1677 & n3635 ) ;
  assign n3637 = n3636 ^ n925 ^ n842 ;
  assign n3638 = n3637 ^ n475 ^ x31 ;
  assign n3640 = n3639 ^ n3638 ^ n1840 ;
  assign n3641 = ( n1511 & n3634 ) | ( n1511 & n3640 ) | ( n3634 & n3640 ) ;
  assign n3642 = ( n3506 & n3633 ) | ( n3506 & ~n3641 ) | ( n3633 & ~n3641 ) ;
  assign n3645 = n3644 ^ n3643 ^ n3642 ;
  assign n3646 = ( ~n2634 & n3628 ) | ( ~n2634 & n3645 ) | ( n3628 & n3645 ) ;
  assign n3647 = ( ~n627 & n736 ) | ( ~n627 & n1595 ) | ( n736 & n1595 ) ;
  assign n3648 = n3647 ^ n1167 ^ x43 ;
  assign n3649 = ( n1040 & n3122 ) | ( n1040 & n3648 ) | ( n3122 & n3648 ) ;
  assign n3650 = ( n411 & n554 ) | ( n411 & ~n1226 ) | ( n554 & ~n1226 ) ;
  assign n3652 = ( x98 & n196 ) | ( x98 & ~n875 ) | ( n196 & ~n875 ) ;
  assign n3651 = ( x2 & ~n708 ) | ( x2 & n2459 ) | ( ~n708 & n2459 ) ;
  assign n3653 = n3652 ^ n3651 ^ n2497 ;
  assign n3654 = ( n677 & n1032 ) | ( n677 & n1436 ) | ( n1032 & n1436 ) ;
  assign n3655 = ( ~n645 & n1571 ) | ( ~n645 & n1971 ) | ( n1571 & n1971 ) ;
  assign n3656 = n3655 ^ n2212 ^ n1384 ;
  assign n3657 = ( ~n381 & n2327 ) | ( ~n381 & n3656 ) | ( n2327 & n3656 ) ;
  assign n3658 = ( n1172 & n3654 ) | ( n1172 & n3657 ) | ( n3654 & n3657 ) ;
  assign n3659 = n3658 ^ n3138 ^ n670 ;
  assign n3660 = ( n3650 & n3653 ) | ( n3650 & n3659 ) | ( n3653 & n3659 ) ;
  assign n3661 = n3660 ^ n3341 ^ n2436 ;
  assign n3662 = ( n1654 & n3649 ) | ( n1654 & n3661 ) | ( n3649 & n3661 ) ;
  assign n3663 = ( n1322 & n1781 ) | ( n1322 & ~n3066 ) | ( n1781 & ~n3066 ) ;
  assign n3665 = ( ~n622 & n1006 ) | ( ~n622 & n1903 ) | ( n1006 & n1903 ) ;
  assign n3664 = n3063 ^ n1543 ^ n1441 ;
  assign n3666 = n3665 ^ n3664 ^ n878 ;
  assign n3667 = n2183 ^ n863 ^ n185 ;
  assign n3668 = ( n404 & ~n799 ) | ( n404 & n1609 ) | ( ~n799 & n1609 ) ;
  assign n3669 = ( ~n526 & n710 ) | ( ~n526 & n712 ) | ( n710 & n712 ) ;
  assign n3670 = ( n912 & n1312 ) | ( n912 & ~n3669 ) | ( n1312 & ~n3669 ) ;
  assign n3671 = ( n332 & n708 ) | ( n332 & n1565 ) | ( n708 & n1565 ) ;
  assign n3672 = ( n3668 & n3670 ) | ( n3668 & ~n3671 ) | ( n3670 & ~n3671 ) ;
  assign n3673 = ( n2787 & ~n3667 ) | ( n2787 & n3672 ) | ( ~n3667 & n3672 ) ;
  assign n3674 = ( ~n312 & n1056 ) | ( ~n312 & n1384 ) | ( n1056 & n1384 ) ;
  assign n3675 = n3674 ^ n1307 ^ n844 ;
  assign n3676 = n3285 ^ n2184 ^ n467 ;
  assign n3677 = ( n2067 & ~n3675 ) | ( n2067 & n3676 ) | ( ~n3675 & n3676 ) ;
  assign n3678 = ( ~n980 & n1243 ) | ( ~n980 & n2376 ) | ( n1243 & n2376 ) ;
  assign n3679 = ( n3673 & n3677 ) | ( n3673 & ~n3678 ) | ( n3677 & ~n3678 ) ;
  assign n3680 = ( n3663 & ~n3666 ) | ( n3663 & n3679 ) | ( ~n3666 & n3679 ) ;
  assign n3681 = ( n787 & n3064 ) | ( n787 & n3220 ) | ( n3064 & n3220 ) ;
  assign n3682 = n1615 ^ n1426 ^ n623 ;
  assign n3683 = ( ~n1292 & n1590 ) | ( ~n1292 & n3682 ) | ( n1590 & n3682 ) ;
  assign n3684 = ( ~n813 & n3681 ) | ( ~n813 & n3683 ) | ( n3681 & n3683 ) ;
  assign n3685 = n3684 ^ n768 ^ n204 ;
  assign n3687 = n2060 ^ n795 ^ n621 ;
  assign n3686 = n887 ^ n762 ^ n696 ;
  assign n3688 = n3687 ^ n3686 ^ n2210 ;
  assign n3689 = ( ~n986 & n1023 ) | ( ~n986 & n1589 ) | ( n1023 & n1589 ) ;
  assign n3690 = n3689 ^ n1490 ^ n1072 ;
  assign n3691 = ( ~n669 & n802 ) | ( ~n669 & n3690 ) | ( n802 & n3690 ) ;
  assign n3692 = ( ~n589 & n3688 ) | ( ~n589 & n3691 ) | ( n3688 & n3691 ) ;
  assign n3693 = ( x7 & n1061 ) | ( x7 & n1471 ) | ( n1061 & n1471 ) ;
  assign n3694 = n3693 ^ n1677 ^ n852 ;
  assign n3695 = ( ~n1205 & n3561 ) | ( ~n1205 & n3694 ) | ( n3561 & n3694 ) ;
  assign n3696 = ( ~n1842 & n2435 ) | ( ~n1842 & n3695 ) | ( n2435 & n3695 ) ;
  assign n3697 = n2355 ^ n1730 ^ n994 ;
  assign n3698 = ( n1441 & n3217 ) | ( n1441 & n3697 ) | ( n3217 & n3697 ) ;
  assign n3699 = n3698 ^ n2437 ^ n1142 ;
  assign n3700 = ( n859 & n2438 ) | ( n859 & n2805 ) | ( n2438 & n2805 ) ;
  assign n3701 = ( ~n533 & n642 ) | ( ~n533 & n1105 ) | ( n642 & n1105 ) ;
  assign n3702 = n3326 ^ n882 ^ n344 ;
  assign n3703 = ( n1643 & n2368 ) | ( n1643 & ~n3629 ) | ( n2368 & ~n3629 ) ;
  assign n3704 = ( n3701 & n3702 ) | ( n3701 & ~n3703 ) | ( n3702 & ~n3703 ) ;
  assign n3705 = n3704 ^ n3632 ^ n1750 ;
  assign n3706 = ( n2654 & n3700 ) | ( n2654 & ~n3705 ) | ( n3700 & ~n3705 ) ;
  assign n3707 = ( n1991 & n3699 ) | ( n1991 & ~n3706 ) | ( n3699 & ~n3706 ) ;
  assign n3708 = ( ~n1510 & n2667 ) | ( ~n1510 & n3707 ) | ( n2667 & n3707 ) ;
  assign n3709 = ( ~n3692 & n3696 ) | ( ~n3692 & n3708 ) | ( n3696 & n3708 ) ;
  assign n3722 = ( x53 & n783 ) | ( x53 & ~n2257 ) | ( n783 & ~n2257 ) ;
  assign n3723 = ( ~n192 & n1256 ) | ( ~n192 & n3169 ) | ( n1256 & n3169 ) ;
  assign n3724 = ( n844 & n3722 ) | ( n844 & ~n3723 ) | ( n3722 & ~n3723 ) ;
  assign n3719 = n720 ^ n522 ^ n301 ;
  assign n3720 = n3719 ^ n3427 ^ n1015 ;
  assign n3721 = n3720 ^ n3522 ^ n522 ;
  assign n3725 = n3724 ^ n3721 ^ n175 ;
  assign n3726 = n3725 ^ n2727 ^ n2488 ;
  assign n3711 = ( ~n435 & n831 ) | ( ~n435 & n2633 ) | ( n831 & n2633 ) ;
  assign n3710 = n3239 ^ n1549 ^ n348 ;
  assign n3712 = n3711 ^ n3710 ^ n923 ;
  assign n3715 = n1570 ^ n1234 ^ n402 ;
  assign n3713 = ( n1218 & ~n1592 ) | ( n1218 & n3165 ) | ( ~n1592 & n3165 ) ;
  assign n3714 = n3713 ^ n1452 ^ n829 ;
  assign n3716 = n3715 ^ n3714 ^ n1959 ;
  assign n3717 = ( ~n2517 & n3712 ) | ( ~n2517 & n3716 ) | ( n3712 & n3716 ) ;
  assign n3718 = n3717 ^ n1878 ^ n1083 ;
  assign n3727 = n3726 ^ n3718 ^ n2953 ;
  assign n3749 = n3531 ^ n2757 ^ n2561 ;
  assign n3750 = n3749 ^ n2336 ^ n1322 ;
  assign n3728 = ( n347 & n708 ) | ( n347 & ~n1079 ) | ( n708 & ~n1079 ) ;
  assign n3729 = n3728 ^ n1239 ^ x25 ;
  assign n3730 = ( ~n154 & n640 ) | ( ~n154 & n932 ) | ( n640 & n932 ) ;
  assign n3731 = ( n1112 & ~n2071 ) | ( n1112 & n2942 ) | ( ~n2071 & n2942 ) ;
  assign n3732 = ( ~n3729 & n3730 ) | ( ~n3729 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3733 = ( ~n140 & n700 ) | ( ~n140 & n1271 ) | ( n700 & n1271 ) ;
  assign n3734 = ( n234 & n655 ) | ( n234 & n1891 ) | ( n655 & n1891 ) ;
  assign n3735 = n3734 ^ n3331 ^ n1164 ;
  assign n3736 = n1451 ^ n1332 ^ n1205 ;
  assign n3737 = n3736 ^ n993 ^ x51 ;
  assign n3738 = ( x33 & n1015 ) | ( x33 & n1219 ) | ( n1015 & n1219 ) ;
  assign n3739 = ( n1884 & n2503 ) | ( n1884 & ~n3738 ) | ( n2503 & ~n3738 ) ;
  assign n3740 = ( n2168 & ~n3737 ) | ( n2168 & n3739 ) | ( ~n3737 & n3739 ) ;
  assign n3741 = n1215 ^ n832 ^ n288 ;
  assign n3742 = ( n443 & n3105 ) | ( n443 & n3741 ) | ( n3105 & n3741 ) ;
  assign n3743 = ( n478 & n1107 ) | ( n478 & n3742 ) | ( n1107 & n3742 ) ;
  assign n3744 = n3743 ^ n3428 ^ n805 ;
  assign n3745 = ( n1628 & n3740 ) | ( n1628 & n3744 ) | ( n3740 & n3744 ) ;
  assign n3746 = ( n3733 & n3735 ) | ( n3733 & n3745 ) | ( n3735 & n3745 ) ;
  assign n3747 = n3746 ^ n2660 ^ n1663 ;
  assign n3748 = ( ~n3105 & n3732 ) | ( ~n3105 & n3747 ) | ( n3732 & n3747 ) ;
  assign n3751 = n3750 ^ n3748 ^ n3191 ;
  assign n3757 = n1691 ^ n209 ^ n137 ;
  assign n3758 = n3757 ^ n2961 ^ n2759 ;
  assign n3752 = ( n656 & n1147 ) | ( n656 & ~n1295 ) | ( n1147 & ~n1295 ) ;
  assign n3753 = n3752 ^ n980 ^ n315 ;
  assign n3754 = n3753 ^ n1661 ^ n1456 ;
  assign n3755 = n3754 ^ n2870 ^ n2620 ;
  assign n3756 = n3755 ^ n3280 ^ n1640 ;
  assign n3759 = n3758 ^ n3756 ^ n1924 ;
  assign n3767 = n2628 ^ n2076 ^ n438 ;
  assign n3766 = ( n717 & ~n1529 ) | ( n717 & n2264 ) | ( ~n1529 & n2264 ) ;
  assign n3765 = n2785 ^ n2600 ^ n2220 ;
  assign n3768 = n3767 ^ n3766 ^ n3765 ;
  assign n3763 = ( n440 & ~n971 ) | ( n440 & n988 ) | ( ~n971 & n988 ) ;
  assign n3761 = ( n336 & n982 ) | ( n336 & ~n1667 ) | ( n982 & ~n1667 ) ;
  assign n3760 = n3440 ^ n1632 ^ n265 ;
  assign n3762 = n3761 ^ n3760 ^ n247 ;
  assign n3764 = n3763 ^ n3762 ^ x47 ;
  assign n3769 = n3768 ^ n3764 ^ n2635 ;
  assign n3814 = ( ~n636 & n1219 ) | ( ~n636 & n1568 ) | ( n1219 & n1568 ) ;
  assign n3810 = n855 ^ n724 ^ x41 ;
  assign n3811 = ( n609 & ~n1321 ) | ( n609 & n3810 ) | ( ~n1321 & n3810 ) ;
  assign n3812 = ( x75 & n2105 ) | ( x75 & n3811 ) | ( n2105 & n3811 ) ;
  assign n3806 = n1209 ^ n471 ^ n179 ;
  assign n3807 = ( ~n211 & n3733 ) | ( ~n211 & n3806 ) | ( n3733 & n3806 ) ;
  assign n3808 = ( ~n2160 & n3315 ) | ( ~n2160 & n3807 ) | ( n3315 & n3807 ) ;
  assign n3809 = ( x34 & ~n2220 ) | ( x34 & n3808 ) | ( ~n2220 & n3808 ) ;
  assign n3813 = n3812 ^ n3809 ^ n1044 ;
  assign n3796 = n3449 ^ n1691 ^ n173 ;
  assign n3797 = n3796 ^ n3347 ^ n1708 ;
  assign n3801 = ( ~n1290 & n1717 ) | ( ~n1290 & n3131 ) | ( n1717 & n3131 ) ;
  assign n3798 = n2068 ^ n1414 ^ n1303 ;
  assign n3799 = n1433 ^ n532 ^ x63 ;
  assign n3800 = ( n1131 & n3798 ) | ( n1131 & ~n3799 ) | ( n3798 & ~n3799 ) ;
  assign n3802 = n3801 ^ n3800 ^ n934 ;
  assign n3803 = ( ~n1919 & n3797 ) | ( ~n1919 & n3802 ) | ( n3797 & n3802 ) ;
  assign n3804 = ( n298 & ~n2665 ) | ( n298 & n3803 ) | ( ~n2665 & n3803 ) ;
  assign n3784 = ( n2876 & ~n3428 ) | ( n2876 & n3496 ) | ( ~n3428 & n3496 ) ;
  assign n3785 = ( ~n191 & n520 ) | ( ~n191 & n694 ) | ( n520 & n694 ) ;
  assign n3786 = n3785 ^ n1389 ^ x58 ;
  assign n3787 = n3488 ^ n780 ^ x38 ;
  assign n3788 = ( n1732 & n3786 ) | ( n1732 & ~n3787 ) | ( n3786 & ~n3787 ) ;
  assign n3789 = n2409 ^ n1059 ^ x97 ;
  assign n3790 = ( n2066 & ~n3024 ) | ( n2066 & n3789 ) | ( ~n3024 & n3789 ) ;
  assign n3791 = ( n565 & n1218 ) | ( n565 & n1707 ) | ( n1218 & n1707 ) ;
  assign n3792 = n3791 ^ n3480 ^ n2931 ;
  assign n3793 = ( ~n564 & n3451 ) | ( ~n564 & n3792 ) | ( n3451 & n3792 ) ;
  assign n3794 = ( ~n1626 & n3790 ) | ( ~n1626 & n3793 ) | ( n3790 & n3793 ) ;
  assign n3795 = ( n3784 & n3788 ) | ( n3784 & n3794 ) | ( n3788 & n3794 ) ;
  assign n3781 = n3341 ^ n1039 ^ n973 ;
  assign n3782 = ( x114 & n2610 ) | ( x114 & ~n3781 ) | ( n2610 & ~n3781 ) ;
  assign n3779 = n2233 ^ n1809 ^ n499 ;
  assign n3777 = n3220 ^ n2036 ^ n463 ;
  assign n3778 = n3777 ^ n2237 ^ n339 ;
  assign n3780 = n3779 ^ n3778 ^ n3199 ;
  assign n3772 = n2182 ^ n955 ^ n548 ;
  assign n3773 = n3772 ^ n1081 ^ n1022 ;
  assign n3774 = ( x23 & n1464 ) | ( x23 & ~n2376 ) | ( n1464 & ~n2376 ) ;
  assign n3775 = ( n3359 & ~n3773 ) | ( n3359 & n3774 ) | ( ~n3773 & n3774 ) ;
  assign n3770 = ( ~n1164 & n1529 ) | ( ~n1164 & n2390 ) | ( n1529 & n2390 ) ;
  assign n3771 = n3770 ^ n2617 ^ n1994 ;
  assign n3776 = n3775 ^ n3771 ^ n818 ;
  assign n3783 = n3782 ^ n3780 ^ n3776 ;
  assign n3805 = n3804 ^ n3795 ^ n3783 ;
  assign n3815 = n3814 ^ n3813 ^ n3805 ;
  assign n3822 = n1563 ^ n430 ^ n257 ;
  assign n3821 = n3801 ^ n1373 ^ n453 ;
  assign n3818 = ( x54 & n482 ) | ( x54 & ~n495 ) | ( n482 & ~n495 ) ;
  assign n3819 = n3818 ^ n2730 ^ n1642 ;
  assign n3816 = n2994 ^ n2586 ^ n1920 ;
  assign n3817 = n3816 ^ n2221 ^ n1607 ;
  assign n3820 = n3819 ^ n3817 ^ n1923 ;
  assign n3823 = n3822 ^ n3821 ^ n3820 ;
  assign n3859 = ( ~x34 & n503 ) | ( ~x34 & n1413 ) | ( n503 & n1413 ) ;
  assign n3860 = ( n278 & ~n1719 ) | ( n278 & n3859 ) | ( ~n1719 & n3859 ) ;
  assign n3861 = n3860 ^ n3331 ^ n327 ;
  assign n3862 = n3861 ^ n2125 ^ n675 ;
  assign n3863 = ( n2000 & ~n3561 ) | ( n2000 & n3862 ) | ( ~n3561 & n3862 ) ;
  assign n3866 = ( ~x1 & n285 ) | ( ~x1 & n1226 ) | ( n285 & n1226 ) ;
  assign n3865 = ( n179 & ~n920 ) | ( n179 & n1229 ) | ( ~n920 & n1229 ) ;
  assign n3867 = n3866 ^ n3865 ^ n2466 ;
  assign n3852 = ( x115 & n1873 ) | ( x115 & n2404 ) | ( n1873 & n2404 ) ;
  assign n3853 = ( x38 & n2102 ) | ( x38 & ~n3852 ) | ( n2102 & ~n3852 ) ;
  assign n3864 = ( n417 & n3342 ) | ( n417 & n3853 ) | ( n3342 & n3853 ) ;
  assign n3868 = n3867 ^ n3864 ^ n2804 ;
  assign n3869 = ( n274 & n312 ) | ( n274 & n1570 ) | ( n312 & n1570 ) ;
  assign n3870 = n3869 ^ n3450 ^ n820 ;
  assign n3871 = ( ~n3863 & n3868 ) | ( ~n3863 & n3870 ) | ( n3868 & n3870 ) ;
  assign n3855 = n3754 ^ n3686 ^ n1898 ;
  assign n3856 = n3855 ^ n1317 ^ n362 ;
  assign n3854 = n3853 ^ n1155 ^ n1121 ;
  assign n3857 = n3856 ^ n3854 ^ n1331 ;
  assign n3849 = n2210 ^ n2208 ^ n953 ;
  assign n3841 = ( n1587 & n1708 ) | ( n1587 & ~n2184 ) | ( n1708 & ~n2184 ) ;
  assign n3842 = ( n3245 & n3723 ) | ( n3245 & n3841 ) | ( n3723 & n3841 ) ;
  assign n3843 = n2417 ^ n1498 ^ n1410 ;
  assign n3844 = ( n1290 & ~n1959 ) | ( n1290 & n3284 ) | ( ~n1959 & n3284 ) ;
  assign n3845 = n3844 ^ n3321 ^ n337 ;
  assign n3846 = ( n1586 & ~n3843 ) | ( n1586 & n3845 ) | ( ~n3843 & n3845 ) ;
  assign n3847 = ( n3739 & n3789 ) | ( n3739 & ~n3846 ) | ( n3789 & ~n3846 ) ;
  assign n3848 = ( n2733 & n3842 ) | ( n2733 & ~n3847 ) | ( n3842 & ~n3847 ) ;
  assign n3835 = n1945 ^ n1197 ^ n277 ;
  assign n3832 = ( ~n268 & n1459 ) | ( ~n268 & n3034 ) | ( n1459 & n3034 ) ;
  assign n3833 = ( n991 & n1050 ) | ( n991 & n3832 ) | ( n1050 & n3832 ) ;
  assign n3831 = n2274 ^ n724 ^ n201 ;
  assign n3834 = n3833 ^ n3831 ^ n2029 ;
  assign n3836 = n3835 ^ n3834 ^ n1137 ;
  assign n3837 = ( ~n1457 & n2341 ) | ( ~n1457 & n3129 ) | ( n2341 & n3129 ) ;
  assign n3838 = ( x76 & n2685 ) | ( x76 & n3837 ) | ( n2685 & n3837 ) ;
  assign n3839 = n3838 ^ n2765 ^ n799 ;
  assign n3840 = ( n2123 & n3836 ) | ( n2123 & ~n3839 ) | ( n3836 & ~n3839 ) ;
  assign n3850 = n3849 ^ n3848 ^ n3840 ;
  assign n3829 = n3537 ^ n1872 ^ n873 ;
  assign n3824 = n1545 ^ n1290 ^ n175 ;
  assign n3825 = ( x60 & n440 ) | ( x60 & ~n2656 ) | ( n440 & ~n2656 ) ;
  assign n3826 = ( n277 & n375 ) | ( n277 & ~n3825 ) | ( n375 & ~n3825 ) ;
  assign n3827 = ( ~x102 & n3824 ) | ( ~x102 & n3826 ) | ( n3824 & n3826 ) ;
  assign n3828 = n3827 ^ n1535 ^ n967 ;
  assign n3830 = n3829 ^ n3828 ^ n2810 ;
  assign n3851 = n3850 ^ n3830 ^ n3009 ;
  assign n3858 = n3857 ^ n3851 ^ n933 ;
  assign n3872 = n3871 ^ n3858 ^ n3448 ;
  assign n3896 = ( ~n814 & n885 ) | ( ~n814 & n1931 ) | ( n885 & n1931 ) ;
  assign n3897 = ( n1231 & n2552 ) | ( n1231 & ~n3896 ) | ( n2552 & ~n3896 ) ;
  assign n3892 = ( ~n1498 & n3436 ) | ( ~n1498 & n3442 ) | ( n3436 & n3442 ) ;
  assign n3891 = n3667 ^ n1871 ^ n872 ;
  assign n3889 = ( x23 & ~n149 ) | ( x23 & n3220 ) | ( ~n149 & n3220 ) ;
  assign n3888 = n2188 ^ n1358 ^ n1203 ;
  assign n3886 = n729 ^ n722 ^ n318 ;
  assign n3887 = n3886 ^ n958 ^ n356 ;
  assign n3890 = n3889 ^ n3888 ^ n3887 ;
  assign n3893 = n3892 ^ n3891 ^ n3890 ;
  assign n3894 = ( n2469 & ~n3186 ) | ( n2469 & n3893 ) | ( ~n3186 & n3893 ) ;
  assign n3895 = n3894 ^ n3182 ^ n2734 ;
  assign n3898 = n3897 ^ n3895 ^ n1977 ;
  assign n3873 = ( n2911 & n2970 ) | ( n2911 & n3345 ) | ( n2970 & n3345 ) ;
  assign n3874 = ( n1043 & n2069 ) | ( n1043 & n3362 ) | ( n2069 & n3362 ) ;
  assign n3875 = n2127 ^ n1267 ^ n380 ;
  assign n3876 = ( n2252 & n3874 ) | ( n2252 & ~n3875 ) | ( n3874 & ~n3875 ) ;
  assign n3877 = n1642 ^ n841 ^ n281 ;
  assign n3878 = ( x23 & n490 ) | ( x23 & ~n3877 ) | ( n490 & ~n3877 ) ;
  assign n3879 = ( n283 & ~n2284 ) | ( n283 & n3878 ) | ( ~n2284 & n3878 ) ;
  assign n3880 = ( ~n402 & n2198 ) | ( ~n402 & n3879 ) | ( n2198 & n3879 ) ;
  assign n3881 = n3880 ^ n1577 ^ n515 ;
  assign n3882 = n3881 ^ n3842 ^ n702 ;
  assign n3883 = ( n2838 & n3581 ) | ( n2838 & ~n3882 ) | ( n3581 & ~n3882 ) ;
  assign n3884 = ( n2924 & n3876 ) | ( n2924 & n3883 ) | ( n3876 & n3883 ) ;
  assign n3885 = ( n712 & n3873 ) | ( n712 & ~n3884 ) | ( n3873 & ~n3884 ) ;
  assign n3899 = n3898 ^ n3885 ^ n976 ;
  assign n3914 = ( ~n170 & n897 ) | ( ~n170 & n3149 ) | ( n897 & n3149 ) ;
  assign n3909 = n2203 ^ n1238 ^ n261 ;
  assign n3910 = n3909 ^ n2101 ^ n594 ;
  assign n3911 = ( n140 & n725 ) | ( n140 & ~n2972 ) | ( n725 & ~n2972 ) ;
  assign n3912 = ( n760 & ~n1181 ) | ( n760 & n3911 ) | ( ~n1181 & n3911 ) ;
  assign n3913 = ( ~n2706 & n3910 ) | ( ~n2706 & n3912 ) | ( n3910 & n3912 ) ;
  assign n3904 = ( x1 & n182 ) | ( x1 & ~n550 ) | ( n182 & ~n550 ) ;
  assign n3905 = n2583 ^ x103 ^ x79 ;
  assign n3906 = ( n3384 & n3904 ) | ( n3384 & ~n3905 ) | ( n3904 & ~n3905 ) ;
  assign n3907 = n3906 ^ n1333 ^ n620 ;
  assign n3903 = n3539 ^ n3273 ^ n633 ;
  assign n3900 = n881 ^ n227 ^ x6 ;
  assign n3901 = n3900 ^ n758 ^ x67 ;
  assign n3902 = ( n875 & n3349 ) | ( n875 & n3901 ) | ( n3349 & n3901 ) ;
  assign n3908 = n3907 ^ n3903 ^ n3902 ;
  assign n3915 = n3914 ^ n3913 ^ n3908 ;
  assign n3916 = ( ~n2190 & n2748 ) | ( ~n2190 & n3597 ) | ( n2748 & n3597 ) ;
  assign n3917 = ( x57 & ~n545 ) | ( x57 & n2432 ) | ( ~n545 & n2432 ) ;
  assign n3918 = n3831 ^ n2871 ^ x35 ;
  assign n3919 = n3918 ^ n3510 ^ n1284 ;
  assign n3920 = ( ~n3175 & n3917 ) | ( ~n3175 & n3919 ) | ( n3917 & n3919 ) ;
  assign n3921 = ( n660 & n1413 ) | ( n660 & ~n2148 ) | ( n1413 & ~n2148 ) ;
  assign n3922 = ( ~n775 & n1953 ) | ( ~n775 & n3921 ) | ( n1953 & n3921 ) ;
  assign n3924 = n3369 ^ n2329 ^ n2030 ;
  assign n3923 = n1945 ^ n1595 ^ n626 ;
  assign n3925 = n3924 ^ n3923 ^ n3157 ;
  assign n3926 = ( ~x49 & n3922 ) | ( ~x49 & n3925 ) | ( n3922 & n3925 ) ;
  assign n3929 = ( n1030 & n1705 ) | ( n1030 & ~n2753 ) | ( n1705 & ~n2753 ) ;
  assign n3930 = n3929 ^ n2939 ^ n1450 ;
  assign n3927 = ( n815 & n1074 ) | ( n815 & ~n1094 ) | ( n1074 & ~n1094 ) ;
  assign n3928 = ( ~n2970 & n3552 ) | ( ~n2970 & n3927 ) | ( n3552 & n3927 ) ;
  assign n3931 = n3930 ^ n3928 ^ n2231 ;
  assign n3939 = n1267 ^ n953 ^ n424 ;
  assign n3940 = n3939 ^ n1646 ^ n756 ;
  assign n3933 = n1607 ^ n622 ^ n217 ;
  assign n3932 = n1134 ^ n1128 ^ n523 ;
  assign n3934 = n3933 ^ n3932 ^ n281 ;
  assign n3935 = n3934 ^ n1047 ^ n260 ;
  assign n3936 = n3935 ^ n1537 ^ n247 ;
  assign n3937 = n3936 ^ n3785 ^ n2111 ;
  assign n3938 = ( n739 & n2352 ) | ( n739 & n3937 ) | ( n2352 & n3937 ) ;
  assign n3941 = n3940 ^ n3938 ^ n2526 ;
  assign n3942 = n3941 ^ n3457 ^ n2117 ;
  assign n3950 = ( n131 & n1598 ) | ( n131 & n2986 ) | ( n1598 & n2986 ) ;
  assign n3951 = ( n198 & n3301 ) | ( n198 & ~n3950 ) | ( n3301 & ~n3950 ) ;
  assign n3952 = n3951 ^ n2023 ^ n726 ;
  assign n3946 = n3186 ^ n2711 ^ n1643 ;
  assign n3947 = ( ~n1493 & n1907 ) | ( ~n1493 & n3946 ) | ( n1907 & n3946 ) ;
  assign n3948 = n3947 ^ n3149 ^ n578 ;
  assign n3944 = ( ~n325 & n1767 ) | ( ~n325 & n3239 ) | ( n1767 & n3239 ) ;
  assign n3943 = ( n2212 & n2965 ) | ( n2212 & ~n3634 ) | ( n2965 & ~n3634 ) ;
  assign n3945 = n3944 ^ n3943 ^ n2298 ;
  assign n3949 = n3948 ^ n3945 ^ n663 ;
  assign n3953 = n3952 ^ n3949 ^ n2591 ;
  assign n3954 = ( n1680 & ~n3942 ) | ( n1680 & n3953 ) | ( ~n3942 & n3953 ) ;
  assign n3955 = ( n3926 & ~n3931 ) | ( n3926 & n3954 ) | ( ~n3931 & n3954 ) ;
  assign n3956 = ( ~n934 & n949 ) | ( ~n934 & n2629 ) | ( n949 & n2629 ) ;
  assign n3957 = n3956 ^ n734 ^ n521 ;
  assign n3958 = n3957 ^ n2662 ^ n1904 ;
  assign n3959 = ( x94 & n1390 ) | ( x94 & n2691 ) | ( n1390 & n2691 ) ;
  assign n3960 = n1263 ^ n1184 ^ n761 ;
  assign n3961 = n3960 ^ n2871 ^ n443 ;
  assign n3962 = ( n2274 & n3959 ) | ( n2274 & ~n3961 ) | ( n3959 & ~n3961 ) ;
  assign n3963 = n3962 ^ n2607 ^ n709 ;
  assign n3965 = n3047 ^ n1142 ^ n917 ;
  assign n3964 = ( n385 & n2758 ) | ( n385 & ~n3281 ) | ( n2758 & ~n3281 ) ;
  assign n3966 = n3965 ^ n3964 ^ n1503 ;
  assign n3967 = ( n3227 & n3494 ) | ( n3227 & n3966 ) | ( n3494 & n3966 ) ;
  assign n3973 = n2633 ^ n1119 ^ x108 ;
  assign n3970 = ( n211 & n557 ) | ( n211 & ~n1155 ) | ( n557 & ~n1155 ) ;
  assign n3971 = n1607 ^ n1566 ^ n872 ;
  assign n3972 = ( n2077 & n3970 ) | ( n2077 & n3971 ) | ( n3970 & n3971 ) ;
  assign n3974 = n3973 ^ n3972 ^ n882 ;
  assign n3975 = n3974 ^ n3178 ^ n965 ;
  assign n3968 = ( ~n2428 & n2917 ) | ( ~n2428 & n3818 ) | ( n2917 & n3818 ) ;
  assign n3969 = n3968 ^ n1578 ^ n1551 ;
  assign n3976 = n3975 ^ n3969 ^ n846 ;
  assign n3977 = n2303 ^ n936 ^ n232 ;
  assign n3978 = ( n944 & n2225 ) | ( n944 & n3977 ) | ( n2225 & n3977 ) ;
  assign n3979 = n1713 ^ n1127 ^ n916 ;
  assign n3980 = ( n270 & n3978 ) | ( n270 & ~n3979 ) | ( n3978 & ~n3979 ) ;
  assign n3981 = ( ~n1505 & n1979 ) | ( ~n1505 & n3980 ) | ( n1979 & n3980 ) ;
  assign n3982 = ( n3967 & ~n3976 ) | ( n3967 & n3981 ) | ( ~n3976 & n3981 ) ;
  assign n3983 = ( ~n3530 & n3963 ) | ( ~n3530 & n3982 ) | ( n3963 & n3982 ) ;
  assign n3989 = n3239 ^ n1417 ^ n768 ;
  assign n3990 = n3450 ^ n3322 ^ n2112 ;
  assign n3991 = ( n3577 & ~n3989 ) | ( n3577 & n3990 ) | ( ~n3989 & n3990 ) ;
  assign n3992 = ( n971 & n3510 ) | ( n971 & ~n3991 ) | ( n3510 & ~n3991 ) ;
  assign n3985 = ( n290 & n1626 ) | ( n290 & ~n3686 ) | ( n1626 & ~n3686 ) ;
  assign n3984 = ( n702 & n859 ) | ( n702 & n1196 ) | ( n859 & n1196 ) ;
  assign n3986 = n3985 ^ n3984 ^ n415 ;
  assign n3987 = ( n176 & n1128 ) | ( n176 & n3986 ) | ( n1128 & n3986 ) ;
  assign n3988 = n3987 ^ n3291 ^ n2190 ;
  assign n3993 = n3992 ^ n3988 ^ n2134 ;
  assign n3994 = n3993 ^ n1492 ^ x96 ;
  assign n3995 = n3007 ^ n2022 ^ n793 ;
  assign n3996 = n3995 ^ n3189 ^ n1074 ;
  assign n3997 = ( ~n1129 & n3203 ) | ( ~n1129 & n3996 ) | ( n3203 & n3996 ) ;
  assign n3998 = n3997 ^ n2108 ^ n218 ;
  assign n4014 = ( n263 & n1536 ) | ( n263 & ~n3896 ) | ( n1536 & ~n3896 ) ;
  assign n4015 = n4014 ^ n1222 ^ n1004 ;
  assign n4010 = n2656 ^ n1744 ^ n1691 ;
  assign n4011 = ( n690 & n1661 ) | ( n690 & ~n4010 ) | ( n1661 & ~n4010 ) ;
  assign n4012 = n3603 ^ n3147 ^ n1769 ;
  assign n4013 = ( n2614 & n4011 ) | ( n2614 & ~n4012 ) | ( n4011 & ~n4012 ) ;
  assign n4016 = n4015 ^ n4013 ^ n2342 ;
  assign n4001 = n1111 ^ n735 ^ x117 ;
  assign n4002 = ( n989 & ~n1647 ) | ( n989 & n4001 ) | ( ~n1647 & n4001 ) ;
  assign n3999 = n3100 ^ n627 ^ x97 ;
  assign n4000 = n3999 ^ n585 ^ n427 ;
  assign n4003 = n4002 ^ n4000 ^ n782 ;
  assign n4004 = n4003 ^ n1635 ^ n310 ;
  assign n4005 = n4004 ^ n2467 ^ n412 ;
  assign n4006 = n3344 ^ n3259 ^ n730 ;
  assign n4007 = n2742 ^ n1076 ^ x40 ;
  assign n4008 = ( n693 & n1404 ) | ( n693 & ~n4007 ) | ( n1404 & ~n4007 ) ;
  assign n4009 = ( n4005 & ~n4006 ) | ( n4005 & n4008 ) | ( ~n4006 & n4008 ) ;
  assign n4017 = n4016 ^ n4009 ^ n2747 ;
  assign n4019 = n4010 ^ n1551 ^ n1223 ;
  assign n4020 = n3320 ^ n1207 ^ n180 ;
  assign n4021 = ( n844 & n4019 ) | ( n844 & ~n4020 ) | ( n4019 & ~n4020 ) ;
  assign n4018 = ( n640 & n2712 ) | ( n640 & n3262 ) | ( n2712 & n3262 ) ;
  assign n4022 = n4021 ^ n4018 ^ n3122 ;
  assign n4032 = ( n2497 & n3361 ) | ( n2497 & ~n3613 ) | ( n3361 & ~n3613 ) ;
  assign n4030 = n2183 ^ n301 ^ n276 ;
  assign n4031 = n4030 ^ n3125 ^ n566 ;
  assign n4023 = n1212 ^ n862 ^ n650 ;
  assign n4024 = ( n363 & ~n2867 ) | ( n363 & n4023 ) | ( ~n2867 & n4023 ) ;
  assign n4025 = n4024 ^ n1125 ^ n894 ;
  assign n4027 = ( n413 & n794 ) | ( n413 & n1499 ) | ( n794 & n1499 ) ;
  assign n4026 = n1561 ^ n1232 ^ n587 ;
  assign n4028 = n4027 ^ n4026 ^ n194 ;
  assign n4029 = ( n875 & n4025 ) | ( n875 & n4028 ) | ( n4025 & n4028 ) ;
  assign n4033 = n4032 ^ n4031 ^ n4029 ;
  assign n4055 = n908 ^ n715 ^ x72 ;
  assign n4053 = n1825 ^ n1630 ^ n625 ;
  assign n4052 = n769 ^ n502 ^ n259 ;
  assign n4054 = n4053 ^ n4052 ^ n3731 ;
  assign n4056 = n4055 ^ n4054 ^ n3503 ;
  assign n4034 = ( ~n775 & n908 ) | ( ~n775 & n2583 ) | ( n908 & n2583 ) ;
  assign n4035 = n3934 ^ n3348 ^ n193 ;
  assign n4036 = n4035 ^ n3381 ^ x83 ;
  assign n4037 = ( n2633 & ~n4034 ) | ( n2633 & n4036 ) | ( ~n4034 & n4036 ) ;
  assign n4038 = n3210 ^ n1169 ^ n828 ;
  assign n4046 = ( n230 & n2546 ) | ( n230 & ~n2773 ) | ( n2546 & ~n2773 ) ;
  assign n4045 = ( n1309 & ~n1768 ) | ( n1309 & n3018 ) | ( ~n1768 & n3018 ) ;
  assign n4044 = n3734 ^ n3041 ^ n1530 ;
  assign n4047 = n4046 ^ n4045 ^ n4044 ;
  assign n4048 = ( n412 & n3205 ) | ( n412 & n4047 ) | ( n3205 & n4047 ) ;
  assign n4049 = ( n1937 & ~n3015 ) | ( n1937 & n4048 ) | ( ~n3015 & n4048 ) ;
  assign n4041 = ( n149 & n1435 ) | ( n149 & ~n3161 ) | ( n1435 & ~n3161 ) ;
  assign n4042 = ( ~n342 & n2071 ) | ( ~n342 & n4041 ) | ( n2071 & n4041 ) ;
  assign n4039 = n2414 ^ n955 ^ n621 ;
  assign n4040 = ( n2479 & ~n3336 ) | ( n2479 & n4039 ) | ( ~n3336 & n4039 ) ;
  assign n4043 = n4042 ^ n4040 ^ n589 ;
  assign n4050 = n4049 ^ n4043 ^ n481 ;
  assign n4051 = ( n4037 & n4038 ) | ( n4037 & ~n4050 ) | ( n4038 & ~n4050 ) ;
  assign n4057 = n4056 ^ n4051 ^ n1514 ;
  assign n4058 = n1589 ^ n994 ^ x75 ;
  assign n4069 = ( ~n348 & n421 ) | ( ~n348 & n1326 ) | ( n421 & n1326 ) ;
  assign n4070 = n4069 ^ n3669 ^ n1016 ;
  assign n4071 = n4070 ^ n2481 ^ n1129 ;
  assign n4072 = ( n1358 & ~n3036 ) | ( n1358 & n3808 ) | ( ~n3036 & n3808 ) ;
  assign n4073 = ( n527 & n4071 ) | ( n527 & n4072 ) | ( n4071 & n4072 ) ;
  assign n4064 = ( x79 & ~n378 ) | ( x79 & n1661 ) | ( ~n378 & n1661 ) ;
  assign n4059 = ( n187 & n2546 ) | ( n187 & n2578 ) | ( n2546 & n2578 ) ;
  assign n4060 = ( ~n550 & n1244 ) | ( ~n550 & n1488 ) | ( n1244 & n1488 ) ;
  assign n4061 = ( n132 & n960 ) | ( n132 & n4060 ) | ( n960 & n4060 ) ;
  assign n4062 = n4061 ^ n1679 ^ n1522 ;
  assign n4063 = ( n1002 & n4059 ) | ( n1002 & n4062 ) | ( n4059 & n4062 ) ;
  assign n4065 = n4064 ^ n4063 ^ n2692 ;
  assign n4066 = n4065 ^ n1470 ^ n1107 ;
  assign n4067 = n4066 ^ n2467 ^ n1852 ;
  assign n4068 = ( n371 & ~n1560 ) | ( n371 & n4067 ) | ( ~n1560 & n4067 ) ;
  assign n4074 = n4073 ^ n4068 ^ n2752 ;
  assign n4075 = ( n1628 & n4058 ) | ( n1628 & n4074 ) | ( n4058 & n4074 ) ;
  assign n4103 = n2136 ^ n1297 ^ n245 ;
  assign n4104 = ( n185 & n3728 ) | ( n185 & n4103 ) | ( n3728 & n4103 ) ;
  assign n4105 = ( n1791 & n3002 ) | ( n1791 & ~n4104 ) | ( n3002 & ~n4104 ) ;
  assign n4101 = ( n1613 & n1736 ) | ( n1613 & n3456 ) | ( n1736 & n3456 ) ;
  assign n4098 = n524 ^ n439 ^ n375 ;
  assign n4099 = ( n601 & n3986 ) | ( n601 & ~n4098 ) | ( n3986 & ~n4098 ) ;
  assign n4100 = ( n2462 & n3517 ) | ( n2462 & n4099 ) | ( n3517 & n4099 ) ;
  assign n4095 = ( x112 & ~n736 ) | ( x112 & n1846 ) | ( ~n736 & n1846 ) ;
  assign n4096 = ( n962 & ~n4030 ) | ( n962 & n4095 ) | ( ~n4030 & n4095 ) ;
  assign n4097 = n4096 ^ n3544 ^ n434 ;
  assign n4102 = n4101 ^ n4100 ^ n4097 ;
  assign n4080 = ( x126 & ~n2803 ) | ( x126 & n3052 ) | ( ~n2803 & n3052 ) ;
  assign n4077 = ( n1279 & n1343 ) | ( n1279 & n2281 ) | ( n1343 & n2281 ) ;
  assign n4078 = ( ~n310 & n3516 ) | ( ~n310 & n4077 ) | ( n3516 & n4077 ) ;
  assign n4076 = n2565 ^ n1476 ^ n1028 ;
  assign n4079 = n4078 ^ n4076 ^ n553 ;
  assign n4081 = n4080 ^ n4079 ^ n2837 ;
  assign n4082 = ( ~n2752 & n3029 ) | ( ~n2752 & n3863 ) | ( n3029 & n3863 ) ;
  assign n4083 = ( n1090 & ~n1804 ) | ( n1090 & n4082 ) | ( ~n1804 & n4082 ) ;
  assign n4084 = n2513 ^ n2433 ^ n971 ;
  assign n4085 = ( n2528 & n2911 ) | ( n2528 & n4084 ) | ( n2911 & n4084 ) ;
  assign n4086 = n3456 ^ n3285 ^ n883 ;
  assign n4089 = n3029 ^ n1083 ^ n487 ;
  assign n4090 = n4089 ^ n1433 ^ n1285 ;
  assign n4087 = ( ~n401 & n988 ) | ( ~n401 & n1730 ) | ( n988 & n1730 ) ;
  assign n4088 = n4087 ^ n2719 ^ n1756 ;
  assign n4091 = n4090 ^ n4088 ^ n2101 ;
  assign n4092 = ( n1776 & n3284 ) | ( n1776 & ~n4091 ) | ( n3284 & ~n4091 ) ;
  assign n4093 = ( n4085 & ~n4086 ) | ( n4085 & n4092 ) | ( ~n4086 & n4092 ) ;
  assign n4094 = ( n4081 & n4083 ) | ( n4081 & n4093 ) | ( n4083 & n4093 ) ;
  assign n4106 = n4105 ^ n4102 ^ n4094 ;
  assign n4115 = n2939 ^ n1356 ^ n1119 ;
  assign n4116 = n4115 ^ n3429 ^ n3263 ;
  assign n4113 = n2087 ^ n1445 ^ n645 ;
  assign n4110 = ( n209 & n1022 ) | ( n209 & ~n2103 ) | ( n1022 & ~n2103 ) ;
  assign n4111 = n4110 ^ n2247 ^ n392 ;
  assign n4109 = ( ~n1378 & n1733 ) | ( ~n1378 & n1875 ) | ( n1733 & n1875 ) ;
  assign n4112 = n4111 ^ n4109 ^ n440 ;
  assign n4107 = n1440 ^ n1422 ^ n1028 ;
  assign n4108 = ( n2300 & n2755 ) | ( n2300 & n4107 ) | ( n2755 & n4107 ) ;
  assign n4114 = n4113 ^ n4112 ^ n4108 ;
  assign n4117 = n4116 ^ n4114 ^ n539 ;
  assign n4118 = ( ~n224 & n326 ) | ( ~n224 & n4117 ) | ( n326 & n4117 ) ;
  assign n4119 = ( n692 & ~n726 ) | ( n692 & n1967 ) | ( ~n726 & n1967 ) ;
  assign n4120 = ( ~n1087 & n2663 ) | ( ~n1087 & n4119 ) | ( n2663 & n4119 ) ;
  assign n4132 = n1485 ^ n829 ^ n349 ;
  assign n4131 = ( n1204 & ~n2094 ) | ( n1204 & n3463 ) | ( ~n2094 & n3463 ) ;
  assign n4133 = n4132 ^ n4131 ^ n480 ;
  assign n4134 = ( n1431 & ~n3351 ) | ( n1431 & n4133 ) | ( ~n3351 & n4133 ) ;
  assign n4130 = n2719 ^ n1811 ^ n1242 ;
  assign n4135 = n4134 ^ n4130 ^ n3162 ;
  assign n4127 = ( n139 & n1515 ) | ( n139 & n2264 ) | ( n1515 & n2264 ) ;
  assign n4128 = n4127 ^ n2793 ^ n1642 ;
  assign n4129 = n4128 ^ n3067 ^ n1973 ;
  assign n4136 = n4135 ^ n4129 ^ n1053 ;
  assign n4123 = n591 ^ n524 ^ n229 ;
  assign n4124 = n4123 ^ n2753 ^ n556 ;
  assign n4125 = ( n259 & n814 ) | ( n259 & n4124 ) | ( n814 & n4124 ) ;
  assign n4121 = ( ~n1360 & n2386 ) | ( ~n1360 & n3853 ) | ( n2386 & n3853 ) ;
  assign n4122 = ( ~n1368 & n3033 ) | ( ~n1368 & n4121 ) | ( n3033 & n4121 ) ;
  assign n4126 = n4125 ^ n4122 ^ n2624 ;
  assign n4137 = n4136 ^ n4126 ^ n809 ;
  assign n4138 = ( ~n2337 & n4120 ) | ( ~n2337 & n4137 ) | ( n4120 & n4137 ) ;
  assign n4139 = n3093 ^ n2449 ^ n2115 ;
  assign n4162 = ( n367 & ~n1009 ) | ( n367 & n1010 ) | ( ~n1009 & n1010 ) ;
  assign n4158 = ( ~n415 & n711 ) | ( ~n415 & n753 ) | ( n711 & n753 ) ;
  assign n4159 = n4158 ^ n3523 ^ n2692 ;
  assign n4160 = ( n2141 & n2341 ) | ( n2141 & ~n4159 ) | ( n2341 & ~n4159 ) ;
  assign n4157 = n2733 ^ n2465 ^ n732 ;
  assign n4161 = n4160 ^ n4157 ^ n1943 ;
  assign n4163 = n4162 ^ n4161 ^ n2347 ;
  assign n4143 = ( x5 & n1633 ) | ( x5 & n2790 ) | ( n1633 & n2790 ) ;
  assign n4144 = n2461 ^ n928 ^ n178 ;
  assign n4145 = n4144 ^ n2059 ^ n511 ;
  assign n4146 = ( n1743 & n2436 ) | ( n1743 & n4145 ) | ( n2436 & n4145 ) ;
  assign n4147 = ( ~n2169 & n4143 ) | ( ~n2169 & n4146 ) | ( n4143 & n4146 ) ;
  assign n4140 = ( x115 & n943 ) | ( x115 & ~n1212 ) | ( n943 & ~n1212 ) ;
  assign n4141 = n2242 ^ n451 ^ x8 ;
  assign n4142 = ( n1845 & n4140 ) | ( n1845 & ~n4141 ) | ( n4140 & ~n4141 ) ;
  assign n4148 = n4147 ^ n4142 ^ n3129 ;
  assign n4149 = ( n3307 & ~n3677 ) | ( n3307 & n4148 ) | ( ~n3677 & n4148 ) ;
  assign n4153 = ( n771 & n1989 ) | ( n771 & ~n2995 ) | ( n1989 & ~n2995 ) ;
  assign n4150 = ( x103 & n179 ) | ( x103 & n1449 ) | ( n179 & n1449 ) ;
  assign n4151 = ( n455 & ~n576 ) | ( n455 & n4077 ) | ( ~n576 & n4077 ) ;
  assign n4152 = ( n3578 & ~n4150 ) | ( n3578 & n4151 ) | ( ~n4150 & n4151 ) ;
  assign n4154 = n4153 ^ n4152 ^ n1839 ;
  assign n4155 = ( ~n881 & n3867 ) | ( ~n881 & n4154 ) | ( n3867 & n4154 ) ;
  assign n4156 = ( n2279 & n4149 ) | ( n2279 & ~n4155 ) | ( n4149 & ~n4155 ) ;
  assign n4164 = n4163 ^ n4156 ^ n570 ;
  assign n4173 = n1585 ^ n619 ^ n543 ;
  assign n4174 = n4173 ^ n1520 ^ n1076 ;
  assign n4175 = ( n732 & ~n1440 ) | ( n732 & n1986 ) | ( ~n1440 & n1986 ) ;
  assign n4176 = ( ~n3147 & n4174 ) | ( ~n3147 & n4175 ) | ( n4174 & n4175 ) ;
  assign n4165 = ( n2502 & n3017 ) | ( n2502 & ~n3634 ) | ( n3017 & ~n3634 ) ;
  assign n4169 = n2492 ^ n2244 ^ n165 ;
  assign n4170 = n4169 ^ n3122 ^ n3017 ;
  assign n4166 = ( ~n516 & n1245 ) | ( ~n516 & n3162 ) | ( n1245 & n3162 ) ;
  assign n4167 = n4166 ^ n2852 ^ n1042 ;
  assign n4168 = n4167 ^ n2088 ^ n1068 ;
  assign n4171 = n4170 ^ n4168 ^ n1942 ;
  assign n4172 = ( n1777 & n4165 ) | ( n1777 & ~n4171 ) | ( n4165 & ~n4171 ) ;
  assign n4177 = n4176 ^ n4172 ^ n984 ;
  assign n4178 = ( ~n2208 & n4009 ) | ( ~n2208 & n4177 ) | ( n4009 & n4177 ) ;
  assign n4192 = ( n434 & n553 ) | ( n434 & n808 ) | ( n553 & n808 ) ;
  assign n4191 = ( ~n285 & n686 ) | ( ~n285 & n1621 ) | ( n686 & n1621 ) ;
  assign n4193 = n4192 ^ n4191 ^ n2482 ;
  assign n4194 = ( n961 & n2870 ) | ( n961 & ~n4193 ) | ( n2870 & ~n4193 ) ;
  assign n4195 = ( n1476 & ~n3706 ) | ( n1476 & n4194 ) | ( ~n3706 & n4194 ) ;
  assign n4179 = n2285 ^ n912 ^ n634 ;
  assign n4180 = n4179 ^ n3417 ^ n907 ;
  assign n4181 = n4180 ^ n3288 ^ n622 ;
  assign n4182 = n4181 ^ n3177 ^ n1261 ;
  assign n4183 = n3207 ^ n386 ^ x118 ;
  assign n4184 = n2023 ^ n1703 ^ n1498 ;
  assign n4185 = n1862 ^ n1836 ^ n536 ;
  assign n4186 = n1392 ^ n1338 ^ n1164 ;
  assign n4187 = ( n4005 & n4185 ) | ( n4005 & n4186 ) | ( n4185 & n4186 ) ;
  assign n4188 = ( n1201 & ~n4184 ) | ( n1201 & n4187 ) | ( ~n4184 & n4187 ) ;
  assign n4189 = ( n3148 & n4183 ) | ( n3148 & n4188 ) | ( n4183 & n4188 ) ;
  assign n4190 = ( n408 & n4182 ) | ( n408 & n4189 ) | ( n4182 & n4189 ) ;
  assign n4196 = n4195 ^ n4190 ^ n3332 ;
  assign n4197 = ( n732 & n836 ) | ( n732 & ~n2333 ) | ( n836 & ~n2333 ) ;
  assign n4198 = ( ~n157 & n867 ) | ( ~n157 & n909 ) | ( n867 & n909 ) ;
  assign n4199 = ( n2263 & ~n4197 ) | ( n2263 & n4198 ) | ( ~n4197 & n4198 ) ;
  assign n4200 = n4199 ^ n3078 ^ n1393 ;
  assign n4201 = n4200 ^ n2981 ^ n2526 ;
  assign n4202 = n751 ^ n409 ^ n232 ;
  assign n4203 = n4202 ^ n2857 ^ n681 ;
  assign n4204 = ( ~n950 & n3985 ) | ( ~n950 & n4090 ) | ( n3985 & n4090 ) ;
  assign n4205 = n4204 ^ n1295 ^ n1015 ;
  assign n4206 = n4205 ^ n3765 ^ n690 ;
  assign n4207 = ( n645 & ~n942 ) | ( n645 & n4206 ) | ( ~n942 & n4206 ) ;
  assign n4208 = ( n1232 & ~n2730 ) | ( n1232 & n4207 ) | ( ~n2730 & n4207 ) ;
  assign n4228 = n2376 ^ n2137 ^ n226 ;
  assign n4224 = ( x62 & n1557 ) | ( x62 & n3476 ) | ( n1557 & n3476 ) ;
  assign n4225 = n4224 ^ n2252 ^ n1948 ;
  assign n4226 = ( n2132 & n2201 ) | ( n2132 & n4225 ) | ( n2201 & n4225 ) ;
  assign n4227 = n4226 ^ n1690 ^ n943 ;
  assign n4229 = n4228 ^ n4227 ^ n509 ;
  assign n4220 = ( n260 & ~n1607 ) | ( n260 & n2027 ) | ( ~n1607 & n2027 ) ;
  assign n4221 = n4220 ^ n3025 ^ n312 ;
  assign n4222 = n4221 ^ n1679 ^ n1521 ;
  assign n4209 = n2409 ^ n1683 ^ n805 ;
  assign n4214 = ( x41 & ~x79 ) | ( x41 & n234 ) | ( ~x79 & n234 ) ;
  assign n4215 = n767 ^ n761 ^ n134 ;
  assign n4216 = ( n1557 & ~n2212 ) | ( n1557 & n4215 ) | ( ~n2212 & n4215 ) ;
  assign n4217 = ( n2639 & ~n4214 ) | ( n2639 & n4216 ) | ( ~n4214 & n4216 ) ;
  assign n4212 = ( n406 & n1281 ) | ( n406 & n2946 ) | ( n1281 & n2946 ) ;
  assign n4210 = n1924 ^ n1464 ^ n453 ;
  assign n4211 = ( n479 & n2485 ) | ( n479 & n4210 ) | ( n2485 & n4210 ) ;
  assign n4213 = n4212 ^ n4211 ^ n129 ;
  assign n4218 = n4217 ^ n4213 ^ n3972 ;
  assign n4219 = ( ~n1870 & n4209 ) | ( ~n1870 & n4218 ) | ( n4209 & n4218 ) ;
  assign n4223 = n4222 ^ n4219 ^ n1304 ;
  assign n4230 = n4229 ^ n4223 ^ n1237 ;
  assign n4231 = n4230 ^ n4092 ^ n1717 ;
  assign n4245 = ( n149 & ~n2058 ) | ( n149 & n3070 ) | ( ~n2058 & n3070 ) ;
  assign n4242 = ( n608 & n3391 ) | ( n608 & n3877 ) | ( n3391 & n3877 ) ;
  assign n4243 = n4242 ^ n3667 ^ n3094 ;
  assign n4244 = ( n2180 & ~n3091 ) | ( n2180 & n4243 ) | ( ~n3091 & n4243 ) ;
  assign n4232 = n2339 ^ n1665 ^ n339 ;
  assign n4233 = ( n2082 & n2376 ) | ( n2082 & ~n4232 ) | ( n2376 & ~n4232 ) ;
  assign n4235 = ( n1093 & n1406 ) | ( n1093 & ~n1486 ) | ( n1406 & ~n1486 ) ;
  assign n4236 = ( n172 & n258 ) | ( n172 & ~n991 ) | ( n258 & ~n991 ) ;
  assign n4237 = ( n392 & n4235 ) | ( n392 & ~n4236 ) | ( n4235 & ~n4236 ) ;
  assign n4238 = n4237 ^ n2007 ^ n292 ;
  assign n4234 = n3190 ^ n1823 ^ n811 ;
  assign n4239 = n4238 ^ n4234 ^ n212 ;
  assign n4240 = ( n406 & ~n4233 ) | ( n406 & n4239 ) | ( ~n4233 & n4239 ) ;
  assign n4241 = ( ~n1596 & n3684 ) | ( ~n1596 & n4240 ) | ( n3684 & n4240 ) ;
  assign n4246 = n4245 ^ n4244 ^ n4241 ;
  assign n4247 = ( ~n1133 & n2156 ) | ( ~n1133 & n3946 ) | ( n2156 & n3946 ) ;
  assign n4248 = ( ~n282 & n455 ) | ( ~n282 & n1110 ) | ( n455 & n1110 ) ;
  assign n4249 = n4248 ^ n1262 ^ x9 ;
  assign n4250 = n4249 ^ n3043 ^ n775 ;
  assign n4251 = ( n536 & n800 ) | ( n536 & n2386 ) | ( n800 & n2386 ) ;
  assign n4252 = ( n4247 & ~n4250 ) | ( n4247 & n4251 ) | ( ~n4250 & n4251 ) ;
  assign n4253 = n2781 ^ n1989 ^ n768 ;
  assign n4254 = n4253 ^ n2244 ^ n376 ;
  assign n4255 = n4254 ^ n1178 ^ n400 ;
  assign n4256 = ( n985 & ~n2023 ) | ( n985 & n3182 ) | ( ~n2023 & n3182 ) ;
  assign n4257 = ( n836 & n960 ) | ( n836 & n3807 ) | ( n960 & n3807 ) ;
  assign n4258 = ( n1590 & n3368 ) | ( n1590 & n4257 ) | ( n3368 & n4257 ) ;
  assign n4259 = ( n1343 & ~n4256 ) | ( n1343 & n4258 ) | ( ~n4256 & n4258 ) ;
  assign n4260 = ( ~n2367 & n3455 ) | ( ~n2367 & n4259 ) | ( n3455 & n4259 ) ;
  assign n4261 = n4260 ^ n3591 ^ n865 ;
  assign n4262 = ( n4252 & n4255 ) | ( n4252 & ~n4261 ) | ( n4255 & ~n4261 ) ;
  assign n4263 = ( n828 & ~n1035 ) | ( n828 & n2173 ) | ( ~n1035 & n2173 ) ;
  assign n4264 = n2941 ^ n1310 ^ n797 ;
  assign n4265 = ( n2315 & n2564 ) | ( n2315 & n4264 ) | ( n2564 & n4264 ) ;
  assign n4266 = n4265 ^ n2021 ^ x115 ;
  assign n4267 = ( n1895 & ~n3194 ) | ( n1895 & n4266 ) | ( ~n3194 & n4266 ) ;
  assign n4268 = ( n2220 & n4263 ) | ( n2220 & n4267 ) | ( n4263 & n4267 ) ;
  assign n4275 = n2195 ^ n1414 ^ n378 ;
  assign n4274 = n1688 ^ n1358 ^ n705 ;
  assign n4269 = n2378 ^ n2278 ^ n822 ;
  assign n4270 = ( n309 & n1088 ) | ( n309 & n4269 ) | ( n1088 & n4269 ) ;
  assign n4271 = ( n1557 & n1571 ) | ( n1557 & ~n4270 ) | ( n1571 & ~n4270 ) ;
  assign n4272 = n4271 ^ n1579 ^ n1525 ;
  assign n4273 = ( n474 & n1293 ) | ( n474 & ~n4272 ) | ( n1293 & ~n4272 ) ;
  assign n4276 = n4275 ^ n4274 ^ n4273 ;
  assign n4277 = n4276 ^ n2760 ^ n1573 ;
  assign n4278 = ( n576 & ~n1353 ) | ( n576 & n2722 ) | ( ~n1353 & n2722 ) ;
  assign n4279 = n4278 ^ n692 ^ x66 ;
  assign n4280 = ( ~n1054 & n2204 ) | ( ~n1054 & n4279 ) | ( n2204 & n4279 ) ;
  assign n4281 = n4146 ^ n3825 ^ n3128 ;
  assign n4282 = ( ~n2141 & n3610 ) | ( ~n2141 & n4281 ) | ( n3610 & n4281 ) ;
  assign n4283 = n3187 ^ n1631 ^ n335 ;
  assign n4284 = ( ~n541 & n1274 ) | ( ~n541 & n4283 ) | ( n1274 & n4283 ) ;
  assign n4285 = n3651 ^ n3109 ^ n2845 ;
  assign n4286 = ( n1266 & n1650 ) | ( n1266 & ~n4285 ) | ( n1650 & ~n4285 ) ;
  assign n4287 = ( n996 & ~n1345 ) | ( n996 & n2721 ) | ( ~n1345 & n2721 ) ;
  assign n4288 = ( ~n1006 & n2384 ) | ( ~n1006 & n4287 ) | ( n2384 & n4287 ) ;
  assign n4289 = ( n4284 & n4286 ) | ( n4284 & ~n4288 ) | ( n4286 & ~n4288 ) ;
  assign n4295 = n3321 ^ n2755 ^ n2492 ;
  assign n4293 = n2416 ^ n1705 ^ n287 ;
  assign n4291 = ( n136 & ~n295 ) | ( n136 & n362 ) | ( ~n295 & n362 ) ;
  assign n4292 = n4291 ^ n2465 ^ n2252 ;
  assign n4294 = n4293 ^ n4292 ^ n1154 ;
  assign n4290 = n3644 ^ n1879 ^ x24 ;
  assign n4296 = n4295 ^ n4294 ^ n4290 ;
  assign n4297 = n3905 ^ n2222 ^ n352 ;
  assign n4298 = ( ~n490 & n1367 ) | ( ~n490 & n1980 ) | ( n1367 & n1980 ) ;
  assign n4299 = n4298 ^ n2012 ^ x67 ;
  assign n4300 = ( n3150 & ~n3835 ) | ( n3150 & n4299 ) | ( ~n3835 & n4299 ) ;
  assign n4301 = ( n3398 & ~n4297 ) | ( n3398 & n4300 ) | ( ~n4297 & n4300 ) ;
  assign n4302 = ( n2506 & n2726 ) | ( n2506 & n4301 ) | ( n2726 & n4301 ) ;
  assign n4303 = ( n4289 & ~n4296 ) | ( n4289 & n4302 ) | ( ~n4296 & n4302 ) ;
  assign n4304 = ( n4280 & n4282 ) | ( n4280 & n4303 ) | ( n4282 & n4303 ) ;
  assign n4315 = n4291 ^ n1028 ^ n738 ;
  assign n4316 = n4315 ^ n3428 ^ n1991 ;
  assign n4312 = n1867 ^ n1355 ^ n762 ;
  assign n4313 = ( n1971 & n3721 ) | ( n1971 & ~n4312 ) | ( n3721 & ~n4312 ) ;
  assign n4310 = n3810 ^ n327 ^ n140 ;
  assign n4306 = ( n1207 & n2083 ) | ( n1207 & ~n3294 ) | ( n2083 & ~n3294 ) ;
  assign n4307 = ( x11 & n2054 ) | ( x11 & ~n4306 ) | ( n2054 & ~n4306 ) ;
  assign n4308 = ( n160 & n237 ) | ( n160 & ~n4307 ) | ( n237 & ~n4307 ) ;
  assign n4309 = n4308 ^ n1899 ^ n1299 ;
  assign n4311 = n4310 ^ n4309 ^ n2144 ;
  assign n4305 = n3004 ^ n1712 ^ x37 ;
  assign n4314 = n4313 ^ n4311 ^ n4305 ;
  assign n4317 = n4316 ^ n4314 ^ n1369 ;
  assign n4318 = n3511 ^ n3448 ^ n940 ;
  assign n4319 = n4318 ^ n2213 ^ n317 ;
  assign n4320 = ( n1876 & ~n3025 ) | ( n1876 & n4319 ) | ( ~n3025 & n4319 ) ;
  assign n4321 = ( n154 & n1028 ) | ( n154 & ~n2682 ) | ( n1028 & ~n2682 ) ;
  assign n4322 = n4321 ^ n4041 ^ n1404 ;
  assign n4327 = ( n676 & n1421 ) | ( n676 & ~n1676 ) | ( n1421 & ~n1676 ) ;
  assign n4328 = n4327 ^ n1467 ^ n1440 ;
  assign n4329 = ( ~n257 & n3824 ) | ( ~n257 & n4328 ) | ( n3824 & n4328 ) ;
  assign n4323 = n1424 ^ n896 ^ n751 ;
  assign n4324 = n4323 ^ n2292 ^ n1609 ;
  assign n4325 = ( n1431 & n2750 ) | ( n1431 & ~n4324 ) | ( n2750 & ~n4324 ) ;
  assign n4326 = ( ~n2068 & n3701 ) | ( ~n2068 & n4325 ) | ( n3701 & n4325 ) ;
  assign n4330 = n4329 ^ n4326 ^ x14 ;
  assign n4331 = ( n2315 & n4287 ) | ( n2315 & ~n4330 ) | ( n4287 & ~n4330 ) ;
  assign n4332 = n3875 ^ n2460 ^ n2419 ;
  assign n4333 = ( ~n4322 & n4331 ) | ( ~n4322 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4334 = ( n1241 & ~n2684 ) | ( n1241 & n3652 ) | ( ~n2684 & n3652 ) ;
  assign n4335 = n1874 ^ n1209 ^ n842 ;
  assign n4336 = n2362 ^ n1219 ^ x35 ;
  assign n4337 = ( n4334 & ~n4335 ) | ( n4334 & n4336 ) | ( ~n4335 & n4336 ) ;
  assign n4338 = n4193 ^ n3281 ^ n2386 ;
  assign n4339 = ( n649 & ~n1005 ) | ( n649 & n4338 ) | ( ~n1005 & n4338 ) ;
  assign n4352 = n1884 ^ n701 ^ n515 ;
  assign n4353 = n4352 ^ n2750 ^ n608 ;
  assign n4351 = ( n181 & ~n730 ) | ( n181 & n3986 ) | ( ~n730 & n3986 ) ;
  assign n4354 = n4353 ^ n4351 ^ n1616 ;
  assign n4348 = ( x107 & ~n535 ) | ( x107 & n3567 ) | ( ~n535 & n3567 ) ;
  assign n4349 = n4348 ^ n1077 ^ n812 ;
  assign n4345 = ( n503 & ~n743 ) | ( n503 & n1834 ) | ( ~n743 & n1834 ) ;
  assign n4346 = ( ~n1517 & n3639 ) | ( ~n1517 & n4345 ) | ( n3639 & n4345 ) ;
  assign n4347 = ( ~n1224 & n3985 ) | ( ~n1224 & n4346 ) | ( n3985 & n4346 ) ;
  assign n4350 = n4349 ^ n4347 ^ n2059 ;
  assign n4343 = n1804 ^ n1274 ^ x85 ;
  assign n4340 = n2793 ^ n2041 ^ n970 ;
  assign n4341 = ( ~n961 & n3694 ) | ( ~n961 & n4340 ) | ( n3694 & n4340 ) ;
  assign n4342 = ( ~n2590 & n3472 ) | ( ~n2590 & n4341 ) | ( n3472 & n4341 ) ;
  assign n4344 = n4343 ^ n4342 ^ n331 ;
  assign n4355 = n4354 ^ n4350 ^ n4344 ;
  assign n4356 = ( ~n2604 & n4339 ) | ( ~n2604 & n4355 ) | ( n4339 & n4355 ) ;
  assign n4376 = ( n336 & ~n2342 ) | ( n336 & n4175 ) | ( ~n2342 & n4175 ) ;
  assign n4377 = ( ~n2990 & n3921 ) | ( ~n2990 & n4376 ) | ( n3921 & n4376 ) ;
  assign n4380 = n2285 ^ n710 ^ n374 ;
  assign n4378 = n2937 ^ n1991 ^ n1730 ;
  assign n4379 = n4378 ^ n3551 ^ n984 ;
  assign n4381 = n4380 ^ n4379 ^ n702 ;
  assign n4383 = ( ~n1451 & n2178 ) | ( ~n1451 & n2339 ) | ( n2178 & n2339 ) ;
  assign n4384 = n2356 ^ n1129 ^ n267 ;
  assign n4385 = ( ~n274 & n657 ) | ( ~n274 & n4384 ) | ( n657 & n4384 ) ;
  assign n4386 = ( n4077 & ~n4383 ) | ( n4077 & n4385 ) | ( ~n4383 & n4385 ) ;
  assign n4382 = ( ~n564 & n1921 ) | ( ~n564 & n2393 ) | ( n1921 & n2393 ) ;
  assign n4387 = n4386 ^ n4382 ^ n3541 ;
  assign n4388 = ( n4377 & n4381 ) | ( n4377 & ~n4387 ) | ( n4381 & ~n4387 ) ;
  assign n4369 = n1534 ^ n1337 ^ n839 ;
  assign n4370 = ( n795 & n2502 ) | ( n795 & ~n4369 ) | ( n2502 & ~n4369 ) ;
  assign n4371 = n2133 ^ n1476 ^ n1447 ;
  assign n4372 = n4371 ^ n2905 ^ n2697 ;
  assign n4373 = ( n3284 & n4370 ) | ( n3284 & ~n4372 ) | ( n4370 & ~n4372 ) ;
  assign n4374 = ( n966 & ~n3063 ) | ( n966 & n4373 ) | ( ~n3063 & n4373 ) ;
  assign n4366 = n3888 ^ n3418 ^ n3303 ;
  assign n4364 = n1400 ^ n887 ^ n297 ;
  assign n4365 = ( n1529 & ~n3073 ) | ( n1529 & n4364 ) | ( ~n3073 & n4364 ) ;
  assign n4367 = n4366 ^ n4365 ^ n1030 ;
  assign n4357 = ( n524 & n3055 ) | ( n524 & ~n4170 ) | ( n3055 & ~n4170 ) ;
  assign n4358 = n2899 ^ n1313 ^ n350 ;
  assign n4359 = ( ~n934 & n1595 ) | ( ~n934 & n3535 ) | ( n1595 & n3535 ) ;
  assign n4360 = n4253 ^ n1554 ^ n1469 ;
  assign n4361 = n3044 ^ n1113 ^ n778 ;
  assign n4362 = ( n4359 & n4360 ) | ( n4359 & ~n4361 ) | ( n4360 & ~n4361 ) ;
  assign n4363 = ( ~n4357 & n4358 ) | ( ~n4357 & n4362 ) | ( n4358 & n4362 ) ;
  assign n4368 = n4367 ^ n4363 ^ n2515 ;
  assign n4375 = n4374 ^ n4368 ^ n1755 ;
  assign n4389 = n4388 ^ n4375 ^ n1491 ;
  assign n4390 = n4389 ^ n3703 ^ n1714 ;
  assign n4391 = n3587 ^ n2490 ^ n2052 ;
  assign n4392 = ( ~n2872 & n3103 ) | ( ~n2872 & n3554 ) | ( n3103 & n3554 ) ;
  assign n4393 = ( n809 & n4060 ) | ( n809 & n4392 ) | ( n4060 & n4392 ) ;
  assign n4394 = n4393 ^ n3135 ^ n1750 ;
  assign n4395 = ( n2620 & n4391 ) | ( n2620 & ~n4394 ) | ( n4391 & ~n4394 ) ;
  assign n4399 = n1350 ^ n1060 ^ n181 ;
  assign n4396 = n1334 ^ n1008 ^ x9 ;
  assign n4397 = n3025 ^ n2676 ^ n1260 ;
  assign n4398 = ( n3198 & n4396 ) | ( n3198 & ~n4397 ) | ( n4396 & ~n4397 ) ;
  assign n4400 = n4399 ^ n4398 ^ n1921 ;
  assign n4401 = n3833 ^ n2793 ^ n533 ;
  assign n4402 = n3999 ^ n2453 ^ x109 ;
  assign n4403 = ( n213 & ~n4232 ) | ( n213 & n4402 ) | ( ~n4232 & n4402 ) ;
  assign n4404 = ( ~n2920 & n4401 ) | ( ~n2920 & n4403 ) | ( n4401 & n4403 ) ;
  assign n4405 = n1549 ^ n555 ^ n324 ;
  assign n4424 = n4024 ^ n262 ^ n215 ;
  assign n4419 = ( ~n189 & n286 ) | ( ~n189 & n4041 ) | ( n286 & n4041 ) ;
  assign n4420 = ( n4045 & n4327 ) | ( n4045 & n4419 ) | ( n4327 & n4419 ) ;
  assign n4417 = ( n320 & n1351 ) | ( n320 & ~n1478 ) | ( n1351 & ~n1478 ) ;
  assign n4418 = n4417 ^ n3837 ^ n2088 ;
  assign n4421 = n4420 ^ n4418 ^ n2202 ;
  assign n4422 = ( ~n2410 & n2541 ) | ( ~n2410 & n4421 ) | ( n2541 & n4421 ) ;
  assign n4423 = ( n203 & ~n510 ) | ( n203 & n4422 ) | ( ~n510 & n4422 ) ;
  assign n4425 = n4424 ^ n4423 ^ n1954 ;
  assign n4416 = ( n1592 & n2359 ) | ( n1592 & ~n2404 ) | ( n2359 & ~n2404 ) ;
  assign n4413 = ( n1660 & n2777 ) | ( n1660 & n3511 ) | ( n2777 & n3511 ) ;
  assign n4411 = ( ~x78 & n1660 ) | ( ~x78 & n3841 ) | ( n1660 & n3841 ) ;
  assign n4407 = n676 ^ n653 ^ x88 ;
  assign n4408 = ( n526 & n1539 ) | ( n526 & n4407 ) | ( n1539 & n4407 ) ;
  assign n4409 = ( n1214 & n2682 ) | ( n1214 & ~n4408 ) | ( n2682 & ~n4408 ) ;
  assign n4410 = n4409 ^ n3122 ^ n1923 ;
  assign n4412 = n4411 ^ n4410 ^ n2386 ;
  assign n4406 = n3331 ^ n2225 ^ n312 ;
  assign n4414 = n4413 ^ n4412 ^ n4406 ;
  assign n4415 = n4414 ^ n4377 ^ n2118 ;
  assign n4426 = n4425 ^ n4416 ^ n4415 ;
  assign n4427 = ( n1191 & ~n4405 ) | ( n1191 & n4426 ) | ( ~n4405 & n4426 ) ;
  assign n4497 = ( n757 & ~n1285 ) | ( n757 & n2852 ) | ( ~n1285 & n2852 ) ;
  assign n4500 = ( ~n1159 & n2569 ) | ( ~n1159 & n3668 ) | ( n2569 & n3668 ) ;
  assign n4498 = ( n481 & ~n2342 ) | ( n481 & n2644 ) | ( ~n2342 & n2644 ) ;
  assign n4499 = ( n407 & n715 ) | ( n407 & ~n4498 ) | ( n715 & ~n4498 ) ;
  assign n4501 = n4500 ^ n4499 ^ n3833 ;
  assign n4502 = ( n466 & n2248 ) | ( n466 & n2518 ) | ( n2248 & n2518 ) ;
  assign n4503 = ( n2952 & ~n4501 ) | ( n2952 & n4502 ) | ( ~n4501 & n4502 ) ;
  assign n4504 = ( n1654 & ~n4497 ) | ( n1654 & n4503 ) | ( ~n4497 & n4503 ) ;
  assign n4491 = n942 ^ n684 ^ n623 ;
  assign n4492 = n4491 ^ n3168 ^ n396 ;
  assign n4493 = ( ~n1371 & n1445 ) | ( ~n1371 & n3455 ) | ( n1445 & n3455 ) ;
  assign n4494 = n3260 ^ n3003 ^ n918 ;
  assign n4495 = ( n4492 & n4493 ) | ( n4492 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4490 = ( n604 & n2056 ) | ( n604 & n3601 ) | ( n2056 & n3601 ) ;
  assign n4487 = ( x37 & ~n726 ) | ( x37 & n848 ) | ( ~n726 & n848 ) ;
  assign n4488 = n4487 ^ n3739 ^ n2418 ;
  assign n4485 = ( n610 & n935 ) | ( n610 & ~n3206 ) | ( n935 & ~n3206 ) ;
  assign n4486 = n4485 ^ n1833 ^ n878 ;
  assign n4482 = n2911 ^ n1610 ^ n1076 ;
  assign n4483 = n4482 ^ x39 ^ x15 ;
  assign n4480 = n2666 ^ n1940 ^ n1147 ;
  assign n4481 = ( n1785 & ~n3111 ) | ( n1785 & n4480 ) | ( ~n3111 & n4480 ) ;
  assign n4476 = ( n618 & n638 ) | ( n618 & n1198 ) | ( n638 & n1198 ) ;
  assign n4477 = n4476 ^ n1828 ^ n1408 ;
  assign n4478 = ( n576 & ~n2308 ) | ( n576 & n2952 ) | ( ~n2308 & n2952 ) ;
  assign n4479 = ( n139 & n4477 ) | ( n139 & n4478 ) | ( n4477 & n4478 ) ;
  assign n4484 = n4483 ^ n4481 ^ n4479 ;
  assign n4489 = n4488 ^ n4486 ^ n4484 ;
  assign n4496 = n4495 ^ n4490 ^ n4489 ;
  assign n4428 = ( n131 & n741 ) | ( n131 & ~n3174 ) | ( n741 & ~n3174 ) ;
  assign n4429 = ( n1237 & ~n3315 ) | ( n1237 & n3495 ) | ( ~n3315 & n3495 ) ;
  assign n4430 = n4429 ^ n4109 ^ n2410 ;
  assign n4431 = n3101 ^ n1258 ^ n569 ;
  assign n4432 = ( n3900 & n4430 ) | ( n3900 & n4431 ) | ( n4430 & n4431 ) ;
  assign n4433 = n4432 ^ n1447 ^ n181 ;
  assign n4472 = n2067 ^ n2012 ^ n146 ;
  assign n4466 = n2752 ^ n858 ^ n684 ;
  assign n4467 = n3540 ^ n1835 ^ n519 ;
  assign n4468 = ( ~n1611 & n4466 ) | ( ~n1611 & n4467 ) | ( n4466 & n4467 ) ;
  assign n4469 = ( n621 & ~n881 ) | ( n621 & n1181 ) | ( ~n881 & n1181 ) ;
  assign n4470 = n4469 ^ n3190 ^ n1775 ;
  assign n4471 = ( n323 & n4468 ) | ( n323 & n4470 ) | ( n4468 & n4470 ) ;
  assign n4473 = n4472 ^ n4471 ^ n2722 ;
  assign n4462 = ( n2207 & ~n3449 ) | ( n2207 & n3874 ) | ( ~n3449 & n3874 ) ;
  assign n4463 = n4462 ^ n3574 ^ n2036 ;
  assign n4459 = n2346 ^ n1810 ^ n1670 ;
  assign n4460 = ( n827 & n3304 ) | ( n827 & n4459 ) | ( n3304 & n4459 ) ;
  assign n4461 = n4460 ^ n2876 ^ n1416 ;
  assign n4464 = n4463 ^ n4461 ^ n3840 ;
  assign n4465 = n4464 ^ n4071 ^ n4026 ;
  assign n4434 = ( n1940 & ~n2138 ) | ( n1940 & n4247 ) | ( ~n2138 & n4247 ) ;
  assign n4435 = ( ~x47 & n2917 ) | ( ~x47 & n4434 ) | ( n2917 & n4434 ) ;
  assign n4436 = n2792 ^ n2473 ^ n2255 ;
  assign n4437 = ( ~n268 & n2859 ) | ( ~n268 & n4225 ) | ( n2859 & n4225 ) ;
  assign n4438 = n4437 ^ n1365 ^ x87 ;
  assign n4439 = ( n3790 & n4436 ) | ( n3790 & n4438 ) | ( n4436 & n4438 ) ;
  assign n4440 = n4439 ^ n3900 ^ n2663 ;
  assign n4441 = ( n848 & n1691 ) | ( n848 & ~n4440 ) | ( n1691 & ~n4440 ) ;
  assign n4449 = ( ~n1324 & n1469 ) | ( ~n1324 & n2209 ) | ( n1469 & n2209 ) ;
  assign n4450 = ( ~n2663 & n2861 ) | ( ~n2663 & n3395 ) | ( n2861 & n3395 ) ;
  assign n4453 = n676 ^ n516 ^ x121 ;
  assign n4451 = n2693 ^ n2283 ^ n962 ;
  assign n4452 = ( n2000 & ~n2505 ) | ( n2000 & n4451 ) | ( ~n2505 & n4451 ) ;
  assign n4454 = n4453 ^ n4452 ^ n1113 ;
  assign n4455 = ( n2220 & ~n3640 ) | ( n2220 & n4454 ) | ( ~n3640 & n4454 ) ;
  assign n4456 = ( n4449 & n4450 ) | ( n4449 & n4455 ) | ( n4450 & n4455 ) ;
  assign n4447 = n3433 ^ n2619 ^ x40 ;
  assign n4448 = ( n129 & n3362 ) | ( n129 & n4447 ) | ( n3362 & n4447 ) ;
  assign n4444 = n627 ^ n301 ^ x50 ;
  assign n4445 = n4444 ^ n1871 ^ n1661 ;
  assign n4442 = ( n447 & n745 ) | ( n447 & n1093 ) | ( n745 & n1093 ) ;
  assign n4443 = ( ~n2409 & n2647 ) | ( ~n2409 & n4442 ) | ( n2647 & n4442 ) ;
  assign n4446 = n4445 ^ n4443 ^ n2356 ;
  assign n4457 = n4456 ^ n4448 ^ n4446 ;
  assign n4458 = ( ~n4435 & n4441 ) | ( ~n4435 & n4457 ) | ( n4441 & n4457 ) ;
  assign n4474 = n4473 ^ n4465 ^ n4458 ;
  assign n4475 = ( n4428 & n4433 ) | ( n4428 & ~n4474 ) | ( n4433 & ~n4474 ) ;
  assign n4505 = n4504 ^ n4496 ^ n4475 ;
  assign n4522 = n3875 ^ n2485 ^ n1605 ;
  assign n4515 = ( n1405 & ~n1946 ) | ( n1405 & n4062 ) | ( ~n1946 & n4062 ) ;
  assign n4516 = n2644 ^ n944 ^ n805 ;
  assign n4517 = ( n219 & ~n928 ) | ( n219 & n4516 ) | ( ~n928 & n4516 ) ;
  assign n4518 = ( n1395 & n3162 ) | ( n1395 & ~n4517 ) | ( n3162 & ~n4517 ) ;
  assign n4519 = n4518 ^ n395 ^ x98 ;
  assign n4520 = ( n3779 & n4515 ) | ( n3779 & ~n4519 ) | ( n4515 & ~n4519 ) ;
  assign n4511 = n1868 ^ n907 ^ n454 ;
  assign n4512 = ( ~x77 & n1248 ) | ( ~x77 & n4511 ) | ( n1248 & n4511 ) ;
  assign n4513 = ( n3020 & n4122 ) | ( n3020 & ~n4512 ) | ( n4122 & ~n4512 ) ;
  assign n4510 = ( ~x53 & n566 ) | ( ~x53 & n1902 ) | ( n566 & n1902 ) ;
  assign n4514 = n4513 ^ n4510 ^ n2210 ;
  assign n4521 = n4520 ^ n4514 ^ n1380 ;
  assign n4506 = n2762 ^ n1351 ^ n473 ;
  assign n4507 = n4506 ^ n2182 ^ n1123 ;
  assign n4508 = ( ~n1973 & n2252 ) | ( ~n1973 & n4507 ) | ( n2252 & n4507 ) ;
  assign n4509 = n4508 ^ n4264 ^ n4247 ;
  assign n4523 = n4522 ^ n4521 ^ n4509 ;
  assign n4526 = ( ~n331 & n3220 ) | ( ~n331 & n4444 ) | ( n3220 & n4444 ) ;
  assign n4525 = n3836 ^ n2056 ^ n471 ;
  assign n4527 = n4526 ^ n4525 ^ n4113 ;
  assign n4524 = ( ~n1087 & n3746 ) | ( ~n1087 & n4406 ) | ( n3746 & n4406 ) ;
  assign n4528 = n4527 ^ n4524 ^ n635 ;
  assign n4531 = ( n1121 & ~n2335 ) | ( n1121 & n3106 ) | ( ~n2335 & n3106 ) ;
  assign n4530 = n2502 ^ n909 ^ x56 ;
  assign n4529 = n3253 ^ n1115 ^ n134 ;
  assign n4532 = n4531 ^ n4530 ^ n4529 ;
  assign n4533 = ( ~n921 & n1483 ) | ( ~n921 & n2175 ) | ( n1483 & n2175 ) ;
  assign n4534 = n4533 ^ n3846 ^ n2388 ;
  assign n4535 = n4205 ^ n1492 ^ n186 ;
  assign n4536 = n2772 ^ n1840 ^ n650 ;
  assign n4537 = n395 ^ n359 ^ n315 ;
  assign n4538 = n4537 ^ n2449 ^ n1808 ;
  assign n4539 = ( n566 & ~n724 ) | ( n566 & n4538 ) | ( ~n724 & n4538 ) ;
  assign n4540 = ( n730 & n3087 ) | ( n730 & n4539 ) | ( n3087 & n4539 ) ;
  assign n4541 = ( n318 & n4536 ) | ( n318 & n4540 ) | ( n4536 & n4540 ) ;
  assign n4542 = ( ~n144 & n1381 ) | ( ~n144 & n4541 ) | ( n1381 & n4541 ) ;
  assign n4543 = n2676 ^ n1427 ^ n785 ;
  assign n4544 = ( n685 & n1380 ) | ( n685 & n2131 ) | ( n1380 & n2131 ) ;
  assign n4545 = ( n267 & n3760 ) | ( n267 & ~n4544 ) | ( n3760 & ~n4544 ) ;
  assign n4546 = ( n802 & n2982 ) | ( n802 & n4545 ) | ( n2982 & n4545 ) ;
  assign n4547 = ( n4542 & n4543 ) | ( n4542 & ~n4546 ) | ( n4543 & ~n4546 ) ;
  assign n4559 = ( n430 & n2684 ) | ( n430 & ~n3527 ) | ( n2684 & ~n3527 ) ;
  assign n4556 = n3327 ^ n1959 ^ n245 ;
  assign n4554 = ( n303 & n397 ) | ( n303 & n4396 ) | ( n397 & n4396 ) ;
  assign n4555 = ( n1591 & ~n4284 ) | ( n1591 & n4554 ) | ( ~n4284 & n4554 ) ;
  assign n4557 = n4556 ^ n4555 ^ n1302 ;
  assign n4553 = n3130 ^ n1669 ^ n1540 ;
  assign n4558 = n4557 ^ n4553 ^ n3914 ;
  assign n4551 = n3879 ^ n2285 ^ n2123 ;
  assign n4549 = ( n1306 & ~n1457 ) | ( n1306 & n3934 ) | ( ~n1457 & n3934 ) ;
  assign n4548 = ( ~x74 & n912 ) | ( ~x74 & n3542 ) | ( n912 & n3542 ) ;
  assign n4550 = n4549 ^ n4548 ^ n533 ;
  assign n4552 = n4551 ^ n4550 ^ n4126 ;
  assign n4560 = n4559 ^ n4558 ^ n4552 ;
  assign n4571 = ( ~x51 & n541 ) | ( ~x51 & n577 ) | ( n541 & n577 ) ;
  assign n4572 = n4571 ^ n547 ^ n522 ;
  assign n4573 = ( n333 & n2111 ) | ( n333 & n4572 ) | ( n2111 & n4572 ) ;
  assign n4561 = ( x31 & n322 ) | ( x31 & n1708 ) | ( n322 & n1708 ) ;
  assign n4562 = ( x53 & ~n963 ) | ( x53 & n1186 ) | ( ~n963 & n1186 ) ;
  assign n4568 = n1801 ^ n1344 ^ n849 ;
  assign n4565 = n3292 ^ n2676 ^ n2639 ;
  assign n4566 = n2779 ^ n1106 ^ x24 ;
  assign n4567 = ( n1644 & n4565 ) | ( n1644 & ~n4566 ) | ( n4565 & ~n4566 ) ;
  assign n4563 = ( n427 & n792 ) | ( n427 & ~n4080 ) | ( n792 & ~n4080 ) ;
  assign n4564 = ( n3691 & n4152 ) | ( n3691 & n4563 ) | ( n4152 & n4563 ) ;
  assign n4569 = n4568 ^ n4567 ^ n4564 ;
  assign n4570 = ( n4561 & n4562 ) | ( n4561 & ~n4569 ) | ( n4562 & ~n4569 ) ;
  assign n4574 = n4573 ^ n4570 ^ n1945 ;
  assign n4575 = ( n2506 & ~n3068 ) | ( n2506 & n4574 ) | ( ~n3068 & n4574 ) ;
  assign n4576 = n2694 ^ n1208 ^ n1177 ;
  assign n4577 = n1542 ^ n1346 ^ n862 ;
  assign n4578 = ( n2634 & n3103 ) | ( n2634 & ~n4577 ) | ( n3103 & ~n4577 ) ;
  assign n4579 = ( n789 & n1263 ) | ( n789 & ~n4328 ) | ( n1263 & ~n4328 ) ;
  assign n4580 = n4579 ^ n3320 ^ n2427 ;
  assign n4581 = ( n4576 & ~n4578 ) | ( n4576 & n4580 ) | ( ~n4578 & n4580 ) ;
  assign n4600 = ( n230 & n1546 ) | ( n230 & n1985 ) | ( n1546 & n1985 ) ;
  assign n4596 = n2141 ^ n1667 ^ n665 ;
  assign n4597 = n4596 ^ n3216 ^ n1520 ;
  assign n4593 = ( n793 & n970 ) | ( n793 & ~n3729 ) | ( n970 & ~n3729 ) ;
  assign n4594 = ( n558 & n2246 ) | ( n558 & n2434 ) | ( n2246 & n2434 ) ;
  assign n4595 = ( ~n954 & n4593 ) | ( ~n954 & n4594 ) | ( n4593 & n4594 ) ;
  assign n4598 = n4597 ^ n4595 ^ n3456 ;
  assign n4591 = ( n809 & n1276 ) | ( n809 & ~n4572 ) | ( n1276 & ~n4572 ) ;
  assign n4590 = ( n2169 & n3169 ) | ( n2169 & ~n3387 ) | ( n3169 & ~n3387 ) ;
  assign n4592 = n4591 ^ n4590 ^ n3890 ;
  assign n4587 = ( ~n1040 & n2087 ) | ( ~n1040 & n2404 ) | ( n2087 & n2404 ) ;
  assign n4588 = ( x101 & ~n1202 ) | ( x101 & n4587 ) | ( ~n1202 & n4587 ) ;
  assign n4583 = ( n324 & n754 ) | ( n324 & n2627 ) | ( n754 & n2627 ) ;
  assign n4584 = n4583 ^ n3763 ^ n2209 ;
  assign n4582 = n2995 ^ n2521 ^ n759 ;
  assign n4585 = n4584 ^ n4582 ^ n2929 ;
  assign n4586 = ( n3355 & n4095 ) | ( n3355 & ~n4585 ) | ( n4095 & ~n4585 ) ;
  assign n4589 = n4588 ^ n4586 ^ n1855 ;
  assign n4599 = n4598 ^ n4592 ^ n4589 ;
  assign n4601 = n4600 ^ n4599 ^ n888 ;
  assign n4627 = n3965 ^ n1124 ^ n437 ;
  assign n4628 = n4627 ^ n1842 ^ n697 ;
  assign n4629 = n4628 ^ n3405 ^ n3384 ;
  assign n4630 = n1301 ^ n223 ^ x95 ;
  assign n4631 = ( ~n2610 & n4629 ) | ( ~n2610 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4624 = ( n158 & n1858 ) | ( n158 & n2639 ) | ( n1858 & n2639 ) ;
  assign n4622 = n3618 ^ n2923 ^ n1609 ;
  assign n4621 = n4334 ^ n3807 ^ n3167 ;
  assign n4623 = n4622 ^ n4621 ^ n860 ;
  assign n4625 = n4624 ^ n4623 ^ x8 ;
  assign n4626 = n4625 ^ n4622 ^ n393 ;
  assign n4602 = n2617 ^ n548 ^ x38 ;
  assign n4608 = ( n239 & n3309 ) | ( n239 & ~n3960 ) | ( n3309 & ~n3960 ) ;
  assign n4604 = n1526 ^ n892 ^ n704 ;
  assign n4605 = n4604 ^ n4113 ^ n1248 ;
  assign n4603 = n3588 ^ n3348 ^ n3024 ;
  assign n4606 = n4605 ^ n4603 ^ n844 ;
  assign n4607 = n4606 ^ n1434 ^ n295 ;
  assign n4609 = n4608 ^ n4607 ^ n1312 ;
  assign n4618 = ( n852 & n2214 ) | ( n852 & n2258 ) | ( n2214 & n2258 ) ;
  assign n4611 = ( x86 & n1599 ) | ( x86 & n1853 ) | ( n1599 & n1853 ) ;
  assign n4612 = n4611 ^ n1707 ^ n841 ;
  assign n4613 = n3362 ^ n2947 ^ n1569 ;
  assign n4614 = n4613 ^ n3189 ^ n2087 ;
  assign n4615 = ( ~x73 & n510 ) | ( ~x73 & n1058 ) | ( n510 & n1058 ) ;
  assign n4616 = n4615 ^ n2926 ^ n1699 ;
  assign n4617 = ( n4612 & ~n4614 ) | ( n4612 & n4616 ) | ( ~n4614 & n4616 ) ;
  assign n4610 = ( x126 & ~n2408 ) | ( x126 & n2776 ) | ( ~n2408 & n2776 ) ;
  assign n4619 = n4618 ^ n4617 ^ n4610 ;
  assign n4620 = ( n4602 & ~n4609 ) | ( n4602 & n4619 ) | ( ~n4609 & n4619 ) ;
  assign n4632 = n4631 ^ n4626 ^ n4620 ;
  assign n4638 = n1212 ^ n943 ^ n873 ;
  assign n4639 = ( n910 & ~n2195 ) | ( n910 & n4638 ) | ( ~n2195 & n4638 ) ;
  assign n4640 = ( n634 & ~n2279 ) | ( n634 & n4639 ) | ( ~n2279 & n4639 ) ;
  assign n4641 = n4640 ^ n1905 ^ n934 ;
  assign n4642 = n4641 ^ n2844 ^ n310 ;
  assign n4634 = n3231 ^ n996 ^ n601 ;
  assign n4635 = n1231 ^ n620 ^ x80 ;
  assign n4636 = ( n4082 & n4634 ) | ( n4082 & ~n4635 ) | ( n4634 & ~n4635 ) ;
  assign n4633 = n4014 ^ n3432 ^ n3044 ;
  assign n4637 = n4636 ^ n4633 ^ n3641 ;
  assign n4643 = n4642 ^ n4637 ^ n2450 ;
  assign n4653 = ( ~n429 & n607 ) | ( ~n429 & n2259 ) | ( n607 & n2259 ) ;
  assign n4651 = ( n883 & n1427 ) | ( n883 & ~n2717 ) | ( n1427 & ~n2717 ) ;
  assign n4652 = n4651 ^ n4573 ^ n1040 ;
  assign n4654 = n4653 ^ n4652 ^ x104 ;
  assign n4650 = n2920 ^ n1945 ^ n538 ;
  assign n4645 = n3406 ^ n3061 ^ n1752 ;
  assign n4644 = n2646 ^ n248 ^ n135 ;
  assign n4646 = n4645 ^ n4644 ^ n869 ;
  assign n4647 = n4646 ^ n3367 ^ n1626 ;
  assign n4648 = n3640 ^ n3085 ^ n2040 ;
  assign n4649 = ( n3596 & n4647 ) | ( n3596 & n4648 ) | ( n4647 & n4648 ) ;
  assign n4655 = n4654 ^ n4650 ^ n4649 ;
  assign n4656 = n4280 ^ n2501 ^ n1101 ;
  assign n4657 = n4656 ^ n3360 ^ n133 ;
  assign n4658 = ( n838 & n1591 ) | ( n838 & n3456 ) | ( n1591 & n3456 ) ;
  assign n4659 = ( n148 & n382 ) | ( n148 & ~n4658 ) | ( n382 & ~n4658 ) ;
  assign n4660 = n4659 ^ n1575 ^ x114 ;
  assign n4661 = n4660 ^ n3676 ^ x55 ;
  assign n4663 = ( ~n904 & n4020 ) | ( ~n904 & n4594 ) | ( n4020 & n4594 ) ;
  assign n4662 = n3588 ^ n2689 ^ x73 ;
  assign n4664 = n4663 ^ n4662 ^ n3779 ;
  assign n4665 = ( n184 & n2177 ) | ( n184 & ~n2433 ) | ( n2177 & ~n2433 ) ;
  assign n4666 = n4665 ^ n2798 ^ n1878 ;
  assign n4667 = ( n792 & ~n3924 ) | ( n792 & n4666 ) | ( ~n3924 & n4666 ) ;
  assign n4668 = ( n4661 & n4664 ) | ( n4661 & n4667 ) | ( n4664 & n4667 ) ;
  assign n4669 = ( ~n560 & n802 ) | ( ~n560 & n2189 ) | ( n802 & n2189 ) ;
  assign n4670 = n4669 ^ n3285 ^ n2167 ;
  assign n4674 = ( ~n165 & n1492 ) | ( ~n165 & n2303 ) | ( n1492 & n2303 ) ;
  assign n4671 = ( ~n414 & n1378 ) | ( ~n414 & n3933 ) | ( n1378 & n3933 ) ;
  assign n4672 = n4671 ^ n2436 ^ n1788 ;
  assign n4673 = ( n1493 & n1965 ) | ( n1493 & n4672 ) | ( n1965 & n4672 ) ;
  assign n4675 = n4674 ^ n4673 ^ n1676 ;
  assign n4676 = ( ~n545 & n2270 ) | ( ~n545 & n4675 ) | ( n2270 & n4675 ) ;
  assign n4677 = ( n355 & ~n4081 ) | ( n355 & n4676 ) | ( ~n4081 & n4676 ) ;
  assign n4678 = n2179 ^ n1043 ^ n940 ;
  assign n4679 = ( n1344 & ~n3613 ) | ( n1344 & n4678 ) | ( ~n3613 & n4678 ) ;
  assign n4680 = n1052 ^ n446 ^ n285 ;
  assign n4681 = ( n393 & n1169 ) | ( n393 & ~n3468 ) | ( n1169 & ~n3468 ) ;
  assign n4682 = ( n410 & n4680 ) | ( n410 & n4681 ) | ( n4680 & n4681 ) ;
  assign n4683 = ( ~n2173 & n4679 ) | ( ~n2173 & n4682 ) | ( n4679 & n4682 ) ;
  assign n4684 = n4683 ^ n3400 ^ n2950 ;
  assign n4685 = ( n4670 & n4677 ) | ( n4670 & ~n4684 ) | ( n4677 & ~n4684 ) ;
  assign n4686 = n1173 ^ n719 ^ n357 ;
  assign n4687 = n4686 ^ n3738 ^ n913 ;
  assign n4688 = ( n138 & n379 ) | ( n138 & ~n4687 ) | ( n379 & ~n4687 ) ;
  assign n4697 = ( ~n1905 & n2161 ) | ( ~n1905 & n4468 ) | ( n2161 & n4468 ) ;
  assign n4689 = ( n896 & n1180 ) | ( n896 & ~n3655 ) | ( n1180 & ~n3655 ) ;
  assign n4690 = n2790 ^ n2718 ^ n1134 ;
  assign n4691 = n4345 ^ n3934 ^ n1321 ;
  assign n4692 = ( ~n613 & n1750 ) | ( ~n613 & n4691 ) | ( n1750 & n4691 ) ;
  assign n4693 = n2886 ^ n647 ^ n230 ;
  assign n4694 = ( n1445 & n2176 ) | ( n1445 & ~n4693 ) | ( n2176 & ~n4693 ) ;
  assign n4695 = ( n4435 & n4692 ) | ( n4435 & ~n4694 ) | ( n4692 & ~n4694 ) ;
  assign n4696 = ( n4689 & n4690 ) | ( n4689 & ~n4695 ) | ( n4690 & ~n4695 ) ;
  assign n4698 = n4697 ^ n4696 ^ n1290 ;
  assign n4711 = ( ~n853 & n2315 ) | ( ~n853 & n2458 ) | ( n2315 & n2458 ) ;
  assign n4712 = ( x22 & n1927 ) | ( x22 & ~n4711 ) | ( n1927 & ~n4711 ) ;
  assign n4702 = n1275 ^ n911 ^ n439 ;
  assign n4703 = ( n1011 & ~n3650 ) | ( n1011 & n4702 ) | ( ~n3650 & n4702 ) ;
  assign n4704 = n3185 ^ n2314 ^ n1497 ;
  assign n4705 = ( ~n251 & n990 ) | ( ~n251 & n1876 ) | ( n990 & n1876 ) ;
  assign n4706 = n4705 ^ n1195 ^ n562 ;
  assign n4707 = ( n1355 & n4704 ) | ( n1355 & ~n4706 ) | ( n4704 & ~n4706 ) ;
  assign n4708 = ( n1215 & n1300 ) | ( n1215 & n4707 ) | ( n1300 & n4707 ) ;
  assign n4709 = ( n965 & n4703 ) | ( n965 & n4708 ) | ( n4703 & n4708 ) ;
  assign n4710 = n4709 ^ n4414 ^ n3434 ;
  assign n4700 = n3463 ^ n1235 ^ n846 ;
  assign n4699 = n3710 ^ n1541 ^ n583 ;
  assign n4701 = n4700 ^ n4699 ^ n4471 ;
  assign n4713 = n4712 ^ n4710 ^ n4701 ;
  assign n4714 = n3070 ^ n2752 ^ n395 ;
  assign n4715 = ( n442 & n1355 ) | ( n442 & ~n4714 ) | ( n1355 & ~n4714 ) ;
  assign n4717 = n4107 ^ n945 ^ n283 ;
  assign n4716 = n3267 ^ n2362 ^ n1031 ;
  assign n4718 = n4717 ^ n4716 ^ n3071 ;
  assign n4719 = ( ~n4713 & n4715 ) | ( ~n4713 & n4718 ) | ( n4715 & n4718 ) ;
  assign n4727 = ( ~n369 & n2182 ) | ( ~n369 & n2298 ) | ( n2182 & n2298 ) ;
  assign n4723 = n2107 ^ n1946 ^ n1402 ;
  assign n4721 = n2574 ^ n1851 ^ n1534 ;
  assign n4722 = ( n894 & ~n902 ) | ( n894 & n4721 ) | ( ~n902 & n4721 ) ;
  assign n4724 = n4723 ^ n4722 ^ n3973 ;
  assign n4725 = n4724 ^ n4325 ^ n1067 ;
  assign n4726 = n4725 ^ n4450 ^ n4256 ;
  assign n4720 = n2327 ^ n739 ^ x119 ;
  assign n4728 = n4727 ^ n4726 ^ n4720 ;
  assign n4729 = ( ~n151 & n530 ) | ( ~n151 & n895 ) | ( n530 & n895 ) ;
  assign n4730 = n4729 ^ n3877 ^ n160 ;
  assign n4731 = n4088 ^ n3836 ^ n3065 ;
  assign n4732 = ( n601 & n946 ) | ( n601 & ~n4731 ) | ( n946 & ~n4731 ) ;
  assign n4733 = n2929 ^ n1968 ^ n137 ;
  assign n4734 = n4733 ^ n2445 ^ n300 ;
  assign n4735 = ( n2010 & n4732 ) | ( n2010 & ~n4734 ) | ( n4732 & ~n4734 ) ;
  assign n4743 = n1851 ^ n582 ^ n168 ;
  assign n4744 = ( n1580 & ~n2320 ) | ( n1580 & n4743 ) | ( ~n2320 & n4743 ) ;
  assign n4745 = n4744 ^ n4233 ^ n1118 ;
  assign n4746 = ( ~n1863 & n4104 ) | ( ~n1863 & n4745 ) | ( n4104 & n4745 ) ;
  assign n4747 = n4746 ^ n3107 ^ n314 ;
  assign n4748 = ( n1728 & n3124 ) | ( n1728 & n4747 ) | ( n3124 & n4747 ) ;
  assign n4749 = ( ~n2431 & n3856 ) | ( ~n2431 & n4748 ) | ( n3856 & n4748 ) ;
  assign n4750 = n3876 ^ n2582 ^ n699 ;
  assign n4751 = ( ~n452 & n3087 ) | ( ~n452 & n4750 ) | ( n3087 & n4750 ) ;
  assign n4752 = n4751 ^ n1941 ^ n1119 ;
  assign n4753 = ( n1775 & ~n4749 ) | ( n1775 & n4752 ) | ( ~n4749 & n4752 ) ;
  assign n4742 = ( n333 & n382 ) | ( n333 & n4429 ) | ( n382 & n4429 ) ;
  assign n4740 = ( n1144 & ~n2849 ) | ( n1144 & n3576 ) | ( ~n2849 & n3576 ) ;
  assign n4738 = ( ~x100 & x116 ) | ( ~x100 & n560 ) | ( x116 & n560 ) ;
  assign n4737 = ( n436 & n701 ) | ( n436 & ~n2501 ) | ( n701 & ~n2501 ) ;
  assign n4736 = n3548 ^ n2142 ^ n895 ;
  assign n4739 = n4738 ^ n4737 ^ n4736 ;
  assign n4741 = n4740 ^ n4739 ^ n409 ;
  assign n4754 = n4753 ^ n4742 ^ n4741 ;
  assign n4773 = ( n171 & n435 ) | ( n171 & n1831 ) | ( n435 & n1831 ) ;
  assign n4769 = ( n146 & n270 ) | ( n146 & ~n522 ) | ( n270 & ~n522 ) ;
  assign n4770 = n4769 ^ n1939 ^ n195 ;
  assign n4771 = n4770 ^ n3271 ^ n202 ;
  assign n4772 = ( n741 & ~n4723 ) | ( n741 & n4771 ) | ( ~n4723 & n4771 ) ;
  assign n4774 = n4773 ^ n4772 ^ n1280 ;
  assign n4775 = ( n449 & n3477 ) | ( n449 & n4774 ) | ( n3477 & n4774 ) ;
  assign n4756 = ( n1594 & n2278 ) | ( n1594 & ~n2454 ) | ( n2278 & ~n2454 ) ;
  assign n4757 = ( n1418 & ~n2928 ) | ( n1418 & n3205 ) | ( ~n2928 & n3205 ) ;
  assign n4758 = ( n2127 & n3304 ) | ( n2127 & ~n3499 ) | ( n3304 & ~n3499 ) ;
  assign n4762 = ( n1459 & n1534 ) | ( n1459 & ~n2944 ) | ( n1534 & ~n2944 ) ;
  assign n4759 = ( ~n470 & n1328 ) | ( ~n470 & n1605 ) | ( n1328 & n1605 ) ;
  assign n4760 = ( n834 & n2427 ) | ( n834 & n3831 ) | ( n2427 & n3831 ) ;
  assign n4761 = ( ~n3147 & n4759 ) | ( ~n3147 & n4760 ) | ( n4759 & n4760 ) ;
  assign n4763 = n4762 ^ n4761 ^ n2337 ;
  assign n4764 = ( n851 & n1350 ) | ( n851 & ~n1512 ) | ( n1350 & ~n1512 ) ;
  assign n4765 = n4764 ^ n4263 ^ n594 ;
  assign n4766 = ( ~n2461 & n4763 ) | ( ~n2461 & n4765 ) | ( n4763 & n4765 ) ;
  assign n4767 = ( n4757 & ~n4758 ) | ( n4757 & n4766 ) | ( ~n4758 & n4766 ) ;
  assign n4768 = ( n1783 & ~n4756 ) | ( n1783 & n4767 ) | ( ~n4756 & n4767 ) ;
  assign n4755 = ( n285 & ~n2865 ) | ( n285 & n3724 ) | ( ~n2865 & n3724 ) ;
  assign n4776 = n4775 ^ n4768 ^ n4755 ;
  assign n4777 = n1263 ^ n863 ^ n271 ;
  assign n4778 = ( n2032 & n2553 ) | ( n2032 & n4777 ) | ( n2553 & n4777 ) ;
  assign n4779 = n4439 ^ n2939 ^ n1002 ;
  assign n4780 = n3930 ^ n2985 ^ n1126 ;
  assign n4781 = ( ~n1376 & n4779 ) | ( ~n1376 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4782 = ( n3106 & ~n4778 ) | ( n3106 & n4781 ) | ( ~n4778 & n4781 ) ;
  assign n4783 = ( n850 & n1836 ) | ( n850 & n3139 ) | ( n1836 & n3139 ) ;
  assign n4784 = n4783 ^ n4525 ^ n3327 ;
  assign n4785 = ( ~n417 & n3929 ) | ( ~n417 & n4784 ) | ( n3929 & n4784 ) ;
  assign n4786 = ( ~n4392 & n4596 ) | ( ~n4392 & n4785 ) | ( n4596 & n4785 ) ;
  assign n4787 = ( n1683 & ~n4162 ) | ( n1683 & n4786 ) | ( ~n4162 & n4786 ) ;
  assign n4788 = ( n1069 & ~n4782 ) | ( n1069 & n4787 ) | ( ~n4782 & n4787 ) ;
  assign n4790 = ( ~n634 & n1090 ) | ( ~n634 & n2762 ) | ( n1090 & n2762 ) ;
  assign n4789 = n3137 ^ n1985 ^ x4 ;
  assign n4791 = n4790 ^ n4789 ^ x79 ;
  assign n4792 = n4791 ^ n3554 ^ n1218 ;
  assign n4793 = ( n1283 & ~n1341 ) | ( n1283 & n1354 ) | ( ~n1341 & n1354 ) ;
  assign n4794 = n4793 ^ n2306 ^ n733 ;
  assign n4795 = n4794 ^ n3479 ^ n2488 ;
  assign n4796 = n3085 ^ n2077 ^ n1680 ;
  assign n4797 = ( n151 & n1243 ) | ( n151 & n2090 ) | ( n1243 & n2090 ) ;
  assign n4798 = ( n767 & n1921 ) | ( n767 & n4797 ) | ( n1921 & n4797 ) ;
  assign n4799 = n4798 ^ n1138 ^ n343 ;
  assign n4800 = ( ~n3735 & n4796 ) | ( ~n3735 & n4799 ) | ( n4796 & n4799 ) ;
  assign n4801 = ( ~n1218 & n4795 ) | ( ~n1218 & n4800 ) | ( n4795 & n4800 ) ;
  assign n4802 = n4801 ^ n2930 ^ n170 ;
  assign n4803 = ( n580 & n897 ) | ( n580 & ~n3731 ) | ( n897 & ~n3731 ) ;
  assign n4804 = ( n639 & n2215 ) | ( n639 & n3016 ) | ( n2215 & n3016 ) ;
  assign n4805 = n4804 ^ n2281 ^ n1215 ;
  assign n4806 = ( n2495 & n4803 ) | ( n2495 & n4805 ) | ( n4803 & n4805 ) ;
  assign n4807 = n4806 ^ n4149 ^ n1067 ;
  assign n4808 = ( ~x74 & n2286 ) | ( ~x74 & n4482 ) | ( n2286 & n4482 ) ;
  assign n4809 = n1902 ^ n1579 ^ n1362 ;
  assign n4810 = ( n641 & ~n2467 ) | ( n641 & n4809 ) | ( ~n2467 & n4809 ) ;
  assign n4811 = n4810 ^ n4159 ^ n3692 ;
  assign n4812 = ( n992 & ~n2177 ) | ( n992 & n3896 ) | ( ~n2177 & n3896 ) ;
  assign n4813 = ( ~n336 & n4811 ) | ( ~n336 & n4812 ) | ( n4811 & n4812 ) ;
  assign n4814 = ( n720 & n3135 ) | ( n720 & n4813 ) | ( n3135 & n4813 ) ;
  assign n4815 = ( n2094 & n4808 ) | ( n2094 & n4814 ) | ( n4808 & n4814 ) ;
  assign n4822 = n1231 ^ n992 ^ x104 ;
  assign n4823 = n4822 ^ n2996 ^ x123 ;
  assign n4824 = n4142 ^ n3212 ^ n2349 ;
  assign n4825 = ( n2719 & n4823 ) | ( n2719 & ~n4824 ) | ( n4823 & ~n4824 ) ;
  assign n4818 = ( n249 & ~n1155 ) | ( n249 & n1486 ) | ( ~n1155 & n1486 ) ;
  assign n4816 = ( n1318 & ~n2244 ) | ( n1318 & n4123 ) | ( ~n2244 & n4123 ) ;
  assign n4817 = n4816 ^ n3824 ^ n980 ;
  assign n4819 = n4818 ^ n4817 ^ n3371 ;
  assign n4820 = n4819 ^ n3828 ^ n531 ;
  assign n4821 = n4820 ^ n3282 ^ n2163 ;
  assign n4826 = n4825 ^ n4821 ^ n2815 ;
  assign n4827 = n2938 ^ n1640 ^ n628 ;
  assign n4828 = n4827 ^ n4556 ^ n954 ;
  assign n4829 = ( n2525 & ~n4257 ) | ( n2525 & n4828 ) | ( ~n4257 & n4828 ) ;
  assign n4830 = ( ~n3986 & n4335 ) | ( ~n3986 & n4829 ) | ( n4335 & n4829 ) ;
  assign n4831 = ( ~n189 & n533 ) | ( ~n189 & n944 ) | ( n533 & n944 ) ;
  assign n4832 = n4831 ^ n4371 ^ n1759 ;
  assign n4833 = n4832 ^ n3010 ^ n707 ;
  assign n4834 = ( n897 & n4705 ) | ( n897 & ~n4756 ) | ( n4705 & ~n4756 ) ;
  assign n4835 = n4834 ^ n1200 ^ n821 ;
  assign n4836 = ( ~n1736 & n4833 ) | ( ~n1736 & n4835 ) | ( n4833 & n4835 ) ;
  assign n4837 = n3811 ^ n1426 ^ n295 ;
  assign n4838 = n4837 ^ n4003 ^ n1046 ;
  assign n4839 = ( n450 & ~n1179 ) | ( n450 & n4838 ) | ( ~n1179 & n4838 ) ;
  assign n4842 = ( n682 & n1567 ) | ( n682 & ~n2113 ) | ( n1567 & ~n2113 ) ;
  assign n4840 = ( n369 & n3547 ) | ( n369 & n4151 ) | ( n3547 & n4151 ) ;
  assign n4841 = ( n900 & n4334 ) | ( n900 & n4840 ) | ( n4334 & n4840 ) ;
  assign n4843 = n4842 ^ n4841 ^ n668 ;
  assign n4844 = ( n3565 & n4839 ) | ( n3565 & n4843 ) | ( n4839 & n4843 ) ;
  assign n4853 = ( n859 & ~n4483 ) | ( n859 & n4760 ) | ( ~n4483 & n4760 ) ;
  assign n4852 = n4796 ^ n3893 ^ n647 ;
  assign n4845 = ( n610 & n1427 ) | ( n610 & n1878 ) | ( n1427 & n1878 ) ;
  assign n4846 = ( n354 & ~n2073 ) | ( n354 & n2798 ) | ( ~n2073 & n2798 ) ;
  assign n4847 = n3237 ^ n1327 ^ n1189 ;
  assign n4848 = ( ~n2068 & n3808 ) | ( ~n2068 & n4847 ) | ( n3808 & n4847 ) ;
  assign n4849 = ( n1130 & n3199 ) | ( n1130 & n4848 ) | ( n3199 & n4848 ) ;
  assign n4850 = n4849 ^ n3261 ^ n2861 ;
  assign n4851 = ( ~n4845 & n4846 ) | ( ~n4845 & n4850 ) | ( n4846 & n4850 ) ;
  assign n4854 = n4853 ^ n4852 ^ n4851 ;
  assign n4855 = ( ~n156 & n201 ) | ( ~n156 & n1495 ) | ( n201 & n1495 ) ;
  assign n4856 = n4855 ^ n3733 ^ n2343 ;
  assign n4857 = n4856 ^ n1368 ^ x66 ;
  assign n4863 = ( ~n502 & n1330 ) | ( ~n502 & n1400 ) | ( n1330 & n1400 ) ;
  assign n4862 = n2699 ^ n2020 ^ n1096 ;
  assign n4864 = n4863 ^ n4862 ^ n1055 ;
  assign n4858 = n2183 ^ n1388 ^ x80 ;
  assign n4859 = ( ~n389 & n942 ) | ( ~n389 & n1876 ) | ( n942 & n1876 ) ;
  assign n4860 = ( n1995 & ~n4858 ) | ( n1995 & n4859 ) | ( ~n4858 & n4859 ) ;
  assign n4861 = n4860 ^ n2796 ^ n977 ;
  assign n4865 = n4864 ^ n4861 ^ n2288 ;
  assign n4873 = n1839 ^ n521 ^ n388 ;
  assign n4874 = n4873 ^ n3946 ^ n3095 ;
  assign n4875 = n4874 ^ n2229 ^ x49 ;
  assign n4870 = n2483 ^ n717 ^ n406 ;
  assign n4871 = ( n2207 & n2616 ) | ( n2207 & n4870 ) | ( n2616 & n4870 ) ;
  assign n4868 = n2407 ^ n1414 ^ n782 ;
  assign n4869 = n4868 ^ n1883 ^ n686 ;
  assign n4872 = n4871 ^ n4869 ^ n784 ;
  assign n4866 = ( n328 & ~n1742 ) | ( n328 & n4248 ) | ( ~n1742 & n4248 ) ;
  assign n4867 = n4866 ^ n2384 ^ n2150 ;
  assign n4876 = n4875 ^ n4872 ^ n4867 ;
  assign n4877 = ( n4857 & n4865 ) | ( n4857 & ~n4876 ) | ( n4865 & ~n4876 ) ;
  assign n4878 = n2777 ^ n1585 ^ n869 ;
  assign n4879 = ( n1831 & n2410 ) | ( n1831 & n4878 ) | ( n2410 & n4878 ) ;
  assign n4880 = ( n262 & ~n676 ) | ( n262 & n4879 ) | ( ~n676 & n4879 ) ;
  assign n4886 = n1659 ^ n1515 ^ x79 ;
  assign n4885 = ( ~n1055 & n3999 ) | ( ~n1055 & n4803 ) | ( n3999 & n4803 ) ;
  assign n4884 = n4761 ^ n2307 ^ n1314 ;
  assign n4887 = n4886 ^ n4885 ^ n4884 ;
  assign n4881 = n4285 ^ n3298 ^ n1053 ;
  assign n4882 = ( n1093 & n3784 ) | ( n1093 & ~n4881 ) | ( n3784 & ~n4881 ) ;
  assign n4883 = n4882 ^ n774 ^ n454 ;
  assign n4888 = n4887 ^ n4883 ^ x65 ;
  assign n4889 = n4888 ^ n3925 ^ x90 ;
  assign n4890 = ( ~n350 & n603 ) | ( ~n350 & n1125 ) | ( n603 & n1125 ) ;
  assign n4891 = ( n1202 & n2067 ) | ( n1202 & ~n3905 ) | ( n2067 & ~n3905 ) ;
  assign n4892 = n4891 ^ n4562 ^ n1598 ;
  assign n4893 = n4892 ^ n1955 ^ n1439 ;
  assign n4894 = n2977 ^ n559 ^ n551 ;
  assign n4895 = ( n1048 & ~n2480 ) | ( n1048 & n4894 ) | ( ~n2480 & n4894 ) ;
  assign n4896 = ( n4890 & n4893 ) | ( n4890 & ~n4895 ) | ( n4893 & ~n4895 ) ;
  assign n4897 = n4738 ^ n3347 ^ n2432 ;
  assign n4898 = ( n886 & n4095 ) | ( n886 & n4897 ) | ( n4095 & n4897 ) ;
  assign n4899 = n4898 ^ n2875 ^ n528 ;
  assign n4903 = n3124 ^ n1218 ^ n954 ;
  assign n4904 = n4903 ^ n2080 ^ n303 ;
  assign n4900 = n3895 ^ n1852 ^ n1450 ;
  assign n4901 = n4900 ^ n1599 ^ n169 ;
  assign n4902 = ( n480 & n4704 ) | ( n480 & n4901 ) | ( n4704 & n4901 ) ;
  assign n4905 = n4904 ^ n4902 ^ n1094 ;
  assign n4906 = ( n1732 & n4899 ) | ( n1732 & n4905 ) | ( n4899 & n4905 ) ;
  assign n4907 = ( n661 & n1355 ) | ( n661 & ~n2243 ) | ( n1355 & ~n2243 ) ;
  assign n4908 = ( n728 & n2280 ) | ( n728 & n4907 ) | ( n2280 & n4907 ) ;
  assign n4909 = n3379 ^ n1712 ^ n1683 ;
  assign n4910 = ( n191 & n3135 ) | ( n191 & ~n4310 ) | ( n3135 & ~n4310 ) ;
  assign n4911 = ( n195 & n883 ) | ( n195 & n4910 ) | ( n883 & n4910 ) ;
  assign n4912 = ( n4908 & n4909 ) | ( n4908 & ~n4911 ) | ( n4909 & ~n4911 ) ;
  assign n4922 = n4358 ^ n1696 ^ n632 ;
  assign n4918 = ( n409 & n695 ) | ( n409 & ~n4797 ) | ( n695 & ~n4797 ) ;
  assign n4919 = n4918 ^ n4672 ^ n1994 ;
  assign n4920 = ( n2464 & n3178 ) | ( n2464 & n4919 ) | ( n3178 & n4919 ) ;
  assign n4913 = ( ~x106 & n2305 ) | ( ~x106 & n4362 ) | ( n2305 & n4362 ) ;
  assign n4914 = ( n1235 & ~n1321 ) | ( n1235 & n2065 ) | ( ~n1321 & n2065 ) ;
  assign n4915 = ( n172 & ~n1040 ) | ( n172 & n4914 ) | ( ~n1040 & n4914 ) ;
  assign n4916 = ( n2302 & n3877 ) | ( n2302 & ~n4915 ) | ( n3877 & ~n4915 ) ;
  assign n4917 = ( n2759 & ~n4913 ) | ( n2759 & n4916 ) | ( ~n4913 & n4916 ) ;
  assign n4921 = n4920 ^ n4917 ^ n1812 ;
  assign n4923 = n4922 ^ n4921 ^ n2258 ;
  assign n4932 = n2794 ^ n1310 ^ n159 ;
  assign n4929 = n4743 ^ n2777 ^ n670 ;
  assign n4930 = ( n1749 & n1897 ) | ( n1749 & n4929 ) | ( n1897 & n4929 ) ;
  assign n4931 = ( n1788 & n2726 ) | ( n1788 & n4930 ) | ( n2726 & n4930 ) ;
  assign n4933 = n4932 ^ n4931 ^ n1564 ;
  assign n4927 = ( ~n571 & n679 ) | ( ~n571 & n1077 ) | ( n679 & n1077 ) ;
  assign n4924 = ( n174 & ~n413 ) | ( n174 & n1213 ) | ( ~n413 & n1213 ) ;
  assign n4925 = n4924 ^ n1288 ^ n1122 ;
  assign n4926 = ( n147 & n3939 ) | ( n147 & ~n4925 ) | ( n3939 & ~n4925 ) ;
  assign n4928 = n4927 ^ n4926 ^ n928 ;
  assign n4934 = n4933 ^ n4928 ^ n2330 ;
  assign n4939 = ( n565 & n2340 ) | ( n565 & n3907 ) | ( n2340 & n3907 ) ;
  assign n4935 = ( n1070 & ~n1605 ) | ( n1070 & n1654 ) | ( ~n1605 & n1654 ) ;
  assign n4936 = ( n1682 & n1874 ) | ( n1682 & n2717 ) | ( n1874 & n2717 ) ;
  assign n4937 = ( n1061 & n3964 ) | ( n1061 & ~n4936 ) | ( n3964 & ~n4936 ) ;
  assign n4938 = ( n1715 & n4935 ) | ( n1715 & ~n4937 ) | ( n4935 & ~n4937 ) ;
  assign n4940 = n4939 ^ n4938 ^ n4588 ;
  assign n4941 = n4940 ^ n2022 ^ n1778 ;
  assign n4942 = n2215 ^ n2161 ^ n941 ;
  assign n4943 = n4942 ^ n4026 ^ n1551 ;
  assign n4944 = n4086 ^ n2692 ^ n1464 ;
  assign n4945 = n4944 ^ n3025 ^ n2974 ;
  assign n4946 = ( n4941 & ~n4943 ) | ( n4941 & n4945 ) | ( ~n4943 & n4945 ) ;
  assign n4947 = n4794 ^ n3945 ^ n2956 ;
  assign n4948 = ( ~n253 & n1494 ) | ( ~n253 & n4947 ) | ( n1494 & n4947 ) ;
  assign n4949 = n3614 ^ n2225 ^ n1486 ;
  assign n4950 = ( ~n149 & n177 ) | ( ~n149 & n1104 ) | ( n177 & n1104 ) ;
  assign n4951 = ( ~n3085 & n3978 ) | ( ~n3085 & n4950 ) | ( n3978 & n4950 ) ;
  assign n4952 = ( ~n2792 & n2939 ) | ( ~n2792 & n4951 ) | ( n2939 & n4951 ) ;
  assign n4953 = n3905 ^ n711 ^ n317 ;
  assign n4954 = ( ~n411 & n1184 ) | ( ~n411 & n4953 ) | ( n1184 & n4953 ) ;
  assign n4955 = ( ~n4949 & n4952 ) | ( ~n4949 & n4954 ) | ( n4952 & n4954 ) ;
  assign n4957 = ( x14 & x85 ) | ( x14 & ~n802 ) | ( x85 & ~n802 ) ;
  assign n4956 = ( n1800 & ~n1906 ) | ( n1800 & n2730 ) | ( ~n1906 & n2730 ) ;
  assign n4958 = n4957 ^ n4956 ^ n1472 ;
  assign n4959 = n2116 ^ n830 ^ n288 ;
  assign n4960 = n4959 ^ n2188 ^ x54 ;
  assign n4961 = ( n1863 & ~n4958 ) | ( n1863 & n4960 ) | ( ~n4958 & n4960 ) ;
  assign n4962 = n4961 ^ n4566 ^ n3647 ;
  assign n4963 = ( ~n1454 & n4955 ) | ( ~n1454 & n4962 ) | ( n4955 & n4962 ) ;
  assign n4964 = ( n1543 & n4948 ) | ( n1543 & ~n4963 ) | ( n4948 & ~n4963 ) ;
  assign n4965 = ( n1758 & n1860 ) | ( n1758 & ~n4572 ) | ( n1860 & ~n4572 ) ;
  assign n4966 = ( n850 & n1052 ) | ( n850 & ~n4554 ) | ( n1052 & ~n4554 ) ;
  assign n4967 = n4966 ^ n909 ^ n608 ;
  assign n4968 = ( n776 & n2041 ) | ( n776 & n4967 ) | ( n2041 & n4967 ) ;
  assign n4969 = ( n4439 & ~n4965 ) | ( n4439 & n4968 ) | ( ~n4965 & n4968 ) ;
  assign n4970 = ( ~n779 & n946 ) | ( ~n779 & n3068 ) | ( n946 & n3068 ) ;
  assign n4971 = ( n850 & ~n3205 ) | ( n850 & n4970 ) | ( ~n3205 & n4970 ) ;
  assign n4972 = ( n3170 & ~n4664 ) | ( n3170 & n4971 ) | ( ~n4664 & n4971 ) ;
  assign n4973 = ( ~n1151 & n2042 ) | ( ~n1151 & n2502 ) | ( n2042 & n2502 ) ;
  assign n4974 = n4973 ^ n4611 ^ n3232 ;
  assign n4975 = ( n2337 & ~n2750 ) | ( n2337 & n4974 ) | ( ~n2750 & n4974 ) ;
  assign n4976 = n4354 ^ n3004 ^ n2733 ;
  assign n4977 = n4976 ^ n1304 ^ n1179 ;
  assign n4978 = ( n3601 & ~n4134 ) | ( n3601 & n4977 ) | ( ~n4134 & n4977 ) ;
  assign n4979 = n3945 ^ n869 ^ n833 ;
  assign n4980 = ( ~n914 & n2793 ) | ( ~n914 & n3686 ) | ( n2793 & n3686 ) ;
  assign n4981 = n4980 ^ n2176 ^ x89 ;
  assign n4982 = n4981 ^ n1705 ^ n780 ;
  assign n4983 = ( n4783 & ~n4979 ) | ( n4783 & n4982 ) | ( ~n4979 & n4982 ) ;
  assign n4984 = ( n215 & n1318 ) | ( n215 & ~n3307 ) | ( n1318 & ~n3307 ) ;
  assign n4985 = n4984 ^ n1216 ^ n1188 ;
  assign n4986 = ( n3849 & n4044 ) | ( n3849 & n4985 ) | ( n4044 & n4985 ) ;
  assign n4987 = ( n330 & n4983 ) | ( n330 & n4986 ) | ( n4983 & n4986 ) ;
  assign n4988 = n4088 ^ n3071 ^ n1016 ;
  assign n4989 = n1358 ^ n621 ^ n191 ;
  assign n4990 = n4989 ^ n3677 ^ n2749 ;
  assign n4991 = n4990 ^ n2484 ^ n2161 ;
  assign n4992 = ( n2488 & n4988 ) | ( n2488 & ~n4991 ) | ( n4988 & ~n4991 ) ;
  assign n4993 = ( ~n2796 & n3921 ) | ( ~n2796 & n4992 ) | ( n3921 & n4992 ) ;
  assign n4994 = n3387 ^ n2236 ^ n1266 ;
  assign n4995 = ( ~n791 & n3620 ) | ( ~n791 & n4039 ) | ( n3620 & n4039 ) ;
  assign n4996 = n4995 ^ n1994 ^ n257 ;
  assign n4997 = n4996 ^ n2903 ^ n1434 ;
  assign n4998 = ( n2428 & n4994 ) | ( n2428 & ~n4997 ) | ( n4994 & ~n4997 ) ;
  assign n4999 = ( n307 & n3805 ) | ( n307 & ~n4998 ) | ( n3805 & ~n4998 ) ;
  assign n5000 = ( n188 & ~n4993 ) | ( n188 & n4999 ) | ( ~n4993 & n4999 ) ;
  assign n5001 = ( n1135 & n3211 ) | ( n1135 & n4816 ) | ( n3211 & n4816 ) ;
  assign n5002 = n5001 ^ n4438 ^ n3414 ;
  assign n5004 = n3690 ^ n3070 ^ x63 ;
  assign n5005 = n5004 ^ n2265 ^ n1947 ;
  assign n5003 = n4220 ^ n1520 ^ n1464 ;
  assign n5006 = n5005 ^ n5003 ^ n2861 ;
  assign n5007 = n5006 ^ n3315 ^ n370 ;
  assign n5008 = ( n2689 & ~n3113 ) | ( n2689 & n5007 ) | ( ~n3113 & n5007 ) ;
  assign n5009 = ( n258 & n1546 ) | ( n258 & n1839 ) | ( n1546 & n1839 ) ;
  assign n5010 = ( ~n1603 & n2834 ) | ( ~n1603 & n5009 ) | ( n2834 & n5009 ) ;
  assign n5011 = ( ~n706 & n5008 ) | ( ~n706 & n5010 ) | ( n5008 & n5010 ) ;
  assign n5012 = ( ~n1018 & n5002 ) | ( ~n1018 & n5011 ) | ( n5002 & n5011 ) ;
  assign n5013 = ( ~n1242 & n1886 ) | ( ~n1242 & n3702 ) | ( n1886 & n3702 ) ;
  assign n5014 = ( n1606 & n4342 ) | ( n1606 & n5013 ) | ( n4342 & n5013 ) ;
  assign n5031 = n435 ^ n309 ^ x6 ;
  assign n5032 = n5031 ^ n3349 ^ n923 ;
  assign n5029 = n4791 ^ n4063 ^ n2879 ;
  assign n5028 = n4382 ^ n1733 ^ n182 ;
  assign n5020 = ( ~n697 & n846 ) | ( ~n697 & n4744 ) | ( n846 & n4744 ) ;
  assign n5022 = ( n568 & ~n1377 ) | ( n568 & n2299 ) | ( ~n1377 & n2299 ) ;
  assign n5023 = n5022 ^ n2641 ^ n717 ;
  assign n5021 = ( n444 & ~n1319 ) | ( n444 & n3970 ) | ( ~n1319 & n3970 ) ;
  assign n5024 = n5023 ^ n5021 ^ n148 ;
  assign n5025 = ( n261 & ~n275 ) | ( n261 & n2094 ) | ( ~n275 & n2094 ) ;
  assign n5026 = ( ~n481 & n4175 ) | ( ~n481 & n5025 ) | ( n4175 & n5025 ) ;
  assign n5027 = ( ~n5020 & n5024 ) | ( ~n5020 & n5026 ) | ( n5024 & n5026 ) ;
  assign n5030 = n5029 ^ n5028 ^ n5027 ;
  assign n5015 = ( n316 & n553 ) | ( n316 & n968 ) | ( n553 & n968 ) ;
  assign n5016 = ( ~n1007 & n1233 ) | ( ~n1007 & n3174 ) | ( n1233 & n3174 ) ;
  assign n5017 = n5016 ^ n2066 ^ n587 ;
  assign n5018 = n3618 ^ n2233 ^ n295 ;
  assign n5019 = ( n5015 & n5017 ) | ( n5015 & n5018 ) | ( n5017 & n5018 ) ;
  assign n5033 = n5032 ^ n5030 ^ n5019 ;
  assign n5034 = n1505 ^ n1025 ^ n931 ;
  assign n5035 = n5034 ^ n850 ^ n228 ;
  assign n5036 = ( n618 & n3532 ) | ( n618 & ~n5035 ) | ( n3532 & ~n5035 ) ;
  assign n5044 = n2126 ^ n1275 ^ n981 ;
  assign n5045 = n5044 ^ n2697 ^ n2361 ;
  assign n5046 = n3829 ^ n1478 ^ n1241 ;
  assign n5047 = ( n291 & n2305 ) | ( n291 & ~n5046 ) | ( n2305 & ~n5046 ) ;
  assign n5051 = n3467 ^ n1066 ^ n200 ;
  assign n5052 = n4224 ^ n2103 ^ n1422 ;
  assign n5053 = n5052 ^ n3950 ^ n2580 ;
  assign n5054 = n3738 ^ n2060 ^ n685 ;
  assign n5055 = n5054 ^ n2642 ^ x43 ;
  assign n5056 = ( n1113 & n2643 ) | ( n1113 & ~n3081 ) | ( n2643 & ~n3081 ) ;
  assign n5057 = ( n1470 & n4122 ) | ( n1470 & n5056 ) | ( n4122 & n5056 ) ;
  assign n5058 = ( n4428 & n5055 ) | ( n4428 & n5057 ) | ( n5055 & n5057 ) ;
  assign n5059 = ( n5051 & ~n5053 ) | ( n5051 & n5058 ) | ( ~n5053 & n5058 ) ;
  assign n5060 = n5059 ^ n3830 ^ n1669 ;
  assign n5048 = ( n598 & n1305 ) | ( n598 & n1633 ) | ( n1305 & n1633 ) ;
  assign n5049 = ( n326 & ~n2211 ) | ( n326 & n2503 ) | ( ~n2211 & n2503 ) ;
  assign n5050 = ( n2265 & n5048 ) | ( n2265 & n5049 ) | ( n5048 & n5049 ) ;
  assign n5061 = n5060 ^ n5050 ^ n1236 ;
  assign n5062 = ( ~n5045 & n5047 ) | ( ~n5045 & n5061 ) | ( n5047 & n5061 ) ;
  assign n5038 = n1641 ^ n233 ^ x38 ;
  assign n5039 = ( n1866 & n3367 ) | ( n1866 & n5038 ) | ( n3367 & n5038 ) ;
  assign n5037 = ( n736 & n1436 ) | ( n736 & n3893 ) | ( n1436 & n3893 ) ;
  assign n5040 = n5039 ^ n5037 ^ n1640 ;
  assign n5041 = n5040 ^ n3816 ^ n225 ;
  assign n5042 = n5041 ^ n4938 ^ n3588 ;
  assign n5043 = n5042 ^ n2497 ^ n1819 ;
  assign n5063 = n5062 ^ n5043 ^ n3913 ;
  assign n5077 = n620 ^ n559 ^ x43 ;
  assign n5078 = n2765 ^ n2309 ^ n2215 ;
  assign n5079 = ( n1589 & n5077 ) | ( n1589 & ~n5078 ) | ( n5077 & ~n5078 ) ;
  assign n5080 = n5079 ^ n1996 ^ n1146 ;
  assign n5081 = ( ~n1444 & n2701 ) | ( ~n1444 & n5080 ) | ( n2701 & n5080 ) ;
  assign n5082 = ( n4286 & ~n4570 ) | ( n4286 & n5081 ) | ( ~n4570 & n5081 ) ;
  assign n5075 = ( n3618 & n4383 ) | ( n3618 & ~n4440 ) | ( n4383 & ~n4440 ) ;
  assign n5072 = ( n2459 & ~n3368 ) | ( n2459 & n3526 ) | ( ~n3368 & n3526 ) ;
  assign n5073 = ( ~n1397 & n2327 ) | ( ~n1397 & n5072 ) | ( n2327 & n5072 ) ;
  assign n5074 = ( ~n613 & n1727 ) | ( ~n613 & n5073 ) | ( n1727 & n5073 ) ;
  assign n5070 = ( n2515 & n3256 ) | ( n2515 & n3650 ) | ( n3256 & n3650 ) ;
  assign n5067 = ( n610 & n795 ) | ( n610 & n2343 ) | ( n795 & n2343 ) ;
  assign n5068 = ( n663 & n3216 ) | ( n663 & n5067 ) | ( n3216 & n5067 ) ;
  assign n5069 = n5068 ^ n4032 ^ n2253 ;
  assign n5064 = ( n641 & n1030 ) | ( n641 & n2145 ) | ( n1030 & n2145 ) ;
  assign n5065 = ( n940 & ~n4169 ) | ( n940 & n4300 ) | ( ~n4169 & n4300 ) ;
  assign n5066 = ( n3921 & n5064 ) | ( n3921 & n5065 ) | ( n5064 & n5065 ) ;
  assign n5071 = n5070 ^ n5069 ^ n5066 ;
  assign n5076 = n5075 ^ n5074 ^ n5071 ;
  assign n5083 = n5082 ^ n5076 ^ n1732 ;
  assign n5084 = ( n3678 & n4783 ) | ( n3678 & n5001 ) | ( n4783 & n5001 ) ;
  assign n5085 = n5084 ^ n3532 ^ n2055 ;
  assign n5086 = n4098 ^ n2339 ^ n726 ;
  assign n5087 = ( n1107 & n2147 ) | ( n1107 & ~n5086 ) | ( n2147 & ~n5086 ) ;
  assign n5088 = n5087 ^ n2629 ^ n2591 ;
  assign n5089 = ( x90 & n2036 ) | ( x90 & ~n2747 ) | ( n2036 & ~n2747 ) ;
  assign n5090 = n4060 ^ n468 ^ n460 ;
  assign n5091 = ( ~n4910 & n5089 ) | ( ~n4910 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5092 = ( n2678 & ~n3401 ) | ( n2678 & n5091 ) | ( ~n3401 & n5091 ) ;
  assign n5093 = ( n244 & ~n891 ) | ( n244 & n5092 ) | ( ~n891 & n5092 ) ;
  assign n5094 = ( ~n2477 & n2570 ) | ( ~n2477 & n5093 ) | ( n2570 & n5093 ) ;
  assign n5095 = n3902 ^ n3634 ^ n2793 ;
  assign n5096 = ( n224 & n644 ) | ( n224 & n5095 ) | ( n644 & n5095 ) ;
  assign n5097 = n3448 ^ n1122 ^ n223 ;
  assign n5098 = n5097 ^ n5077 ^ n1188 ;
  assign n5114 = ( x39 & ~n361 ) | ( x39 & n655 ) | ( ~n361 & n655 ) ;
  assign n5102 = ( ~n887 & n1524 ) | ( ~n887 & n2527 ) | ( n1524 & n2527 ) ;
  assign n5099 = n1504 ^ n443 ^ x98 ;
  assign n5100 = ( ~n583 & n1565 ) | ( ~n583 & n5099 ) | ( n1565 & n5099 ) ;
  assign n5101 = n5100 ^ n3699 ^ n1554 ;
  assign n5103 = n5102 ^ n5101 ^ n3956 ;
  assign n5104 = ( n2402 & n3758 ) | ( n2402 & n3904 ) | ( n3758 & n3904 ) ;
  assign n5110 = n3017 ^ n1191 ^ n914 ;
  assign n5108 = ( n480 & n1285 ) | ( n480 & ~n3124 ) | ( n1285 & ~n3124 ) ;
  assign n5109 = ( n1037 & n1148 ) | ( n1037 & ~n5108 ) | ( n1148 & ~n5108 ) ;
  assign n5105 = ( n1063 & n1448 ) | ( n1063 & n3799 ) | ( n1448 & n3799 ) ;
  assign n5106 = ( x53 & n3648 ) | ( x53 & ~n5105 ) | ( n3648 & ~n5105 ) ;
  assign n5107 = ( n780 & n1537 ) | ( n780 & ~n5106 ) | ( n1537 & ~n5106 ) ;
  assign n5111 = n5110 ^ n5109 ^ n5107 ;
  assign n5112 = ( n340 & n1095 ) | ( n340 & ~n5111 ) | ( n1095 & ~n5111 ) ;
  assign n5113 = ( n5103 & ~n5104 ) | ( n5103 & n5112 ) | ( ~n5104 & n5112 ) ;
  assign n5115 = n5114 ^ n5113 ^ n4703 ;
  assign n5131 = n4711 ^ n4197 ^ n1120 ;
  assign n5138 = ( n238 & n356 ) | ( n238 & n378 ) | ( n356 & n378 ) ;
  assign n5135 = n1290 ^ n1155 ^ n459 ;
  assign n5136 = n5135 ^ n1344 ^ n386 ;
  assign n5133 = ( ~n813 & n2428 ) | ( ~n813 & n4010 ) | ( n2428 & n4010 ) ;
  assign n5132 = n4089 ^ n2460 ^ n292 ;
  assign n5134 = n5133 ^ n5132 ^ n3011 ;
  assign n5137 = n5136 ^ n5134 ^ n2610 ;
  assign n5139 = n5138 ^ n5137 ^ n3067 ;
  assign n5140 = n5139 ^ n3139 ^ n1284 ;
  assign n5141 = ( ~n1379 & n2724 ) | ( ~n1379 & n3874 ) | ( n2724 & n3874 ) ;
  assign n5142 = n5141 ^ n2246 ^ n1312 ;
  assign n5143 = ( x56 & n2564 ) | ( x56 & n5142 ) | ( n2564 & n5142 ) ;
  assign n5144 = ( n5131 & ~n5140 ) | ( n5131 & n5143 ) | ( ~n5140 & n5143 ) ;
  assign n5128 = n1980 ^ n1174 ^ n264 ;
  assign n5129 = ( n505 & n3343 ) | ( n505 & n5128 ) | ( n3343 & n5128 ) ;
  assign n5126 = n1664 ^ n1378 ^ n596 ;
  assign n5124 = n2233 ^ n1400 ^ n1347 ;
  assign n5123 = n3656 ^ n3090 ^ n1371 ;
  assign n5121 = ( x29 & ~n3731 ) | ( x29 & n3777 ) | ( ~n3731 & n3777 ) ;
  assign n5118 = n1776 ^ n1098 ^ n211 ;
  assign n5119 = n5118 ^ n2343 ^ n2065 ;
  assign n5120 = n5119 ^ n4309 ^ n3446 ;
  assign n5122 = n5121 ^ n5120 ^ n3265 ;
  assign n5125 = n5124 ^ n5123 ^ n5122 ;
  assign n5127 = n5126 ^ n5125 ^ n4035 ;
  assign n5130 = n5129 ^ n5127 ^ n2504 ;
  assign n5116 = ( ~n856 & n1653 ) | ( ~n856 & n2225 ) | ( n1653 & n2225 ) ;
  assign n5117 = ( ~n2069 & n3405 ) | ( ~n2069 & n5116 ) | ( n3405 & n5116 ) ;
  assign n5145 = n5144 ^ n5130 ^ n5117 ;
  assign n5146 = n1504 ^ n853 ^ n635 ;
  assign n5147 = ( ~n772 & n2395 ) | ( ~n772 & n5146 ) | ( n2395 & n5146 ) ;
  assign n5148 = n5147 ^ n4009 ^ n437 ;
  assign n5149 = n2528 ^ n544 ^ n377 ;
  assign n5150 = n2007 ^ n1144 ^ n872 ;
  assign n5151 = n5150 ^ n5025 ^ n3229 ;
  assign n5154 = ( x13 & x14 ) | ( x13 & n1831 ) | ( x14 & n1831 ) ;
  assign n5152 = n3590 ^ n782 ^ n468 ;
  assign n5153 = n5152 ^ n3628 ^ n1109 ;
  assign n5155 = n5154 ^ n5153 ^ n826 ;
  assign n5156 = ( ~n5149 & n5151 ) | ( ~n5149 & n5155 ) | ( n5151 & n5155 ) ;
  assign n5157 = n4613 ^ n3654 ^ n388 ;
  assign n5158 = n5157 ^ n3706 ^ n1865 ;
  assign n5186 = n4041 ^ n1106 ^ n1091 ;
  assign n5159 = ( n509 & n4030 ) | ( n509 & n4291 ) | ( n4030 & n4291 ) ;
  assign n5160 = ( n244 & n1184 ) | ( n244 & ~n1346 ) | ( n1184 & ~n1346 ) ;
  assign n5161 = n5160 ^ n2403 ^ n1878 ;
  assign n5162 = ( ~n186 & n5159 ) | ( ~n186 & n5161 ) | ( n5159 & n5161 ) ;
  assign n5163 = ( n1536 & n3340 ) | ( n1536 & ~n5162 ) | ( n3340 & ~n5162 ) ;
  assign n5164 = ( n1783 & n1889 ) | ( n1783 & n5163 ) | ( n1889 & n5163 ) ;
  assign n5165 = ( n1287 & n3535 ) | ( n1287 & n5164 ) | ( n3535 & n5164 ) ;
  assign n5178 = ( ~n675 & n922 ) | ( ~n675 & n1047 ) | ( n922 & n1047 ) ;
  assign n5179 = ( n492 & n1081 ) | ( n492 & n5178 ) | ( n1081 & n5178 ) ;
  assign n5177 = n4224 ^ n2282 ^ n575 ;
  assign n5180 = n5179 ^ n5177 ^ n601 ;
  assign n5181 = ( n941 & ~n2569 ) | ( n941 & n5180 ) | ( ~n2569 & n5180 ) ;
  assign n5170 = n2201 ^ n1568 ^ n417 ;
  assign n5171 = n5170 ^ n2214 ^ n2059 ;
  assign n5172 = n5171 ^ n510 ^ x85 ;
  assign n5169 = n2902 ^ n1278 ^ n443 ;
  assign n5173 = n5172 ^ n5169 ^ n2932 ;
  assign n5174 = ( n205 & n1410 ) | ( n205 & ~n3638 ) | ( n1410 & ~n3638 ) ;
  assign n5175 = n3811 ^ n2912 ^ n186 ;
  assign n5176 = ( ~n5173 & n5174 ) | ( ~n5173 & n5175 ) | ( n5174 & n5175 ) ;
  assign n5182 = n5181 ^ n5176 ^ n3742 ;
  assign n5183 = n5182 ^ n3640 ^ x15 ;
  assign n5166 = ( ~n417 & n2407 ) | ( ~n417 & n5160 ) | ( n2407 & n5160 ) ;
  assign n5167 = n5166 ^ n3670 ^ n502 ;
  assign n5168 = n5167 ^ n3729 ^ x55 ;
  assign n5184 = n5183 ^ n5168 ^ n4771 ;
  assign n5185 = ( n954 & n5165 ) | ( n954 & ~n5184 ) | ( n5165 & ~n5184 ) ;
  assign n5187 = n5186 ^ n5185 ^ n1028 ;
  assign n5188 = ( n1939 & n1951 ) | ( n1939 & ~n5187 ) | ( n1951 & ~n5187 ) ;
  assign n5190 = ( n797 & ~n1672 ) | ( n797 & n2093 ) | ( ~n1672 & n2093 ) ;
  assign n5191 = n5190 ^ n4603 ^ n477 ;
  assign n5189 = ( ~n428 & n1845 ) | ( ~n428 & n2764 ) | ( n1845 & n2764 ) ;
  assign n5192 = n5191 ^ n5189 ^ n1466 ;
  assign n5193 = ( n185 & n321 ) | ( n185 & n644 ) | ( n321 & n644 ) ;
  assign n5194 = n4159 ^ n3234 ^ n928 ;
  assign n5195 = ( n2697 & ~n5193 ) | ( n2697 & n5194 ) | ( ~n5193 & n5194 ) ;
  assign n5196 = n5195 ^ n4743 ^ n2604 ;
  assign n5199 = n4863 ^ n1362 ^ n814 ;
  assign n5197 = ( n261 & n1378 ) | ( n261 & ~n2971 ) | ( n1378 & ~n2971 ) ;
  assign n5198 = n5197 ^ n5124 ^ n1791 ;
  assign n5200 = n5199 ^ n5198 ^ n2058 ;
  assign n5201 = ( n4640 & n5196 ) | ( n4640 & n5200 ) | ( n5196 & n5200 ) ;
  assign n5227 = n2040 ^ n296 ^ n292 ;
  assign n5231 = n2968 ^ n2034 ^ n349 ;
  assign n5229 = n4248 ^ n1420 ^ n472 ;
  assign n5230 = ( ~n1091 & n4216 ) | ( ~n1091 & n5229 ) | ( n4216 & n5229 ) ;
  assign n5232 = n5231 ^ n5230 ^ n653 ;
  assign n5233 = n5232 ^ n1931 ^ n1025 ;
  assign n5228 = n4185 ^ n3802 ^ n236 ;
  assign n5234 = n5233 ^ n5228 ^ n4169 ;
  assign n5236 = n1781 ^ n365 ^ n130 ;
  assign n5235 = n2066 ^ n1392 ^ n791 ;
  assign n5237 = n5236 ^ n5235 ^ n1683 ;
  assign n5238 = ( n1238 & n2787 ) | ( n1238 & n4482 ) | ( n2787 & n4482 ) ;
  assign n5239 = ( n561 & n5237 ) | ( n561 & ~n5238 ) | ( n5237 & ~n5238 ) ;
  assign n5240 = ( n3458 & n4297 ) | ( n3458 & n5239 ) | ( n4297 & n5239 ) ;
  assign n5241 = ( n5227 & ~n5234 ) | ( n5227 & n5240 ) | ( ~n5234 & n5240 ) ;
  assign n5208 = n4818 ^ n1669 ^ n1488 ;
  assign n5209 = n5208 ^ n4150 ^ n2741 ;
  assign n5210 = n3086 ^ n365 ^ n359 ;
  assign n5211 = ( x0 & n446 ) | ( x0 & ~n2126 ) | ( n446 & ~n2126 ) ;
  assign n5212 = n4216 ^ n1008 ^ n168 ;
  assign n5219 = ( n2838 & n4542 ) | ( n2838 & ~n5001 ) | ( n4542 & ~n5001 ) ;
  assign n5216 = ( ~n374 & n2437 ) | ( ~n374 & n3000 ) | ( n2437 & n3000 ) ;
  assign n5213 = n1359 ^ n1065 ^ n519 ;
  assign n5214 = ( n2079 & n2460 ) | ( n2079 & n5213 ) | ( n2460 & n5213 ) ;
  assign n5215 = n5214 ^ n3644 ^ n426 ;
  assign n5217 = n5216 ^ n5215 ^ n2000 ;
  assign n5218 = n5217 ^ n4848 ^ n4563 ;
  assign n5220 = n5219 ^ n5218 ^ n2103 ;
  assign n5221 = ( x25 & n5212 ) | ( x25 & n5220 ) | ( n5212 & n5220 ) ;
  assign n5222 = ( n751 & n5211 ) | ( n751 & n5221 ) | ( n5211 & n5221 ) ;
  assign n5223 = ( ~n1310 & n5210 ) | ( ~n1310 & n5222 ) | ( n5210 & n5222 ) ;
  assign n5224 = ( n3041 & n4420 ) | ( n3041 & ~n5223 ) | ( n4420 & ~n5223 ) ;
  assign n5225 = ( ~n2085 & n5209 ) | ( ~n2085 & n5224 ) | ( n5209 & n5224 ) ;
  assign n5226 = ( ~n676 & n3675 ) | ( ~n676 & n5225 ) | ( n3675 & n5225 ) ;
  assign n5202 = ( ~n1712 & n3062 ) | ( ~n1712 & n4124 ) | ( n3062 & n4124 ) ;
  assign n5203 = ( n787 & n2403 ) | ( n787 & n2676 ) | ( n2403 & n2676 ) ;
  assign n5204 = n4596 ^ n4371 ^ n390 ;
  assign n5205 = ( n2148 & ~n5203 ) | ( n2148 & n5204 ) | ( ~n5203 & n5204 ) ;
  assign n5206 = n5205 ^ n1628 ^ n1458 ;
  assign n5207 = ( n4935 & n5202 ) | ( n4935 & ~n5206 ) | ( n5202 & ~n5206 ) ;
  assign n5242 = n5241 ^ n5226 ^ n5207 ;
  assign n5247 = ( n729 & n1681 ) | ( n729 & ~n1735 ) | ( n1681 & ~n1735 ) ;
  assign n5245 = ( n510 & ~n871 ) | ( n510 & n2128 ) | ( ~n871 & n2128 ) ;
  assign n5243 = ( n209 & n464 ) | ( n209 & ~n5178 ) | ( n464 & ~n5178 ) ;
  assign n5244 = ( n1052 & ~n3427 ) | ( n1052 & n5243 ) | ( ~n3427 & n5243 ) ;
  assign n5246 = n5245 ^ n5244 ^ n619 ;
  assign n5248 = n5247 ^ n5246 ^ x95 ;
  assign n5249 = ( ~n568 & n2295 ) | ( ~n568 & n5248 ) | ( n2295 & n5248 ) ;
  assign n5250 = ( ~n3231 & n4098 ) | ( ~n3231 & n5249 ) | ( n4098 & n5249 ) ;
  assign n5263 = n3362 ^ n1789 ^ n839 ;
  assign n5264 = n4293 ^ n4271 ^ n587 ;
  assign n5265 = ( n2555 & n3339 ) | ( n2555 & n4379 ) | ( n3339 & n4379 ) ;
  assign n5266 = ( n5263 & ~n5264 ) | ( n5263 & n5265 ) | ( ~n5264 & n5265 ) ;
  assign n5259 = ( n574 & ~n2439 ) | ( n574 & n3765 ) | ( ~n2439 & n3765 ) ;
  assign n5260 = n5259 ^ n4810 ^ n2393 ;
  assign n5261 = n5260 ^ n4158 ^ n2246 ;
  assign n5258 = ( x104 & n3555 ) | ( x104 & ~n4437 ) | ( n3555 & ~n4437 ) ;
  assign n5262 = n5261 ^ n5258 ^ n158 ;
  assign n5251 = n2698 ^ n2419 ^ n460 ;
  assign n5252 = n5251 ^ n3781 ^ n3189 ;
  assign n5253 = ( n2169 & n4122 ) | ( n2169 & n5252 ) | ( n4122 & n5252 ) ;
  assign n5254 = ( ~n713 & n746 ) | ( ~n713 & n3476 ) | ( n746 & n3476 ) ;
  assign n5255 = n5254 ^ n4046 ^ n3111 ;
  assign n5256 = ( n2595 & ~n5253 ) | ( n2595 & n5255 ) | ( ~n5253 & n5255 ) ;
  assign n5257 = n5256 ^ n3678 ^ n1812 ;
  assign n5267 = n5266 ^ n5262 ^ n5257 ;
  assign n5268 = n5267 ^ n4869 ^ n142 ;
  assign n5274 = n1935 ^ n1728 ^ n515 ;
  assign n5275 = ( n642 & n4847 ) | ( n642 & ~n5274 ) | ( n4847 & ~n5274 ) ;
  assign n5273 = n5044 ^ n2220 ^ n668 ;
  assign n5269 = n2244 ^ n1353 ^ n524 ;
  assign n5270 = n5269 ^ n5089 ^ n4168 ;
  assign n5271 = n5270 ^ n5065 ^ n534 ;
  assign n5272 = ( n2643 & n2741 ) | ( n2643 & n5271 ) | ( n2741 & n5271 ) ;
  assign n5276 = n5275 ^ n5273 ^ n5272 ;
  assign n5277 = ( ~n1096 & n2220 ) | ( ~n1096 & n5276 ) | ( n2220 & n5276 ) ;
  assign n5280 = n5025 ^ n786 ^ n266 ;
  assign n5281 = ( n893 & n1101 ) | ( n893 & n5280 ) | ( n1101 & n5280 ) ;
  assign n5282 = ( n4165 & ~n4646 ) | ( n4165 & n5281 ) | ( ~n4646 & n5281 ) ;
  assign n5287 = ( x72 & ~n2419 ) | ( x72 & n3677 ) | ( ~n2419 & n3677 ) ;
  assign n5283 = n2574 ^ n1694 ^ n1074 ;
  assign n5284 = ( n1501 & ~n2186 ) | ( n1501 & n5283 ) | ( ~n2186 & n5283 ) ;
  assign n5285 = ( n1052 & n3892 ) | ( n1052 & n5284 ) | ( n3892 & n5284 ) ;
  assign n5286 = ( n718 & n2280 ) | ( n718 & n5285 ) | ( n2280 & n5285 ) ;
  assign n5288 = n5287 ^ n5286 ^ n1277 ;
  assign n5289 = ( n2341 & ~n5282 ) | ( n2341 & n5288 ) | ( ~n5282 & n5288 ) ;
  assign n5278 = ( ~n2000 & n2328 ) | ( ~n2000 & n2814 ) | ( n2328 & n2814 ) ;
  assign n5279 = n5278 ^ n3438 ^ n2338 ;
  assign n5290 = n5289 ^ n5279 ^ n2994 ;
  assign n5298 = n3978 ^ n1216 ^ n490 ;
  assign n5293 = ( n1385 & n2501 ) | ( n1385 & n4002 ) | ( n2501 & n4002 ) ;
  assign n5294 = n3318 ^ n1134 ^ n303 ;
  assign n5295 = ( n599 & ~n5293 ) | ( n599 & n5294 ) | ( ~n5293 & n5294 ) ;
  assign n5296 = n5295 ^ n3810 ^ n2883 ;
  assign n5297 = n5296 ^ n2660 ^ n154 ;
  assign n5291 = n4174 ^ n3946 ^ n526 ;
  assign n5292 = ( n141 & ~n3057 ) | ( n141 & n5291 ) | ( ~n3057 & n5291 ) ;
  assign n5299 = n5298 ^ n5297 ^ n5292 ;
  assign n5300 = ( n2845 & ~n4968 ) | ( n2845 & n5299 ) | ( ~n4968 & n5299 ) ;
  assign n5335 = n3256 ^ n2745 ^ n1860 ;
  assign n5331 = n5280 ^ n1343 ^ n1254 ;
  assign n5332 = n5331 ^ n2874 ^ n918 ;
  assign n5333 = ( ~n782 & n2876 ) | ( ~n782 & n5332 ) | ( n2876 & n5332 ) ;
  assign n5329 = n4628 ^ n2542 ^ n409 ;
  assign n5313 = n2662 ^ n1748 ^ n516 ;
  assign n5330 = n5329 ^ n5313 ^ n3545 ;
  assign n5334 = n5333 ^ n5330 ^ n2896 ;
  assign n5336 = n5335 ^ n5334 ^ n799 ;
  assign n5326 = ( n545 & n3430 ) | ( n545 & n3431 ) | ( n3430 & n3431 ) ;
  assign n5327 = n5326 ^ n4058 ^ n3454 ;
  assign n5301 = ( n1295 & ~n3457 ) | ( n1295 & n5052 ) | ( ~n3457 & n5052 ) ;
  assign n5302 = n5301 ^ n2131 ^ n524 ;
  assign n5303 = n4796 ^ n3323 ^ n213 ;
  assign n5304 = ( n1838 & n3467 ) | ( n1838 & n3886 ) | ( n3467 & n3886 ) ;
  assign n5305 = ( n2338 & n4055 ) | ( n2338 & n5304 ) | ( n4055 & n5304 ) ;
  assign n5306 = ( n2119 & n2704 ) | ( n2119 & ~n5305 ) | ( n2704 & ~n5305 ) ;
  assign n5307 = n5306 ^ n2008 ^ n724 ;
  assign n5308 = n5307 ^ n5306 ^ n2343 ;
  assign n5309 = ( n215 & ~n1630 ) | ( n215 & n4595 ) | ( ~n1630 & n4595 ) ;
  assign n5317 = ( n992 & n1390 ) | ( n992 & ~n1626 ) | ( n1390 & ~n1626 ) ;
  assign n5316 = n3406 ^ n2366 ^ n1836 ;
  assign n5312 = ( x100 & n2429 ) | ( x100 & n3741 ) | ( n2429 & n3741 ) ;
  assign n5314 = n5313 ^ n5312 ^ n1661 ;
  assign n5310 = ( n1571 & n2712 ) | ( n1571 & n3535 ) | ( n2712 & n3535 ) ;
  assign n5311 = ( x34 & ~n2904 ) | ( x34 & n5310 ) | ( ~n2904 & n5310 ) ;
  assign n5315 = n5314 ^ n5311 ^ n1999 ;
  assign n5318 = n5317 ^ n5316 ^ n5315 ;
  assign n5319 = ( n3996 & n4225 ) | ( n3996 & n5318 ) | ( n4225 & n5318 ) ;
  assign n5320 = ( n3154 & n5309 ) | ( n3154 & n5319 ) | ( n5309 & n5319 ) ;
  assign n5321 = ( ~n1298 & n1486 ) | ( ~n1298 & n3834 ) | ( n1486 & n3834 ) ;
  assign n5322 = ( x0 & ~n1909 ) | ( x0 & n5321 ) | ( ~n1909 & n5321 ) ;
  assign n5323 = ( ~n762 & n3611 ) | ( ~n762 & n5322 ) | ( n3611 & n5322 ) ;
  assign n5324 = ( ~n5308 & n5320 ) | ( ~n5308 & n5323 ) | ( n5320 & n5323 ) ;
  assign n5325 = ( n5302 & ~n5303 ) | ( n5302 & n5324 ) | ( ~n5303 & n5324 ) ;
  assign n5328 = n5327 ^ n5325 ^ n2926 ;
  assign n5337 = n5336 ^ n5328 ^ n415 ;
  assign n5338 = n5337 ^ n2976 ^ n1264 ;
  assign n5353 = ( x9 & n2248 ) | ( x9 & n3556 ) | ( n2248 & n3556 ) ;
  assign n5354 = ( ~n974 & n4942 ) | ( ~n974 & n5353 ) | ( n4942 & n5353 ) ;
  assign n5349 = n4325 ^ n3425 ^ n2141 ;
  assign n5350 = ( x116 & n415 ) | ( x116 & ~n2296 ) | ( n415 & ~n2296 ) ;
  assign n5351 = n5350 ^ n1784 ^ n814 ;
  assign n5352 = ( n5123 & ~n5349 ) | ( n5123 & n5351 ) | ( ~n5349 & n5351 ) ;
  assign n5342 = n2697 ^ n1028 ^ n895 ;
  assign n5343 = n5342 ^ n4669 ^ n1807 ;
  assign n5340 = ( n168 & ~n1170 ) | ( n168 & n1507 ) | ( ~n1170 & n1507 ) ;
  assign n5339 = n1143 ^ n895 ^ n360 ;
  assign n5341 = n5340 ^ n5339 ^ n3255 ;
  assign n5344 = n5343 ^ n5341 ^ n2115 ;
  assign n5345 = n1343 ^ n725 ^ n650 ;
  assign n5346 = n5345 ^ n1999 ^ n1005 ;
  assign n5347 = ( n3118 & n3275 ) | ( n3118 & n5346 ) | ( n3275 & n5346 ) ;
  assign n5348 = ( n1504 & ~n5344 ) | ( n1504 & n5347 ) | ( ~n5344 & n5347 ) ;
  assign n5355 = n5354 ^ n5352 ^ n5348 ;
  assign n5356 = n4439 ^ n2375 ^ n1208 ;
  assign n5357 = ( n1980 & n3088 ) | ( n1980 & n5356 ) | ( n3088 & n5356 ) ;
  assign n5358 = n3644 ^ n645 ^ n303 ;
  assign n5359 = ( n819 & n4760 ) | ( n819 & n5358 ) | ( n4760 & n5358 ) ;
  assign n5360 = n5359 ^ n4706 ^ n3432 ;
  assign n5361 = ( ~n291 & n5357 ) | ( ~n291 & n5360 ) | ( n5357 & n5360 ) ;
  assign n5362 = ( n1227 & n5047 ) | ( n1227 & ~n5361 ) | ( n5047 & ~n5361 ) ;
  assign n5363 = ( n657 & n1923 ) | ( n657 & n2448 ) | ( n1923 & n2448 ) ;
  assign n5364 = ( n1173 & ~n4519 ) | ( n1173 & n5363 ) | ( ~n4519 & n5363 ) ;
  assign n5365 = ( ~n1827 & n5362 ) | ( ~n1827 & n5364 ) | ( n5362 & n5364 ) ;
  assign n5366 = ( ~n3511 & n4005 ) | ( ~n3511 & n4256 ) | ( n4005 & n4256 ) ;
  assign n5377 = n5175 ^ n4711 ^ n3657 ;
  assign n5372 = ( n371 & n3503 ) | ( n371 & n3729 ) | ( n3503 & n3729 ) ;
  assign n5373 = n5372 ^ n2939 ^ n608 ;
  assign n5374 = ( ~n2631 & n3767 ) | ( ~n2631 & n4429 ) | ( n3767 & n4429 ) ;
  assign n5375 = ( n493 & n549 ) | ( n493 & n3557 ) | ( n549 & n3557 ) ;
  assign n5376 = ( ~n5373 & n5374 ) | ( ~n5373 & n5375 ) | ( n5374 & n5375 ) ;
  assign n5378 = n5377 ^ n5376 ^ n2126 ;
  assign n5367 = n2204 ^ n712 ^ x33 ;
  assign n5368 = n5367 ^ n3196 ^ n1774 ;
  assign n5369 = ( n440 & n2608 ) | ( n440 & ~n5368 ) | ( n2608 & ~n5368 ) ;
  assign n5370 = n5369 ^ n4297 ^ n1312 ;
  assign n5371 = n5370 ^ n2897 ^ n1472 ;
  assign n5379 = n5378 ^ n5371 ^ n2229 ;
  assign n5380 = ( n2183 & ~n2512 ) | ( n2183 & n3157 ) | ( ~n2512 & n3157 ) ;
  assign n5385 = ( n1709 & n1938 ) | ( n1709 & ~n4526 ) | ( n1938 & ~n4526 ) ;
  assign n5386 = n5385 ^ n2701 ^ n861 ;
  assign n5384 = n4447 ^ n3105 ^ n1362 ;
  assign n5381 = ( n805 & ~n1900 ) | ( n805 & n2701 ) | ( ~n1900 & n2701 ) ;
  assign n5382 = n5381 ^ n1786 ^ n262 ;
  assign n5383 = n5382 ^ n3511 ^ n1947 ;
  assign n5387 = n5386 ^ n5384 ^ n5383 ;
  assign n5388 = ( ~n1893 & n5380 ) | ( ~n1893 & n5387 ) | ( n5380 & n5387 ) ;
  assign n5389 = ( n5366 & n5379 ) | ( n5366 & n5388 ) | ( n5379 & n5388 ) ;
  assign n5407 = ( n1073 & ~n1727 ) | ( n1073 & n5314 ) | ( ~n1727 & n5314 ) ;
  assign n5410 = ( n923 & n3904 ) | ( n923 & ~n4951 ) | ( n3904 & ~n4951 ) ;
  assign n5408 = ( n1182 & n4334 ) | ( n1182 & ~n5179 ) | ( n4334 & ~n5179 ) ;
  assign n5409 = n5408 ^ n2681 ^ n1940 ;
  assign n5411 = n5410 ^ n5409 ^ n872 ;
  assign n5412 = ( n1512 & n5407 ) | ( n1512 & n5411 ) | ( n5407 & n5411 ) ;
  assign n5403 = n1551 ^ n507 ^ n144 ;
  assign n5404 = ( ~n396 & n3792 ) | ( ~n396 & n5403 ) | ( n3792 & n5403 ) ;
  assign n5400 = ( ~n727 & n1062 ) | ( ~n727 & n1367 ) | ( n1062 & n1367 ) ;
  assign n5401 = ( n231 & n2977 ) | ( n231 & n5400 ) | ( n2977 & n5400 ) ;
  assign n5402 = n5401 ^ n4428 ^ n1668 ;
  assign n5405 = n5404 ^ n5402 ^ n1829 ;
  assign n5406 = n5405 ^ n4368 ^ n1111 ;
  assign n5390 = ( n627 & n1805 ) | ( n627 & n2848 ) | ( n1805 & n2848 ) ;
  assign n5391 = n5390 ^ n3757 ^ x96 ;
  assign n5392 = n5391 ^ n2862 ^ n739 ;
  assign n5393 = n4227 ^ n3477 ^ n3139 ;
  assign n5394 = ( n1807 & ~n5392 ) | ( n1807 & n5393 ) | ( ~n5392 & n5393 ) ;
  assign n5395 = ( ~n1251 & n5054 ) | ( ~n1251 & n5394 ) | ( n5054 & n5394 ) ;
  assign n5396 = n2313 ^ n1691 ^ n1567 ;
  assign n5397 = n4369 ^ n2429 ^ n2060 ;
  assign n5398 = ( n187 & n5396 ) | ( n187 & n5397 ) | ( n5396 & n5397 ) ;
  assign n5399 = ( n1460 & n5395 ) | ( n1460 & n5398 ) | ( n5395 & n5398 ) ;
  assign n5413 = n5412 ^ n5406 ^ n5399 ;
  assign n5414 = n3567 ^ n964 ^ n719 ;
  assign n5415 = n5414 ^ n3326 ^ n675 ;
  assign n5416 = ( x62 & n725 ) | ( x62 & ~n3124 ) | ( n725 & ~n3124 ) ;
  assign n5417 = ( n818 & n872 ) | ( n818 & ~n5416 ) | ( n872 & ~n5416 ) ;
  assign n5418 = ( ~n1254 & n5415 ) | ( ~n1254 & n5417 ) | ( n5415 & n5417 ) ;
  assign n5419 = n5418 ^ n3825 ^ n640 ;
  assign n5420 = ( n2687 & n3426 ) | ( n2687 & ~n4607 ) | ( n3426 & ~n4607 ) ;
  assign n5421 = n5319 ^ n3530 ^ n3027 ;
  assign n5422 = n5421 ^ n3681 ^ x47 ;
  assign n5423 = ( n5419 & n5420 ) | ( n5419 & ~n5422 ) | ( n5420 & ~n5422 ) ;
  assign n5428 = ( x92 & n423 ) | ( x92 & ~n922 ) | ( n423 & ~n922 ) ;
  assign n5426 = ( n1209 & ~n1612 ) | ( n1209 & n1710 ) | ( ~n1612 & n1710 ) ;
  assign n5424 = ( x27 & ~n1841 ) | ( x27 & n2309 ) | ( ~n1841 & n2309 ) ;
  assign n5425 = n5424 ^ n4428 ^ n1016 ;
  assign n5427 = n5426 ^ n5425 ^ n2201 ;
  assign n5429 = n5428 ^ n5427 ^ n3100 ;
  assign n5430 = n5429 ^ n3873 ^ n3098 ;
  assign n5431 = ( n2102 & n3404 ) | ( n2102 & n4091 ) | ( n3404 & n4091 ) ;
  assign n5432 = ( ~n1341 & n2374 ) | ( ~n1341 & n3187 ) | ( n2374 & n3187 ) ;
  assign n5433 = ( n2162 & ~n4805 ) | ( n2162 & n5432 ) | ( ~n4805 & n5432 ) ;
  assign n5436 = ( n1703 & n1936 ) | ( n1703 & n2183 ) | ( n1936 & n2183 ) ;
  assign n5435 = n2521 ^ n1769 ^ n1048 ;
  assign n5434 = ( n2204 & n2220 ) | ( n2204 & n4571 ) | ( n2220 & n4571 ) ;
  assign n5437 = n5436 ^ n5435 ^ n5434 ;
  assign n5438 = ( n1623 & n3110 ) | ( n1623 & ~n5437 ) | ( n3110 & ~n5437 ) ;
  assign n5439 = n3314 ^ n1132 ^ n652 ;
  assign n5440 = ( n148 & n746 ) | ( n148 & ~n5439 ) | ( n746 & ~n5439 ) ;
  assign n5441 = ( n571 & ~n3168 ) | ( n571 & n5341 ) | ( ~n3168 & n5341 ) ;
  assign n5442 = ( n3399 & ~n5440 ) | ( n3399 & n5441 ) | ( ~n5440 & n5441 ) ;
  assign n5443 = ( n5433 & n5438 ) | ( n5433 & n5442 ) | ( n5438 & n5442 ) ;
  assign n5450 = ( ~n550 & n886 ) | ( ~n550 & n2365 ) | ( n886 & n2365 ) ;
  assign n5451 = n5450 ^ n1451 ^ n955 ;
  assign n5448 = ( ~n848 & n1426 ) | ( ~n848 & n2050 ) | ( n1426 & n2050 ) ;
  assign n5449 = n5448 ^ n2491 ^ n2209 ;
  assign n5446 = ( ~n137 & n2367 ) | ( ~n137 & n3305 ) | ( n2367 & n3305 ) ;
  assign n5444 = ( n706 & n970 ) | ( n706 & ~n3002 ) | ( n970 & ~n3002 ) ;
  assign n5445 = ( n1682 & ~n4110 ) | ( n1682 & n5444 ) | ( ~n4110 & n5444 ) ;
  assign n5447 = n5446 ^ n5445 ^ x121 ;
  assign n5452 = n5451 ^ n5449 ^ n5447 ;
  assign n5453 = ( n4463 & n4669 ) | ( n4463 & ~n5452 ) | ( n4669 & ~n5452 ) ;
  assign n5456 = n1464 ^ n1333 ^ n148 ;
  assign n5457 = ( n3944 & n4174 ) | ( n3944 & ~n5456 ) | ( n4174 & ~n5456 ) ;
  assign n5454 = ( n1279 & ~n3582 ) | ( n1279 & n5067 ) | ( ~n3582 & n5067 ) ;
  assign n5455 = ( ~n1180 & n1359 ) | ( ~n1180 & n5454 ) | ( n1359 & n5454 ) ;
  assign n5458 = n5457 ^ n5455 ^ n2161 ;
  assign n5480 = ( n2236 & n3581 ) | ( n2236 & n3973 ) | ( n3581 & n3973 ) ;
  assign n5476 = ( ~n447 & n3490 ) | ( ~n447 & n4460 ) | ( n3490 & n4460 ) ;
  assign n5477 = n5476 ^ n1350 ^ n1249 ;
  assign n5470 = n632 ^ n310 ^ n291 ;
  assign n5471 = n5470 ^ n2764 ^ n1971 ;
  assign n5472 = n2419 ^ n2037 ^ n906 ;
  assign n5473 = ( ~n536 & n5471 ) | ( ~n536 & n5472 ) | ( n5471 & n5472 ) ;
  assign n5474 = n5473 ^ n5408 ^ n437 ;
  assign n5475 = n5474 ^ n1864 ^ n718 ;
  assign n5478 = n5477 ^ n5475 ^ n755 ;
  assign n5479 = ( ~n648 & n3796 ) | ( ~n648 & n5478 ) | ( n3796 & n5478 ) ;
  assign n5466 = ( n1179 & n2208 ) | ( n1179 & n2621 ) | ( n2208 & n2621 ) ;
  assign n5467 = n3429 ^ n2389 ^ n1070 ;
  assign n5468 = ( n3490 & ~n5466 ) | ( n3490 & n5467 ) | ( ~n5466 & n5467 ) ;
  assign n5459 = n4027 ^ n2685 ^ n255 ;
  assign n5460 = ( ~n1184 & n2993 ) | ( ~n1184 & n4039 ) | ( n2993 & n4039 ) ;
  assign n5461 = ( n1180 & n1206 ) | ( n1180 & n5460 ) | ( n1206 & n5460 ) ;
  assign n5462 = n5461 ^ n1002 ^ n984 ;
  assign n5463 = n5462 ^ n1481 ^ n651 ;
  assign n5464 = n5463 ^ n1946 ^ n381 ;
  assign n5465 = ( ~n1157 & n5459 ) | ( ~n1157 & n5464 ) | ( n5459 & n5464 ) ;
  assign n5469 = n5468 ^ n5465 ^ n3632 ;
  assign n5481 = n5480 ^ n5479 ^ n5469 ;
  assign n5489 = n1355 ^ n1184 ^ n263 ;
  assign n5487 = ( ~n1751 & n2734 ) | ( ~n1751 & n4585 ) | ( n2734 & n4585 ) ;
  assign n5485 = n2101 ^ n1686 ^ n823 ;
  assign n5484 = n5179 ^ n1861 ^ n800 ;
  assign n5482 = ( n142 & ~n748 ) | ( n142 & n889 ) | ( ~n748 & n889 ) ;
  assign n5483 = n5482 ^ n4613 ^ n4373 ;
  assign n5486 = n5485 ^ n5484 ^ n5483 ;
  assign n5488 = n5487 ^ n5486 ^ n465 ;
  assign n5490 = n5489 ^ n5488 ^ n3600 ;
  assign n5497 = n2859 ^ n2831 ^ n1204 ;
  assign n5498 = ( n334 & n4501 ) | ( n334 & n5497 ) | ( n4501 & n5497 ) ;
  assign n5491 = n1619 ^ n1595 ^ x40 ;
  assign n5492 = n5491 ^ n3835 ^ n1582 ;
  assign n5493 = n3936 ^ n1667 ^ x127 ;
  assign n5494 = ( n3703 & ~n5492 ) | ( n3703 & n5493 ) | ( ~n5492 & n5493 ) ;
  assign n5495 = ( ~n1922 & n2339 ) | ( ~n1922 & n5494 ) | ( n2339 & n5494 ) ;
  assign n5496 = ( ~n1774 & n2176 ) | ( ~n1774 & n5495 ) | ( n2176 & n5495 ) ;
  assign n5499 = n5498 ^ n5496 ^ n2241 ;
  assign n5501 = ( ~x41 & n1685 ) | ( ~x41 & n2698 ) | ( n1685 & n2698 ) ;
  assign n5500 = n4257 ^ n3704 ^ n335 ;
  assign n5502 = n5501 ^ n5500 ^ n771 ;
  assign n5504 = n2621 ^ n2527 ^ n652 ;
  assign n5505 = ( x88 & ~n250 ) | ( x88 & n5504 ) | ( ~n250 & n5504 ) ;
  assign n5503 = n3457 ^ n3454 ^ n3191 ;
  assign n5506 = n5505 ^ n5503 ^ n5386 ;
  assign n5507 = ( n775 & n5502 ) | ( n775 & n5506 ) | ( n5502 & n5506 ) ;
  assign n5508 = n3855 ^ n3676 ^ n900 ;
  assign n5509 = n5508 ^ n4142 ^ n2256 ;
  assign n5514 = n4383 ^ n2070 ^ x77 ;
  assign n5515 = ( n4586 & ~n4855 ) | ( n4586 & n5514 ) | ( ~n4855 & n5514 ) ;
  assign n5510 = ( n645 & n1005 ) | ( n645 & n4135 ) | ( n1005 & n4135 ) ;
  assign n5511 = n3714 ^ n2203 ^ n210 ;
  assign n5512 = ( n400 & n5510 ) | ( n400 & ~n5511 ) | ( n5510 & ~n5511 ) ;
  assign n5513 = n5512 ^ n690 ^ x120 ;
  assign n5516 = n5515 ^ n5513 ^ n3104 ;
  assign n5517 = ( n5212 & n5509 ) | ( n5212 & ~n5516 ) | ( n5509 & ~n5516 ) ;
  assign n5521 = ( x106 & ~n803 ) | ( x106 & n1829 ) | ( ~n803 & n1829 ) ;
  assign n5522 = n5521 ^ n3619 ^ n1226 ;
  assign n5520 = ( n166 & n4010 ) | ( n166 & n4379 ) | ( n4010 & n4379 ) ;
  assign n5518 = ( n1136 & n1535 ) | ( n1136 & ~n1698 ) | ( n1535 & ~n1698 ) ;
  assign n5519 = n5518 ^ n2525 ^ x6 ;
  assign n5523 = n5522 ^ n5520 ^ n5519 ;
  assign n5529 = n2051 ^ n433 ^ n353 ;
  assign n5528 = ( ~x34 & n294 ) | ( ~x34 & n1052 ) | ( n294 & n1052 ) ;
  assign n5530 = n5529 ^ n5528 ^ n2668 ;
  assign n5526 = ( n345 & n972 ) | ( n345 & n4957 ) | ( n972 & n4957 ) ;
  assign n5527 = ( n1368 & n2505 ) | ( n1368 & n5526 ) | ( n2505 & n5526 ) ;
  assign n5531 = n5530 ^ n5527 ^ n931 ;
  assign n5524 = n4364 ^ n2719 ^ n227 ;
  assign n5525 = ( n1276 & n2523 ) | ( n1276 & ~n5524 ) | ( n2523 & ~n5524 ) ;
  assign n5532 = n5531 ^ n5525 ^ n3007 ;
  assign n5533 = n1327 ^ n811 ^ n692 ;
  assign n5534 = n5533 ^ n1887 ^ n1561 ;
  assign n5535 = n3729 ^ n1328 ^ x91 ;
  assign n5536 = ( ~n806 & n932 ) | ( ~n806 & n5178 ) | ( n932 & n5178 ) ;
  assign n5537 = ( n3921 & n4095 ) | ( n3921 & n5536 ) | ( n4095 & n5536 ) ;
  assign n5538 = n3971 ^ n2274 ^ n709 ;
  assign n5539 = ( n780 & n2748 ) | ( n780 & ~n5538 ) | ( n2748 & ~n5538 ) ;
  assign n5540 = ( x12 & ~n4834 ) | ( x12 & n5539 ) | ( ~n4834 & n5539 ) ;
  assign n5541 = n4055 ^ n3543 ^ n2608 ;
  assign n5542 = ( n809 & n5540 ) | ( n809 & n5541 ) | ( n5540 & n5541 ) ;
  assign n5543 = ( n926 & n2771 ) | ( n926 & ~n5542 ) | ( n2771 & ~n5542 ) ;
  assign n5559 = n4769 ^ n707 ^ x90 ;
  assign n5558 = n1273 ^ n1098 ^ n239 ;
  assign n5560 = n5559 ^ n5558 ^ n2438 ;
  assign n5554 = n3294 ^ n769 ^ n631 ;
  assign n5555 = ( n1651 & n2837 ) | ( n1651 & n5554 ) | ( n2837 & n5554 ) ;
  assign n5556 = n3495 ^ n3412 ^ n917 ;
  assign n5557 = ( ~n2313 & n5555 ) | ( ~n2313 & n5556 ) | ( n5555 & n5556 ) ;
  assign n5544 = ( n413 & n1490 ) | ( n413 & ~n2400 ) | ( n1490 & ~n2400 ) ;
  assign n5545 = n1967 ^ n260 ^ n214 ;
  assign n5546 = n1781 ^ n676 ^ n495 ;
  assign n5547 = ( x107 & n511 ) | ( x107 & ~n2256 ) | ( n511 & ~n2256 ) ;
  assign n5548 = n5547 ^ n1436 ^ n812 ;
  assign n5549 = ( n804 & ~n5546 ) | ( n804 & n5548 ) | ( ~n5546 & n5548 ) ;
  assign n5550 = ( n3742 & n3807 ) | ( n3742 & ~n5549 ) | ( n3807 & ~n5549 ) ;
  assign n5551 = ( n275 & n5545 ) | ( n275 & ~n5550 ) | ( n5545 & ~n5550 ) ;
  assign n5552 = ( ~n3109 & n3778 ) | ( ~n3109 & n5551 ) | ( n3778 & n5551 ) ;
  assign n5553 = ( ~n968 & n5544 ) | ( ~n968 & n5552 ) | ( n5544 & n5552 ) ;
  assign n5561 = n5560 ^ n5557 ^ n5553 ;
  assign n5562 = ( ~n1439 & n1452 ) | ( ~n1439 & n5561 ) | ( n1452 & n5561 ) ;
  assign n5563 = ( x20 & ~n473 ) | ( x20 & n3810 ) | ( ~n473 & n3810 ) ;
  assign n5564 = ( x58 & ~n982 ) | ( x58 & n5563 ) | ( ~n982 & n5563 ) ;
  assign n5565 = ( ~n308 & n1246 ) | ( ~n308 & n2137 ) | ( n1246 & n2137 ) ;
  assign n5566 = n4299 ^ n825 ^ n466 ;
  assign n5567 = ( n3806 & ~n5565 ) | ( n3806 & n5566 ) | ( ~n5565 & n5566 ) ;
  assign n5568 = ( x52 & n5564 ) | ( x52 & ~n5567 ) | ( n5564 & ~n5567 ) ;
  assign n5575 = ( n632 & n1450 ) | ( n632 & ~n2175 ) | ( n1450 & ~n2175 ) ;
  assign n5570 = n5038 ^ n2280 ^ n239 ;
  assign n5571 = ( n1752 & n2244 ) | ( n1752 & ~n5570 ) | ( n2244 & ~n5570 ) ;
  assign n5572 = n5571 ^ n3050 ^ n428 ;
  assign n5569 = ( n1216 & n3503 ) | ( n1216 & n4265 ) | ( n3503 & n4265 ) ;
  assign n5573 = n5572 ^ n5569 ^ n1510 ;
  assign n5574 = n5573 ^ n1206 ^ n680 ;
  assign n5576 = n5575 ^ n5574 ^ n2307 ;
  assign n5589 = ( x37 & n263 ) | ( x37 & ~n4459 ) | ( n263 & ~n4459 ) ;
  assign n5590 = ( ~n1563 & n3056 ) | ( ~n1563 & n5589 ) | ( n3056 & n5589 ) ;
  assign n5585 = ( n790 & n3906 ) | ( n790 & ~n4407 ) | ( n3906 & ~n4407 ) ;
  assign n5586 = ( n1873 & ~n3504 ) | ( n1873 & n5585 ) | ( ~n3504 & n5585 ) ;
  assign n5581 = n3845 ^ n3196 ^ n2080 ;
  assign n5582 = ( n454 & n3552 ) | ( n454 & ~n5581 ) | ( n3552 & ~n5581 ) ;
  assign n5583 = ( n2527 & n3115 ) | ( n2527 & n5582 ) | ( n3115 & n5582 ) ;
  assign n5584 = n5583 ^ n4445 ^ n1016 ;
  assign n5587 = n5586 ^ n5584 ^ n2929 ;
  assign n5579 = ( n726 & n1967 ) | ( n726 & n3052 ) | ( n1967 & n3052 ) ;
  assign n5580 = n5579 ^ n4123 ^ n1738 ;
  assign n5577 = n3303 ^ n2593 ^ n281 ;
  assign n5578 = ( ~x51 & n4098 ) | ( ~x51 & n5577 ) | ( n4098 & n5577 ) ;
  assign n5588 = n5587 ^ n5580 ^ n5578 ;
  assign n5591 = n5590 ^ n5588 ^ n899 ;
  assign n5592 = n1303 ^ n1166 ^ x36 ;
  assign n5593 = ( ~n1069 & n2859 ) | ( ~n1069 & n5592 ) | ( n2859 & n5592 ) ;
  assign n5594 = ( ~n965 & n2054 ) | ( ~n965 & n2504 ) | ( n2054 & n2504 ) ;
  assign n5595 = n2686 ^ n1630 ^ n942 ;
  assign n5596 = n5414 ^ n3100 ^ n1902 ;
  assign n5597 = ( n358 & n5595 ) | ( n358 & n5596 ) | ( n5595 & n5596 ) ;
  assign n5598 = ( n1991 & ~n5594 ) | ( n1991 & n5597 ) | ( ~n5594 & n5597 ) ;
  assign n5599 = ( n4047 & n5593 ) | ( n4047 & ~n5598 ) | ( n5593 & ~n5598 ) ;
  assign n5600 = n3566 ^ n3029 ^ n1843 ;
  assign n5601 = ( ~n834 & n1110 ) | ( ~n834 & n5600 ) | ( n1110 & n5600 ) ;
  assign n5602 = n5601 ^ n5405 ^ n791 ;
  assign n5603 = n3818 ^ n2408 ^ n1019 ;
  assign n5604 = ( ~n173 & n1916 ) | ( ~n173 & n3000 ) | ( n1916 & n3000 ) ;
  assign n5605 = ( n2621 & n4212 ) | ( n2621 & n5604 ) | ( n4212 & n5604 ) ;
  assign n5606 = ( n4219 & n5603 ) | ( n4219 & n5605 ) | ( n5603 & n5605 ) ;
  assign n5608 = ( n457 & ~n916 ) | ( n457 & n1744 ) | ( ~n916 & n1744 ) ;
  assign n5609 = ( n2365 & ~n4659 ) | ( n2365 & n5608 ) | ( ~n4659 & n5608 ) ;
  assign n5610 = n5609 ^ n3177 ^ n1727 ;
  assign n5607 = ( n2413 & ~n4447 ) | ( n2413 & n4717 ) | ( ~n4447 & n4717 ) ;
  assign n5611 = n5610 ^ n5607 ^ n5207 ;
  assign n5617 = ( ~n2300 & n3137 ) | ( ~n2300 & n3494 ) | ( n3137 & n3494 ) ;
  assign n5618 = n5617 ^ n3116 ^ n1430 ;
  assign n5615 = ( n1770 & n1932 ) | ( n1770 & n3808 ) | ( n1932 & n3808 ) ;
  assign n5616 = n5615 ^ n3537 ^ n2045 ;
  assign n5612 = ( n523 & ~n2870 ) | ( n523 & n4279 ) | ( ~n2870 & n4279 ) ;
  assign n5613 = ( n1792 & ~n4318 ) | ( n1792 & n4326 ) | ( ~n4318 & n4326 ) ;
  assign n5614 = ( x20 & n5612 ) | ( x20 & n5613 ) | ( n5612 & n5613 ) ;
  assign n5619 = n5618 ^ n5616 ^ n5614 ;
  assign n5623 = n5136 ^ n1893 ^ n987 ;
  assign n5624 = n5623 ^ n4891 ^ n1049 ;
  assign n5625 = ( n395 & n1404 ) | ( n395 & n3272 ) | ( n1404 & n3272 ) ;
  assign n5626 = ( ~n2308 & n5624 ) | ( ~n2308 & n5625 ) | ( n5624 & n5625 ) ;
  assign n5627 = n5626 ^ n1486 ^ n192 ;
  assign n5628 = ( n699 & n3944 ) | ( n699 & n5627 ) | ( n3944 & n5627 ) ;
  assign n5621 = ( n1486 & ~n1703 ) | ( n1486 & n5120 ) | ( ~n1703 & n5120 ) ;
  assign n5620 = ( n365 & n652 ) | ( n365 & n5312 ) | ( n652 & n5312 ) ;
  assign n5622 = n5621 ^ n5620 ^ n2438 ;
  assign n5629 = n5628 ^ n5622 ^ n898 ;
  assign n5630 = ( ~n2603 & n4345 ) | ( ~n2603 & n5274 ) | ( n4345 & n5274 ) ;
  assign n5631 = ( ~x74 & n2064 ) | ( ~x74 & n3933 ) | ( n2064 & n3933 ) ;
  assign n5632 = n5449 ^ n1436 ^ x39 ;
  assign n5633 = ( ~n464 & n4408 ) | ( ~n464 & n5632 ) | ( n4408 & n5632 ) ;
  assign n5634 = n5583 ^ n1840 ^ x118 ;
  assign n5635 = n5634 ^ n2210 ^ n2071 ;
  assign n5636 = ( ~n313 & n5633 ) | ( ~n313 & n5635 ) | ( n5633 & n5635 ) ;
  assign n5637 = ( n5630 & n5631 ) | ( n5630 & ~n5636 ) | ( n5631 & ~n5636 ) ;
  assign n5638 = ( n772 & ~n3131 ) | ( n772 & n3757 ) | ( ~n3131 & n3757 ) ;
  assign n5639 = n3240 ^ n2495 ^ x67 ;
  assign n5640 = n5023 ^ n4902 ^ n4346 ;
  assign n5641 = ( n5638 & n5639 ) | ( n5638 & ~n5640 ) | ( n5639 & ~n5640 ) ;
  assign n5642 = ( n676 & ~n2496 ) | ( n676 & n4914 ) | ( ~n2496 & n4914 ) ;
  assign n5644 = ( ~n1274 & n2993 ) | ( ~n1274 & n5023 ) | ( n2993 & n5023 ) ;
  assign n5643 = ( ~n338 & n412 ) | ( ~n338 & n3517 ) | ( n412 & n3517 ) ;
  assign n5645 = n5644 ^ n5643 ^ n4541 ;
  assign n5646 = ( ~n2831 & n5642 ) | ( ~n2831 & n5645 ) | ( n5642 & n5645 ) ;
  assign n5647 = ( n152 & ~n229 ) | ( n152 & n1468 ) | ( ~n229 & n1468 ) ;
  assign n5648 = ( n2654 & ~n3636 ) | ( n2654 & n5647 ) | ( ~n3636 & n5647 ) ;
  assign n5652 = ( x4 & n485 ) | ( x4 & n3946 ) | ( n485 & n3946 ) ;
  assign n5649 = ( n472 & n1197 ) | ( n472 & n5377 ) | ( n1197 & n5377 ) ;
  assign n5650 = n5649 ^ n1180 ^ n867 ;
  assign n5651 = ( n2254 & ~n3034 ) | ( n2254 & n5650 ) | ( ~n3034 & n5650 ) ;
  assign n5653 = n5652 ^ n5651 ^ n4316 ;
  assign n5654 = n5653 ^ n2954 ^ n1536 ;
  assign n5655 = ( n2203 & n5648 ) | ( n2203 & n5654 ) | ( n5648 & n5654 ) ;
  assign n5656 = ( ~n3252 & n5646 ) | ( ~n3252 & n5655 ) | ( n5646 & n5655 ) ;
  assign n5657 = ( n285 & ~n2782 ) | ( n285 & n2793 ) | ( ~n2782 & n2793 ) ;
  assign n5658 = n5657 ^ n5273 ^ n525 ;
  assign n5664 = n3506 ^ n891 ^ n614 ;
  assign n5659 = n2757 ^ n1904 ^ n215 ;
  assign n5660 = ( n387 & n607 ) | ( n387 & n975 ) | ( n607 & n975 ) ;
  assign n5661 = ( ~n257 & n287 ) | ( ~n257 & n4439 ) | ( n287 & n4439 ) ;
  assign n5662 = ( ~n1925 & n5660 ) | ( ~n1925 & n5661 ) | ( n5660 & n5661 ) ;
  assign n5663 = ( n2228 & n5659 ) | ( n2228 & n5662 ) | ( n5659 & n5662 ) ;
  assign n5665 = n5664 ^ n5663 ^ n2372 ;
  assign n5666 = ( n323 & ~n3857 ) | ( n323 & n5665 ) | ( ~n3857 & n5665 ) ;
  assign n5667 = ( n519 & n5343 ) | ( n519 & ~n5666 ) | ( n5343 & ~n5666 ) ;
  assign n5670 = ( n2659 & ~n3585 ) | ( n2659 & n4199 ) | ( ~n3585 & n4199 ) ;
  assign n5668 = n4582 ^ n4069 ^ n483 ;
  assign n5669 = n5668 ^ n4901 ^ n3050 ;
  assign n5671 = n5670 ^ n5669 ^ n5212 ;
  assign n5672 = n5671 ^ n4755 ^ n2545 ;
  assign n5673 = ( n2034 & n3779 ) | ( n2034 & n5165 ) | ( n3779 & n5165 ) ;
  assign n5684 = n1937 ^ n1496 ^ n1112 ;
  assign n5685 = ( n1815 & n5426 ) | ( n1815 & n5684 ) | ( n5426 & n5684 ) ;
  assign n5686 = ( n2330 & n3839 ) | ( n2330 & n5685 ) | ( n3839 & n5685 ) ;
  assign n5682 = n864 ^ n795 ^ n618 ;
  assign n5683 = ( n1183 & ~n1879 ) | ( n1183 & n5682 ) | ( ~n1879 & n5682 ) ;
  assign n5687 = n5686 ^ n5683 ^ n4181 ;
  assign n5680 = n3892 ^ n3782 ^ n3397 ;
  assign n5676 = ( ~x51 & n1483 ) | ( ~x51 & n3413 ) | ( n1483 & n3413 ) ;
  assign n5677 = ( n580 & n2968 ) | ( n580 & ~n5676 ) | ( n2968 & ~n5676 ) ;
  assign n5678 = ( ~n469 & n2286 ) | ( ~n469 & n5677 ) | ( n2286 & n5677 ) ;
  assign n5674 = ( n486 & n3606 ) | ( n486 & n5392 ) | ( n3606 & n5392 ) ;
  assign n5675 = n5674 ^ n4799 ^ n159 ;
  assign n5679 = n5678 ^ n5675 ^ n4257 ;
  assign n5681 = n5680 ^ n5679 ^ n2575 ;
  assign n5688 = n5687 ^ n5681 ^ n1632 ;
  assign n5689 = ( n2535 & n3433 ) | ( n2535 & n4079 ) | ( n3433 & n4079 ) ;
  assign n5690 = ( ~n1839 & n3394 ) | ( ~n1839 & n4078 ) | ( n3394 & n4078 ) ;
  assign n5691 = n5690 ^ n5592 ^ n557 ;
  assign n5692 = ( n2621 & n5689 ) | ( n2621 & n5691 ) | ( n5689 & n5691 ) ;
  assign n5693 = ( ~n195 & n3600 ) | ( ~n195 & n5692 ) | ( n3600 & n5692 ) ;
  assign n5695 = ( n2007 & n3313 ) | ( n2007 & n5259 ) | ( n3313 & n5259 ) ;
  assign n5696 = ( ~n2389 & n3341 ) | ( ~n2389 & n5695 ) | ( n3341 & n5695 ) ;
  assign n5694 = n5308 ^ n2976 ^ n1426 ;
  assign n5697 = n5696 ^ n5694 ^ n4538 ;
  assign n5706 = n3019 ^ n1448 ^ n1218 ;
  assign n5704 = ( n658 & ~n959 ) | ( n658 & n4084 ) | ( ~n959 & n4084 ) ;
  assign n5705 = n5704 ^ n2375 ^ n1287 ;
  assign n5698 = n4705 ^ n873 ^ n272 ;
  assign n5699 = ( n511 & ~n4084 ) | ( n511 & n5698 ) | ( ~n4084 & n5698 ) ;
  assign n5700 = n3627 ^ n1903 ^ n1434 ;
  assign n5701 = ( x119 & n1145 ) | ( x119 & n5700 ) | ( n1145 & n5700 ) ;
  assign n5702 = ( x18 & n4327 ) | ( x18 & ~n5701 ) | ( n4327 & ~n5701 ) ;
  assign n5703 = ( ~n3800 & n5699 ) | ( ~n3800 & n5702 ) | ( n5699 & n5702 ) ;
  assign n5707 = n5706 ^ n5705 ^ n5703 ;
  assign n5709 = ( n979 & n1355 ) | ( n979 & ~n3198 ) | ( n1355 & ~n3198 ) ;
  assign n5708 = n4506 ^ n993 ^ x103 ;
  assign n5710 = n5709 ^ n5708 ^ n716 ;
  assign n5711 = ( n419 & ~n5411 ) | ( n419 & n5710 ) | ( ~n5411 & n5710 ) ;
  assign n5715 = n5312 ^ n4891 ^ n3961 ;
  assign n5716 = ( ~n1130 & n2871 ) | ( ~n1130 & n5715 ) | ( n2871 & n5715 ) ;
  assign n5712 = n3912 ^ n3180 ^ n547 ;
  assign n5713 = ( ~x83 & n3296 ) | ( ~x83 & n5712 ) | ( n3296 & n5712 ) ;
  assign n5714 = n5713 ^ n4081 ^ n3620 ;
  assign n5717 = n5716 ^ n5714 ^ n4091 ;
  assign n5727 = n2409 ^ n2157 ^ n327 ;
  assign n5732 = n2719 ^ n780 ^ n418 ;
  assign n5733 = n5732 ^ n4014 ^ n3812 ;
  assign n5728 = ( n614 & n1408 ) | ( n614 & ~n2303 ) | ( n1408 & ~n2303 ) ;
  assign n5729 = ( n2472 & ~n3463 ) | ( n2472 & n4026 ) | ( ~n3463 & n4026 ) ;
  assign n5730 = n5729 ^ n1699 ^ n524 ;
  assign n5731 = ( n242 & n5728 ) | ( n242 & n5730 ) | ( n5728 & n5730 ) ;
  assign n5734 = n5733 ^ n5731 ^ n3688 ;
  assign n5735 = ( ~n980 & n5727 ) | ( ~n980 & n5734 ) | ( n5727 & n5734 ) ;
  assign n5736 = n5735 ^ n4799 ^ x52 ;
  assign n5719 = n3331 ^ n3167 ^ n263 ;
  assign n5720 = ( n2262 & n4410 ) | ( n2262 & ~n5719 ) | ( n4410 & ~n5719 ) ;
  assign n5724 = n1688 ^ n1316 ^ n265 ;
  assign n5721 = ( ~n630 & n698 ) | ( ~n630 & n3062 ) | ( n698 & n3062 ) ;
  assign n5722 = ( n1208 & n1854 ) | ( n1208 & n5721 ) | ( n1854 & n5721 ) ;
  assign n5723 = n5722 ^ n5152 ^ n3964 ;
  assign n5725 = n5724 ^ n5723 ^ x16 ;
  assign n5726 = ( n4257 & n5720 ) | ( n4257 & n5725 ) | ( n5720 & n5725 ) ;
  assign n5737 = n5736 ^ n5726 ^ n5477 ;
  assign n5718 = ( ~n2230 & n2914 ) | ( ~n2230 & n3735 ) | ( n2914 & n3735 ) ;
  assign n5738 = n5737 ^ n5718 ^ n327 ;
  assign n5739 = n742 ^ n262 ^ x65 ;
  assign n5740 = n5739 ^ n5024 ^ n2006 ;
  assign n5741 = ( n957 & n3000 ) | ( n957 & n4061 ) | ( n3000 & n4061 ) ;
  assign n5742 = ( x115 & n464 ) | ( x115 & ~n4369 ) | ( n464 & ~n4369 ) ;
  assign n5743 = n5742 ^ n2753 ^ n2208 ;
  assign n5744 = n5743 ^ n1580 ^ n138 ;
  assign n5745 = n2525 ^ n2097 ^ n1650 ;
  assign n5746 = n5745 ^ n3139 ^ n1197 ;
  assign n5747 = ( n1874 & n5744 ) | ( n1874 & ~n5746 ) | ( n5744 & ~n5746 ) ;
  assign n5748 = ( n5004 & n5741 ) | ( n5004 & n5747 ) | ( n5741 & n5747 ) ;
  assign n5749 = ( n2619 & n4930 ) | ( n2619 & ~n5748 ) | ( n4930 & ~n5748 ) ;
  assign n5750 = ( n1303 & n3557 ) | ( n1303 & ~n5749 ) | ( n3557 & ~n5749 ) ;
  assign n5751 = ( ~n944 & n5740 ) | ( ~n944 & n5750 ) | ( n5740 & n5750 ) ;
  assign n5752 = ( n4540 & ~n5456 ) | ( n4540 & n5751 ) | ( ~n5456 & n5751 ) ;
  assign n5753 = ( n2091 & n2310 ) | ( n2091 & ~n3051 ) | ( n2310 & ~n3051 ) ;
  assign n5754 = n4731 ^ n1844 ^ n1214 ;
  assign n5755 = ( n3720 & ~n5253 ) | ( n3720 & n5754 ) | ( ~n5253 & n5754 ) ;
  assign n5756 = ( ~n1837 & n5753 ) | ( ~n1837 & n5755 ) | ( n5753 & n5755 ) ;
  assign n5757 = ( n1298 & n3631 ) | ( n1298 & ~n4439 ) | ( n3631 & ~n4439 ) ;
  assign n5758 = ( n328 & n2688 ) | ( n328 & ~n5757 ) | ( n2688 & ~n5757 ) ;
  assign n5759 = n3972 ^ n3437 ^ n1387 ;
  assign n5760 = ( n1546 & n5758 ) | ( n1546 & n5759 ) | ( n5758 & n5759 ) ;
  assign n5763 = ( n381 & ~n2529 ) | ( n381 & n5743 ) | ( ~n2529 & n5743 ) ;
  assign n5761 = ( ~n410 & n962 ) | ( ~n410 & n1839 ) | ( n962 & n1839 ) ;
  assign n5762 = ( n2749 & n3305 ) | ( n2749 & n5761 ) | ( n3305 & n5761 ) ;
  assign n5764 = n5763 ^ n5762 ^ n3414 ;
  assign n5765 = n4364 ^ n4030 ^ n2274 ;
  assign n5766 = n5765 ^ n2538 ^ n453 ;
  assign n5767 = ( n464 & n535 ) | ( n464 & ~n3641 ) | ( n535 & ~n3641 ) ;
  assign n5768 = n5767 ^ n3551 ^ n2377 ;
  assign n5769 = n5451 ^ n5031 ^ n3220 ;
  assign n5770 = n5769 ^ n3991 ^ n705 ;
  assign n5771 = n5770 ^ n3589 ^ n1146 ;
  assign n5772 = ( n2058 & n5768 ) | ( n2058 & ~n5771 ) | ( n5768 & ~n5771 ) ;
  assign n5773 = ( n1072 & n1238 ) | ( n1072 & ~n2677 ) | ( n1238 & ~n2677 ) ;
  assign n5774 = ( n2127 & n3317 ) | ( n2127 & ~n5773 ) | ( n3317 & ~n5773 ) ;
  assign n5775 = ( n1196 & n1801 ) | ( n1196 & n3179 ) | ( n1801 & n3179 ) ;
  assign n5776 = ( n2878 & n2924 ) | ( n2878 & ~n5775 ) | ( n2924 & ~n5775 ) ;
  assign n5777 = ( n724 & ~n5774 ) | ( n724 & n5776 ) | ( ~n5774 & n5776 ) ;
  assign n5778 = ( ~n5766 & n5772 ) | ( ~n5766 & n5777 ) | ( n5772 & n5777 ) ;
  assign n5781 = ( n1441 & n1715 ) | ( n1441 & ~n4526 ) | ( n1715 & ~n4526 ) ;
  assign n5782 = n2030 ^ n815 ^ n315 ;
  assign n5783 = ( ~n5091 & n5781 ) | ( ~n5091 & n5782 ) | ( n5781 & n5782 ) ;
  assign n5787 = n3204 ^ n2579 ^ n853 ;
  assign n5784 = ( n3372 & n3401 ) | ( n3372 & ~n4561 ) | ( n3401 & ~n4561 ) ;
  assign n5785 = ( n2075 & ~n5700 ) | ( n2075 & n5784 ) | ( ~n5700 & n5784 ) ;
  assign n5786 = ( n2628 & n4600 ) | ( n2628 & ~n5785 ) | ( n4600 & ~n5785 ) ;
  assign n5788 = n5787 ^ n5786 ^ n3198 ;
  assign n5789 = ( n5368 & n5783 ) | ( n5368 & ~n5788 ) | ( n5783 & ~n5788 ) ;
  assign n5779 = ( ~n1639 & n1650 ) | ( ~n1639 & n4340 ) | ( n1650 & n4340 ) ;
  assign n5780 = n5779 ^ n4047 ^ n440 ;
  assign n5790 = n5789 ^ n5780 ^ n408 ;
  assign n5810 = ( n1361 & ~n1694 ) | ( n1361 & n2422 ) | ( ~n1694 & n2422 ) ;
  assign n5811 = ( n694 & n3691 ) | ( n694 & ~n5810 ) | ( n3691 & ~n5810 ) ;
  assign n5795 = ( n2434 & n2462 ) | ( n2434 & n2518 ) | ( n2462 & n2518 ) ;
  assign n5800 = n871 ^ n636 ^ n261 ;
  assign n5801 = ( n3107 & ~n3742 ) | ( n3107 & n5800 ) | ( ~n3742 & n5800 ) ;
  assign n5802 = n5801 ^ n4783 ^ n1456 ;
  assign n5797 = n5097 ^ n3911 ^ n343 ;
  assign n5798 = ( n2759 & n5020 ) | ( n2759 & ~n5797 ) | ( n5020 & ~n5797 ) ;
  assign n5799 = n5798 ^ n3151 ^ n407 ;
  assign n5796 = n866 ^ n660 ^ n195 ;
  assign n5803 = n5802 ^ n5799 ^ n5796 ;
  assign n5804 = ( n2412 & n5795 ) | ( n2412 & n5803 ) | ( n5795 & n5803 ) ;
  assign n5805 = ( n1007 & n3116 ) | ( n1007 & n3918 ) | ( n3116 & n3918 ) ;
  assign n5806 = n5805 ^ n1731 ^ n905 ;
  assign n5807 = n3729 ^ n1429 ^ n1345 ;
  assign n5808 = ( n1990 & n3638 ) | ( n1990 & n5807 ) | ( n3638 & n5807 ) ;
  assign n5809 = ( n5804 & n5806 ) | ( n5804 & ~n5808 ) | ( n5806 & ~n5808 ) ;
  assign n5791 = ( ~n1343 & n2597 ) | ( ~n1343 & n3837 ) | ( n2597 & n3837 ) ;
  assign n5792 = n5791 ^ n3628 ^ n1765 ;
  assign n5793 = ( n1791 & ~n4508 ) | ( n1791 & n5792 ) | ( ~n4508 & n5792 ) ;
  assign n5794 = n5793 ^ n5605 ^ n219 ;
  assign n5812 = n5811 ^ n5809 ^ n5794 ;
  assign n5813 = n3844 ^ n2296 ^ n2009 ;
  assign n5814 = n4976 ^ n4827 ^ n1036 ;
  assign n5815 = ( ~n3818 & n5034 ) | ( ~n3818 & n5814 ) | ( n5034 & n5814 ) ;
  assign n5816 = ( n220 & n3876 ) | ( n220 & n4973 ) | ( n3876 & n4973 ) ;
  assign n5817 = n5816 ^ n5017 ^ n4466 ;
  assign n5818 = n5783 ^ n4054 ^ n1953 ;
  assign n5819 = n5818 ^ n4569 ^ n185 ;
  assign n5820 = ( n5815 & n5817 ) | ( n5815 & ~n5819 ) | ( n5817 & ~n5819 ) ;
  assign n5821 = ( n2671 & n5813 ) | ( n2671 & n5820 ) | ( n5813 & n5820 ) ;
  assign n5826 = n4966 ^ n2929 ^ n2321 ;
  assign n5822 = n1942 ^ n859 ^ n570 ;
  assign n5823 = n4312 ^ n1554 ^ n1220 ;
  assign n5824 = n5823 ^ n2490 ^ x52 ;
  assign n5825 = ( n4996 & n5822 ) | ( n4996 & n5824 ) | ( n5822 & n5824 ) ;
  assign n5827 = n5826 ^ n5825 ^ n4256 ;
  assign n5828 = ( n3352 & ~n5174 ) | ( n3352 & n5827 ) | ( ~n5174 & n5827 ) ;
  assign n5851 = n2269 ^ n2016 ^ n1455 ;
  assign n5849 = ( n652 & n2680 ) | ( n652 & n5210 ) | ( n2680 & n5210 ) ;
  assign n5847 = n4082 ^ n2957 ^ n2202 ;
  assign n5840 = ( ~n1201 & n1387 ) | ( ~n1201 & n2373 ) | ( n1387 & n2373 ) ;
  assign n5842 = ( n144 & n506 ) | ( n144 & ~n1186 ) | ( n506 & ~n1186 ) ;
  assign n5843 = n5842 ^ n3042 ^ n2804 ;
  assign n5841 = ( n326 & ~n581 ) | ( n326 & n2044 ) | ( ~n581 & n2044 ) ;
  assign n5844 = n5843 ^ n5841 ^ n4385 ;
  assign n5829 = ( x109 & ~n581 ) | ( x109 & n5170 ) | ( ~n581 & n5170 ) ;
  assign n5830 = n5829 ^ n4495 ^ n1874 ;
  assign n5845 = n5830 ^ n5441 ^ n4732 ;
  assign n5846 = ( n5840 & n5844 ) | ( n5840 & n5845 ) | ( n5844 & n5845 ) ;
  assign n5848 = n5847 ^ n5846 ^ n3568 ;
  assign n5850 = n5849 ^ n5848 ^ n1932 ;
  assign n5836 = ( ~n1080 & n4428 ) | ( ~n1080 & n5482 ) | ( n4428 & n5482 ) ;
  assign n5835 = ( n610 & n1719 ) | ( n610 & n4053 ) | ( n1719 & n4053 ) ;
  assign n5837 = n5836 ^ n5835 ^ n289 ;
  assign n5838 = ( x67 & n4602 ) | ( x67 & n5837 ) | ( n4602 & n5837 ) ;
  assign n5832 = n2322 ^ n1659 ^ n180 ;
  assign n5833 = ( ~n5511 & n5567 ) | ( ~n5511 & n5832 ) | ( n5567 & n5832 ) ;
  assign n5831 = n5830 ^ n4634 ^ n1483 ;
  assign n5834 = n5833 ^ n5831 ^ n3283 ;
  assign n5839 = n5838 ^ n5834 ^ n4122 ;
  assign n5852 = n5851 ^ n5850 ^ n5839 ;
  assign n5853 = n2896 ^ n893 ^ x47 ;
  assign n5854 = n5853 ^ n3525 ^ n822 ;
  assign n5855 = n5854 ^ n4444 ^ n2998 ;
  assign n5856 = ( ~n1323 & n5502 ) | ( ~n1323 & n5855 ) | ( n5502 & n5855 ) ;
  assign n5870 = n3881 ^ n1716 ^ n1396 ;
  assign n5871 = n5870 ^ n2439 ^ n301 ;
  assign n5868 = n3644 ^ n753 ^ x35 ;
  assign n5869 = ( n924 & ~n3682 ) | ( n924 & n5868 ) | ( ~n3682 & n5868 ) ;
  assign n5866 = n4680 ^ n1087 ^ n849 ;
  assign n5863 = ( ~n252 & n2243 ) | ( ~n252 & n4364 ) | ( n2243 & n4364 ) ;
  assign n5864 = n5863 ^ n3126 ^ n904 ;
  assign n5861 = ( x77 & n289 ) | ( x77 & n1374 ) | ( n289 & n1374 ) ;
  assign n5862 = n5861 ^ n3889 ^ n649 ;
  assign n5858 = n2408 ^ n844 ^ n493 ;
  assign n5859 = n5858 ^ n2255 ^ n1449 ;
  assign n5857 = ( n540 & ~n1206 ) | ( n540 & n2849 ) | ( ~n1206 & n2849 ) ;
  assign n5860 = n5859 ^ n5857 ^ n5199 ;
  assign n5865 = n5864 ^ n5862 ^ n5860 ;
  assign n5867 = n5866 ^ n5865 ^ n777 ;
  assign n5872 = n5871 ^ n5869 ^ n5867 ;
  assign n5873 = ( n1886 & ~n5500 ) | ( n1886 & n5872 ) | ( ~n5500 & n5872 ) ;
  assign n5874 = n5873 ^ n3455 ^ n1814 ;
  assign n5875 = ( n2712 & n5856 ) | ( n2712 & ~n5874 ) | ( n5856 & ~n5874 ) ;
  assign n5876 = n1164 ^ n782 ^ n674 ;
  assign n5877 = n5876 ^ n5375 ^ n4808 ;
  assign n5878 = ( n1207 & n2791 ) | ( n1207 & ~n4120 ) | ( n2791 & ~n4120 ) ;
  assign n5880 = ( n840 & ~n1157 ) | ( n840 & n3807 ) | ( ~n1157 & n3807 ) ;
  assign n5879 = ( n1100 & n2897 ) | ( n1100 & ~n3478 ) | ( n2897 & ~n3478 ) ;
  assign n5881 = n5880 ^ n5879 ^ n2620 ;
  assign n5882 = n5881 ^ n4104 ^ n2856 ;
  assign n5883 = n5725 ^ n1076 ^ n796 ;
  assign n5884 = ( n1202 & ~n1446 ) | ( n1202 & n3648 ) | ( ~n1446 & n3648 ) ;
  assign n5885 = n5884 ^ n2020 ^ n616 ;
  assign n5886 = n5885 ^ n4260 ^ n2910 ;
  assign n5887 = ( ~n4605 & n5883 ) | ( ~n4605 & n5886 ) | ( n5883 & n5886 ) ;
  assign n5888 = ( n816 & n5882 ) | ( n816 & ~n5887 ) | ( n5882 & ~n5887 ) ;
  assign n5893 = n5859 ^ n4495 ^ n3957 ;
  assign n5889 = n5851 ^ n5417 ^ n3139 ;
  assign n5890 = ( n1689 & n3922 ) | ( n1689 & n4832 ) | ( n3922 & n4832 ) ;
  assign n5891 = ( ~n2414 & n5889 ) | ( ~n2414 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5892 = n5891 ^ n4240 ^ n1601 ;
  assign n5894 = n5893 ^ n5892 ^ n180 ;
  assign n5904 = n5210 ^ n3186 ^ n2308 ;
  assign n5902 = ( n802 & ~n2186 ) | ( n802 & n4419 ) | ( ~n2186 & n4419 ) ;
  assign n5903 = n5902 ^ n1796 ^ n780 ;
  assign n5899 = n3207 ^ n2779 ^ n288 ;
  assign n5900 = n5899 ^ n5434 ^ n2428 ;
  assign n5895 = ( n392 & ~n2151 ) | ( n392 & n3999 ) | ( ~n2151 & n3999 ) ;
  assign n5896 = n4953 ^ n2200 ^ n818 ;
  assign n5897 = ( n1978 & n5895 ) | ( n1978 & ~n5896 ) | ( n5895 & ~n5896 ) ;
  assign n5898 = n5897 ^ n3190 ^ n2900 ;
  assign n5901 = n5900 ^ n5898 ^ n210 ;
  assign n5905 = n5904 ^ n5903 ^ n5901 ;
  assign n5906 = ( n2072 & ~n3151 ) | ( n2072 & n5905 ) | ( ~n3151 & n5905 ) ;
  assign n5907 = n5906 ^ n602 ^ n131 ;
  assign n5909 = n4453 ^ n1247 ^ n862 ;
  assign n5908 = n4518 ^ n3585 ^ n2832 ;
  assign n5910 = n5909 ^ n5908 ^ n699 ;
  assign n5913 = ( ~n784 & n1018 ) | ( ~n784 & n3043 ) | ( n1018 & n3043 ) ;
  assign n5911 = n3174 ^ n1672 ^ n520 ;
  assign n5912 = n5911 ^ n1925 ^ x118 ;
  assign n5914 = n5913 ^ n5912 ^ n1943 ;
  assign n5915 = n3691 ^ n2483 ^ n2160 ;
  assign n5916 = ( ~n743 & n5914 ) | ( ~n743 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5917 = n5916 ^ n1912 ^ x106 ;
  assign n5918 = n4080 ^ n3211 ^ n1776 ;
  assign n5919 = ( ~x119 & n1844 ) | ( ~x119 & n2218 ) | ( n1844 & n2218 ) ;
  assign n5920 = ( n3417 & n5918 ) | ( n3417 & ~n5919 ) | ( n5918 & ~n5919 ) ;
  assign n5921 = ( n504 & ~n1539 ) | ( n504 & n2116 ) | ( ~n1539 & n2116 ) ;
  assign n5922 = ( n197 & n1179 ) | ( n197 & ~n5921 ) | ( n1179 & ~n5921 ) ;
  assign n5923 = n4310 ^ n2047 ^ n1331 ;
  assign n5924 = ( n5208 & ~n5922 ) | ( n5208 & n5923 ) | ( ~n5922 & n5923 ) ;
  assign n5925 = ( n562 & n5920 ) | ( n562 & ~n5924 ) | ( n5920 & ~n5924 ) ;
  assign n5926 = n4080 ^ n1551 ^ n369 ;
  assign n5927 = ( ~n354 & n1525 ) | ( ~n354 & n5926 ) | ( n1525 & n5926 ) ;
  assign n5928 = ( ~n2163 & n5729 ) | ( ~n2163 & n5927 ) | ( n5729 & n5927 ) ;
  assign n5929 = ( n2256 & n4767 ) | ( n2256 & n5928 ) | ( n4767 & n5928 ) ;
  assign n5959 = n1707 ^ n1162 ^ n257 ;
  assign n5952 = n2778 ^ n1452 ^ n1202 ;
  assign n5953 = n5952 ^ n3182 ^ n1832 ;
  assign n5954 = n1593 ^ n984 ^ n446 ;
  assign n5955 = n5954 ^ n1706 ^ n177 ;
  assign n5956 = ( ~n5396 & n5953 ) | ( ~n5396 & n5955 ) | ( n5953 & n5955 ) ;
  assign n5957 = n5956 ^ n5728 ^ n4279 ;
  assign n5958 = n5957 ^ n4818 ^ n1767 ;
  assign n5930 = n5247 ^ n2530 ^ n486 ;
  assign n5931 = n5930 ^ n750 ^ x77 ;
  assign n5932 = ( n3452 & n4351 ) | ( n3452 & ~n5931 ) | ( n4351 & ~n5931 ) ;
  assign n5933 = n5266 ^ n359 ^ n140 ;
  assign n5948 = n5372 ^ n4257 ^ n845 ;
  assign n5949 = n5948 ^ n5177 ^ n2650 ;
  assign n5942 = n4633 ^ n4365 ^ n262 ;
  assign n5944 = ( n359 & ~n865 ) | ( n359 & n3734 ) | ( ~n865 & n3734 ) ;
  assign n5943 = ( ~n2337 & n4039 ) | ( ~n2337 & n5342 ) | ( n4039 & n5342 ) ;
  assign n5945 = n5944 ^ n5943 ^ n3840 ;
  assign n5946 = n4221 ^ n2732 ^ n819 ;
  assign n5947 = ( ~n5942 & n5945 ) | ( ~n5942 & n5946 ) | ( n5945 & n5946 ) ;
  assign n5937 = ( n235 & ~n434 ) | ( n235 & n2087 ) | ( ~n434 & n2087 ) ;
  assign n5938 = ( n835 & n1302 ) | ( n835 & n5937 ) | ( n1302 & n5937 ) ;
  assign n5939 = n5938 ^ n2575 ^ n2314 ;
  assign n5940 = ( n3742 & n5126 ) | ( n3742 & n5939 ) | ( n5126 & n5939 ) ;
  assign n5934 = n5624 ^ n2322 ^ n264 ;
  assign n5935 = ( ~n3588 & n3861 ) | ( ~n3588 & n5934 ) | ( n3861 & n5934 ) ;
  assign n5936 = n5935 ^ n4790 ^ n4238 ;
  assign n5941 = n5940 ^ n5936 ^ n3974 ;
  assign n5950 = n5949 ^ n5947 ^ n5941 ;
  assign n5951 = ( ~n5932 & n5933 ) | ( ~n5932 & n5950 ) | ( n5933 & n5950 ) ;
  assign n5960 = n5959 ^ n5958 ^ n5951 ;
  assign n5961 = ( x11 & n730 ) | ( x11 & n5367 ) | ( n730 & n5367 ) ;
  assign n5962 = n5961 ^ n3095 ^ n1224 ;
  assign n5963 = n4499 ^ n4380 ^ n353 ;
  assign n5964 = ( n5617 & n5962 ) | ( n5617 & ~n5963 ) | ( n5962 & ~n5963 ) ;
  assign n5966 = n1259 ^ n635 ^ n493 ;
  assign n5965 = ( ~n502 & n954 ) | ( ~n502 & n5739 ) | ( n954 & n5739 ) ;
  assign n5967 = n5966 ^ n5965 ^ n1951 ;
  assign n5975 = ( ~n1647 & n3002 ) | ( ~n1647 & n4143 ) | ( n3002 & n4143 ) ;
  assign n5972 = n5657 ^ n2001 ^ n660 ;
  assign n5973 = n5972 ^ n1685 ^ n1318 ;
  assign n5974 = ( n2140 & ~n4927 ) | ( n2140 & n5973 ) | ( ~n4927 & n5973 ) ;
  assign n5968 = n1232 ^ n752 ^ n421 ;
  assign n5969 = ( ~n435 & n2864 ) | ( ~n435 & n5968 ) | ( n2864 & n5968 ) ;
  assign n5970 = n5969 ^ n3404 ^ n3332 ;
  assign n5971 = n5970 ^ n5322 ^ n743 ;
  assign n5976 = n5975 ^ n5974 ^ n5971 ;
  assign n5977 = ( n134 & ~n5967 ) | ( n134 & n5976 ) | ( ~n5967 & n5976 ) ;
  assign n5983 = ( n3523 & n3552 ) | ( n3523 & ~n5169 ) | ( n3552 & ~n5169 ) ;
  assign n5979 = n3048 ^ n2465 ^ n544 ;
  assign n5980 = n5979 ^ n775 ^ n696 ;
  assign n5978 = n4544 ^ n3022 ^ n2903 ;
  assign n5981 = n5980 ^ n5978 ^ n4628 ;
  assign n5982 = n5981 ^ n5327 ^ n1989 ;
  assign n5984 = n5983 ^ n5982 ^ n1642 ;
  assign n5985 = ( ~n1646 & n3363 ) | ( ~n1646 & n5984 ) | ( n3363 & n5984 ) ;
  assign n5986 = ( ~n227 & n1224 ) | ( ~n227 & n5985 ) | ( n1224 & n5985 ) ;
  assign n5991 = ( ~n326 & n717 ) | ( ~n326 & n1058 ) | ( n717 & n1058 ) ;
  assign n5987 = ( x71 & ~n1072 ) | ( x71 & n1435 ) | ( ~n1072 & n1435 ) ;
  assign n5988 = n5987 ^ n4678 ^ n1336 ;
  assign n5989 = n5988 ^ n1426 ^ n1273 ;
  assign n5990 = ( n921 & n2234 ) | ( n921 & n5989 ) | ( n2234 & n5989 ) ;
  assign n5992 = n5991 ^ n5990 ^ n4082 ;
  assign n5993 = n3730 ^ n2566 ^ n1935 ;
  assign n5994 = ( ~n1473 & n3045 ) | ( ~n1473 & n5993 ) | ( n3045 & n5993 ) ;
  assign n5995 = n5994 ^ n2465 ^ n1338 ;
  assign n5999 = n2214 ^ n1707 ^ n1083 ;
  assign n5997 = n4274 ^ n3231 ^ n1077 ;
  assign n5996 = ( n638 & ~n899 ) | ( n638 & n2517 ) | ( ~n899 & n2517 ) ;
  assign n5998 = n5997 ^ n5996 ^ n3081 ;
  assign n6000 = n5999 ^ n5998 ^ n2406 ;
  assign n6005 = ( ~n768 & n3035 ) | ( ~n768 & n5489 ) | ( n3035 & n5489 ) ;
  assign n6001 = ( n2268 & ~n3614 ) | ( n2268 & n5861 ) | ( ~n3614 & n5861 ) ;
  assign n6002 = ( n669 & n696 ) | ( n669 & n2097 ) | ( n696 & n2097 ) ;
  assign n6003 = n6002 ^ n713 ^ n309 ;
  assign n6004 = ( n3446 & n6001 ) | ( n3446 & ~n6003 ) | ( n6001 & ~n6003 ) ;
  assign n6006 = n6005 ^ n6004 ^ n1103 ;
  assign n6007 = ( n435 & ~n987 ) | ( n435 & n1354 ) | ( ~n987 & n1354 ) ;
  assign n6008 = n3061 ^ n2368 ^ n706 ;
  assign n6009 = n6008 ^ n4083 ^ n669 ;
  assign n6010 = ( ~n3835 & n3978 ) | ( ~n3835 & n6009 ) | ( n3978 & n6009 ) ;
  assign n6023 = ( x120 & n568 ) | ( x120 & n1101 ) | ( n568 & n1101 ) ;
  assign n6024 = ( n1006 & n3088 ) | ( n1006 & ~n6023 ) | ( n3088 & ~n6023 ) ;
  assign n6025 = ( ~n1350 & n3341 ) | ( ~n1350 & n6024 ) | ( n3341 & n6024 ) ;
  assign n6026 = n6025 ^ n5408 ^ n1316 ;
  assign n6011 = ( n658 & n2297 ) | ( n658 & n3567 ) | ( n2297 & n3567 ) ;
  assign n6015 = ( n1454 & ~n1471 ) | ( n1454 & n2419 ) | ( ~n1471 & n2419 ) ;
  assign n6012 = n4604 ^ n714 ^ n264 ;
  assign n6013 = ( n1499 & n1950 ) | ( n1499 & n6012 ) | ( n1950 & n6012 ) ;
  assign n6014 = n6013 ^ n3601 ^ n652 ;
  assign n6016 = n6015 ^ n6014 ^ n1176 ;
  assign n6017 = ( ~x78 & n443 ) | ( ~x78 & n1156 ) | ( n443 & n1156 ) ;
  assign n6018 = n6017 ^ n940 ^ n191 ;
  assign n6019 = ( n712 & n1460 ) | ( n712 & ~n6018 ) | ( n1460 & ~n6018 ) ;
  assign n6020 = ( ~n987 & n2023 ) | ( ~n987 & n6019 ) | ( n2023 & n6019 ) ;
  assign n6021 = ( n951 & ~n4865 ) | ( n951 & n6020 ) | ( ~n4865 & n6020 ) ;
  assign n6022 = ( n6011 & n6016 ) | ( n6011 & n6021 ) | ( n6016 & n6021 ) ;
  assign n6027 = n6026 ^ n6022 ^ n5479 ;
  assign n6045 = n4091 ^ n3587 ^ n3150 ;
  assign n6048 = ( n1561 & n1621 ) | ( n1561 & n2150 ) | ( n1621 & n2150 ) ;
  assign n6046 = ( n1450 & n1570 ) | ( n1450 & ~n2247 ) | ( n1570 & ~n2247 ) ;
  assign n6047 = ( n734 & ~n1334 ) | ( n734 & n6046 ) | ( ~n1334 & n6046 ) ;
  assign n6049 = n6048 ^ n6047 ^ n463 ;
  assign n6050 = ( n2914 & n6045 ) | ( n2914 & n6049 ) | ( n6045 & n6049 ) ;
  assign n6043 = n2218 ^ n404 ^ n135 ;
  assign n6042 = n3688 ^ n3005 ^ x114 ;
  assign n6044 = n6043 ^ n6042 ^ x120 ;
  assign n6051 = n6050 ^ n6044 ^ n4798 ;
  assign n6036 = ( n1089 & n1507 ) | ( n1089 & n4798 ) | ( n1507 & n4798 ) ;
  assign n6037 = ( n660 & n1143 ) | ( n660 & ~n2550 ) | ( n1143 & ~n2550 ) ;
  assign n6038 = ( n4809 & n6036 ) | ( n4809 & n6037 ) | ( n6036 & n6037 ) ;
  assign n6039 = ( n2023 & n4847 ) | ( n2023 & ~n6038 ) | ( n4847 & ~n6038 ) ;
  assign n6032 = n3359 ^ n3203 ^ n533 ;
  assign n6033 = ( n3084 & n5570 ) | ( n3084 & n6032 ) | ( n5570 & n6032 ) ;
  assign n6034 = n6033 ^ n5254 ^ n3677 ;
  assign n6028 = ( n1115 & n2438 ) | ( n1115 & ~n3152 ) | ( n2438 & ~n3152 ) ;
  assign n6029 = ( n4087 & ~n4710 ) | ( n4087 & n5190 ) | ( ~n4710 & n5190 ) ;
  assign n6030 = n6029 ^ n5734 ^ n1935 ;
  assign n6031 = ( ~n340 & n6028 ) | ( ~n340 & n6030 ) | ( n6028 & n6030 ) ;
  assign n6035 = n6034 ^ n6031 ^ n5713 ;
  assign n6040 = n6039 ^ n6035 ^ n2996 ;
  assign n6041 = n6040 ^ n4513 ^ n617 ;
  assign n6052 = n6051 ^ n6041 ^ n4866 ;
  assign n6060 = ( ~n2206 & n5062 ) | ( ~n2206 & n5263 ) | ( n5062 & n5263 ) ;
  assign n6056 = ( n311 & ~n1212 ) | ( n311 & n5326 ) | ( ~n1212 & n5326 ) ;
  assign n6054 = ( n451 & ~n641 ) | ( n451 & n5203 ) | ( ~n641 & n5203 ) ;
  assign n6055 = ( n402 & ~n979 ) | ( n402 & n6054 ) | ( ~n979 & n6054 ) ;
  assign n6057 = n6056 ^ n6055 ^ n869 ;
  assign n6058 = n6057 ^ n2023 ^ n800 ;
  assign n6053 = ( ~n227 & n2577 ) | ( ~n227 & n2702 ) | ( n2577 & n2702 ) ;
  assign n6059 = n6058 ^ n6053 ^ n286 ;
  assign n6061 = n6060 ^ n6059 ^ n2890 ;
  assign n6068 = ( ~x20 & n1179 ) | ( ~x20 & n1783 ) | ( n1179 & n1783 ) ;
  assign n6069 = n6068 ^ n3701 ^ n932 ;
  assign n6070 = n6069 ^ n4748 ^ n2957 ;
  assign n6071 = n6070 ^ n4722 ^ n3396 ;
  assign n6065 = ( n1832 & n4525 ) | ( n1832 & n5741 ) | ( n4525 & n5741 ) ;
  assign n6066 = n6065 ^ n4307 ^ n172 ;
  assign n6072 = n6071 ^ n6066 ^ n4842 ;
  assign n6063 = ( ~n1766 & n2008 ) | ( ~n1766 & n3043 ) | ( n2008 & n3043 ) ;
  assign n6062 = n4833 ^ n4108 ^ n1762 ;
  assign n6064 = n6063 ^ n6062 ^ n255 ;
  assign n6067 = n6066 ^ n6064 ^ n5383 ;
  assign n6073 = n6072 ^ n6067 ^ n1200 ;
  assign n6074 = n4145 ^ n2674 ^ n2355 ;
  assign n6075 = ( n805 & n1124 ) | ( n805 & ~n5134 ) | ( n1124 & ~n5134 ) ;
  assign n6076 = ( n2323 & ~n2528 ) | ( n2323 & n6075 ) | ( ~n2528 & n6075 ) ;
  assign n6077 = ( ~n3852 & n4659 ) | ( ~n3852 & n6076 ) | ( n4659 & n6076 ) ;
  assign n6078 = ( n2711 & n6074 ) | ( n2711 & ~n6077 ) | ( n6074 & ~n6077 ) ;
  assign n6085 = ( n690 & n1661 ) | ( n690 & ~n5259 ) | ( n1661 & ~n5259 ) ;
  assign n6086 = ( n412 & ~n5539 ) | ( n412 & n6085 ) | ( ~n5539 & n6085 ) ;
  assign n6082 = ( n607 & ~n1103 ) | ( n607 & n3634 ) | ( ~n1103 & n3634 ) ;
  assign n6083 = n6082 ^ n3835 ^ n2059 ;
  assign n6084 = ( n610 & n6028 ) | ( n610 & n6083 ) | ( n6028 & n6083 ) ;
  assign n6087 = n6086 ^ n6084 ^ n5480 ;
  assign n6079 = n4873 ^ n1284 ^ n278 ;
  assign n6080 = n6079 ^ n372 ^ n337 ;
  assign n6081 = n6080 ^ n6005 ^ n4300 ;
  assign n6088 = n6087 ^ n6081 ^ n3007 ;
  assign n6089 = n6088 ^ n5255 ^ n3690 ;
  assign n6090 = n6089 ^ n4388 ^ n1039 ;
  assign n6091 = ( ~n3893 & n4455 ) | ( ~n3893 & n6090 ) | ( n4455 & n6090 ) ;
  assign n6092 = ( ~n969 & n2454 ) | ( ~n969 & n2627 ) | ( n2454 & n2627 ) ;
  assign n6093 = n6092 ^ n2910 ^ n643 ;
  assign n6094 = n2228 ^ n717 ^ n502 ;
  assign n6095 = n6094 ^ n3861 ^ n2111 ;
  assign n6096 = ( n5454 & n6093 ) | ( n5454 & n6095 ) | ( n6093 & n6095 ) ;
  assign n6106 = n5449 ^ n3450 ^ n2649 ;
  assign n6107 = ( n202 & ~n1960 ) | ( n202 & n6106 ) | ( ~n1960 & n6106 ) ;
  assign n6108 = n6107 ^ n5396 ^ n1329 ;
  assign n6109 = ( ~n4087 & n4927 ) | ( ~n4087 & n6108 ) | ( n4927 & n6108 ) ;
  assign n6110 = n6109 ^ n5186 ^ n4361 ;
  assign n6097 = n3475 ^ n2837 ^ n1315 ;
  assign n6098 = n4583 ^ n3939 ^ n3652 ;
  assign n6099 = ( n2677 & n5009 ) | ( n2677 & ~n6098 ) | ( n5009 & ~n6098 ) ;
  assign n6100 = ( ~n157 & n2124 ) | ( ~n157 & n2311 ) | ( n2124 & n2311 ) ;
  assign n6101 = n5784 ^ n2758 ^ n367 ;
  assign n6102 = ( ~n1550 & n2248 ) | ( ~n1550 & n3502 ) | ( n2248 & n3502 ) ;
  assign n6103 = ( ~n420 & n6101 ) | ( ~n420 & n6102 ) | ( n6101 & n6102 ) ;
  assign n6104 = ( ~n5026 & n6100 ) | ( ~n5026 & n6103 ) | ( n6100 & n6103 ) ;
  assign n6105 = ( n6097 & ~n6099 ) | ( n6097 & n6104 ) | ( ~n6099 & n6104 ) ;
  assign n6111 = n6110 ^ n6105 ^ n6001 ;
  assign n6112 = ( n290 & n6096 ) | ( n290 & n6111 ) | ( n6096 & n6111 ) ;
  assign n6113 = ( n2234 & ~n3540 ) | ( n2234 & n4384 ) | ( ~n3540 & n4384 ) ;
  assign n6114 = ( n155 & n1659 ) | ( n155 & n6113 ) | ( n1659 & n6113 ) ;
  assign n6115 = ( n2204 & ~n3349 ) | ( n2204 & n6114 ) | ( ~n3349 & n6114 ) ;
  assign n6119 = ( n584 & ~n5304 ) | ( n584 & n5939 ) | ( ~n5304 & n5939 ) ;
  assign n6120 = n3878 ^ n1261 ^ n650 ;
  assign n6121 = ( n181 & n2395 ) | ( n181 & ~n6120 ) | ( n2395 & ~n6120 ) ;
  assign n6122 = ( n1680 & n6119 ) | ( n1680 & ~n6121 ) | ( n6119 & ~n6121 ) ;
  assign n6117 = ( ~n1667 & n1679 ) | ( ~n1667 & n3505 ) | ( n1679 & n3505 ) ;
  assign n6116 = ( n624 & ~n2383 ) | ( n624 & n3563 ) | ( ~n2383 & n3563 ) ;
  assign n6118 = n6117 ^ n6116 ^ n5162 ;
  assign n6123 = n6122 ^ n6118 ^ n3699 ;
  assign n6124 = ( ~x121 & n4226 ) | ( ~x121 & n5171 ) | ( n4226 & n5171 ) ;
  assign n6125 = ( n2400 & n5861 ) | ( n2400 & n6124 ) | ( n5861 & n6124 ) ;
  assign n6126 = ( n3071 & n4101 ) | ( n3071 & ~n6125 ) | ( n4101 & ~n6125 ) ;
  assign n6129 = n3911 ^ n3843 ^ n365 ;
  assign n6127 = ( ~n934 & n2300 ) | ( ~n934 & n3950 ) | ( n2300 & n3950 ) ;
  assign n6128 = n6127 ^ n1349 ^ n852 ;
  assign n6130 = n6129 ^ n6128 ^ n5801 ;
  assign n6131 = ( n1730 & n2781 ) | ( n1730 & n6130 ) | ( n2781 & n6130 ) ;
  assign n6132 = n5031 ^ n1589 ^ n643 ;
  assign n6133 = ( ~x126 & n2050 ) | ( ~x126 & n6132 ) | ( n2050 & n6132 ) ;
  assign n6134 = ( ~n1503 & n2256 ) | ( ~n1503 & n6133 ) | ( n2256 & n6133 ) ;
  assign n6135 = n6134 ^ n4967 ^ n527 ;
  assign n6136 = n6135 ^ n3391 ^ n204 ;
  assign n6137 = n6136 ^ n5308 ^ n2467 ;
  assign n6138 = ( n6126 & ~n6131 ) | ( n6126 & n6137 ) | ( ~n6131 & n6137 ) ;
  assign n6139 = ( n6115 & n6123 ) | ( n6115 & ~n6138 ) | ( n6123 & ~n6138 ) ;
  assign n6140 = ( n401 & n1306 ) | ( n401 & ~n2323 ) | ( n1306 & ~n2323 ) ;
  assign n6141 = n6140 ^ n1651 ^ n443 ;
  assign n6142 = n6141 ^ n4216 ^ n1915 ;
  assign n6143 = n6142 ^ n3791 ^ x0 ;
  assign n6144 = ( n2067 & n3247 ) | ( n2067 & n6143 ) | ( n3247 & n6143 ) ;
  assign n6150 = n2133 ^ n1708 ^ n133 ;
  assign n6145 = ( ~n272 & n506 ) | ( ~n272 & n1128 ) | ( n506 & n1128 ) ;
  assign n6146 = ( n1028 & n2773 ) | ( n1028 & ~n4401 ) | ( n2773 & ~n4401 ) ;
  assign n6147 = ( n4627 & n6145 ) | ( n4627 & n6146 ) | ( n6145 & n6146 ) ;
  assign n6148 = n6147 ^ n2259 ^ n1696 ;
  assign n6149 = ( ~n301 & n5661 ) | ( ~n301 & n6148 ) | ( n5661 & n6148 ) ;
  assign n6151 = n6150 ^ n6149 ^ n1624 ;
  assign n6152 = ( n132 & n300 ) | ( n132 & n2222 ) | ( n300 & n2222 ) ;
  assign n6176 = ( ~n765 & n1266 ) | ( ~n765 & n3614 ) | ( n1266 & n3614 ) ;
  assign n6175 = ( n328 & n1664 ) | ( n328 & n1928 ) | ( n1664 & n1928 ) ;
  assign n6173 = n2498 ^ n1197 ^ n464 ;
  assign n6174 = ( ~n4318 & n5994 ) | ( ~n4318 & n6173 ) | ( n5994 & n6173 ) ;
  assign n6177 = n6176 ^ n6175 ^ n6174 ;
  assign n6168 = n5968 ^ n3426 ^ n2531 ;
  assign n6169 = n1265 ^ n357 ^ n300 ;
  assign n6170 = ( n810 & ~n6168 ) | ( n810 & n6169 ) | ( ~n6168 & n6169 ) ;
  assign n6171 = n6170 ^ n4831 ^ n334 ;
  assign n6172 = n6171 ^ n871 ^ x66 ;
  assign n6159 = n3516 ^ n2730 ^ n881 ;
  assign n6160 = ( n846 & n1336 ) | ( n846 & ~n3379 ) | ( n1336 & ~n3379 ) ;
  assign n6161 = n6160 ^ n3869 ^ n3182 ;
  assign n6162 = n1411 ^ n913 ^ n678 ;
  assign n6163 = ( n3577 & ~n3781 ) | ( n3577 & n5009 ) | ( ~n3781 & n5009 ) ;
  assign n6164 = ( n236 & n6162 ) | ( n236 & n6163 ) | ( n6162 & n6163 ) ;
  assign n6165 = ( n6159 & n6161 ) | ( n6159 & ~n6164 ) | ( n6161 & ~n6164 ) ;
  assign n6166 = n6165 ^ n3628 ^ n2049 ;
  assign n6156 = ( ~n421 & n755 ) | ( ~n421 & n862 ) | ( n755 & n862 ) ;
  assign n6157 = n6156 ^ n2733 ^ n1043 ;
  assign n6155 = n2162 ^ n158 ^ n157 ;
  assign n6153 = ( n1094 & ~n1950 ) | ( n1094 & n5008 ) | ( ~n1950 & n5008 ) ;
  assign n6154 = ( n3009 & n3225 ) | ( n3009 & ~n6153 ) | ( n3225 & ~n6153 ) ;
  assign n6158 = n6157 ^ n6155 ^ n6154 ;
  assign n6167 = n6166 ^ n6158 ^ n1611 ;
  assign n6178 = n6177 ^ n6172 ^ n6167 ;
  assign n6179 = n6178 ^ n5291 ^ n285 ;
  assign n6180 = ( n2968 & n5264 ) | ( n2968 & ~n6179 ) | ( n5264 & ~n6179 ) ;
  assign n6181 = ( n507 & ~n1288 ) | ( n507 & n1708 ) | ( ~n1288 & n1708 ) ;
  assign n6182 = ( n3147 & ~n4656 ) | ( n3147 & n6181 ) | ( ~n4656 & n6181 ) ;
  assign n6183 = n2757 ^ n1767 ^ n1179 ;
  assign n6184 = n5594 ^ n4638 ^ n242 ;
  assign n6187 = ( ~n836 & n2549 ) | ( ~n836 & n3342 ) | ( n2549 & n3342 ) ;
  assign n6188 = ( n952 & n4158 ) | ( n952 & n6187 ) | ( n4158 & n6187 ) ;
  assign n6189 = ( n896 & n2356 ) | ( n896 & ~n6188 ) | ( n2356 & ~n6188 ) ;
  assign n6190 = n6189 ^ n1115 ^ n488 ;
  assign n6186 = ( n227 & n2816 ) | ( n227 & n3416 ) | ( n2816 & n3416 ) ;
  assign n6185 = n2708 ^ n1443 ^ n873 ;
  assign n6191 = n6190 ^ n6186 ^ n6185 ;
  assign n6192 = ( n6183 & n6184 ) | ( n6183 & n6191 ) | ( n6184 & n6191 ) ;
  assign n6193 = ( n2565 & n3394 ) | ( n2565 & n4215 ) | ( n3394 & n4215 ) ;
  assign n6194 = n6193 ^ n5135 ^ n1765 ;
  assign n6195 = n3381 ^ n1680 ^ n703 ;
  assign n6196 = ( ~n1836 & n5230 ) | ( ~n1836 & n6195 ) | ( n5230 & n6195 ) ;
  assign n6197 = ( n1612 & n4504 ) | ( n1612 & n6196 ) | ( n4504 & n6196 ) ;
  assign n6198 = ( n1039 & n6194 ) | ( n1039 & ~n6197 ) | ( n6194 & ~n6197 ) ;
  assign n6199 = ( n544 & n2509 ) | ( n544 & n4459 ) | ( n2509 & n4459 ) ;
  assign n6200 = n4402 ^ n1507 ^ n849 ;
  assign n6201 = n6200 ^ n5132 ^ n1899 ;
  assign n6202 = n2892 ^ n744 ^ n702 ;
  assign n6203 = n6202 ^ n5714 ^ n1594 ;
  assign n6204 = ( n1310 & n6201 ) | ( n1310 & ~n6203 ) | ( n6201 & ~n6203 ) ;
  assign n6205 = ( ~n4992 & n6199 ) | ( ~n4992 & n6204 ) | ( n6199 & n6204 ) ;
  assign n6206 = ( n2702 & ~n2826 ) | ( n2702 & n5039 ) | ( ~n2826 & n5039 ) ;
  assign n6207 = ( n1320 & ~n1659 ) | ( n1320 & n1973 ) | ( ~n1659 & n1973 ) ;
  assign n6208 = n812 ^ n149 ^ x85 ;
  assign n6209 = n6208 ^ n3338 ^ n690 ;
  assign n6210 = n6209 ^ n1795 ^ n822 ;
  assign n6211 = ( n1950 & ~n2634 ) | ( n1950 & n5784 ) | ( ~n2634 & n5784 ) ;
  assign n6212 = n6211 ^ n1493 ^ n911 ;
  assign n6213 = n6212 ^ n4793 ^ n4527 ;
  assign n6214 = ( x1 & n6210 ) | ( x1 & n6213 ) | ( n6210 & n6213 ) ;
  assign n6215 = ( n223 & ~n723 ) | ( n223 & n1253 ) | ( ~n723 & n1253 ) ;
  assign n6216 = ( n1363 & ~n6214 ) | ( n1363 & n6215 ) | ( ~n6214 & n6215 ) ;
  assign n6217 = ( n940 & n3242 ) | ( n940 & n3977 ) | ( n3242 & n3977 ) ;
  assign n6218 = n1074 ^ n970 ^ n873 ;
  assign n6219 = n6218 ^ n1498 ^ n762 ;
  assign n6220 = n6219 ^ n3686 ^ n316 ;
  assign n6221 = ( n1568 & n2355 ) | ( n1568 & n2377 ) | ( n2355 & n2377 ) ;
  assign n6222 = n2639 ^ n1974 ^ n1363 ;
  assign n6223 = n6222 ^ n4370 ^ n2156 ;
  assign n6224 = ( n2174 & ~n6221 ) | ( n2174 & n6223 ) | ( ~n6221 & n6223 ) ;
  assign n6225 = ( n1442 & ~n3016 ) | ( n1442 & n6224 ) | ( ~n3016 & n6224 ) ;
  assign n6226 = n2702 ^ n2616 ^ n783 ;
  assign n6227 = n5899 ^ n5037 ^ n3123 ;
  assign n6228 = n3392 ^ n2724 ^ n590 ;
  assign n6229 = ( ~n6226 & n6227 ) | ( ~n6226 & n6228 ) | ( n6227 & n6228 ) ;
  assign n6230 = ( n6220 & ~n6225 ) | ( n6220 & n6229 ) | ( ~n6225 & n6229 ) ;
  assign n6231 = ( n3987 & n6217 ) | ( n3987 & ~n6230 ) | ( n6217 & ~n6230 ) ;
  assign n6232 = ( n6207 & n6216 ) | ( n6207 & ~n6231 ) | ( n6216 & ~n6231 ) ;
  assign n6233 = ( ~n5209 & n6206 ) | ( ~n5209 & n6232 ) | ( n6206 & n6232 ) ;
  assign n6241 = n3265 ^ n1306 ^ n714 ;
  assign n6237 = ( n404 & n1959 ) | ( n404 & n2489 ) | ( n1959 & n2489 ) ;
  assign n6238 = ( x124 & n3426 ) | ( x124 & n4665 ) | ( n3426 & n4665 ) ;
  assign n6239 = ( n2385 & n6237 ) | ( n2385 & n6238 ) | ( n6237 & n6238 ) ;
  assign n6235 = n5293 ^ n2583 ^ n1151 ;
  assign n6234 = n4903 ^ n1691 ^ n1485 ;
  assign n6236 = n6235 ^ n6234 ^ n4626 ;
  assign n6240 = n6239 ^ n6236 ^ n5477 ;
  assign n6242 = n6241 ^ n6240 ^ n1708 ;
  assign n6245 = ( n764 & n3893 ) | ( n764 & n5785 ) | ( n3893 & n5785 ) ;
  assign n6246 = n6245 ^ n960 ^ n140 ;
  assign n6243 = n968 ^ n811 ^ n243 ;
  assign n6244 = ( n2396 & ~n5016 ) | ( n2396 & n6243 ) | ( ~n5016 & n6243 ) ;
  assign n6247 = n6246 ^ n6244 ^ n1751 ;
  assign n6248 = ( n1523 & n4214 ) | ( n1523 & n6247 ) | ( n4214 & n6247 ) ;
  assign n6249 = ( ~n2433 & n6015 ) | ( ~n2433 & n6248 ) | ( n6015 & n6248 ) ;
  assign n6250 = n2806 ^ n769 ^ n176 ;
  assign n6251 = n5544 ^ n3161 ^ n2948 ;
  assign n6253 = n6113 ^ n3660 ^ n834 ;
  assign n6252 = ( ~n2607 & n5178 ) | ( ~n2607 & n5547 ) | ( n5178 & n5547 ) ;
  assign n6254 = n6253 ^ n6252 ^ n2281 ;
  assign n6255 = ( n6250 & n6251 ) | ( n6250 & ~n6254 ) | ( n6251 & ~n6254 ) ;
  assign n6256 = n6048 ^ n2124 ^ n375 ;
  assign n6257 = n4793 ^ n2852 ^ n798 ;
  assign n6258 = ( n1680 & n1709 ) | ( n1680 & n6257 ) | ( n1709 & n6257 ) ;
  assign n6259 = n2516 ^ n785 ^ n758 ;
  assign n6260 = ( n2920 & ~n3698 ) | ( n2920 & n6259 ) | ( ~n3698 & n6259 ) ;
  assign n6261 = ( n6256 & ~n6258 ) | ( n6256 & n6260 ) | ( ~n6258 & n6260 ) ;
  assign n6283 = ( n1373 & ~n4269 ) | ( n1373 & n4571 ) | ( ~n4269 & n4571 ) ;
  assign n6284 = ( n1337 & n3181 ) | ( n1337 & ~n6283 ) | ( n3181 & ~n6283 ) ;
  assign n6285 = n6284 ^ n4064 ^ n1404 ;
  assign n6280 = n3585 ^ n2397 ^ n1718 ;
  assign n6281 = n6280 ^ n3553 ^ x96 ;
  assign n6282 = ( n2381 & n2782 ) | ( n2381 & n6281 ) | ( n2782 & n6281 ) ;
  assign n6277 = ( ~x26 & n1508 ) | ( ~x26 & n2409 ) | ( n1508 & n2409 ) ;
  assign n6276 = ( n1098 & n1142 ) | ( n1098 & n2419 ) | ( n1142 & n2419 ) ;
  assign n6278 = n6277 ^ n6276 ^ n5408 ;
  assign n6268 = ( ~n215 & n2687 ) | ( ~n215 & n5450 ) | ( n2687 & n5450 ) ;
  assign n6270 = ( n3130 & n3451 ) | ( n3130 & n4927 ) | ( n3451 & n4927 ) ;
  assign n6271 = n6270 ^ n4452 ^ n3893 ;
  assign n6272 = n6271 ^ n5881 ^ n2355 ;
  assign n6269 = ( n827 & n4280 ) | ( n827 & n5918 ) | ( n4280 & n5918 ) ;
  assign n6273 = n6272 ^ n6269 ^ n6048 ;
  assign n6274 = ( n2849 & n6268 ) | ( n2849 & ~n6273 ) | ( n6268 & ~n6273 ) ;
  assign n6275 = n6274 ^ n2830 ^ n1236 ;
  assign n6265 = n3866 ^ n2461 ^ n806 ;
  assign n6266 = n6265 ^ n1201 ^ n529 ;
  assign n6262 = ( n272 & ~n3446 ) | ( n272 & n3542 ) | ( ~n3446 & n3542 ) ;
  assign n6263 = ( n952 & ~n5100 ) | ( n952 & n6262 ) | ( ~n5100 & n6262 ) ;
  assign n6264 = ( n2908 & n5459 ) | ( n2908 & ~n6263 ) | ( n5459 & ~n6263 ) ;
  assign n6267 = n6266 ^ n6264 ^ n3581 ;
  assign n6279 = n6278 ^ n6275 ^ n6267 ;
  assign n6286 = n6285 ^ n6282 ^ n6279 ;
  assign n6287 = ( ~n1033 & n2617 ) | ( ~n1033 & n3723 ) | ( n2617 & n3723 ) ;
  assign n6288 = n6287 ^ n5112 ^ n178 ;
  assign n6289 = ( ~n1400 & n3989 ) | ( ~n1400 & n6288 ) | ( n3989 & n6288 ) ;
  assign n6290 = ( n1894 & ~n4758 ) | ( n1894 & n6289 ) | ( ~n4758 & n6289 ) ;
  assign n6294 = n890 ^ n724 ^ n292 ;
  assign n6291 = ( n1354 & n1731 ) | ( n1354 & ~n1855 ) | ( n1731 & ~n1855 ) ;
  assign n6292 = n2355 ^ n1593 ^ x92 ;
  assign n6293 = ( n444 & n6291 ) | ( n444 & ~n6292 ) | ( n6291 & ~n6292 ) ;
  assign n6295 = n6294 ^ n6293 ^ n5100 ;
  assign n6296 = ( n1488 & n2545 ) | ( n1488 & n6295 ) | ( n2545 & n6295 ) ;
  assign n6297 = ( n3752 & ~n5510 ) | ( n3752 & n6296 ) | ( ~n5510 & n6296 ) ;
  assign n6298 = ( ~n436 & n2656 ) | ( ~n436 & n6297 ) | ( n2656 & n6297 ) ;
  assign n6299 = n6298 ^ n3834 ^ n2404 ;
  assign n6300 = ( n697 & n935 ) | ( n697 & n1977 ) | ( n935 & n1977 ) ;
  assign n6301 = ( n535 & ~n3069 ) | ( n535 & n6300 ) | ( ~n3069 & n6300 ) ;
  assign n6302 = n6301 ^ n2110 ^ n716 ;
  assign n6303 = n3691 ^ n1144 ^ n764 ;
  assign n6304 = ( n593 & n4756 ) | ( n593 & ~n6303 ) | ( n4756 & ~n6303 ) ;
  assign n6305 = ( n1259 & n6302 ) | ( n1259 & ~n6304 ) | ( n6302 & ~n6304 ) ;
  assign n6306 = n6305 ^ n4113 ^ n1917 ;
  assign n6307 = ( n651 & n6299 ) | ( n651 & ~n6306 ) | ( n6299 & ~n6306 ) ;
  assign n6308 = n3574 ^ n2813 ^ n1689 ;
  assign n6309 = ( n1883 & n2569 ) | ( n1883 & n4053 ) | ( n2569 & n4053 ) ;
  assign n6310 = n4797 ^ n3752 ^ n373 ;
  assign n6311 = ( n2462 & n3929 ) | ( n2462 & ~n6310 ) | ( n3929 & ~n6310 ) ;
  assign n6312 = ( n6308 & ~n6309 ) | ( n6308 & n6311 ) | ( ~n6309 & n6311 ) ;
  assign n6313 = n3999 ^ n703 ^ n428 ;
  assign n6314 = ( ~n341 & n2840 ) | ( ~n341 & n6313 ) | ( n2840 & n6313 ) ;
  assign n6315 = ( ~n1016 & n2569 ) | ( ~n1016 & n3219 ) | ( n2569 & n3219 ) ;
  assign n6316 = n6315 ^ n573 ^ n178 ;
  assign n6317 = ( ~x18 & n1912 ) | ( ~x18 & n6316 ) | ( n1912 & n6316 ) ;
  assign n6318 = n6317 ^ n5038 ^ n2164 ;
  assign n6319 = n5706 ^ n4308 ^ n531 ;
  assign n6320 = n1631 ^ n904 ^ n652 ;
  assign n6321 = n5970 ^ n5067 ^ n2948 ;
  assign n6322 = ( n1859 & n6320 ) | ( n1859 & ~n6321 ) | ( n6320 & ~n6321 ) ;
  assign n6323 = ( n2701 & n3380 ) | ( n2701 & n3770 ) | ( n3380 & n3770 ) ;
  assign n6327 = n3896 ^ n3814 ^ n900 ;
  assign n6328 = n6327 ^ n5926 ^ n5575 ;
  assign n6324 = ( n406 & n726 ) | ( n406 & ~n4235 ) | ( n726 & ~n4235 ) ;
  assign n6325 = ( ~n2226 & n3785 ) | ( ~n2226 & n6324 ) | ( n3785 & n6324 ) ;
  assign n6326 = n6325 ^ n5373 ^ n2125 ;
  assign n6329 = n6328 ^ n6326 ^ n1880 ;
  assign n6330 = ( n622 & ~n6323 ) | ( n622 & n6329 ) | ( ~n6323 & n6329 ) ;
  assign n6331 = ( n6319 & ~n6322 ) | ( n6319 & n6330 ) | ( ~n6322 & n6330 ) ;
  assign n6332 = ( ~n6314 & n6318 ) | ( ~n6314 & n6331 ) | ( n6318 & n6331 ) ;
  assign n6333 = n2502 ^ n1695 ^ n271 ;
  assign n6334 = n6333 ^ n2152 ^ n1654 ;
  assign n6335 = ( n1261 & ~n2464 ) | ( n1261 & n6334 ) | ( ~n2464 & n6334 ) ;
  assign n6336 = n6335 ^ n4293 ^ n162 ;
  assign n6337 = ( n565 & n1754 ) | ( n565 & n6336 ) | ( n1754 & n6336 ) ;
  assign n6343 = ( n1079 & n2116 ) | ( n1079 & n2697 ) | ( n2116 & n2697 ) ;
  assign n6344 = ( n1241 & n3713 ) | ( n1241 & ~n6343 ) | ( n3713 & ~n6343 ) ;
  assign n6345 = ( ~n635 & n3584 ) | ( ~n635 & n6344 ) | ( n3584 & n6344 ) ;
  assign n6346 = ( ~n2881 & n5401 ) | ( ~n2881 & n6345 ) | ( n5401 & n6345 ) ;
  assign n6340 = ( n330 & n344 ) | ( n330 & ~n501 ) | ( n344 & ~n501 ) ;
  assign n6338 = n6276 ^ n3704 ^ n805 ;
  assign n6339 = ( ~n2850 & n3672 ) | ( ~n2850 & n6338 ) | ( n3672 & n6338 ) ;
  assign n6341 = n6340 ^ n6339 ^ n4350 ;
  assign n6342 = n6341 ^ n5762 ^ n465 ;
  assign n6347 = n6346 ^ n6342 ^ n1401 ;
  assign n6348 = ( ~n2809 & n6337 ) | ( ~n2809 & n6347 ) | ( n6337 & n6347 ) ;
  assign n6349 = ( n6312 & ~n6332 ) | ( n6312 & n6348 ) | ( ~n6332 & n6348 ) ;
  assign n6350 = n3284 ^ n2896 ^ n599 ;
  assign n6351 = ( n1136 & ~n3016 ) | ( n1136 & n6350 ) | ( ~n3016 & n6350 ) ;
  assign n6352 = n5213 ^ n4191 ^ n630 ;
  assign n6353 = ( n4141 & n6351 ) | ( n4141 & n6352 ) | ( n6351 & n6352 ) ;
  assign n6354 = n6353 ^ n3388 ^ n1654 ;
  assign n6356 = n2046 ^ n1478 ^ n784 ;
  assign n6357 = ( n1724 & n5586 ) | ( n1724 & ~n6356 ) | ( n5586 & ~n6356 ) ;
  assign n6358 = n6357 ^ n3323 ^ n2089 ;
  assign n6359 = ( x112 & n1929 ) | ( x112 & ~n6358 ) | ( n1929 & ~n6358 ) ;
  assign n6360 = n4700 ^ n3051 ^ n1814 ;
  assign n6361 = n6360 ^ n5243 ^ n3897 ;
  assign n6362 = ( ~n1054 & n6359 ) | ( ~n1054 & n6361 ) | ( n6359 & n6361 ) ;
  assign n6363 = ( n834 & ~n1208 ) | ( n834 & n6362 ) | ( ~n1208 & n6362 ) ;
  assign n6355 = ( n424 & ~n4649 ) | ( n424 & n5508 ) | ( ~n4649 & n5508 ) ;
  assign n6364 = n6363 ^ n6355 ^ n580 ;
  assign n6373 = ( n437 & n2104 ) | ( n437 & n3543 ) | ( n2104 & n3543 ) ;
  assign n6371 = n5571 ^ n2766 ^ n1433 ;
  assign n6372 = ( n1437 & n4858 ) | ( n1437 & ~n6371 ) | ( n4858 & ~n6371 ) ;
  assign n6365 = n2561 ^ n2257 ^ n341 ;
  assign n6366 = n6365 ^ n3321 ^ n1371 ;
  assign n6367 = n6366 ^ n3437 ^ n2127 ;
  assign n6368 = ( n591 & ~n3438 ) | ( n591 & n5313 ) | ( ~n3438 & n5313 ) ;
  assign n6369 = n6368 ^ n3282 ^ n3115 ;
  assign n6370 = ( ~n4137 & n6367 ) | ( ~n4137 & n6369 ) | ( n6367 & n6369 ) ;
  assign n6374 = n6373 ^ n6372 ^ n6370 ;
  assign n6375 = n4501 ^ n3451 ^ n1271 ;
  assign n6376 = ( n1010 & n1310 ) | ( n1010 & ~n6375 ) | ( n1310 & ~n6375 ) ;
  assign n6377 = ( ~n2473 & n5003 ) | ( ~n2473 & n6376 ) | ( n5003 & n6376 ) ;
  assign n6378 = n6377 ^ n6239 ^ n318 ;
  assign n6380 = ( n537 & n730 ) | ( n537 & n3956 ) | ( n730 & n3956 ) ;
  assign n6381 = n4272 ^ n2768 ^ n501 ;
  assign n6382 = n6381 ^ n6058 ^ n2041 ;
  assign n6383 = ( n1492 & ~n6380 ) | ( n1492 & n6382 ) | ( ~n6380 & n6382 ) ;
  assign n6379 = n4600 ^ n2698 ^ n2468 ;
  assign n6384 = n6383 ^ n6379 ^ n4144 ;
  assign n6385 = ( n283 & n836 ) | ( n283 & ~n6384 ) | ( n836 & ~n6384 ) ;
  assign n6388 = ( n443 & ~n1105 ) | ( n443 & n4095 ) | ( ~n1105 & n4095 ) ;
  assign n6386 = n1449 ^ n1165 ^ n521 ;
  assign n6387 = ( n1829 & n2697 ) | ( n1829 & ~n6386 ) | ( n2697 & ~n6386 ) ;
  assign n6389 = n6388 ^ n6387 ^ n1371 ;
  assign n6396 = ( ~n1185 & n2753 ) | ( ~n1185 & n4493 ) | ( n2753 & n4493 ) ;
  assign n6397 = ( n1206 & ~n4588 ) | ( n1206 & n6396 ) | ( ~n4588 & n6396 ) ;
  assign n6390 = n3375 ^ n2303 ^ n1124 ;
  assign n6391 = ( ~n1432 & n3262 ) | ( ~n1432 & n6390 ) | ( n3262 & n6390 ) ;
  assign n6392 = n6063 ^ n4598 ^ n850 ;
  assign n6393 = ( n753 & n2128 ) | ( n753 & ~n3618 ) | ( n2128 & ~n3618 ) ;
  assign n6394 = n6393 ^ n2300 ^ n1166 ;
  assign n6395 = ( ~n6391 & n6392 ) | ( ~n6391 & n6394 ) | ( n6392 & n6394 ) ;
  assign n6398 = n6397 ^ n6395 ^ n6271 ;
  assign n6404 = n932 ^ n292 ^ n237 ;
  assign n6405 = ( n2132 & n2459 ) | ( n2132 & n6404 ) | ( n2459 & n6404 ) ;
  assign n6403 = n3846 ^ n3307 ^ n1986 ;
  assign n6406 = n6405 ^ n6403 ^ n1605 ;
  assign n6399 = ( ~n1383 & n1622 ) | ( ~n1383 & n4283 ) | ( n1622 & n4283 ) ;
  assign n6400 = ( ~n476 & n796 ) | ( ~n476 & n1113 ) | ( n796 & n1113 ) ;
  assign n6401 = ( n2734 & n3471 ) | ( n2734 & ~n3628 ) | ( n3471 & ~n3628 ) ;
  assign n6402 = ( n6399 & n6400 ) | ( n6399 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6407 = n6406 ^ n6402 ^ n1570 ;
  assign n6408 = n4449 ^ n4168 ^ n1510 ;
  assign n6411 = n3071 ^ n2203 ^ n268 ;
  assign n6409 = n1465 ^ n731 ^ n293 ;
  assign n6410 = ( n771 & n4043 ) | ( n771 & ~n6409 ) | ( n4043 & ~n6409 ) ;
  assign n6412 = n6411 ^ n6410 ^ n3720 ;
  assign n6413 = ( n1465 & n6408 ) | ( n1465 & n6412 ) | ( n6408 & n6412 ) ;
  assign n6414 = n1599 ^ n782 ^ n767 ;
  assign n6415 = n6414 ^ n814 ^ n183 ;
  assign n6416 = ( ~n4661 & n5390 ) | ( ~n4661 & n6415 ) | ( n5390 & n6415 ) ;
  assign n6417 = n6416 ^ n2521 ^ n1789 ;
  assign n6418 = ( x42 & ~n2149 ) | ( x42 & n6417 ) | ( ~n2149 & n6417 ) ;
  assign n6419 = ( n216 & n3524 ) | ( n216 & n6124 ) | ( n3524 & n6124 ) ;
  assign n6420 = ( n2621 & n6226 ) | ( n2621 & n6419 ) | ( n6226 & n6419 ) ;
  assign n6421 = ( n784 & ~n3907 ) | ( n784 & n6420 ) | ( ~n3907 & n6420 ) ;
  assign n6422 = n6421 ^ n6122 ^ n5997 ;
  assign n6423 = n6422 ^ n3110 ^ n2536 ;
  assign n6424 = n3960 ^ n3478 ^ n329 ;
  assign n6435 = ( n1129 & n3431 ) | ( n1129 & ~n4492 ) | ( n3431 & ~n4492 ) ;
  assign n6431 = n3077 ^ n1501 ^ n1373 ;
  assign n6432 = ( n1286 & ~n1360 ) | ( n1286 & n3519 ) | ( ~n1360 & n3519 ) ;
  assign n6433 = ( n1544 & n1576 ) | ( n1544 & n6432 ) | ( n1576 & n6432 ) ;
  assign n6434 = ( ~n1462 & n6431 ) | ( ~n1462 & n6433 ) | ( n6431 & n6433 ) ;
  assign n6425 = ( n214 & ~n2845 ) | ( n214 & n6063 ) | ( ~n2845 & n6063 ) ;
  assign n6426 = ( n2139 & ~n3009 ) | ( n2139 & n6425 ) | ( ~n3009 & n6425 ) ;
  assign n6427 = n859 ^ n486 ^ n481 ;
  assign n6428 = ( n598 & n2433 ) | ( n598 & ~n6427 ) | ( n2433 & ~n6427 ) ;
  assign n6429 = ( n1268 & ~n3675 ) | ( n1268 & n6428 ) | ( ~n3675 & n6428 ) ;
  assign n6430 = ( ~n1246 & n6426 ) | ( ~n1246 & n6429 ) | ( n6426 & n6429 ) ;
  assign n6436 = n6435 ^ n6434 ^ n6430 ;
  assign n6437 = ( n5515 & n6424 ) | ( n5515 & ~n6436 ) | ( n6424 & ~n6436 ) ;
  assign n6438 = ( n474 & n6423 ) | ( n474 & ~n6437 ) | ( n6423 & ~n6437 ) ;
  assign n6447 = n3068 ^ n2260 ^ n946 ;
  assign n6448 = ( n1386 & n4228 ) | ( n1386 & n6447 ) | ( n4228 & n6447 ) ;
  assign n6439 = ( n509 & n2111 ) | ( n509 & n2195 ) | ( n2111 & n2195 ) ;
  assign n6440 = n6439 ^ n5403 ^ n3151 ;
  assign n6441 = n6440 ^ n1313 ^ n312 ;
  assign n6443 = ( n2411 & n2732 ) | ( n2411 & ~n3891 ) | ( n2732 & ~n3891 ) ;
  assign n6444 = n6443 ^ n3442 ^ n463 ;
  assign n6442 = ( n841 & n2147 ) | ( n841 & n3700 ) | ( n2147 & n3700 ) ;
  assign n6445 = n6444 ^ n6442 ^ n1589 ;
  assign n6446 = ( n5678 & ~n6441 ) | ( n5678 & n6445 ) | ( ~n6441 & n6445 ) ;
  assign n6449 = n6448 ^ n6446 ^ n4029 ;
  assign n6450 = n2489 ^ n2181 ^ n1915 ;
  assign n6453 = ( n241 & n2550 ) | ( n241 & ~n2945 ) | ( n2550 & ~n2945 ) ;
  assign n6451 = n2132 ^ n278 ^ x77 ;
  assign n6452 = ( n1394 & ~n3844 ) | ( n1394 & n6451 ) | ( ~n3844 & n6451 ) ;
  assign n6454 = n6453 ^ n6452 ^ n866 ;
  assign n6455 = ( n4149 & n6450 ) | ( n4149 & ~n6454 ) | ( n6450 & ~n6454 ) ;
  assign n6456 = ( ~n1929 & n2797 ) | ( ~n1929 & n6291 ) | ( n2797 & n6291 ) ;
  assign n6457 = n6427 ^ n4671 ^ n748 ;
  assign n6458 = ( n1097 & ~n1137 ) | ( n1097 & n6457 ) | ( ~n1137 & n6457 ) ;
  assign n6459 = ( n1034 & n6456 ) | ( n1034 & n6458 ) | ( n6456 & n6458 ) ;
  assign n6474 = n5742 ^ n4364 ^ n1729 ;
  assign n6462 = n3516 ^ n2232 ^ n1851 ;
  assign n6463 = ( ~n1054 & n1524 ) | ( ~n1054 & n5706 ) | ( n1524 & n5706 ) ;
  assign n6464 = ( n5375 & n6462 ) | ( n5375 & n6463 ) | ( n6462 & n6463 ) ;
  assign n6465 = n6464 ^ n3824 ^ n1192 ;
  assign n6460 = n3905 ^ n2563 ^ n1499 ;
  assign n6461 = ( ~n2567 & n2872 ) | ( ~n2567 & n6460 ) | ( n2872 & n6460 ) ;
  assign n6466 = n6465 ^ n6461 ^ n2349 ;
  assign n6467 = ( x74 & n431 ) | ( x74 & ~n1945 ) | ( n431 & ~n1945 ) ;
  assign n6468 = n6467 ^ n2643 ^ n1134 ;
  assign n6469 = ( n4173 & n5235 ) | ( n4173 & n6468 ) | ( n5235 & n6468 ) ;
  assign n6470 = ( ~x72 & n2755 ) | ( ~x72 & n6469 ) | ( n2755 & n6469 ) ;
  assign n6471 = n6470 ^ n5745 ^ n1526 ;
  assign n6472 = n6471 ^ n6291 ^ n2538 ;
  assign n6473 = ( n2783 & ~n6466 ) | ( n2783 & n6472 ) | ( ~n6466 & n6472 ) ;
  assign n6475 = n6474 ^ n6473 ^ n4332 ;
  assign n6476 = ( n1108 & ~n6335 ) | ( n1108 & n6475 ) | ( ~n6335 & n6475 ) ;
  assign n6477 = ( n858 & ~n2201 ) | ( n858 & n3830 ) | ( ~n2201 & n3830 ) ;
  assign n6478 = n5536 ^ n902 ^ n723 ;
  assign n6479 = ( n2793 & n3265 ) | ( n2793 & n4607 ) | ( n3265 & n4607 ) ;
  assign n6480 = ( ~x109 & n3210 ) | ( ~x109 & n3855 ) | ( n3210 & n3855 ) ;
  assign n6481 = ( ~n806 & n1425 ) | ( ~n806 & n6480 ) | ( n1425 & n6480 ) ;
  assign n6491 = ( ~n284 & n4582 ) | ( ~n284 & n5131 ) | ( n4582 & n5131 ) ;
  assign n6492 = ( n2792 & n6175 ) | ( n2792 & n6491 ) | ( n6175 & n6491 ) ;
  assign n6482 = n3470 ^ n1759 ^ n234 ;
  assign n6483 = ( n1391 & n2937 ) | ( n1391 & ~n6482 ) | ( n2937 & ~n6482 ) ;
  assign n6484 = n6483 ^ n5919 ^ n1102 ;
  assign n6485 = ( n1942 & n2660 ) | ( n1942 & n3924 ) | ( n2660 & n3924 ) ;
  assign n6487 = ( n1776 & n3301 ) | ( n1776 & n3576 ) | ( n3301 & n3576 ) ;
  assign n6486 = ( n2762 & n2933 ) | ( n2762 & ~n5004 ) | ( n2933 & ~n5004 ) ;
  assign n6488 = n6487 ^ n6486 ^ n3755 ;
  assign n6489 = ( n5860 & n6485 ) | ( n5860 & n6488 ) | ( n6485 & n6488 ) ;
  assign n6490 = ( ~n3030 & n6484 ) | ( ~n3030 & n6489 ) | ( n6484 & n6489 ) ;
  assign n6493 = n6492 ^ n6490 ^ n856 ;
  assign n6494 = n5734 ^ n5437 ^ n244 ;
  assign n6495 = n4265 ^ n3441 ^ n2050 ;
  assign n6497 = n2821 ^ n2550 ^ n1069 ;
  assign n6496 = ( n2387 & ~n3447 ) | ( n2387 & n3620 ) | ( ~n3447 & n3620 ) ;
  assign n6498 = n6497 ^ n6496 ^ n2285 ;
  assign n6499 = n6498 ^ n3150 ^ n2149 ;
  assign n6500 = ( n1786 & n2596 ) | ( n1786 & ~n2934 ) | ( n2596 & ~n2934 ) ;
  assign n6501 = ( ~n1179 & n6499 ) | ( ~n1179 & n6500 ) | ( n6499 & n6500 ) ;
  assign n6502 = n6501 ^ n3129 ^ n293 ;
  assign n6503 = ( ~n2556 & n6495 ) | ( ~n2556 & n6502 ) | ( n6495 & n6502 ) ;
  assign n6504 = ( ~x122 & n993 ) | ( ~x122 & n1341 ) | ( n993 & n1341 ) ;
  assign n6507 = n5046 ^ n3767 ^ n579 ;
  assign n6505 = ( ~n228 & n4284 ) | ( ~n228 & n6409 ) | ( n4284 & n6409 ) ;
  assign n6506 = n6505 ^ n3616 ^ n166 ;
  assign n6508 = n6507 ^ n6506 ^ n1981 ;
  assign n6509 = n2542 ^ n1789 ^ n225 ;
  assign n6510 = n6509 ^ n2749 ^ n197 ;
  assign n6511 = ( n265 & ~n1602 ) | ( n265 & n1934 ) | ( ~n1602 & n1934 ) ;
  assign n6512 = n6511 ^ n4451 ^ n966 ;
  assign n6517 = ( n2394 & n3542 ) | ( n2394 & n4870 ) | ( n3542 & n4870 ) ;
  assign n6513 = ( n376 & n1580 ) | ( n376 & n4153 ) | ( n1580 & n4153 ) ;
  assign n6514 = ( n1594 & n3652 ) | ( n1594 & n6513 ) | ( n3652 & n6513 ) ;
  assign n6515 = n6514 ^ n6235 ^ n3544 ;
  assign n6516 = n6515 ^ n6268 ^ n5968 ;
  assign n6518 = n6517 ^ n6516 ^ n5935 ;
  assign n6519 = n6518 ^ n3571 ^ n2115 ;
  assign n6520 = ( n615 & ~n2321 ) | ( n615 & n3418 ) | ( ~n2321 & n3418 ) ;
  assign n6521 = ( n938 & n2507 ) | ( n938 & ~n4712 ) | ( n2507 & ~n4712 ) ;
  assign n6522 = ( n3206 & n6520 ) | ( n3206 & n6521 ) | ( n6520 & n6521 ) ;
  assign n6523 = ( n6512 & n6519 ) | ( n6512 & n6522 ) | ( n6519 & n6522 ) ;
  assign n6524 = ( n2186 & n3918 ) | ( n2186 & n5528 ) | ( n3918 & n5528 ) ;
  assign n6525 = n6524 ^ n3792 ^ n2273 ;
  assign n6526 = n6300 ^ n1475 ^ n266 ;
  assign n6527 = n6526 ^ n3073 ^ n270 ;
  assign n6528 = ( ~n1301 & n6525 ) | ( ~n1301 & n6527 ) | ( n6525 & n6527 ) ;
  assign n6534 = n1118 ^ n859 ^ x33 ;
  assign n6529 = ( ~n2210 & n3836 ) | ( ~n2210 & n4014 ) | ( n3836 & n4014 ) ;
  assign n6530 = ( ~n1078 & n1275 ) | ( ~n1078 & n2512 ) | ( n1275 & n2512 ) ;
  assign n6531 = ( n2501 & ~n4417 ) | ( n2501 & n6530 ) | ( ~n4417 & n6530 ) ;
  assign n6532 = ( n978 & n5628 ) | ( n978 & n6531 ) | ( n5628 & n6531 ) ;
  assign n6533 = ( ~n4853 & n6529 ) | ( ~n4853 & n6532 ) | ( n6529 & n6532 ) ;
  assign n6535 = n6534 ^ n6533 ^ n2361 ;
  assign n6536 = n4218 ^ n2182 ^ n1787 ;
  assign n6537 = n4378 ^ n1989 ^ n563 ;
  assign n6538 = n6537 ^ n4180 ^ n3842 ;
  assign n6550 = n3368 ^ n1805 ^ n473 ;
  assign n6539 = ( n610 & n2813 ) | ( n610 & n4345 ) | ( n2813 & n4345 ) ;
  assign n6540 = ( ~x82 & n399 ) | ( ~x82 & n1138 ) | ( n399 & n1138 ) ;
  assign n6541 = n2898 ^ n2784 ^ n791 ;
  assign n6542 = n6541 ^ n3316 ^ n1228 ;
  assign n6543 = n6542 ^ n1983 ^ n1666 ;
  assign n6544 = ( n1562 & n6540 ) | ( n1562 & n6543 ) | ( n6540 & n6543 ) ;
  assign n6545 = ( n1310 & n1392 ) | ( n1310 & n2674 ) | ( n1392 & n2674 ) ;
  assign n6546 = n6545 ^ n1546 ^ n1353 ;
  assign n6547 = n6546 ^ n4253 ^ n1461 ;
  assign n6548 = ( n2734 & n3900 ) | ( n2734 & n6547 ) | ( n3900 & n6547 ) ;
  assign n6549 = ( n6539 & n6544 ) | ( n6539 & n6548 ) | ( n6544 & n6548 ) ;
  assign n6551 = n6550 ^ n6549 ^ n5725 ;
  assign n6557 = ( ~n850 & n2713 ) | ( ~n850 & n2863 ) | ( n2713 & n2863 ) ;
  assign n6554 = ( n249 & n3846 ) | ( n249 & n4180 ) | ( n3846 & n4180 ) ;
  assign n6555 = ( ~n625 & n4272 ) | ( ~n625 & n6554 ) | ( n4272 & n6554 ) ;
  assign n6556 = ( n3452 & n3540 ) | ( n3452 & n6555 ) | ( n3540 & n6555 ) ;
  assign n6558 = n6557 ^ n6556 ^ n1009 ;
  assign n6552 = n4595 ^ n3639 ^ n3634 ;
  assign n6553 = ( ~n2633 & n3952 ) | ( ~n2633 & n6552 ) | ( n3952 & n6552 ) ;
  assign n6559 = n6558 ^ n6553 ^ n968 ;
  assign n6560 = n6559 ^ n4217 ^ n3576 ;
  assign n6561 = n5966 ^ n5057 ^ n1366 ;
  assign n6562 = ( n3455 & n5252 ) | ( n3455 & ~n6561 ) | ( n5252 & ~n6561 ) ;
  assign n6563 = n6562 ^ n5590 ^ n441 ;
  assign n6566 = n2459 ^ n2407 ^ n1455 ;
  assign n6565 = n5306 ^ n3272 ^ n1801 ;
  assign n6564 = ( ~n2162 & n3985 ) | ( ~n2162 & n4724 ) | ( n3985 & n4724 ) ;
  assign n6567 = n6566 ^ n6565 ^ n6564 ;
  assign n6574 = n6268 ^ n3608 ^ n2346 ;
  assign n6571 = n4432 ^ n3876 ^ n1830 ;
  assign n6572 = n6571 ^ n2820 ^ n2199 ;
  assign n6568 = n4269 ^ n3126 ^ n2487 ;
  assign n6569 = n6568 ^ n2070 ^ n1881 ;
  assign n6570 = n6569 ^ n2755 ^ n219 ;
  assign n6573 = n6572 ^ n6570 ^ n950 ;
  assign n6575 = n6574 ^ n6573 ^ n3762 ;
  assign n6579 = ( n661 & n2920 ) | ( n661 & n5260 ) | ( n2920 & n5260 ) ;
  assign n6576 = ( n2687 & n4816 ) | ( n2687 & n5909 ) | ( n4816 & n5909 ) ;
  assign n6577 = ( x120 & ~n5835 ) | ( x120 & n6576 ) | ( ~n5835 & n6576 ) ;
  assign n6578 = n6577 ^ n6200 ^ n5970 ;
  assign n6580 = n6579 ^ n6578 ^ n5026 ;
  assign n6581 = n3045 ^ n1454 ^ n333 ;
  assign n6582 = ( ~n1763 & n2409 ) | ( ~n1763 & n6581 ) | ( n2409 & n6581 ) ;
  assign n6583 = ( ~n892 & n6580 ) | ( ~n892 & n6582 ) | ( n6580 & n6582 ) ;
  assign n6584 = n6583 ^ n3096 ^ n1601 ;
  assign n6585 = ( n2333 & n6575 ) | ( n2333 & n6584 ) | ( n6575 & n6584 ) ;
  assign n6586 = ( n6171 & n6567 ) | ( n6171 & n6585 ) | ( n6567 & n6585 ) ;
  assign n6587 = ( n3094 & ~n6563 ) | ( n3094 & n6586 ) | ( ~n6563 & n6586 ) ;
  assign n6588 = n3577 ^ n1270 ^ n1176 ;
  assign n6593 = ( x116 & ~n279 ) | ( x116 & n5410 ) | ( ~n279 & n5410 ) ;
  assign n6594 = n6593 ^ n5787 ^ n691 ;
  assign n6589 = n3651 ^ n1434 ^ x104 ;
  assign n6590 = n6589 ^ n4759 ^ n677 ;
  assign n6591 = n5151 ^ n2499 ^ n407 ;
  assign n6592 = ( ~n4548 & n6590 ) | ( ~n4548 & n6591 ) | ( n6590 & n6591 ) ;
  assign n6595 = n6594 ^ n6592 ^ x110 ;
  assign n6596 = ( n3918 & n6588 ) | ( n3918 & n6595 ) | ( n6588 & n6595 ) ;
  assign n6597 = n4411 ^ n564 ^ n444 ;
  assign n6598 = ( n536 & n2050 ) | ( n536 & n5893 ) | ( n2050 & n5893 ) ;
  assign n6599 = ( n1541 & ~n1778 ) | ( n1541 & n6598 ) | ( ~n1778 & n6598 ) ;
  assign n6600 = ( x102 & n603 ) | ( x102 & n1285 ) | ( n603 & n1285 ) ;
  assign n6601 = ( ~n2937 & n5550 ) | ( ~n2937 & n6600 ) | ( n5550 & n6600 ) ;
  assign n6602 = n3482 ^ n3301 ^ n2934 ;
  assign n6603 = n6602 ^ n1292 ^ n226 ;
  assign n6604 = ( n1762 & n6601 ) | ( n1762 & n6603 ) | ( n6601 & n6603 ) ;
  assign n6605 = ( n1196 & n1384 ) | ( n1196 & n1545 ) | ( n1384 & n1545 ) ;
  assign n6606 = ( n4577 & n6604 ) | ( n4577 & n6605 ) | ( n6604 & n6605 ) ;
  assign n6607 = ( ~n2044 & n4226 ) | ( ~n2044 & n5912 ) | ( n4226 & n5912 ) ;
  assign n6608 = n6607 ^ n5831 ^ n5793 ;
  assign n6609 = ( n446 & ~n2163 ) | ( n446 & n2792 ) | ( ~n2163 & n2792 ) ;
  assign n6610 = n6609 ^ n3739 ^ n2241 ;
  assign n6611 = n6610 ^ n5621 ^ n1868 ;
  assign n6612 = ( n1099 & ~n4683 ) | ( n1099 & n6611 ) | ( ~n4683 & n6611 ) ;
  assign n6613 = n6612 ^ n3927 ^ n1644 ;
  assign n6614 = n4977 ^ n3457 ^ x123 ;
  assign n6617 = n2852 ^ n870 ^ n515 ;
  assign n6615 = ( n1471 & n1959 ) | ( n1471 & n2684 ) | ( n1959 & n2684 ) ;
  assign n6616 = n6615 ^ n4907 ^ n1122 ;
  assign n6618 = n6617 ^ n6616 ^ n5118 ;
  assign n6619 = n6618 ^ n2328 ^ x88 ;
  assign n6620 = n6619 ^ n3433 ^ n1154 ;
  assign n6621 = ( n452 & n527 ) | ( n452 & n6620 ) | ( n527 & n6620 ) ;
  assign n6622 = ( ~n1766 & n6614 ) | ( ~n1766 & n6621 ) | ( n6614 & n6621 ) ;
  assign n6623 = n2399 ^ n1621 ^ n278 ;
  assign n6624 = n6623 ^ n6573 ^ n2835 ;
  assign n6625 = n6624 ^ n3429 ^ n1095 ;
  assign n6626 = ( n1719 & ~n6622 ) | ( n1719 & n6625 ) | ( ~n6622 & n6625 ) ;
  assign n6627 = ( n328 & ~n1884 ) | ( n328 & n2971 ) | ( ~n1884 & n2971 ) ;
  assign n6628 = n6627 ^ n3307 ^ n777 ;
  assign n6629 = ( n654 & n1356 ) | ( n654 & n2346 ) | ( n1356 & n2346 ) ;
  assign n6631 = ( n1239 & n1476 ) | ( n1239 & n6124 ) | ( n1476 & n6124 ) ;
  assign n6632 = ( n983 & n1121 ) | ( n983 & ~n6631 ) | ( n1121 & ~n6631 ) ;
  assign n6633 = n2633 ^ n617 ^ n419 ;
  assign n6634 = ( n275 & n3952 ) | ( n275 & n6633 ) | ( n3952 & n6633 ) ;
  assign n6635 = ( n358 & n6632 ) | ( n358 & ~n6634 ) | ( n6632 & ~n6634 ) ;
  assign n6630 = ( ~n665 & n1047 ) | ( ~n665 & n4544 ) | ( n1047 & n4544 ) ;
  assign n6636 = n6635 ^ n6630 ^ n373 ;
  assign n6637 = ( n3529 & n6629 ) | ( n3529 & ~n6636 ) | ( n6629 & ~n6636 ) ;
  assign n6643 = ( ~n1123 & n2007 ) | ( ~n1123 & n6432 ) | ( n2007 & n6432 ) ;
  assign n6640 = n1948 ^ n1179 ^ n805 ;
  assign n6641 = n4132 ^ n1476 ^ n1320 ;
  assign n6642 = ( n3703 & ~n6640 ) | ( n3703 & n6641 ) | ( ~n6640 & n6641 ) ;
  assign n6638 = ( n2978 & ~n3430 ) | ( n2978 & n4220 ) | ( ~n3430 & n4220 ) ;
  assign n6639 = ( ~n3964 & n4731 ) | ( ~n3964 & n6638 ) | ( n4731 & n6638 ) ;
  assign n6644 = n6643 ^ n6642 ^ n6639 ;
  assign n6645 = n2938 ^ n2227 ^ n1076 ;
  assign n6646 = n2924 ^ n2573 ^ n653 ;
  assign n6647 = ( n1810 & n6645 ) | ( n1810 & ~n6646 ) | ( n6645 & ~n6646 ) ;
  assign n6648 = n2682 ^ n1846 ^ n1266 ;
  assign n6649 = n6648 ^ n3686 ^ n2079 ;
  assign n6650 = n5539 ^ n4109 ^ n2839 ;
  assign n6651 = n5124 ^ n2549 ^ n399 ;
  assign n6652 = ( n3108 & n3635 ) | ( n3108 & ~n6651 ) | ( n3635 & ~n6651 ) ;
  assign n6653 = ( x58 & n6650 ) | ( x58 & n6652 ) | ( n6650 & n6652 ) ;
  assign n6654 = n6653 ^ n3471 ^ n3239 ;
  assign n6659 = ( n217 & n1751 ) | ( n217 & ~n5416 ) | ( n1751 & ~n5416 ) ;
  assign n6660 = n6659 ^ n4842 ^ n413 ;
  assign n6655 = n4372 ^ n2450 ^ n1447 ;
  assign n6656 = ( n1852 & n4088 ) | ( n1852 & n4191 ) | ( n4088 & n4191 ) ;
  assign n6657 = n6656 ^ n2346 ^ n1562 ;
  assign n6658 = ( ~n2649 & n6655 ) | ( ~n2649 & n6657 ) | ( n6655 & n6657 ) ;
  assign n6661 = n6660 ^ n6658 ^ n4079 ;
  assign n6662 = ( n6649 & n6654 ) | ( n6649 & ~n6661 ) | ( n6654 & ~n6661 ) ;
  assign n6663 = ( n3708 & n6237 ) | ( n3708 & n6350 ) | ( n6237 & n6350 ) ;
  assign n6664 = ( x110 & n3752 ) | ( x110 & n4822 ) | ( n3752 & n4822 ) ;
  assign n6665 = ( n1274 & n2421 ) | ( n1274 & ~n6664 ) | ( n2421 & ~n6664 ) ;
  assign n6668 = n3753 ^ n3667 ^ n1896 ;
  assign n6666 = n4777 ^ n2410 ^ n1917 ;
  assign n6667 = ( n2594 & n2734 ) | ( n2594 & ~n6666 ) | ( n2734 & ~n6666 ) ;
  assign n6669 = n6668 ^ n6667 ^ n6367 ;
  assign n6670 = ( n448 & n4564 ) | ( n448 & n5045 ) | ( n4564 & n5045 ) ;
  assign n6671 = ( ~n3419 & n4365 ) | ( ~n3419 & n5269 ) | ( n4365 & n5269 ) ;
  assign n6672 = ( n1647 & ~n6670 ) | ( n1647 & n6671 ) | ( ~n6670 & n6671 ) ;
  assign n6673 = ( n2668 & n5140 ) | ( n2668 & ~n6672 ) | ( n5140 & ~n6672 ) ;
  assign n6674 = ( n1026 & n6669 ) | ( n1026 & ~n6673 ) | ( n6669 & ~n6673 ) ;
  assign n6675 = ( ~n5021 & n6665 ) | ( ~n5021 & n6674 ) | ( n6665 & n6674 ) ;
  assign n6676 = ( n2275 & ~n3525 ) | ( n2275 & n3877 ) | ( ~n3525 & n3877 ) ;
  assign n6677 = n6676 ^ n4204 ^ n2204 ;
  assign n6678 = ( n1417 & n2453 ) | ( n1417 & ~n2520 ) | ( n2453 & ~n2520 ) ;
  assign n6679 = ( ~n3269 & n6337 ) | ( ~n3269 & n6678 ) | ( n6337 & n6678 ) ;
  assign n6680 = ( n985 & ~n1307 ) | ( n985 & n1459 ) | ( ~n1307 & n1459 ) ;
  assign n6681 = ( n633 & n920 ) | ( n633 & n1994 ) | ( n920 & n1994 ) ;
  assign n6682 = ( x80 & ~n3601 ) | ( x80 & n6681 ) | ( ~n3601 & n6681 ) ;
  assign n6683 = ( ~n3016 & n6680 ) | ( ~n3016 & n6682 ) | ( n6680 & n6682 ) ;
  assign n6704 = ( n3861 & ~n3930 ) | ( n3861 & n4143 ) | ( ~n3930 & n4143 ) ;
  assign n6705 = n6704 ^ n5493 ^ n1127 ;
  assign n6696 = n2506 ^ n783 ^ n235 ;
  assign n6697 = n6696 ^ n377 ^ n284 ;
  assign n6698 = n6697 ^ n1029 ^ n279 ;
  assign n6699 = ( n730 & n751 ) | ( n730 & ~n3491 ) | ( n751 & ~n3491 ) ;
  assign n6700 = n6699 ^ n2982 ^ n2000 ;
  assign n6701 = n6700 ^ n6509 ^ n812 ;
  assign n6702 = ( n1073 & n1922 ) | ( n1073 & ~n6701 ) | ( n1922 & ~n6701 ) ;
  assign n6703 = ( ~n5446 & n6698 ) | ( ~n5446 & n6702 ) | ( n6698 & n6702 ) ;
  assign n6684 = ( n2266 & ~n3557 ) | ( n2266 & n6156 ) | ( ~n3557 & n6156 ) ;
  assign n6685 = ( n1048 & n2139 ) | ( n1048 & n3834 ) | ( n2139 & n3834 ) ;
  assign n6686 = ( n1520 & ~n3398 ) | ( n1520 & n6685 ) | ( ~n3398 & n6685 ) ;
  assign n6687 = ( n173 & n6684 ) | ( n173 & n6686 ) | ( n6684 & n6686 ) ;
  assign n6688 = n4274 ^ n2258 ^ n152 ;
  assign n6689 = ( n2355 & ~n5160 ) | ( n2355 & n6688 ) | ( ~n5160 & n6688 ) ;
  assign n6690 = n6689 ^ n1857 ^ n172 ;
  assign n6691 = n6690 ^ n2475 ^ n203 ;
  assign n6692 = n6691 ^ n3799 ^ n1659 ;
  assign n6693 = n6692 ^ n4382 ^ n365 ;
  assign n6694 = n6693 ^ n5470 ^ n2671 ;
  assign n6695 = ( n413 & ~n6687 ) | ( n413 & n6694 ) | ( ~n6687 & n6694 ) ;
  assign n6706 = n6705 ^ n6703 ^ n6695 ;
  assign n6707 = n6706 ^ n6105 ^ n3603 ;
  assign n6708 = n3736 ^ n3229 ^ n1001 ;
  assign n6709 = ( n223 & ~n3218 ) | ( n223 & n5895 ) | ( ~n3218 & n5895 ) ;
  assign n6710 = ( n1642 & ~n1924 ) | ( n1642 & n6709 ) | ( ~n1924 & n6709 ) ;
  assign n6711 = ( n312 & n599 ) | ( n312 & n2201 ) | ( n599 & n2201 ) ;
  assign n6712 = n6711 ^ n989 ^ x55 ;
  assign n6713 = ( n1211 & n3488 ) | ( n1211 & n6712 ) | ( n3488 & n6712 ) ;
  assign n6715 = ( n1851 & n1936 ) | ( n1851 & ~n4253 ) | ( n1936 & ~n4253 ) ;
  assign n6714 = n2956 ^ n511 ^ x13 ;
  assign n6716 = n6715 ^ n6714 ^ n362 ;
  assign n6717 = ( n533 & n6713 ) | ( n533 & n6716 ) | ( n6713 & n6716 ) ;
  assign n6718 = ( n6708 & n6710 ) | ( n6708 & n6717 ) | ( n6710 & n6717 ) ;
  assign n6719 = ( n1874 & ~n2506 ) | ( n1874 & n5344 ) | ( ~n2506 & n5344 ) ;
  assign n6720 = ( n536 & n4656 ) | ( n536 & ~n6681 ) | ( n4656 & ~n6681 ) ;
  assign n6721 = ( n2140 & n6719 ) | ( n2140 & n6720 ) | ( n6719 & n6720 ) ;
  assign n6722 = ( ~n418 & n1475 ) | ( ~n418 & n3478 ) | ( n1475 & n3478 ) ;
  assign n6723 = n4721 ^ n1907 ^ n386 ;
  assign n6724 = n318 ^ x76 ^ x48 ;
  assign n6725 = n6724 ^ n2278 ^ n2051 ;
  assign n6726 = n5073 ^ n5055 ^ n4935 ;
  assign n6727 = ( n1370 & n6725 ) | ( n1370 & n6726 ) | ( n6725 & n6726 ) ;
  assign n6728 = ( ~n4228 & n4775 ) | ( ~n4228 & n6727 ) | ( n4775 & n6727 ) ;
  assign n6729 = ( n6722 & ~n6723 ) | ( n6722 & n6728 ) | ( ~n6723 & n6728 ) ;
  assign n6730 = n6358 ^ n4745 ^ n1843 ;
  assign n6734 = ( ~n2422 & n5152 ) | ( ~n2422 & n5460 ) | ( n5152 & n5460 ) ;
  assign n6732 = ( n418 & n2671 ) | ( n418 & ~n5179 ) | ( n2671 & ~n5179 ) ;
  assign n6731 = n5123 ^ n3421 ^ n293 ;
  assign n6733 = n6732 ^ n6731 ^ n1017 ;
  assign n6735 = n6734 ^ n6733 ^ n4319 ;
  assign n6743 = n4061 ^ n2541 ^ n2224 ;
  assign n6741 = n6444 ^ n5409 ^ n673 ;
  assign n6742 = n6741 ^ n6124 ^ n1526 ;
  assign n6737 = n4269 ^ n1284 ^ n773 ;
  assign n6738 = n6737 ^ n2898 ^ n1222 ;
  assign n6736 = ( n3029 & ~n3785 ) | ( n3029 & n3863 ) | ( ~n3785 & n3863 ) ;
  assign n6739 = n6738 ^ n6736 ^ n3061 ;
  assign n6740 = n6739 ^ n4316 ^ n309 ;
  assign n6744 = n6743 ^ n6742 ^ n6740 ;
  assign n6747 = ( n134 & ~n1344 ) | ( n134 & n3091 ) | ( ~n1344 & n3091 ) ;
  assign n6745 = ( n1961 & n5371 ) | ( n1961 & ~n6468 ) | ( n5371 & ~n6468 ) ;
  assign n6746 = n6745 ^ n6266 ^ n425 ;
  assign n6748 = n6747 ^ n6746 ^ n6042 ;
  assign n6749 = ( n629 & ~n5798 ) | ( n629 & n6748 ) | ( ~n5798 & n6748 ) ;
  assign n6750 = ( n6735 & ~n6744 ) | ( n6735 & n6749 ) | ( ~n6744 & n6749 ) ;
  assign n6751 = ( x73 & n258 ) | ( x73 & n999 ) | ( n258 & n999 ) ;
  assign n6755 = ( n282 & ~n3213 ) | ( n282 & n3486 ) | ( ~n3213 & n3486 ) ;
  assign n6753 = n2760 ^ n1452 ^ n144 ;
  assign n6752 = n6708 ^ n564 ^ n253 ;
  assign n6754 = n6753 ^ n6752 ^ n3003 ;
  assign n6756 = n6755 ^ n6754 ^ n2008 ;
  assign n6759 = n3634 ^ n2305 ^ n1020 ;
  assign n6760 = n6759 ^ n2884 ^ x121 ;
  assign n6761 = ( n1478 & n2677 ) | ( n1478 & n6760 ) | ( n2677 & n6760 ) ;
  assign n6757 = ( n473 & n1037 ) | ( n473 & ~n4449 ) | ( n1037 & ~n4449 ) ;
  assign n6758 = ( n2912 & ~n4870 ) | ( n2912 & n6757 ) | ( ~n4870 & n6757 ) ;
  assign n6762 = n6761 ^ n6758 ^ n3524 ;
  assign n6763 = ( n6751 & n6756 ) | ( n6751 & n6762 ) | ( n6756 & n6762 ) ;
  assign n6764 = ( ~n3160 & n3704 ) | ( ~n3160 & n5886 ) | ( n3704 & n5886 ) ;
  assign n6773 = n5131 ^ n4512 ^ n2034 ;
  assign n6765 = n6753 ^ n5757 ^ n1141 ;
  assign n6766 = ( n1345 & n1756 ) | ( n1345 & n3906 ) | ( n1756 & n3906 ) ;
  assign n6767 = ( ~n1527 & n2297 ) | ( ~n1527 & n2972 ) | ( n2297 & n2972 ) ;
  assign n6768 = n3600 ^ n1569 ^ n895 ;
  assign n6769 = ( n1891 & n6767 ) | ( n1891 & ~n6768 ) | ( n6767 & ~n6768 ) ;
  assign n6770 = ( n497 & n6766 ) | ( n497 & ~n6769 ) | ( n6766 & ~n6769 ) ;
  assign n6771 = ( ~n2787 & n3039 ) | ( ~n2787 & n6770 ) | ( n3039 & n6770 ) ;
  assign n6772 = ( n6188 & ~n6765 ) | ( n6188 & n6771 ) | ( ~n6765 & n6771 ) ;
  assign n6774 = n6773 ^ n6772 ^ n5264 ;
  assign n6776 = n6643 ^ n5236 ^ n1186 ;
  assign n6777 = ( ~n129 & n5835 ) | ( ~n129 & n6776 ) | ( n5835 & n6776 ) ;
  assign n6775 = ( n2275 & n4860 ) | ( n2275 & n5893 ) | ( n4860 & n5893 ) ;
  assign n6778 = n6777 ^ n6775 ^ n4718 ;
  assign n6779 = n5993 ^ n5449 ^ n891 ;
  assign n6780 = ( n1667 & n4233 ) | ( n1667 & n5550 ) | ( n4233 & n5550 ) ;
  assign n6781 = ( n1465 & n5221 ) | ( n1465 & ~n6780 ) | ( n5221 & ~n6780 ) ;
  assign n6782 = n4822 ^ n3762 ^ n2572 ;
  assign n6790 = n6769 ^ n4712 ^ n1202 ;
  assign n6791 = n6790 ^ n6678 ^ n4469 ;
  assign n6792 = ( n3742 & n5080 ) | ( n3742 & n6791 ) | ( n5080 & n6791 ) ;
  assign n6793 = ( n1239 & n1551 ) | ( n1239 & ~n4095 ) | ( n1551 & ~n4095 ) ;
  assign n6794 = n6793 ^ n2473 ^ n2415 ;
  assign n6795 = n6794 ^ n1913 ^ n1908 ;
  assign n6796 = ( ~n3710 & n6792 ) | ( ~n3710 & n6795 ) | ( n6792 & n6795 ) ;
  assign n6786 = ( n2125 & n2660 ) | ( n2125 & ~n2662 ) | ( n2660 & ~n2662 ) ;
  assign n6787 = n6786 ^ n4940 ^ n788 ;
  assign n6783 = n4204 ^ n4123 ^ n2295 ;
  assign n6784 = n2782 ^ n2194 ^ n1200 ;
  assign n6785 = ( ~n5439 & n6783 ) | ( ~n5439 & n6784 ) | ( n6783 & n6784 ) ;
  assign n6788 = n6787 ^ n6785 ^ n1973 ;
  assign n6789 = ( ~n901 & n3720 ) | ( ~n901 & n6788 ) | ( n3720 & n6788 ) ;
  assign n6797 = n6796 ^ n6789 ^ n6046 ;
  assign n6798 = n2547 ^ n782 ^ n369 ;
  assign n6799 = n6798 ^ n6111 ^ n4627 ;
  assign n6800 = ( n2688 & n5989 ) | ( n2688 & n6799 ) | ( n5989 & n6799 ) ;
  assign n6801 = n1887 ^ n591 ^ n519 ;
  assign n6802 = ( n998 & n1310 ) | ( n998 & ~n4678 ) | ( n1310 & ~n4678 ) ;
  assign n6803 = ( n348 & ~n3327 ) | ( n348 & n6802 ) | ( ~n3327 & n6802 ) ;
  assign n6804 = ( n2115 & n2839 ) | ( n2115 & n6803 ) | ( n2839 & n6803 ) ;
  assign n6805 = n6804 ^ n4232 ^ n3203 ;
  assign n6810 = ( n2951 & n3903 ) | ( n2951 & n4858 ) | ( n3903 & n4858 ) ;
  assign n6807 = n4890 ^ n4827 ^ n4578 ;
  assign n6806 = ( n577 & ~n1541 ) | ( n577 & n2661 ) | ( ~n1541 & n2661 ) ;
  assign n6808 = n6807 ^ n6806 ^ n975 ;
  assign n6809 = n6808 ^ n1908 ^ n547 ;
  assign n6811 = n6810 ^ n6809 ^ n5081 ;
  assign n6812 = n6811 ^ n3436 ^ n3064 ;
  assign n6813 = ( n6801 & n6805 ) | ( n6801 & n6812 ) | ( n6805 & n6812 ) ;
  assign n6820 = n3990 ^ n3341 ^ n312 ;
  assign n6816 = ( n170 & n333 ) | ( n170 & n525 ) | ( n333 & n525 ) ;
  assign n6817 = ( ~n1404 & n1955 ) | ( ~n1404 & n3542 ) | ( n1955 & n3542 ) ;
  assign n6818 = n6817 ^ n301 ^ x29 ;
  assign n6819 = ( n3312 & n6816 ) | ( n3312 & n6818 ) | ( n6816 & n6818 ) ;
  assign n6814 = n3669 ^ n2315 ^ n2206 ;
  assign n6815 = ( n1657 & n2039 ) | ( n1657 & ~n6814 ) | ( n2039 & ~n6814 ) ;
  assign n6821 = n6820 ^ n6819 ^ n6815 ;
  assign n6825 = n2373 ^ n2067 ^ n811 ;
  assign n6823 = ( n2692 & n3228 ) | ( n2692 & ~n6343 ) | ( n3228 & ~n6343 ) ;
  assign n6822 = n4562 ^ n2656 ^ n2019 ;
  assign n6824 = n6823 ^ n6822 ^ n2291 ;
  assign n6826 = n6825 ^ n6824 ^ n1073 ;
  assign n6827 = ( n1100 & n2218 ) | ( n1100 & n6826 ) | ( n2218 & n6826 ) ;
  assign n6838 = ( ~x67 & n730 ) | ( ~x67 & n3528 ) | ( n730 & n3528 ) ;
  assign n6835 = n1692 ^ n846 ^ n529 ;
  assign n6836 = n6835 ^ n538 ^ n235 ;
  assign n6837 = n6836 ^ n5131 ^ n2547 ;
  assign n6839 = n6838 ^ n6837 ^ n4191 ;
  assign n6828 = ( ~n1492 & n2315 ) | ( ~n1492 & n3540 ) | ( n2315 & n3540 ) ;
  assign n6829 = ( ~x122 & n3486 ) | ( ~x122 & n6828 ) | ( n3486 & n6828 ) ;
  assign n6830 = ( n906 & n2856 ) | ( n906 & n5245 ) | ( n2856 & n5245 ) ;
  assign n6831 = n6830 ^ n5785 ^ n3455 ;
  assign n6832 = ( n2090 & n2771 ) | ( n2090 & ~n6831 ) | ( n2771 & ~n6831 ) ;
  assign n6833 = ( n553 & n6829 ) | ( n553 & ~n6832 ) | ( n6829 & ~n6832 ) ;
  assign n6834 = ( n2787 & n6591 ) | ( n2787 & ~n6833 ) | ( n6591 & ~n6833 ) ;
  assign n6840 = n6839 ^ n6834 ^ n5160 ;
  assign n6841 = ( ~n3062 & n4163 ) | ( ~n3062 & n4875 ) | ( n4163 & n4875 ) ;
  assign n6846 = ( n177 & ~n657 ) | ( n177 & n1879 ) | ( ~n657 & n1879 ) ;
  assign n6842 = ( n1664 & ~n2619 ) | ( n1664 & n4804 ) | ( ~n2619 & n4804 ) ;
  assign n6843 = ( x87 & n4259 ) | ( x87 & n6842 ) | ( n4259 & n6842 ) ;
  assign n6844 = ( ~n2942 & n5803 ) | ( ~n2942 & n6843 ) | ( n5803 & n6843 ) ;
  assign n6845 = ( n3861 & ~n3972 ) | ( n3861 & n6844 ) | ( ~n3972 & n6844 ) ;
  assign n6847 = n6846 ^ n6845 ^ n4467 ;
  assign n6848 = n1985 ^ n1782 ^ n1712 ;
  assign n6849 = n3906 ^ n1868 ^ x104 ;
  assign n6850 = n6849 ^ n6258 ^ n3860 ;
  assign n6851 = ( n2874 & ~n6848 ) | ( n2874 & n6850 ) | ( ~n6848 & n6850 ) ;
  assign n6852 = ( n2365 & ~n2918 ) | ( n2365 & n5432 ) | ( ~n2918 & n5432 ) ;
  assign n6853 = ( ~n2708 & n5391 ) | ( ~n2708 & n6852 ) | ( n5391 & n6852 ) ;
  assign n6854 = n2376 ^ n1413 ^ n817 ;
  assign n6855 = n6854 ^ n2778 ^ n1241 ;
  assign n6856 = n6855 ^ n1142 ^ x106 ;
  assign n6857 = n6856 ^ n3424 ^ n654 ;
  assign n6858 = ( n285 & n6853 ) | ( n285 & ~n6857 ) | ( n6853 & ~n6857 ) ;
  assign n6887 = n5972 ^ n4544 ^ n429 ;
  assign n6859 = ( n258 & ~n2082 ) | ( n258 & n5254 ) | ( ~n2082 & n5254 ) ;
  assign n6860 = n6859 ^ n3111 ^ n632 ;
  assign n6861 = ( n3859 & n4612 ) | ( n3859 & ~n6860 ) | ( n4612 & ~n6860 ) ;
  assign n6862 = ( ~n734 & n1298 ) | ( ~n734 & n5390 ) | ( n1298 & n5390 ) ;
  assign n6867 = ( x99 & n1448 ) | ( x99 & ~n1697 ) | ( n1448 & ~n1697 ) ;
  assign n6863 = n3576 ^ n2305 ^ n387 ;
  assign n6864 = n2628 ^ n2138 ^ n763 ;
  assign n6865 = ( ~n819 & n950 ) | ( ~n819 & n6864 ) | ( n950 & n6864 ) ;
  assign n6866 = ( n5937 & n6863 ) | ( n5937 & n6865 ) | ( n6863 & n6865 ) ;
  assign n6868 = n6867 ^ n6866 ^ n2433 ;
  assign n6869 = ( ~n437 & n6862 ) | ( ~n437 & n6868 ) | ( n6862 & n6868 ) ;
  assign n6870 = n6869 ^ n2915 ^ n1484 ;
  assign n6871 = ( ~n3459 & n6861 ) | ( ~n3459 & n6870 ) | ( n6861 & n6870 ) ;
  assign n6872 = n2014 ^ n1870 ^ x104 ;
  assign n6873 = ( ~n520 & n1213 ) | ( ~n520 & n3476 ) | ( n1213 & n3476 ) ;
  assign n6874 = ( ~n544 & n3285 ) | ( ~n544 & n6873 ) | ( n3285 & n6873 ) ;
  assign n6875 = n5460 ^ n1337 ^ n810 ;
  assign n6876 = n6875 ^ n5999 ^ n1077 ;
  assign n6877 = ( n6872 & ~n6874 ) | ( n6872 & n6876 ) | ( ~n6874 & n6876 ) ;
  assign n6880 = n5193 ^ n1892 ^ n839 ;
  assign n6881 = ( n178 & ~n1336 ) | ( n178 & n6880 ) | ( ~n1336 & n6880 ) ;
  assign n6882 = n6881 ^ n3062 ^ n1346 ;
  assign n6883 = n6882 ^ n1380 ^ n879 ;
  assign n6879 = n6256 ^ n5624 ^ n3869 ;
  assign n6878 = n5128 ^ n4958 ^ n4909 ;
  assign n6884 = n6883 ^ n6879 ^ n6878 ;
  assign n6885 = ( n1906 & ~n5553 ) | ( n1906 & n6884 ) | ( ~n5553 & n6884 ) ;
  assign n6886 = ( n6871 & ~n6877 ) | ( n6871 & n6885 ) | ( ~n6877 & n6885 ) ;
  assign n6888 = n6887 ^ n6886 ^ n5691 ;
  assign n6899 = ( n1485 & ~n1932 ) | ( n1485 & n5404 ) | ( ~n1932 & n5404 ) ;
  assign n6896 = n3665 ^ n1720 ^ n868 ;
  assign n6897 = ( x50 & ~n1750 ) | ( x50 & n2504 ) | ( ~n1750 & n2504 ) ;
  assign n6898 = ( ~x46 & n6896 ) | ( ~x46 & n6897 ) | ( n6896 & n6897 ) ;
  assign n6892 = ( n1006 & ~n5467 ) | ( n1006 & n5586 ) | ( ~n5467 & n5586 ) ;
  assign n6889 = ( n976 & n5526 ) | ( n976 & n6336 ) | ( n5526 & n6336 ) ;
  assign n6890 = ( n319 & n3645 ) | ( n319 & n6889 ) | ( n3645 & n6889 ) ;
  assign n6891 = n6890 ^ n5401 ^ n4679 ;
  assign n6893 = n6892 ^ n6891 ^ n5285 ;
  assign n6894 = n6893 ^ n5860 ^ n3372 ;
  assign n6895 = n6894 ^ n4174 ^ n3821 ;
  assign n6900 = n6899 ^ n6898 ^ n6895 ;
  assign n6902 = ( ~n1386 & n4003 ) | ( ~n1386 & n4725 ) | ( n4003 & n4725 ) ;
  assign n6901 = ( n833 & n1544 ) | ( n833 & ~n4469 ) | ( n1544 & ~n4469 ) ;
  assign n6903 = n6902 ^ n6901 ^ n2901 ;
  assign n6904 = ( n1005 & n2066 ) | ( n1005 & ~n3876 ) | ( n2066 & ~n3876 ) ;
  assign n6905 = ( n1102 & n1525 ) | ( n1102 & n6807 ) | ( n1525 & n6807 ) ;
  assign n6906 = ( ~n3023 & n6904 ) | ( ~n3023 & n6905 ) | ( n6904 & n6905 ) ;
  assign n6907 = n6906 ^ n1609 ^ n873 ;
  assign n6908 = n6907 ^ n2445 ^ n2340 ;
  assign n6909 = ( n1523 & n3332 ) | ( n1523 & n5315 ) | ( n3332 & n5315 ) ;
  assign n6913 = n4989 ^ n4352 ^ n2183 ;
  assign n6914 = n6913 ^ n2489 ^ n1823 ;
  assign n6910 = n1938 ^ n1025 ^ n993 ;
  assign n6911 = ( n1527 & n1812 ) | ( n1527 & n6910 ) | ( n1812 & n6910 ) ;
  assign n6912 = ( n3757 & n5953 ) | ( n3757 & n6911 ) | ( n5953 & n6911 ) ;
  assign n6915 = n6914 ^ n6912 ^ n206 ;
  assign n6916 = n6915 ^ n5694 ^ n2633 ;
  assign n6920 = ( n1213 & n1366 ) | ( n1213 & ~n4744 ) | ( n1366 & ~n4744 ) ;
  assign n6919 = n5702 ^ n2772 ^ n2664 ;
  assign n6917 = n4110 ^ n2579 ^ n1467 ;
  assign n6918 = n6917 ^ n1006 ^ n649 ;
  assign n6921 = n6920 ^ n6919 ^ n6918 ;
  assign n6922 = ( ~n552 & n2176 ) | ( ~n552 & n4027 ) | ( n2176 & n4027 ) ;
  assign n6923 = n6922 ^ n4128 ^ n2650 ;
  assign n6928 = n2253 ^ n1379 ^ n1023 ;
  assign n6929 = n6928 ^ n1944 ^ n1620 ;
  assign n6927 = n6206 ^ n4360 ^ n401 ;
  assign n6924 = ( n2051 & ~n2702 ) | ( n2051 & n3483 ) | ( ~n2702 & n3483 ) ;
  assign n6925 = ( n1697 & n3454 ) | ( n1697 & ~n6924 ) | ( n3454 & ~n6924 ) ;
  assign n6926 = ( n1293 & n5689 ) | ( n1293 & n6925 ) | ( n5689 & n6925 ) ;
  assign n6930 = n6929 ^ n6927 ^ n6926 ;
  assign n6931 = ( ~n3029 & n6923 ) | ( ~n3029 & n6930 ) | ( n6923 & n6930 ) ;
  assign n6932 = n4463 ^ n2501 ^ n1950 ;
  assign n6933 = n6932 ^ n4293 ^ n250 ;
  assign n6934 = n6933 ^ n5914 ^ n1748 ;
  assign n6935 = ( ~n1901 & n3057 ) | ( ~n1901 & n4293 ) | ( n3057 & n4293 ) ;
  assign n6936 = ( ~n617 & n1430 ) | ( ~n617 & n6935 ) | ( n1430 & n6935 ) ;
  assign n6937 = n6864 ^ n2413 ^ n971 ;
  assign n6938 = ( x60 & n6936 ) | ( x60 & ~n6937 ) | ( n6936 & ~n6937 ) ;
  assign n6939 = ( x58 & n2090 ) | ( x58 & n4147 ) | ( n2090 & n4147 ) ;
  assign n6940 = ( n2481 & n4248 ) | ( n2481 & ~n6467 ) | ( n4248 & ~n6467 ) ;
  assign n6941 = n6940 ^ n5456 ^ n720 ;
  assign n6944 = n5456 ^ n1641 ^ x61 ;
  assign n6945 = n6944 ^ n4511 ^ n1011 ;
  assign n6946 = ( n270 & ~n906 ) | ( n270 & n1716 ) | ( ~n906 & n1716 ) ;
  assign n6947 = ( ~n2210 & n5912 ) | ( ~n2210 & n6946 ) | ( n5912 & n6946 ) ;
  assign n6948 = ( ~n2167 & n6945 ) | ( ~n2167 & n6947 ) | ( n6945 & n6947 ) ;
  assign n6943 = ( n1220 & n1671 ) | ( n1220 & ~n4937 ) | ( n1671 & ~n4937 ) ;
  assign n6942 = n6444 ^ n5357 ^ n4096 ;
  assign n6949 = n6948 ^ n6943 ^ n6942 ;
  assign n6950 = ( n2220 & ~n5101 ) | ( n2220 & n6949 ) | ( ~n5101 & n6949 ) ;
  assign n6951 = ( n4376 & ~n6941 ) | ( n4376 & n6950 ) | ( ~n6941 & n6950 ) ;
  assign n6952 = ( n845 & n4283 ) | ( n845 & ~n5739 ) | ( n4283 & ~n5739 ) ;
  assign n6953 = n3632 ^ n3483 ^ n177 ;
  assign n6954 = ( n1893 & n5007 ) | ( n1893 & ~n6953 ) | ( n5007 & ~n6953 ) ;
  assign n6959 = n5079 ^ n1354 ^ n691 ;
  assign n6960 = ( n2413 & n6163 ) | ( n2413 & ~n6959 ) | ( n6163 & ~n6959 ) ;
  assign n6956 = ( n2777 & n3552 ) | ( n2777 & n4967 ) | ( n3552 & n4967 ) ;
  assign n6955 = ( n3938 & n4996 ) | ( n3938 & n5189 ) | ( n4996 & n5189 ) ;
  assign n6957 = n6956 ^ n6955 ^ n1046 ;
  assign n6958 = n6957 ^ n4653 ^ n2626 ;
  assign n6961 = n6960 ^ n6958 ^ n2164 ;
  assign n6962 = ( ~n6952 & n6954 ) | ( ~n6952 & n6961 ) | ( n6954 & n6961 ) ;
  assign n6963 = n5372 ^ n4850 ^ n1159 ;
  assign n6964 = ( ~n4991 & n6902 ) | ( ~n4991 & n6963 ) | ( n6902 & n6963 ) ;
  assign n6965 = ( n289 & ~n1737 ) | ( n289 & n3057 ) | ( ~n1737 & n3057 ) ;
  assign n6966 = ( n4434 & n6959 ) | ( n4434 & n6965 ) | ( n6959 & n6965 ) ;
  assign n6967 = n6966 ^ n3320 ^ n2001 ;
  assign n6968 = n6967 ^ n4282 ^ n1180 ;
  assign n6969 = ( ~n1201 & n6964 ) | ( ~n1201 & n6968 ) | ( n6964 & n6968 ) ;
  assign n6984 = ( n1352 & n3827 ) | ( n1352 & n6106 ) | ( n3827 & n6106 ) ;
  assign n6982 = n4049 ^ n2035 ^ n178 ;
  assign n6980 = n3209 ^ n1893 ^ n1400 ;
  assign n6981 = n6980 ^ n2489 ^ n482 ;
  assign n6983 = n6982 ^ n6981 ^ n3521 ;
  assign n6970 = n4536 ^ n3869 ^ n3292 ;
  assign n6971 = ( n1105 & n1149 ) | ( n1105 & n5235 ) | ( n1149 & n5235 ) ;
  assign n6972 = ( n3017 & n4045 ) | ( n3017 & ~n6971 ) | ( n4045 & ~n6971 ) ;
  assign n6973 = ( ~n560 & n4452 ) | ( ~n560 & n5235 ) | ( n4452 & n5235 ) ;
  assign n6974 = n6973 ^ n6823 ^ n4804 ;
  assign n6975 = ( n3472 & ~n6972 ) | ( n3472 & n6974 ) | ( ~n6972 & n6974 ) ;
  assign n6976 = ( n219 & n1407 ) | ( n219 & ~n6975 ) | ( n1407 & ~n6975 ) ;
  assign n6977 = n6976 ^ n1782 ^ n648 ;
  assign n6978 = ( x8 & n4052 ) | ( x8 & ~n6977 ) | ( n4052 & ~n6977 ) ;
  assign n6979 = ( n2776 & ~n6970 ) | ( n2776 & n6978 ) | ( ~n6970 & n6978 ) ;
  assign n6985 = n6984 ^ n6983 ^ n6979 ;
  assign n6990 = n2294 ^ n1896 ^ n1764 ;
  assign n6986 = ( ~n1315 & n2148 ) | ( ~n1315 & n3906 ) | ( n2148 & n3906 ) ;
  assign n6987 = n6986 ^ n5461 ^ n2164 ;
  assign n6988 = ( n2420 & n5605 ) | ( n2420 & ~n6987 ) | ( n5605 & ~n6987 ) ;
  assign n6989 = n6988 ^ n5842 ^ n4379 ;
  assign n6991 = n6990 ^ n6989 ^ n388 ;
  assign n6992 = ( n179 & n3172 ) | ( n179 & ~n6387 ) | ( n3172 & ~n6387 ) ;
  assign n6993 = ( n365 & n6991 ) | ( n365 & n6992 ) | ( n6991 & n6992 ) ;
  assign n6994 = ( n392 & n5502 ) | ( n392 & ~n6547 ) | ( n5502 & ~n6547 ) ;
  assign n6995 = n3186 ^ n1046 ^ n564 ;
  assign n6996 = ( n3962 & n6836 ) | ( n3962 & ~n6995 ) | ( n6836 & ~n6995 ) ;
  assign n6997 = ( ~n2118 & n6994 ) | ( ~n2118 & n6996 ) | ( n6994 & n6996 ) ;
  assign n6998 = ( n213 & n5030 ) | ( n213 & n6997 ) | ( n5030 & n6997 ) ;
  assign n6999 = ( n3985 & ~n4209 ) | ( n3985 & n6020 ) | ( ~n4209 & n6020 ) ;
  assign n7000 = ( ~n2561 & n5006 ) | ( ~n2561 & n6999 ) | ( n5006 & n6999 ) ;
  assign n7001 = n6045 ^ n5659 ^ n3547 ;
  assign n7002 = ( n2663 & ~n7000 ) | ( n2663 & n7001 ) | ( ~n7000 & n7001 ) ;
  assign n7003 = n7002 ^ n6617 ^ n2569 ;
  assign n7004 = ( ~n1597 & n2088 ) | ( ~n1597 & n2971 ) | ( n2088 & n2971 ) ;
  assign n7005 = ( n1309 & n6245 ) | ( n1309 & n7004 ) | ( n6245 & n7004 ) ;
  assign n7006 = n7005 ^ n5710 ^ x104 ;
  assign n7007 = ( ~n505 & n835 ) | ( ~n505 & n1740 ) | ( n835 & n1740 ) ;
  assign n7008 = ( n726 & ~n1133 ) | ( n726 & n1608 ) | ( ~n1133 & n1608 ) ;
  assign n7009 = n7008 ^ n6759 ^ n3419 ;
  assign n7010 = ( n1225 & n7007 ) | ( n1225 & n7009 ) | ( n7007 & n7009 ) ;
  assign n7011 = ( n3228 & ~n4608 ) | ( n3228 & n7010 ) | ( ~n4608 & n7010 ) ;
  assign n7012 = ( n6157 & n7006 ) | ( n6157 & ~n7011 ) | ( n7006 & ~n7011 ) ;
  assign n7013 = ( n2138 & ~n7003 ) | ( n2138 & n7012 ) | ( ~n7003 & n7012 ) ;
  assign n7014 = n6002 ^ n4958 ^ n3965 ;
  assign n7015 = n3617 ^ n2247 ^ n1876 ;
  assign n7016 = n1844 ^ n808 ^ n188 ;
  assign n7017 = ( n208 & n3801 ) | ( n208 & n7016 ) | ( n3801 & n7016 ) ;
  assign n7018 = ( ~n6424 & n7015 ) | ( ~n6424 & n7017 ) | ( n7015 & n7017 ) ;
  assign n7019 = ( n5501 & n7014 ) | ( n5501 & ~n7018 ) | ( n7014 & ~n7018 ) ;
  assign n7020 = n7019 ^ n6815 ^ n4845 ;
  assign n7021 = ( n3447 & n3725 ) | ( n3447 & n7020 ) | ( n3725 & n7020 ) ;
  assign n7026 = n5397 ^ n3428 ^ n419 ;
  assign n7027 = n7026 ^ n6798 ^ n891 ;
  assign n7022 = n5997 ^ n4315 ^ n963 ;
  assign n7023 = ( n543 & ~n2334 ) | ( n543 & n7022 ) | ( ~n2334 & n7022 ) ;
  assign n7024 = n7023 ^ n5357 ^ n506 ;
  assign n7025 = n7024 ^ n3635 ^ n2270 ;
  assign n7028 = n7027 ^ n7025 ^ n1351 ;
  assign n7029 = n7028 ^ n5225 ^ n3776 ;
  assign n7032 = n3115 ^ n724 ^ n612 ;
  assign n7033 = ( n200 & n3093 ) | ( n200 & n7032 ) | ( n3093 & n7032 ) ;
  assign n7030 = n3723 ^ n2448 ^ n341 ;
  assign n7031 = ( n466 & n2913 ) | ( n466 & n7030 ) | ( n2913 & n7030 ) ;
  assign n7034 = n7033 ^ n7031 ^ n1848 ;
  assign n7035 = n4111 ^ n1591 ^ n1244 ;
  assign n7045 = ( n1295 & n2886 ) | ( n1295 & n6862 ) | ( n2886 & n6862 ) ;
  assign n7040 = ( n255 & ~n345 ) | ( n255 & n901 ) | ( ~n345 & n901 ) ;
  assign n7041 = ( n1105 & n2527 ) | ( n1105 & n6697 ) | ( n2527 & n6697 ) ;
  assign n7042 = ( n1503 & n5034 ) | ( n1503 & n7041 ) | ( n5034 & n7041 ) ;
  assign n7043 = ( n2528 & ~n7040 ) | ( n2528 & n7042 ) | ( ~n7040 & n7042 ) ;
  assign n7039 = ( x35 & n1996 ) | ( x35 & n3591 ) | ( n1996 & n3591 ) ;
  assign n7044 = n7043 ^ n7039 ^ n1920 ;
  assign n7036 = n4470 ^ n1966 ^ n1549 ;
  assign n7037 = ( n2268 & ~n2688 ) | ( n2268 & n6905 ) | ( ~n2688 & n6905 ) ;
  assign n7038 = ( n4718 & n7036 ) | ( n4718 & ~n7037 ) | ( n7036 & ~n7037 ) ;
  assign n7046 = n7045 ^ n7044 ^ n7038 ;
  assign n7047 = ( n7034 & n7035 ) | ( n7034 & n7046 ) | ( n7035 & n7046 ) ;
  assign n7049 = ( n131 & n1503 ) | ( n131 & n2072 ) | ( n1503 & n2072 ) ;
  assign n7048 = ( n608 & n3131 ) | ( n608 & ~n3505 ) | ( n3131 & ~n3505 ) ;
  assign n7050 = n7049 ^ n7048 ^ n2415 ;
  assign n7051 = ( ~x28 & n3653 ) | ( ~x28 & n3904 ) | ( n3653 & n3904 ) ;
  assign n7052 = n7051 ^ n4193 ^ n2516 ;
  assign n7053 = n5128 ^ n4354 ^ n1393 ;
  assign n7054 = ( n813 & n7052 ) | ( n813 & ~n7053 ) | ( n7052 & ~n7053 ) ;
  assign n7055 = n4163 ^ n2824 ^ n1559 ;
  assign n7056 = ( ~n6640 & n7054 ) | ( ~n6640 & n7055 ) | ( n7054 & n7055 ) ;
  assign n7059 = ( n503 & n722 ) | ( n503 & n2634 ) | ( n722 & n2634 ) ;
  assign n7060 = n7059 ^ n1765 ^ n1691 ;
  assign n7057 = ( n737 & n5632 ) | ( n737 & ~n5864 ) | ( n5632 & ~n5864 ) ;
  assign n7058 = ( n2468 & n6274 ) | ( n2468 & ~n7057 ) | ( n6274 & ~n7057 ) ;
  assign n7061 = n7060 ^ n7058 ^ x126 ;
  assign n7062 = ( n7050 & n7056 ) | ( n7050 & n7061 ) | ( n7056 & n7061 ) ;
  assign n7063 = n6546 ^ n4224 ^ n1213 ;
  assign n7064 = n7063 ^ n2326 ^ n138 ;
  assign n7067 = ( n2167 & n3971 ) | ( n2167 & n4169 ) | ( n3971 & n4169 ) ;
  assign n7068 = n7067 ^ n5459 ^ n4298 ;
  assign n7065 = n6206 ^ n3647 ^ n2898 ;
  assign n7066 = ( n1820 & ~n4563 ) | ( n1820 & n7065 ) | ( ~n4563 & n7065 ) ;
  assign n7069 = n7068 ^ n7066 ^ n7032 ;
  assign n7070 = n2403 ^ n918 ^ n170 ;
  assign n7071 = n2393 ^ n1741 ^ n618 ;
  assign n7072 = ( n3774 & ~n7070 ) | ( n3774 & n7071 ) | ( ~n7070 & n7071 ) ;
  assign n7073 = ( n2627 & ~n4187 ) | ( n2627 & n7072 ) | ( ~n4187 & n7072 ) ;
  assign n7074 = ( n334 & ~n2719 ) | ( n334 & n3494 ) | ( ~n2719 & n3494 ) ;
  assign n7075 = n7074 ^ n6329 ^ n4950 ;
  assign n7076 = ( n3519 & n3669 ) | ( n3519 & ~n5715 ) | ( n3669 & ~n5715 ) ;
  assign n7077 = n7076 ^ n2760 ^ n177 ;
  assign n7078 = n5053 ^ n5020 ^ n2649 ;
  assign n7079 = ( n2317 & ~n7077 ) | ( n2317 & n7078 ) | ( ~n7077 & n7078 ) ;
  assign n7080 = n5183 ^ n5118 ^ n3960 ;
  assign n7081 = ( n1129 & n1223 ) | ( n1129 & ~n3189 ) | ( n1223 & ~n3189 ) ;
  assign n7082 = ( n1586 & ~n2543 ) | ( n1586 & n6871 ) | ( ~n2543 & n6871 ) ;
  assign n7083 = ( n1653 & n1869 ) | ( n1653 & n4639 ) | ( n1869 & n4639 ) ;
  assign n7084 = n3874 ^ n1370 ^ n959 ;
  assign n7086 = n3326 ^ n833 ^ n646 ;
  assign n7085 = ( n899 & n1659 ) | ( n899 & n1697 ) | ( n1659 & n1697 ) ;
  assign n7087 = n7086 ^ n7085 ^ n2516 ;
  assign n7088 = ( n7083 & ~n7084 ) | ( n7083 & n7087 ) | ( ~n7084 & n7087 ) ;
  assign n7089 = n7051 ^ n4612 ^ n576 ;
  assign n7090 = n3804 ^ n2205 ^ n1675 ;
  assign n7091 = n3265 ^ n2988 ^ n1664 ;
  assign n7092 = ( ~n849 & n7090 ) | ( ~n849 & n7091 ) | ( n7090 & n7091 ) ;
  assign n7093 = n7092 ^ n4012 ^ n1473 ;
  assign n7094 = n7093 ^ n1178 ^ n1119 ;
  assign n7095 = ( ~n7088 & n7089 ) | ( ~n7088 & n7094 ) | ( n7089 & n7094 ) ;
  assign n7099 = n1656 ^ n508 ^ n374 ;
  assign n7097 = ( ~n1052 & n1611 ) | ( ~n1052 & n4451 ) | ( n1611 & n4451 ) ;
  assign n7098 = ( n640 & n6033 ) | ( n640 & ~n7097 ) | ( n6033 & ~n7097 ) ;
  assign n7096 = n2744 ^ n1880 ^ x80 ;
  assign n7100 = n7099 ^ n7098 ^ n7096 ;
  assign n7101 = ( n5348 & ~n7095 ) | ( n5348 & n7100 ) | ( ~n7095 & n7100 ) ;
  assign n7108 = n1080 ^ n835 ^ n702 ;
  assign n7109 = n7108 ^ n1874 ^ n1040 ;
  assign n7110 = n7109 ^ n2937 ^ n1739 ;
  assign n7105 = ( n414 & n3323 ) | ( n414 & ~n4140 ) | ( n3323 & ~n4140 ) ;
  assign n7106 = n7105 ^ n5110 ^ n4000 ;
  assign n7107 = ( n1514 & n2202 ) | ( n1514 & n7106 ) | ( n2202 & n7106 ) ;
  assign n7102 = n6583 ^ n6405 ^ n3952 ;
  assign n7103 = n7102 ^ n4327 ^ n2906 ;
  assign n7104 = n7103 ^ n6666 ^ n5690 ;
  assign n7111 = n7110 ^ n7107 ^ n7104 ;
  assign n7112 = ( n818 & n892 ) | ( n818 & ~n1819 ) | ( n892 & ~n1819 ) ;
  assign n7113 = ( n1440 & n4747 ) | ( n1440 & n7112 ) | ( n4747 & n7112 ) ;
  assign n7114 = n2632 ^ n874 ^ n285 ;
  assign n7115 = ( n735 & ~n908 ) | ( n735 & n1090 ) | ( ~n908 & n1090 ) ;
  assign n7116 = ( n4675 & n7114 ) | ( n4675 & n7115 ) | ( n7114 & n7115 ) ;
  assign n7120 = n3702 ^ n2347 ^ n2247 ;
  assign n7117 = ( ~n1181 & n1502 ) | ( ~n1181 & n7015 ) | ( n1502 & n7015 ) ;
  assign n7118 = ( x37 & n690 ) | ( x37 & ~n7117 ) | ( n690 & ~n7117 ) ;
  assign n7119 = ( n1683 & ~n3706 ) | ( n1683 & n7118 ) | ( ~n3706 & n7118 ) ;
  assign n7121 = n7120 ^ n7119 ^ n2412 ;
  assign n7122 = ( n7113 & ~n7116 ) | ( n7113 & n7121 ) | ( ~n7116 & n7121 ) ;
  assign n7124 = n6773 ^ n1149 ^ n288 ;
  assign n7125 = n7124 ^ n1135 ^ n603 ;
  assign n7123 = ( n1393 & n1612 ) | ( n1393 & n4762 ) | ( n1612 & n4762 ) ;
  assign n7126 = n7125 ^ n7123 ^ n5259 ;
  assign n7127 = n7126 ^ n6953 ^ n193 ;
  assign n7128 = ( n4016 & n6085 ) | ( n4016 & ~n6555 ) | ( n6085 & ~n6555 ) ;
  assign n7136 = ( n194 & n740 ) | ( n194 & ~n899 ) | ( n740 & ~n899 ) ;
  assign n7137 = ( n321 & n1609 ) | ( n321 & n7136 ) | ( n1609 & n7136 ) ;
  assign n7134 = n2910 ^ n1179 ^ n1068 ;
  assign n7132 = ( ~n2282 & n2948 ) | ( ~n2282 & n3041 ) | ( n2948 & n3041 ) ;
  assign n7133 = ( n2880 & n5582 ) | ( n2880 & n7132 ) | ( n5582 & n7132 ) ;
  assign n7130 = ( n1530 & n4593 ) | ( n1530 & ~n6658 ) | ( n4593 & ~n6658 ) ;
  assign n7131 = n7130 ^ n6270 ^ n1798 ;
  assign n7135 = n7134 ^ n7133 ^ n7131 ;
  assign n7129 = n4241 ^ n3710 ^ x67 ;
  assign n7138 = n7137 ^ n7135 ^ n7129 ;
  assign n7139 = n5189 ^ n2568 ^ x92 ;
  assign n7140 = ( ~n424 & n1273 ) | ( ~n424 & n2711 ) | ( n1273 & n2711 ) ;
  assign n7141 = n7140 ^ n6367 ^ n4472 ;
  assign n7154 = ( n754 & n1242 ) | ( n754 & n6645 ) | ( n1242 & n6645 ) ;
  assign n7152 = n1594 ^ n485 ^ x83 ;
  assign n7150 = ( n288 & ~n957 ) | ( n288 & n1817 ) | ( ~n957 & n1817 ) ;
  assign n7151 = n7150 ^ n6018 ^ n1657 ;
  assign n7153 = n7152 ^ n7151 ^ n6561 ;
  assign n7155 = n7154 ^ n7153 ^ n3310 ;
  assign n7148 = n4861 ^ n4092 ^ n3247 ;
  assign n7149 = n7148 ^ n5489 ^ n3467 ;
  assign n7145 = ( ~n545 & n935 ) | ( ~n545 & n3345 ) | ( n935 & n3345 ) ;
  assign n7146 = n7145 ^ n2597 ^ n2055 ;
  assign n7143 = ( n219 & n1279 ) | ( n219 & n2354 ) | ( n1279 & n2354 ) ;
  assign n7144 = n7143 ^ n2869 ^ x79 ;
  assign n7142 = n6017 ^ n2973 ^ n897 ;
  assign n7147 = n7146 ^ n7144 ^ n7142 ;
  assign n7156 = n7155 ^ n7149 ^ n7147 ;
  assign n7157 = n7156 ^ n5598 ^ n2460 ;
  assign n7158 = ( n683 & ~n703 ) | ( n683 & n2358 ) | ( ~n703 & n2358 ) ;
  assign n7159 = ( n410 & n5314 ) | ( n410 & ~n6012 ) | ( n5314 & ~n6012 ) ;
  assign n7160 = ( ~n5484 & n7158 ) | ( ~n5484 & n7159 ) | ( n7158 & n7159 ) ;
  assign n7161 = n7160 ^ n3418 ^ n1146 ;
  assign n7162 = ( n2141 & n2482 ) | ( n2141 & ~n5377 ) | ( n2482 & ~n5377 ) ;
  assign n7163 = ( ~n3100 & n6784 ) | ( ~n3100 & n7162 ) | ( n6784 & n7162 ) ;
  assign n7164 = ( n456 & n1300 ) | ( n456 & n2241 ) | ( n1300 & n2241 ) ;
  assign n7165 = n5734 ^ n5727 ^ n239 ;
  assign n7166 = ( n6162 & n7164 ) | ( n6162 & ~n7165 ) | ( n7164 & ~n7165 ) ;
  assign n7167 = ( n7161 & n7163 ) | ( n7161 & ~n7166 ) | ( n7163 & ~n7166 ) ;
  assign n7168 = ( ~n385 & n927 ) | ( ~n385 & n1315 ) | ( n927 & n1315 ) ;
  assign n7169 = n7168 ^ n3738 ^ n1112 ;
  assign n7170 = n3832 ^ n1066 ^ n159 ;
  assign n7171 = ( n6019 & ~n6534 ) | ( n6019 & n7170 ) | ( ~n6534 & n7170 ) ;
  assign n7172 = ( n4536 & n6700 ) | ( n4536 & ~n7171 ) | ( n6700 & ~n7171 ) ;
  assign n7173 = n6773 ^ n2025 ^ n1054 ;
  assign n7174 = n5963 ^ n4461 ^ n395 ;
  assign n7175 = ( n4056 & n7173 ) | ( n4056 & n7174 ) | ( n7173 & n7174 ) ;
  assign n7176 = ( n6955 & ~n7172 ) | ( n6955 & n7175 ) | ( ~n7172 & n7175 ) ;
  assign n7177 = ( n2611 & n5581 ) | ( n2611 & n5700 ) | ( n5581 & n5700 ) ;
  assign n7178 = n7177 ^ n3633 ^ n1413 ;
  assign n7179 = ( n7169 & n7176 ) | ( n7169 & ~n7178 ) | ( n7176 & ~n7178 ) ;
  assign n7187 = ( n922 & n2622 ) | ( n922 & ~n4144 ) | ( n2622 & ~n4144 ) ;
  assign n7188 = ( ~n956 & n1152 ) | ( ~n956 & n2282 ) | ( n1152 & n2282 ) ;
  assign n7189 = n7188 ^ n5765 ^ n5538 ;
  assign n7190 = ( n271 & n3861 ) | ( n271 & n6315 ) | ( n3861 & n6315 ) ;
  assign n7191 = n7190 ^ n4265 ^ n742 ;
  assign n7192 = ( ~n7187 & n7189 ) | ( ~n7187 & n7191 ) | ( n7189 & n7191 ) ;
  assign n7184 = n3093 ^ n2250 ^ x59 ;
  assign n7180 = ( x116 & n794 ) | ( x116 & ~n1222 ) | ( n794 & ~n1222 ) ;
  assign n7181 = ( n1418 & n1988 ) | ( n1418 & ~n7180 ) | ( n1988 & ~n7180 ) ;
  assign n7182 = ( n3181 & n4200 ) | ( n3181 & n7181 ) | ( n4200 & n7181 ) ;
  assign n7183 = n7182 ^ n4332 ^ x0 ;
  assign n7185 = n7184 ^ n7183 ^ n5180 ;
  assign n7186 = n7185 ^ n6107 ^ n237 ;
  assign n7193 = n7192 ^ n7186 ^ n5175 ;
  assign n7194 = ( n190 & n1047 ) | ( n190 & ~n6798 ) | ( n1047 & ~n6798 ) ;
  assign n7195 = ( n1059 & n4973 ) | ( n1059 & n6320 ) | ( n4973 & n6320 ) ;
  assign n7199 = n3651 ^ n2760 ^ x49 ;
  assign n7197 = ( n3528 & ~n3952 ) | ( n3528 & n4793 ) | ( ~n3952 & n4793 ) ;
  assign n7196 = n6594 ^ n3593 ^ n1211 ;
  assign n7198 = n7197 ^ n7196 ^ n1481 ;
  assign n7200 = n7199 ^ n7198 ^ n619 ;
  assign n7201 = ( n7194 & n7195 ) | ( n7194 & ~n7200 ) | ( n7195 & ~n7200 ) ;
  assign n7202 = n7201 ^ n2671 ^ n393 ;
  assign n7203 = n7202 ^ n6412 ^ n1231 ;
  assign n7207 = n3481 ^ n3152 ^ n3025 ;
  assign n7204 = n3812 ^ n964 ^ n907 ;
  assign n7205 = ( n3288 & n4256 ) | ( n3288 & ~n7204 ) | ( n4256 & ~n7204 ) ;
  assign n7206 = ( n4517 & ~n5373 ) | ( n4517 & n7205 ) | ( ~n5373 & n7205 ) ;
  assign n7208 = n7207 ^ n7206 ^ n1905 ;
  assign n7210 = ( n1911 & ~n2495 ) | ( n1911 & n3648 ) | ( ~n2495 & n3648 ) ;
  assign n7211 = ( n2138 & ~n2161 ) | ( n2138 & n7210 ) | ( ~n2161 & n7210 ) ;
  assign n7209 = n3733 ^ n3719 ^ n619 ;
  assign n7212 = n7211 ^ n7209 ^ n4873 ;
  assign n7213 = ( n137 & ~n761 ) | ( n137 & n7212 ) | ( ~n761 & n7212 ) ;
  assign n7225 = ( n762 & n1929 ) | ( n762 & n6046 ) | ( n1929 & n6046 ) ;
  assign n7226 = n7225 ^ n4611 ^ n2879 ;
  assign n7214 = n3860 ^ n2241 ^ n1133 ;
  assign n7215 = n7214 ^ n893 ^ n594 ;
  assign n7216 = n7215 ^ n4424 ^ n1511 ;
  assign n7217 = ( n476 & n584 ) | ( n476 & ~n1461 ) | ( n584 & ~n1461 ) ;
  assign n7218 = n7217 ^ n2480 ^ n816 ;
  assign n7219 = n7218 ^ n5952 ^ n4382 ;
  assign n7220 = n7219 ^ n4808 ^ n3249 ;
  assign n7221 = n7220 ^ n3198 ^ x110 ;
  assign n7222 = n6711 ^ n5164 ^ n915 ;
  assign n7223 = ( n7216 & n7221 ) | ( n7216 & ~n7222 ) | ( n7221 & ~n7222 ) ;
  assign n7224 = n7223 ^ n2994 ^ n2278 ;
  assign n7227 = n7226 ^ n7224 ^ n1828 ;
  assign n7228 = n4900 ^ n544 ^ n323 ;
  assign n7229 = ( x84 & n678 ) | ( x84 & n1917 ) | ( n678 & n1917 ) ;
  assign n7230 = ( n1987 & ~n2958 ) | ( n1987 & n7229 ) | ( ~n2958 & n7229 ) ;
  assign n7231 = n7017 ^ n748 ^ n515 ;
  assign n7232 = n7231 ^ n751 ^ n703 ;
  assign n7233 = ( n7228 & n7230 ) | ( n7228 & ~n7232 ) | ( n7230 & ~n7232 ) ;
  assign n7234 = n6512 ^ n4597 ^ n3742 ;
  assign n7235 = ( n2610 & ~n3388 ) | ( n2610 & n5583 ) | ( ~n3388 & n5583 ) ;
  assign n7236 = ( ~x92 & n3593 ) | ( ~x92 & n7235 ) | ( n3593 & n7235 ) ;
  assign n7237 = ( n383 & n2137 ) | ( n383 & ~n7189 ) | ( n2137 & ~n7189 ) ;
  assign n7242 = n2315 ^ n1354 ^ n636 ;
  assign n7243 = ( ~n2252 & n6826 ) | ( ~n2252 & n7242 ) | ( n6826 & n7242 ) ;
  assign n7238 = ( n704 & n1376 ) | ( n704 & n2649 ) | ( n1376 & n2649 ) ;
  assign n7239 = ( n2236 & n3655 ) | ( n2236 & n7238 ) | ( n3655 & n7238 ) ;
  assign n7240 = ( n3495 & ~n5109 ) | ( n3495 & n7239 ) | ( ~n5109 & n7239 ) ;
  assign n7241 = n7240 ^ n5312 ^ n4332 ;
  assign n7244 = n7243 ^ n7241 ^ n2537 ;
  assign n7245 = ( n2202 & n2241 ) | ( n2202 & ~n3476 ) | ( n2241 & ~n3476 ) ;
  assign n7246 = ( ~n166 & n185 ) | ( ~n166 & n7245 ) | ( n185 & n7245 ) ;
  assign n7247 = n7246 ^ n3071 ^ n871 ;
  assign n7248 = ( n411 & ~n5252 ) | ( n411 & n7247 ) | ( ~n5252 & n7247 ) ;
  assign n7249 = ( ~n4539 & n6243 ) | ( ~n4539 & n7248 ) | ( n6243 & n7248 ) ;
  assign n7252 = ( n1982 & ~n2115 ) | ( n1982 & n2484 ) | ( ~n2115 & n2484 ) ;
  assign n7253 = ( n612 & n2264 ) | ( n612 & n7252 ) | ( n2264 & n7252 ) ;
  assign n7250 = n4918 ^ n737 ^ n681 ;
  assign n7251 = n7250 ^ n3298 ^ n1501 ;
  assign n7254 = n7253 ^ n7251 ^ n2292 ;
  assign n7255 = n2948 ^ n1625 ^ n1273 ;
  assign n7256 = ( n575 & ~n3960 ) | ( n575 & n5263 ) | ( ~n3960 & n5263 ) ;
  assign n7257 = ( n258 & n7255 ) | ( n258 & ~n7256 ) | ( n7255 & ~n7256 ) ;
  assign n7258 = ( n2773 & n7254 ) | ( n2773 & ~n7257 ) | ( n7254 & ~n7257 ) ;
  assign n7259 = n3928 ^ n3858 ^ n2459 ;
  assign n7264 = ( n416 & n459 ) | ( n416 & n2487 ) | ( n459 & n2487 ) ;
  assign n7265 = ( n1081 & n3752 ) | ( n1081 & ~n7264 ) | ( n3752 & ~n7264 ) ;
  assign n7266 = ( n1954 & n2022 ) | ( n1954 & n7265 ) | ( n2022 & n7265 ) ;
  assign n7260 = n6080 ^ n5440 ^ n620 ;
  assign n7261 = n7260 ^ n1363 ^ n695 ;
  assign n7262 = ( ~n955 & n988 ) | ( ~n955 & n7261 ) | ( n988 & n7261 ) ;
  assign n7263 = ( n293 & n2260 ) | ( n293 & n7262 ) | ( n2260 & n7262 ) ;
  assign n7267 = n7266 ^ n7263 ^ n1962 ;
  assign n7268 = n7267 ^ n6016 ^ n4237 ;
  assign n7269 = ( x8 & n2006 ) | ( x8 & n4840 ) | ( n2006 & n4840 ) ;
  assign n7270 = n7269 ^ n1207 ^ n988 ;
  assign n7271 = ( ~n2399 & n3678 ) | ( ~n2399 & n5425 ) | ( n3678 & n5425 ) ;
  assign n7276 = ( n523 & n2051 ) | ( n523 & n3048 ) | ( n2051 & n3048 ) ;
  assign n7277 = n7276 ^ n3969 ^ n3781 ;
  assign n7274 = ( n1869 & n1990 ) | ( n1869 & ~n5785 ) | ( n1990 & ~n5785 ) ;
  assign n7272 = ( n1206 & n2248 ) | ( n1206 & n3150 ) | ( n2248 & n3150 ) ;
  assign n7273 = n7272 ^ n3757 ^ n905 ;
  assign n7275 = n7274 ^ n7273 ^ n6568 ;
  assign n7278 = n7277 ^ n7275 ^ n1149 ;
  assign n7279 = ( n7270 & n7271 ) | ( n7270 & ~n7278 ) | ( n7271 & ~n7278 ) ;
  assign n7280 = ( n552 & ~n3728 ) | ( n552 & n4112 ) | ( ~n3728 & n4112 ) ;
  assign n7281 = n7280 ^ n3655 ^ n3493 ;
  assign n7282 = n5966 ^ n4255 ^ n3319 ;
  assign n7283 = ( n6123 & ~n7281 ) | ( n6123 & n7282 ) | ( ~n7281 & n7282 ) ;
  assign n7284 = n7283 ^ n2826 ^ n1419 ;
  assign n7285 = ( n356 & n2663 ) | ( n356 & n4495 ) | ( n2663 & n4495 ) ;
  assign n7286 = n7285 ^ n5197 ^ n3563 ;
  assign n7287 = n4543 ^ n886 ^ x42 ;
  assign n7288 = n4868 ^ n3211 ^ n3045 ;
  assign n7289 = ( x16 & n202 ) | ( x16 & ~n7288 ) | ( n202 & ~n7288 ) ;
  assign n7290 = ( n3114 & ~n7287 ) | ( n3114 & n7289 ) | ( ~n7287 & n7289 ) ;
  assign n7291 = ( n3549 & n5525 ) | ( n3549 & n6367 ) | ( n5525 & n6367 ) ;
  assign n7292 = ( ~n818 & n2548 ) | ( ~n818 & n4484 ) | ( n2548 & n4484 ) ;
  assign n7293 = ( n2399 & n2664 ) | ( n2399 & ~n7292 ) | ( n2664 & ~n7292 ) ;
  assign n7294 = ( n4595 & n5594 ) | ( n4595 & n6936 ) | ( n5594 & n6936 ) ;
  assign n7296 = ( x2 & n1668 ) | ( x2 & ~n3581 ) | ( n1668 & ~n3581 ) ;
  assign n7297 = n7296 ^ n3806 ^ n1753 ;
  assign n7298 = n7297 ^ n3601 ^ n2916 ;
  assign n7295 = n1753 ^ n1644 ^ n1440 ;
  assign n7299 = n7298 ^ n7295 ^ n581 ;
  assign n7300 = n4092 ^ n2685 ^ n521 ;
  assign n7301 = n7300 ^ n3589 ^ n2886 ;
  assign n7302 = ( ~n2601 & n5754 ) | ( ~n2601 & n7301 ) | ( n5754 & n7301 ) ;
  assign n7303 = n7302 ^ n1910 ^ n958 ;
  assign n7304 = ( n7294 & n7299 ) | ( n7294 & ~n7303 ) | ( n7299 & ~n7303 ) ;
  assign n7305 = ( n454 & n1712 ) | ( n454 & n7304 ) | ( n1712 & n7304 ) ;
  assign n7306 = ( n2609 & n3219 ) | ( n2609 & n5173 ) | ( n3219 & n5173 ) ;
  assign n7307 = ( ~n1074 & n3863 ) | ( ~n1074 & n7306 ) | ( n3863 & n7306 ) ;
  assign n7308 = ( n2445 & ~n3864 ) | ( n2445 & n7307 ) | ( ~n3864 & n7307 ) ;
  assign n7309 = n7308 ^ n6484 ^ n3820 ;
  assign n7333 = n6723 ^ n4531 ^ n1867 ;
  assign n7334 = ( ~n2033 & n2391 ) | ( ~n2033 & n5724 ) | ( n2391 & n5724 ) ;
  assign n7335 = ( n442 & ~n3722 ) | ( n442 & n7334 ) | ( ~n3722 & n7334 ) ;
  assign n7336 = n6094 ^ n2588 ^ n667 ;
  assign n7337 = n7336 ^ n5791 ^ n2225 ;
  assign n7338 = ( n793 & ~n3345 ) | ( n793 & n7337 ) | ( ~n3345 & n7337 ) ;
  assign n7339 = ( n5432 & n7335 ) | ( n5432 & n7338 ) | ( n7335 & n7338 ) ;
  assign n7340 = ( n6258 & n7333 ) | ( n6258 & ~n7339 ) | ( n7333 & ~n7339 ) ;
  assign n7311 = n2370 ^ n1099 ^ n1078 ;
  assign n7312 = ( x80 & n2996 ) | ( x80 & n7311 ) | ( n2996 & n7311 ) ;
  assign n7313 = n7312 ^ n3553 ^ n2552 ;
  assign n7310 = ( x6 & n182 ) | ( x6 & n460 ) | ( n182 & n460 ) ;
  assign n7314 = n7313 ^ n7310 ^ n1835 ;
  assign n7315 = n7314 ^ n1981 ^ x74 ;
  assign n7316 = ( ~n4260 & n6161 ) | ( ~n4260 & n7315 ) | ( n6161 & n7315 ) ;
  assign n7317 = n6651 ^ n1629 ^ n1450 ;
  assign n7318 = n7317 ^ n6316 ^ n1452 ;
  assign n7319 = n6193 ^ n4723 ^ n1072 ;
  assign n7320 = n7319 ^ n1532 ^ n1044 ;
  assign n7322 = ( n588 & n3181 ) | ( n588 & n6589 ) | ( n3181 & n6589 ) ;
  assign n7323 = n7322 ^ n5961 ^ n1770 ;
  assign n7324 = ( ~n688 & n1030 ) | ( ~n688 & n7323 ) | ( n1030 & n7323 ) ;
  assign n7321 = ( n932 & ~n1968 ) | ( n932 & n4833 ) | ( ~n1968 & n4833 ) ;
  assign n7325 = n7324 ^ n7321 ^ n2249 ;
  assign n7326 = ( x59 & n2222 ) | ( x59 & n3124 ) | ( n2222 & n3124 ) ;
  assign n7327 = ( x11 & n719 ) | ( x11 & ~n7326 ) | ( n719 & ~n7326 ) ;
  assign n7328 = ( ~n1312 & n1910 ) | ( ~n1312 & n7327 ) | ( n1910 & n7327 ) ;
  assign n7329 = n7328 ^ n3785 ^ n669 ;
  assign n7330 = ( n7320 & n7325 ) | ( n7320 & n7329 ) | ( n7325 & n7329 ) ;
  assign n7331 = ( n7316 & ~n7318 ) | ( n7316 & n7330 ) | ( ~n7318 & n7330 ) ;
  assign n7332 = ( n5958 & ~n7120 ) | ( n5958 & n7331 ) | ( ~n7120 & n7331 ) ;
  assign n7341 = n7340 ^ n7332 ^ n5862 ;
  assign n7342 = ( ~n474 & n3886 ) | ( ~n474 & n5544 ) | ( n3886 & n5544 ) ;
  assign n7343 = n5515 ^ n5383 ^ n202 ;
  assign n7344 = n3463 ^ n1691 ^ n603 ;
  assign n7345 = ( n1868 & n3710 ) | ( n1868 & ~n7344 ) | ( n3710 & ~n7344 ) ;
  assign n7346 = ( n2385 & n6615 ) | ( n2385 & ~n7345 ) | ( n6615 & ~n7345 ) ;
  assign n7347 = ( n2929 & ~n4084 ) | ( n2929 & n4542 ) | ( ~n4084 & n4542 ) ;
  assign n7348 = ( x2 & n2371 ) | ( x2 & n7347 ) | ( n2371 & n7347 ) ;
  assign n7349 = ( n1994 & n5004 ) | ( n1994 & n7348 ) | ( n5004 & n7348 ) ;
  assign n7350 = ( n4490 & ~n7346 ) | ( n4490 & n7349 ) | ( ~n7346 & n7349 ) ;
  assign n7351 = ( n7342 & ~n7343 ) | ( n7342 & n7350 ) | ( ~n7343 & n7350 ) ;
  assign n7352 = ( n2449 & n2985 ) | ( n2449 & ~n5409 ) | ( n2985 & ~n5409 ) ;
  assign n7353 = ( n2049 & ~n2972 ) | ( n2049 & n5110 ) | ( ~n2972 & n5110 ) ;
  assign n7354 = n7353 ^ n7322 ^ n5233 ;
  assign n7355 = ( n2214 & ~n5769 ) | ( n2214 & n7354 ) | ( ~n5769 & n7354 ) ;
  assign n7356 = n7355 ^ n3969 ^ n823 ;
  assign n7364 = n6798 ^ n2293 ^ n2109 ;
  assign n7357 = n1171 ^ n378 ^ x26 ;
  assign n7358 = ( n1005 & n6127 ) | ( n1005 & ~n7253 ) | ( n6127 & ~n7253 ) ;
  assign n7359 = n3606 ^ n1136 ^ n970 ;
  assign n7360 = ( n7357 & n7358 ) | ( n7357 & ~n7359 ) | ( n7358 & ~n7359 ) ;
  assign n7361 = ( n229 & n2092 ) | ( n229 & ~n5104 ) | ( n2092 & ~n5104 ) ;
  assign n7362 = n7361 ^ n335 ^ n311 ;
  assign n7363 = ( ~n7008 & n7360 ) | ( ~n7008 & n7362 ) | ( n7360 & n7362 ) ;
  assign n7365 = n7364 ^ n7363 ^ n6458 ;
  assign n7366 = ( n7352 & ~n7356 ) | ( n7352 & n7365 ) | ( ~n7356 & n7365 ) ;
  assign n7370 = n5281 ^ n1593 ^ n722 ;
  assign n7371 = ( ~x50 & n5161 ) | ( ~x50 & n7370 ) | ( n5161 & n7370 ) ;
  assign n7367 = ( ~n848 & n1619 ) | ( ~n848 & n2040 ) | ( n1619 & n2040 ) ;
  assign n7368 = ( n1455 & n2906 ) | ( n1455 & n3874 ) | ( n2906 & n3874 ) ;
  assign n7369 = ( n997 & n7367 ) | ( n997 & n7368 ) | ( n7367 & n7368 ) ;
  assign n7372 = n7371 ^ n7369 ^ n2306 ;
  assign n7373 = ( ~n1132 & n1930 ) | ( ~n1132 & n4275 ) | ( n1930 & n4275 ) ;
  assign n7380 = ( n849 & ~n1742 ) | ( n849 & n2491 ) | ( ~n1742 & n2491 ) ;
  assign n7381 = n7380 ^ n3842 ^ n729 ;
  assign n7374 = n4459 ^ n648 ^ n541 ;
  assign n7375 = ( n1753 & ~n2248 ) | ( n1753 & n7374 ) | ( ~n2248 & n7374 ) ;
  assign n7376 = ( n1886 & n6187 ) | ( n1886 & n7229 ) | ( n6187 & n7229 ) ;
  assign n7377 = n4918 ^ n1150 ^ n807 ;
  assign n7378 = ( n226 & ~n1513 ) | ( n226 & n7377 ) | ( ~n1513 & n7377 ) ;
  assign n7379 = ( n7375 & ~n7376 ) | ( n7375 & n7378 ) | ( ~n7376 & n7378 ) ;
  assign n7382 = n7381 ^ n7379 ^ n1131 ;
  assign n7383 = ( ~n338 & n2297 ) | ( ~n338 & n4897 ) | ( n2297 & n4897 ) ;
  assign n7384 = n7383 ^ n5685 ^ n3153 ;
  assign n7385 = n7384 ^ n1480 ^ n559 ;
  assign n7386 = ( n7188 & ~n7382 ) | ( n7188 & n7385 ) | ( ~n7382 & n7385 ) ;
  assign n7387 = n7386 ^ n3898 ^ n3360 ;
  assign n7399 = ( n3062 & ~n4717 ) | ( n3062 & n6635 ) | ( ~n4717 & n6635 ) ;
  assign n7395 = n7358 ^ n4952 ^ x122 ;
  assign n7396 = n7395 ^ n1402 ^ n974 ;
  assign n7394 = ( n5579 & n6300 ) | ( n5579 & n7124 ) | ( n6300 & n7124 ) ;
  assign n7397 = n7396 ^ n7394 ^ n1564 ;
  assign n7388 = n5682 ^ n1998 ^ n829 ;
  assign n7389 = ( n1437 & ~n3574 ) | ( n1437 & n7388 ) | ( ~n3574 & n7388 ) ;
  assign n7390 = ( ~n1854 & n4194 ) | ( ~n1854 & n7301 ) | ( n4194 & n7301 ) ;
  assign n7391 = ( ~n4224 & n4336 ) | ( ~n4224 & n7390 ) | ( n4336 & n7390 ) ;
  assign n7392 = ( n5227 & n7389 ) | ( n5227 & n7391 ) | ( n7389 & n7391 ) ;
  assign n7393 = ( n2160 & n6219 ) | ( n2160 & ~n7392 ) | ( n6219 & ~n7392 ) ;
  assign n7398 = n7397 ^ n7393 ^ n3244 ;
  assign n7400 = n7399 ^ n7398 ^ n209 ;
  assign n7401 = ( n232 & ~n1056 ) | ( n232 & n3131 ) | ( ~n1056 & n3131 ) ;
  assign n7402 = n7401 ^ n4325 ^ n3991 ;
  assign n7403 = ( n1059 & n2978 ) | ( n1059 & n3977 ) | ( n2978 & n3977 ) ;
  assign n7404 = ( ~n1604 & n7402 ) | ( ~n1604 & n7403 ) | ( n7402 & n7403 ) ;
  assign n7414 = n3837 ^ n2305 ^ n1262 ;
  assign n7410 = n2524 ^ n1719 ^ n196 ;
  assign n7411 = ( n4743 & n5805 ) | ( n4743 & ~n7410 ) | ( n5805 & ~n7410 ) ;
  assign n7412 = ( ~n3669 & n6116 ) | ( ~n3669 & n7411 ) | ( n6116 & n7411 ) ;
  assign n7413 = ( n772 & n3134 ) | ( n772 & n7412 ) | ( n3134 & n7412 ) ;
  assign n7405 = n2419 ^ n1114 ^ n988 ;
  assign n7406 = ( n1936 & n5955 ) | ( n1936 & ~n7405 ) | ( n5955 & ~n7405 ) ;
  assign n7407 = ( n4491 & n7015 ) | ( n4491 & n7406 ) | ( n7015 & n7406 ) ;
  assign n7408 = ( x77 & n137 ) | ( x77 & n7407 ) | ( n137 & n7407 ) ;
  assign n7409 = n7408 ^ n3675 ^ x90 ;
  assign n7415 = n7414 ^ n7413 ^ n7409 ;
  assign n7416 = ( n536 & ~n2162 ) | ( n536 & n5372 ) | ( ~n2162 & n5372 ) ;
  assign n7417 = ( n203 & n7061 ) | ( n203 & ~n7416 ) | ( n7061 & ~n7416 ) ;
  assign n7428 = n1875 ^ n999 ^ n526 ;
  assign n7424 = n6986 ^ n4936 ^ n2455 ;
  assign n7425 = n7424 ^ n6627 ^ n5401 ;
  assign n7426 = n7425 ^ n7322 ^ n4915 ;
  assign n7427 = n7426 ^ n4343 ^ n2105 ;
  assign n7429 = n7428 ^ n7427 ^ n3513 ;
  assign n7420 = n4805 ^ n2557 ^ n1496 ;
  assign n7419 = n6054 ^ n2913 ^ x32 ;
  assign n7421 = n7420 ^ n7419 ^ n1026 ;
  assign n7422 = n7421 ^ n3714 ^ n1475 ;
  assign n7418 = n5397 ^ n1510 ^ n963 ;
  assign n7423 = n7422 ^ n7418 ^ n3791 ;
  assign n7430 = n7429 ^ n7423 ^ n3914 ;
  assign n7434 = n2698 ^ n1697 ^ n520 ;
  assign n7435 = ( ~n2441 & n5445 ) | ( ~n2441 & n7434 ) | ( n5445 & n7434 ) ;
  assign n7432 = n4793 ^ n1170 ^ n1146 ;
  assign n7433 = n7432 ^ n3676 ^ n2124 ;
  assign n7436 = n7435 ^ n7433 ^ n1910 ;
  assign n7431 = n6802 ^ n3557 ^ n3317 ;
  assign n7437 = n7436 ^ n7431 ^ n6161 ;
  assign n7438 = ( n5069 & n6235 ) | ( n5069 & n7437 ) | ( n6235 & n7437 ) ;
  assign n7439 = ( ~n1932 & n3466 ) | ( ~n1932 & n7438 ) | ( n3466 & n7438 ) ;
  assign n7440 = ( ~n3552 & n6069 ) | ( ~n3552 & n7354 ) | ( n6069 & n7354 ) ;
  assign n7441 = n6213 ^ n3085 ^ n1553 ;
  assign n7442 = ( n5384 & n5936 ) | ( n5384 & ~n7441 ) | ( n5936 & ~n7441 ) ;
  assign n7443 = n7015 ^ n3449 ^ n488 ;
  assign n7444 = ( ~n2883 & n6084 ) | ( ~n2883 & n6450 ) | ( n6084 & n6450 ) ;
  assign n7445 = ( ~n2252 & n7443 ) | ( ~n2252 & n7444 ) | ( n7443 & n7444 ) ;
  assign n7446 = ( n479 & n1418 ) | ( n479 & n7445 ) | ( n1418 & n7445 ) ;
  assign n7447 = ( n2282 & n3267 ) | ( n2282 & n4931 ) | ( n3267 & n4931 ) ;
  assign n7448 = n7447 ^ n2453 ^ x102 ;
  assign n7449 = ( n457 & n872 ) | ( n457 & n2522 ) | ( n872 & n2522 ) ;
  assign n7450 = ( n4552 & ~n5151 ) | ( n4552 & n7449 ) | ( ~n5151 & n7449 ) ;
  assign n7451 = n7450 ^ n7104 ^ n1772 ;
  assign n7457 = ( n631 & ~n1027 ) | ( n631 & n2060 ) | ( ~n1027 & n2060 ) ;
  assign n7458 = ( n801 & n4232 ) | ( n801 & ~n5652 ) | ( n4232 & ~n5652 ) ;
  assign n7459 = ( n2516 & n7457 ) | ( n2516 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7460 = ( n1824 & n2131 ) | ( n1824 & ~n7459 ) | ( n2131 & ~n7459 ) ;
  assign n7461 = ( n1634 & n5664 ) | ( n1634 & ~n7460 ) | ( n5664 & ~n7460 ) ;
  assign n7452 = n2240 ^ n2027 ^ n1426 ;
  assign n7453 = ( n2954 & ~n3196 ) | ( n2954 & n3650 ) | ( ~n3196 & n3650 ) ;
  assign n7454 = n7453 ^ n621 ^ n583 ;
  assign n7455 = ( ~n5922 & n7452 ) | ( ~n5922 & n7454 ) | ( n7452 & n7454 ) ;
  assign n7456 = ( n4938 & n5350 ) | ( n4938 & n7455 ) | ( n5350 & n7455 ) ;
  assign n7462 = n7461 ^ n7456 ^ n1828 ;
  assign n7465 = ( n970 & n2314 ) | ( n970 & ~n3905 ) | ( n2314 & ~n3905 ) ;
  assign n7466 = n7465 ^ n2205 ^ n2011 ;
  assign n7463 = n7425 ^ n6609 ^ n2581 ;
  assign n7464 = ( n768 & ~n2441 ) | ( n768 & n7463 ) | ( ~n2441 & n7463 ) ;
  assign n7467 = n7466 ^ n7464 ^ n5222 ;
  assign n7473 = n6959 ^ n1076 ^ n307 ;
  assign n7471 = ( n344 & ~n6208 ) | ( n344 & n6836 ) | ( ~n6208 & n6836 ) ;
  assign n7472 = n7471 ^ n6609 ^ n1375 ;
  assign n7470 = ( n1441 & ~n1624 ) | ( n1441 & n3132 ) | ( ~n1624 & n3132 ) ;
  assign n7474 = n7473 ^ n7472 ^ n7470 ;
  assign n7475 = ( ~n1080 & n6875 ) | ( ~n1080 & n7474 ) | ( n6875 & n7474 ) ;
  assign n7476 = n7475 ^ n3271 ^ x110 ;
  assign n7469 = n3528 ^ n2354 ^ n2112 ;
  assign n7468 = n2057 ^ n1723 ^ n340 ;
  assign n7477 = n7476 ^ n7469 ^ n7468 ;
  assign n7478 = ( n2435 & n4855 ) | ( n2435 & ~n5302 ) | ( n4855 & ~n5302 ) ;
  assign n7479 = ( n3374 & n5008 ) | ( n3374 & ~n7190 ) | ( n5008 & ~n7190 ) ;
  assign n7480 = n6724 ^ n1629 ^ n129 ;
  assign n7481 = n7480 ^ n5840 ^ n557 ;
  assign n7482 = n7481 ^ n2948 ^ n1162 ;
  assign n7483 = n7482 ^ n4929 ^ n1258 ;
  assign n7484 = ( n1363 & n7479 ) | ( n1363 & n7483 ) | ( n7479 & n7483 ) ;
  assign n7485 = n7484 ^ n6189 ^ n4494 ;
  assign n7486 = ( n4029 & n6265 ) | ( n4029 & ~n7485 ) | ( n6265 & ~n7485 ) ;
  assign n7487 = n7486 ^ n6947 ^ n5857 ;
  assign n7488 = n6798 ^ n4270 ^ n1578 ;
  assign n7489 = n7488 ^ n3763 ^ n482 ;
  assign n7490 = ( n2154 & n2416 ) | ( n2154 & ~n7489 ) | ( n2416 & ~n7489 ) ;
  assign n7491 = n7490 ^ n5044 ^ n2578 ;
  assign n7492 = n7491 ^ n1803 ^ n215 ;
  assign n7494 = n1838 ^ n612 ^ x120 ;
  assign n7493 = n2547 ^ n2073 ^ n487 ;
  assign n7495 = n7494 ^ n7493 ^ n4347 ;
  assign n7496 = ( n2536 & n6071 ) | ( n2536 & n7495 ) | ( n6071 & n7495 ) ;
  assign n7497 = n1785 ^ n1749 ^ n509 ;
  assign n7498 = ( n151 & n2660 ) | ( n151 & ~n4549 ) | ( n2660 & ~n4549 ) ;
  assign n7499 = n7498 ^ n3382 ^ n3367 ;
  assign n7500 = n7499 ^ n2918 ^ n412 ;
  assign n7501 = ( ~n506 & n7497 ) | ( ~n506 & n7500 ) | ( n7497 & n7500 ) ;
  assign n7502 = ( ~n3765 & n5334 ) | ( ~n3765 & n7501 ) | ( n5334 & n7501 ) ;
  assign n7503 = n7502 ^ n5221 ^ n311 ;
  assign n7504 = n7503 ^ n5262 ^ n4481 ;
  assign n7510 = n3087 ^ n2874 ^ n1012 ;
  assign n7511 = ( n422 & n2263 ) | ( n422 & ~n7510 ) | ( n2263 & ~n7510 ) ;
  assign n7509 = n3839 ^ n2508 ^ n1087 ;
  assign n7512 = n7511 ^ n7509 ^ n3856 ;
  assign n7513 = n7512 ^ n1659 ^ n589 ;
  assign n7505 = n2028 ^ n1676 ^ n937 ;
  assign n7506 = ( n3481 & n4152 ) | ( n3481 & ~n7505 ) | ( n4152 & ~n7505 ) ;
  assign n7507 = ( n4265 & n6201 ) | ( n4265 & n7506 ) | ( n6201 & n7506 ) ;
  assign n7508 = ( n3273 & n4905 ) | ( n3273 & ~n7507 ) | ( n4905 & ~n7507 ) ;
  assign n7514 = n7513 ^ n7508 ^ n5342 ;
  assign n7517 = n7509 ^ n3130 ^ n1531 ;
  assign n7518 = ( ~n2314 & n7180 ) | ( ~n2314 & n7517 ) | ( n7180 & n7517 ) ;
  assign n7515 = ( n366 & n1624 ) | ( n366 & n2793 ) | ( n1624 & n2793 ) ;
  assign n7516 = ( n2480 & n7323 ) | ( n2480 & n7515 ) | ( n7323 & n7515 ) ;
  assign n7519 = n7518 ^ n7516 ^ n4614 ;
  assign n7520 = n3240 ^ n3004 ^ n1411 ;
  assign n7521 = ( n1010 & ~n2861 ) | ( n1010 & n7520 ) | ( ~n2861 & n7520 ) ;
  assign n7523 = ( x1 & n1323 ) | ( x1 & n2208 ) | ( n1323 & n2208 ) ;
  assign n7522 = n3364 ^ n2121 ^ n528 ;
  assign n7524 = n7523 ^ n7522 ^ n5104 ;
  assign n7525 = n5403 ^ n356 ^ n281 ;
  assign n7526 = n7525 ^ n5460 ^ n1722 ;
  assign n7527 = ( n3196 & n4738 ) | ( n3196 & ~n7526 ) | ( n4738 & ~n7526 ) ;
  assign n7528 = ( n2098 & n5090 ) | ( n2098 & ~n7189 ) | ( n5090 & ~n7189 ) ;
  assign n7530 = n7070 ^ n2139 ^ n1293 ;
  assign n7531 = n7530 ^ n5135 ^ n592 ;
  assign n7532 = n7531 ^ n4915 ^ n1792 ;
  assign n7529 = ( n813 & ~n3832 ) | ( n813 & n4743 ) | ( ~n3832 & n4743 ) ;
  assign n7533 = n7532 ^ n7529 ^ n3281 ;
  assign n7534 = ( ~n6097 & n7528 ) | ( ~n6097 & n7533 ) | ( n7528 & n7533 ) ;
  assign n7535 = ( n1925 & n2311 ) | ( n1925 & ~n7534 ) | ( n2311 & ~n7534 ) ;
  assign n7537 = ( n342 & n1832 ) | ( n342 & n2448 ) | ( n1832 & n2448 ) ;
  assign n7538 = n7537 ^ n2848 ^ n2476 ;
  assign n7536 = ( ~n1915 & n3150 ) | ( ~n1915 & n6940 ) | ( n3150 & n6940 ) ;
  assign n7539 = n7538 ^ n7536 ^ n1766 ;
  assign n7540 = ( n2720 & n3167 ) | ( n2720 & ~n7539 ) | ( n3167 & ~n7539 ) ;
  assign n7544 = n2389 ^ n1923 ^ n1001 ;
  assign n7545 = ( n3808 & ~n6905 ) | ( n3808 & n7544 ) | ( ~n6905 & n7544 ) ;
  assign n7541 = n3110 ^ n3007 ^ n1424 ;
  assign n7542 = n7541 ^ n3073 ^ n229 ;
  assign n7543 = ( n2093 & ~n4746 ) | ( n2093 & n7542 ) | ( ~n4746 & n7542 ) ;
  assign n7546 = n7545 ^ n7543 ^ n4514 ;
  assign n7547 = ( n202 & n1473 ) | ( n202 & ~n2201 ) | ( n1473 & ~n2201 ) ;
  assign n7548 = n4926 ^ n1995 ^ n433 ;
  assign n7549 = ( ~n4559 & n5105 ) | ( ~n4559 & n7548 ) | ( n5105 & n7548 ) ;
  assign n7550 = n7549 ^ n2577 ^ n1740 ;
  assign n7551 = n3775 ^ n2466 ^ n540 ;
  assign n7552 = ( n2407 & ~n4217 ) | ( n2407 & n7551 ) | ( ~n4217 & n7551 ) ;
  assign n7553 = ( ~n7547 & n7550 ) | ( ~n7547 & n7552 ) | ( n7550 & n7552 ) ;
  assign n7554 = n3294 ^ n2399 ^ n2370 ;
  assign n7555 = n7554 ^ n5904 ^ n2550 ;
  assign n7556 = n7555 ^ n4259 ^ n4105 ;
  assign n7557 = n2565 ^ n293 ^ n259 ;
  assign n7558 = ( ~n2430 & n3814 ) | ( ~n2430 & n7557 ) | ( n3814 & n7557 ) ;
  assign n7559 = ( n1696 & n7124 ) | ( n1696 & ~n7558 ) | ( n7124 & ~n7558 ) ;
  assign n7560 = n7559 ^ n5557 ^ n4002 ;
  assign n7561 = n5059 ^ n3246 ^ n2168 ;
  assign n7562 = ( n1670 & n3058 ) | ( n1670 & n5698 ) | ( n3058 & n5698 ) ;
  assign n7563 = ( ~n5317 & n5952 ) | ( ~n5317 & n7562 ) | ( n5952 & n7562 ) ;
  assign n7564 = ( n726 & n2975 ) | ( n726 & ~n7563 ) | ( n2975 & ~n7563 ) ;
  assign n7565 = ( n5527 & n7561 ) | ( n5527 & ~n7564 ) | ( n7561 & ~n7564 ) ;
  assign n7566 = ( n164 & n951 ) | ( n164 & n4069 ) | ( n951 & n4069 ) ;
  assign n7567 = ( ~n7560 & n7565 ) | ( ~n7560 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7568 = ( n5893 & n7556 ) | ( n5893 & ~n7567 ) | ( n7556 & ~n7567 ) ;
  assign n7569 = ( x20 & n282 ) | ( x20 & n2591 ) | ( n282 & n2591 ) ;
  assign n7570 = ( n1586 & ~n2346 ) | ( n1586 & n5428 ) | ( ~n2346 & n5428 ) ;
  assign n7571 = n7570 ^ n5628 ^ n2633 ;
  assign n7572 = n7388 ^ n6396 ^ n777 ;
  assign n7573 = ( n7569 & n7571 ) | ( n7569 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = ( n609 & n780 ) | ( n609 & ~n918 ) | ( n780 & ~n918 ) ;
  assign n7575 = n7574 ^ n3362 ^ n1065 ;
  assign n7577 = ( n2520 & ~n3217 ) | ( n2520 & n5293 ) | ( ~n3217 & n5293 ) ;
  assign n7576 = ( n828 & n1190 ) | ( n828 & ~n2203 ) | ( n1190 & ~n2203 ) ;
  assign n7578 = n7577 ^ n7576 ^ n2029 ;
  assign n7579 = n7578 ^ n5061 ^ n601 ;
  assign n7580 = ( n7573 & n7575 ) | ( n7573 & n7579 ) | ( n7575 & n7579 ) ;
  assign n7582 = ( n1544 & ~n2450 ) | ( n1544 & n2685 ) | ( ~n2450 & n2685 ) ;
  assign n7583 = n7582 ^ n5826 ^ n3039 ;
  assign n7581 = ( ~n3095 & n5436 ) | ( ~n3095 & n6859 ) | ( n5436 & n6859 ) ;
  assign n7584 = n7583 ^ n7581 ^ n3740 ;
  assign n7585 = ( n738 & ~n1197 ) | ( n738 & n2711 ) | ( ~n1197 & n2711 ) ;
  assign n7586 = n982 ^ n720 ^ n195 ;
  assign n7587 = ( n1377 & n7585 ) | ( n1377 & ~n7586 ) | ( n7585 & ~n7586 ) ;
  assign n7588 = n7180 ^ n2622 ^ x64 ;
  assign n7589 = n3624 ^ n2913 ^ n172 ;
  assign n7590 = ( ~n2400 & n7588 ) | ( ~n2400 & n7589 ) | ( n7588 & n7589 ) ;
  assign n7591 = n5245 ^ n559 ^ n346 ;
  assign n7592 = ( ~n3445 & n7590 ) | ( ~n3445 & n7591 ) | ( n7590 & n7591 ) ;
  assign n7598 = n1857 ^ n1674 ^ n532 ;
  assign n7599 = ( ~n227 & n569 ) | ( ~n227 & n7598 ) | ( n569 & n7598 ) ;
  assign n7600 = n7599 ^ n5670 ^ n771 ;
  assign n7601 = n7600 ^ n1716 ^ n562 ;
  assign n7593 = n5178 ^ n3523 ^ n2011 ;
  assign n7594 = ( n999 & ~n1542 ) | ( n999 & n7593 ) | ( ~n1542 & n7593 ) ;
  assign n7595 = n6028 ^ n5381 ^ n3699 ;
  assign n7596 = ( n1743 & n7594 ) | ( n1743 & n7595 ) | ( n7594 & n7595 ) ;
  assign n7597 = ( n3385 & n6411 ) | ( n3385 & n7596 ) | ( n6411 & n7596 ) ;
  assign n7602 = n7601 ^ n7597 ^ n5529 ;
  assign n7603 = ( n1773 & n5661 ) | ( n1773 & ~n7602 ) | ( n5661 & ~n7602 ) ;
  assign n7604 = ( n5493 & n7592 ) | ( n5493 & ~n7603 ) | ( n7592 & ~n7603 ) ;
  assign n7605 = n7604 ^ n6447 ^ n4021 ;
  assign n7609 = n3689 ^ n3137 ^ n1434 ;
  assign n7610 = n7609 ^ n3414 ^ n1339 ;
  assign n7611 = n7610 ^ n3181 ^ n1721 ;
  assign n7606 = n3306 ^ n1031 ^ n360 ;
  assign n7607 = ( n1781 & n4232 ) | ( n1781 & n4384 ) | ( n4232 & n4384 ) ;
  assign n7608 = ( n356 & n7606 ) | ( n356 & ~n7607 ) | ( n7606 & ~n7607 ) ;
  assign n7612 = n7611 ^ n7608 ^ n902 ;
  assign n7613 = ( n1379 & n1991 ) | ( n1379 & ~n5979 ) | ( n1991 & ~n5979 ) ;
  assign n7614 = ( x65 & ~n5210 ) | ( x65 & n6212 ) | ( ~n5210 & n6212 ) ;
  assign n7615 = ( n2882 & n4187 ) | ( n2882 & n7614 ) | ( n4187 & n7614 ) ;
  assign n7616 = n7615 ^ n2119 ^ n461 ;
  assign n7617 = ( ~n7612 & n7613 ) | ( ~n7612 & n7616 ) | ( n7613 & n7616 ) ;
  assign n7618 = n6651 ^ n3934 ^ n675 ;
  assign n7619 = n7618 ^ n274 ^ n191 ;
  assign n7624 = ( n700 & n4918 ) | ( n700 & n5090 ) | ( n4918 & n5090 ) ;
  assign n7621 = ( n433 & n2322 ) | ( n433 & n2418 ) | ( n2322 & n2418 ) ;
  assign n7620 = n4089 ^ n2687 ^ n915 ;
  assign n7622 = n7621 ^ n7620 ^ n414 ;
  assign n7623 = n7622 ^ n6844 ^ n1266 ;
  assign n7625 = n7624 ^ n7623 ^ n2473 ;
  assign n7626 = ( ~n6817 & n7619 ) | ( ~n6817 & n7625 ) | ( n7619 & n7625 ) ;
  assign n7632 = n2939 ^ n1857 ^ n1041 ;
  assign n7633 = n7632 ^ n7004 ^ n5787 ;
  assign n7634 = ( n1559 & ~n6175 ) | ( n1559 & n7633 ) | ( ~n6175 & n7633 ) ;
  assign n7635 = n6049 ^ n5909 ^ n2343 ;
  assign n7636 = ( n5125 & n7634 ) | ( n5125 & n7635 ) | ( n7634 & n7635 ) ;
  assign n7630 = ( n1438 & ~n3299 ) | ( n1438 & n5213 ) | ( ~n3299 & n5213 ) ;
  assign n7631 = n7630 ^ n4647 ^ n746 ;
  assign n7628 = ( n2467 & n3323 ) | ( n2467 & n4123 ) | ( n3323 & n4123 ) ;
  assign n7627 = n7482 ^ n4835 ^ n2738 ;
  assign n7629 = n7628 ^ n7627 ^ n4041 ;
  assign n7637 = n7636 ^ n7631 ^ n7629 ;
  assign n7638 = ( n1196 & n1345 ) | ( n1196 & n5055 ) | ( n1345 & n5055 ) ;
  assign n7639 = n7638 ^ n5005 ^ n4671 ;
  assign n7640 = n3496 ^ n2386 ^ x117 ;
  assign n7641 = n2527 ^ n1766 ^ n814 ;
  assign n7642 = n7641 ^ n2109 ^ n966 ;
  assign n7643 = ( ~n4587 & n6419 ) | ( ~n4587 & n7642 ) | ( n6419 & n7642 ) ;
  assign n7644 = ( ~n7216 & n7640 ) | ( ~n7216 & n7643 ) | ( n7640 & n7643 ) ;
  assign n7645 = ( n923 & n6280 ) | ( n923 & ~n7185 ) | ( n6280 & ~n7185 ) ;
  assign n7646 = n7598 ^ n2083 ^ n1177 ;
  assign n7649 = n3081 ^ n1192 ^ n448 ;
  assign n7650 = ( n3774 & n3798 ) | ( n3774 & n7649 ) | ( n3798 & n7649 ) ;
  assign n7648 = n3392 ^ n321 ^ n212 ;
  assign n7647 = ( x124 & n4275 ) | ( x124 & n7517 ) | ( n4275 & n7517 ) ;
  assign n7651 = n7650 ^ n7648 ^ n7647 ;
  assign n7652 = ( n1629 & ~n7646 ) | ( n1629 & n7651 ) | ( ~n7646 & n7651 ) ;
  assign n7653 = n5664 ^ n4416 ^ n4169 ;
  assign n7654 = ( n2648 & n3985 ) | ( n2648 & ~n4793 ) | ( n3985 & ~n4793 ) ;
  assign n7655 = ( n2656 & n3454 ) | ( n2656 & ~n7654 ) | ( n3454 & ~n7654 ) ;
  assign n7656 = ( ~n5379 & n6895 ) | ( ~n5379 & n7655 ) | ( n6895 & n7655 ) ;
  assign n7658 = n2778 ^ n1356 ^ n311 ;
  assign n7657 = ( n501 & n1424 ) | ( n501 & ~n6054 ) | ( n1424 & ~n6054 ) ;
  assign n7659 = n7658 ^ n7657 ^ n2768 ;
  assign n7660 = n7659 ^ n3438 ^ n422 ;
  assign n7661 = n7660 ^ n7618 ^ n6649 ;
  assign n7662 = n6312 ^ n6277 ^ n4286 ;
  assign n7663 = n6889 ^ n5132 ^ n1326 ;
  assign n7664 = ( n998 & n1974 ) | ( n998 & n7663 ) | ( n1974 & n7663 ) ;
  assign n7665 = n5418 ^ n3545 ^ n1260 ;
  assign n7666 = n7665 ^ n829 ^ n639 ;
  assign n7667 = n6640 ^ n1804 ^ n362 ;
  assign n7668 = n3100 ^ n141 ^ x97 ;
  assign n7669 = ( n4566 & ~n7667 ) | ( n4566 & n7668 ) | ( ~n7667 & n7668 ) ;
  assign n7670 = n7669 ^ n7589 ^ n5967 ;
  assign n7671 = n5044 ^ n3600 ^ n2211 ;
  assign n7672 = ( n1636 & ~n4498 ) | ( n1636 & n7671 ) | ( ~n4498 & n7671 ) ;
  assign n7673 = n7672 ^ n6487 ^ x115 ;
  assign n7674 = ( n1830 & n7670 ) | ( n1830 & n7673 ) | ( n7670 & n7673 ) ;
  assign n7675 = ( n4187 & ~n7666 ) | ( n4187 & n7674 ) | ( ~n7666 & n7674 ) ;
  assign n7676 = ( n6668 & n7664 ) | ( n6668 & n7675 ) | ( n7664 & n7675 ) ;
  assign n7679 = n6386 ^ n5497 ^ n750 ;
  assign n7680 = n7679 ^ n7270 ^ n1921 ;
  assign n7681 = ( n2872 & ~n3808 ) | ( n2872 & n7680 ) | ( ~n3808 & n7680 ) ;
  assign n7677 = n2461 ^ n980 ^ n730 ;
  assign n7678 = n7677 ^ n3674 ^ n2385 ;
  assign n7682 = n7681 ^ n7678 ^ n6277 ;
  assign n7688 = ( n2240 & ~n3740 ) | ( n2240 & n5316 ) | ( ~n3740 & n5316 ) ;
  assign n7689 = ( n493 & n3050 ) | ( n493 & ~n7688 ) | ( n3050 & ~n7688 ) ;
  assign n7685 = ( n937 & ~n2861 ) | ( n937 & n4382 ) | ( ~n2861 & n4382 ) ;
  assign n7686 = ( ~n1585 & n4414 ) | ( ~n1585 & n7685 ) | ( n4414 & n7685 ) ;
  assign n7687 = ( n5101 & ~n7593 ) | ( n5101 & n7686 ) | ( ~n7593 & n7686 ) ;
  assign n7683 = n4953 ^ n1239 ^ n249 ;
  assign n7684 = n7683 ^ n1284 ^ n1219 ;
  assign n7690 = n7689 ^ n7687 ^ n7684 ;
  assign n7691 = n7619 ^ n4907 ^ n4613 ;
  assign n7704 = n3831 ^ n2764 ^ n232 ;
  assign n7701 = ( ~n497 & n1901 ) | ( ~n497 & n5659 ) | ( n1901 & n5659 ) ;
  assign n7700 = ( n2440 & n3446 ) | ( n2440 & n5131 ) | ( n3446 & n5131 ) ;
  assign n7702 = n7701 ^ n7700 ^ n2657 ;
  assign n7697 = ( n2460 & ~n2553 ) | ( n2460 & n5682 ) | ( ~n2553 & n5682 ) ;
  assign n7698 = n7697 ^ n7481 ^ n170 ;
  assign n7699 = ( n3499 & n5699 ) | ( n3499 & ~n7698 ) | ( n5699 & ~n7698 ) ;
  assign n7703 = n7702 ^ n7699 ^ n328 ;
  assign n7705 = n7704 ^ n7703 ^ n1772 ;
  assign n7692 = n4953 ^ n2096 ^ n1661 ;
  assign n7693 = n7692 ^ n6356 ^ n1833 ;
  assign n7694 = ( n3166 & n3832 ) | ( n3166 & ~n5725 ) | ( n3832 & ~n5725 ) ;
  assign n7695 = ( n2532 & n3408 ) | ( n2532 & n7694 ) | ( n3408 & n7694 ) ;
  assign n7696 = ( n6193 & n7693 ) | ( n6193 & n7695 ) | ( n7693 & n7695 ) ;
  assign n7706 = n7705 ^ n7696 ^ n6240 ;
  assign n7707 = n6591 ^ n4364 ^ n695 ;
  assign n7708 = ( n599 & n7356 ) | ( n599 & ~n7707 ) | ( n7356 & ~n7707 ) ;
  assign n7709 = n5131 ^ n3645 ^ n3107 ;
  assign n7710 = n7709 ^ n4649 ^ n3149 ;
  assign n7717 = ( ~x42 & n3029 ) | ( ~x42 & n5805 ) | ( n3029 & n5805 ) ;
  assign n7711 = n3781 ^ n645 ^ x13 ;
  assign n7712 = ( n461 & ~n3307 ) | ( n461 & n5665 ) | ( ~n3307 & n5665 ) ;
  assign n7713 = ( n2584 & ~n3054 ) | ( n2584 & n7712 ) | ( ~n3054 & n7712 ) ;
  assign n7714 = n7713 ^ n7642 ^ n7425 ;
  assign n7715 = ( n199 & n4717 ) | ( n199 & ~n7714 ) | ( n4717 & ~n7714 ) ;
  assign n7716 = ( n4656 & ~n7711 ) | ( n4656 & n7715 ) | ( ~n7711 & n7715 ) ;
  assign n7718 = n7717 ^ n7716 ^ n2949 ;
  assign n7720 = ( n2488 & ~n3029 ) | ( n2488 & n3807 ) | ( ~n3029 & n3807 ) ;
  assign n7719 = ( n2964 & n3944 ) | ( n2964 & ~n5571 ) | ( n3944 & ~n5571 ) ;
  assign n7721 = n7720 ^ n7719 ^ n3149 ;
  assign n7732 = ( n445 & n4301 ) | ( n445 & n5853 ) | ( n4301 & n5853 ) ;
  assign n7727 = n3341 ^ n2995 ^ n1749 ;
  assign n7724 = ( n251 & n964 ) | ( n251 & n1624 ) | ( n964 & n1624 ) ;
  assign n7723 = ( n989 & ~n1099 ) | ( n989 & n3773 ) | ( ~n1099 & n3773 ) ;
  assign n7725 = n7724 ^ n7723 ^ n3165 ;
  assign n7726 = ( n1969 & ~n3047 ) | ( n1969 & n7725 ) | ( ~n3047 & n7725 ) ;
  assign n7722 = n4976 ^ n3903 ^ n1117 ;
  assign n7728 = n7727 ^ n7726 ^ n7722 ;
  assign n7729 = ( n2190 & n7683 ) | ( n2190 & n7728 ) | ( n7683 & n7728 ) ;
  assign n7730 = n7680 ^ n5556 ^ n2832 ;
  assign n7731 = ( n1236 & ~n7729 ) | ( n1236 & n7730 ) | ( ~n7729 & n7730 ) ;
  assign n7733 = n7732 ^ n7731 ^ n2306 ;
  assign n7734 = ( n447 & n639 ) | ( n447 & ~n704 ) | ( n639 & ~n704 ) ;
  assign n7735 = n7734 ^ n6277 ^ n5865 ;
  assign n7736 = n7672 ^ n3591 ^ n3363 ;
  assign n7737 = n6339 ^ n5607 ^ n2971 ;
  assign n7738 = ( x40 & ~n7736 ) | ( x40 & n7737 ) | ( ~n7736 & n7737 ) ;
  assign n7739 = ( n1147 & ~n4218 ) | ( n1147 & n7738 ) | ( ~n4218 & n7738 ) ;
  assign n7740 = n5511 ^ n4053 ^ n3085 ;
  assign n7741 = ( n3644 & n5560 ) | ( n3644 & n7242 ) | ( n5560 & n7242 ) ;
  assign n7742 = ( n4624 & n5573 ) | ( n4624 & n7741 ) | ( n5573 & n7741 ) ;
  assign n7743 = n7380 ^ n5842 ^ n4624 ;
  assign n7744 = ( n3755 & n7697 ) | ( n3755 & n7743 ) | ( n7697 & n7743 ) ;
  assign n7745 = n5514 ^ n4853 ^ n2039 ;
  assign n7746 = ( ~n176 & n2158 ) | ( ~n176 & n6709 ) | ( n2158 & n6709 ) ;
  assign n7747 = ( ~n7646 & n7745 ) | ( ~n7646 & n7746 ) | ( n7745 & n7746 ) ;
  assign n7748 = n7747 ^ n5857 ^ n718 ;
  assign n7749 = ( n555 & n7744 ) | ( n555 & ~n7748 ) | ( n7744 & ~n7748 ) ;
  assign n7753 = ( ~x124 & n4270 ) | ( ~x124 & n5739 ) | ( n4270 & n5739 ) ;
  assign n7754 = n7753 ^ n2126 ^ x92 ;
  assign n7755 = n7754 ^ n6429 ^ n1642 ;
  assign n7756 = n7755 ^ n6798 ^ n2821 ;
  assign n7751 = n3349 ^ n1725 ^ x15 ;
  assign n7750 = n6136 ^ n3042 ^ n2519 ;
  assign n7752 = n7751 ^ n7750 ^ n1595 ;
  assign n7757 = n7756 ^ n7752 ^ n2632 ;
  assign n7763 = n3314 ^ n2327 ^ n807 ;
  assign n7764 = n7763 ^ n2943 ^ x119 ;
  assign n7759 = ( n1133 & n1269 ) | ( n1133 & n3130 ) | ( n1269 & n3130 ) ;
  assign n7760 = n4638 ^ n1289 ^ n393 ;
  assign n7761 = ( n3273 & n7759 ) | ( n3273 & n7760 ) | ( n7759 & n7760 ) ;
  assign n7762 = n7761 ^ n6620 ^ n3647 ;
  assign n7758 = n7726 ^ n5963 ^ n1874 ;
  assign n7765 = n7764 ^ n7762 ^ n7758 ;
  assign n7769 = ( x121 & n181 ) | ( x121 & n445 ) | ( n181 & n445 ) ;
  assign n7770 = ( ~n1828 & n3774 ) | ( ~n1828 & n7769 ) | ( n3774 & n7769 ) ;
  assign n7767 = ( ~n205 & n2614 ) | ( ~n205 & n5895 ) | ( n2614 & n5895 ) ;
  assign n7766 = n7049 ^ n5831 ^ n3745 ;
  assign n7768 = n7767 ^ n7766 ^ n2072 ;
  assign n7771 = n7770 ^ n7768 ^ n1736 ;
  assign n7772 = ( n1638 & n3204 ) | ( n1638 & n7051 ) | ( n3204 & n7051 ) ;
  assign n7782 = n2007 ^ n1946 ^ n827 ;
  assign n7783 = n7782 ^ n5970 ^ n5312 ;
  assign n7779 = ( n979 & n2764 ) | ( n979 & ~n2769 ) | ( n2764 & ~n2769 ) ;
  assign n7780 = ( n2589 & n3261 ) | ( n2589 & ~n5385 ) | ( n3261 & ~n5385 ) ;
  assign n7781 = ( n6771 & n7779 ) | ( n6771 & n7780 ) | ( n7779 & n7780 ) ;
  assign n7776 = ( n903 & ~n2073 ) | ( n903 & n2387 ) | ( ~n2073 & n2387 ) ;
  assign n7777 = ( ~n235 & n3393 ) | ( ~n235 & n7776 ) | ( n3393 & n7776 ) ;
  assign n7775 = n7015 ^ n3184 ^ n1088 ;
  assign n7773 = n3972 ^ n925 ^ n881 ;
  assign n7774 = n7773 ^ n3601 ^ n3340 ;
  assign n7778 = n7777 ^ n7775 ^ n7774 ;
  assign n7784 = n7783 ^ n7781 ^ n7778 ;
  assign n7785 = ( n5168 & ~n7772 ) | ( n5168 & n7784 ) | ( ~n7772 & n7784 ) ;
  assign n7786 = n6882 ^ n6090 ^ n4771 ;
  assign n7798 = ( n2461 & ~n2735 ) | ( n2461 & n6443 ) | ( ~n2735 & n6443 ) ;
  assign n7799 = ( ~n1241 & n6623 ) | ( ~n1241 & n7798 ) | ( n6623 & n7798 ) ;
  assign n7796 = n6588 ^ n5030 ^ n2281 ;
  assign n7794 = n3740 ^ n2674 ^ n2521 ;
  assign n7792 = ( n809 & n2373 ) | ( n809 & ~n5228 ) | ( n2373 & ~n5228 ) ;
  assign n7793 = ( ~n4624 & n5782 ) | ( ~n4624 & n7792 ) | ( n5782 & n7792 ) ;
  assign n7795 = n7794 ^ n7793 ^ n5219 ;
  assign n7790 = ( n705 & n1781 ) | ( n705 & ~n3628 ) | ( n1781 & ~n3628 ) ;
  assign n7788 = n2855 ^ n2333 ^ n1153 ;
  assign n7787 = ( n1682 & n4971 ) | ( n1682 & n6030 ) | ( n4971 & n6030 ) ;
  assign n7789 = n7788 ^ n7787 ^ n7732 ;
  assign n7791 = n7790 ^ n7789 ^ n461 ;
  assign n7797 = n7796 ^ n7795 ^ n7791 ;
  assign n7800 = n7799 ^ n7797 ^ n6070 ;
  assign n7801 = n4198 ^ n3833 ^ n1298 ;
  assign n7802 = ( n2560 & ~n6170 ) | ( n2560 & n7801 ) | ( ~n6170 & n7801 ) ;
  assign n7803 = ( ~n3581 & n4060 ) | ( ~n3581 & n7802 ) | ( n4060 & n7802 ) ;
  assign n7804 = n7803 ^ n7299 ^ n7044 ;
  assign n7805 = ( n6630 & n6794 ) | ( n6630 & ~n7804 ) | ( n6794 & ~n7804 ) ;
  assign n7806 = ( n1545 & ~n1677 ) | ( n1545 & n7805 ) | ( ~n1677 & n7805 ) ;
  assign n7823 = ( n1076 & n2110 ) | ( n1076 & ~n3230 ) | ( n2110 & ~n3230 ) ;
  assign n7824 = ( n990 & ~n2791 ) | ( n990 & n3576 ) | ( ~n2791 & n3576 ) ;
  assign n7825 = ( n4974 & ~n5710 ) | ( n4974 & n7824 ) | ( ~n5710 & n7824 ) ;
  assign n7826 = ( n4499 & ~n7823 ) | ( n4499 & n7825 ) | ( ~n7823 & n7825 ) ;
  assign n7827 = ( n2015 & ~n2886 ) | ( n2015 & n7826 ) | ( ~n2886 & n7826 ) ;
  assign n7807 = n3256 ^ n1952 ^ n794 ;
  assign n7808 = ( n343 & ~n2101 ) | ( n343 & n7807 ) | ( ~n2101 & n7807 ) ;
  assign n7809 = n7808 ^ n2468 ^ n775 ;
  assign n7810 = ( n516 & n3938 ) | ( n516 & n4463 ) | ( n3938 & n4463 ) ;
  assign n7811 = n7810 ^ n4340 ^ n3711 ;
  assign n7812 = n5232 ^ n2508 ^ n2462 ;
  assign n7813 = n7812 ^ n6317 ^ n1072 ;
  assign n7814 = n5680 ^ n923 ^ n198 ;
  assign n7815 = n7814 ^ n5720 ^ n1434 ;
  assign n7816 = ( n4545 & n6292 ) | ( n4545 & ~n7815 ) | ( n6292 & ~n7815 ) ;
  assign n7817 = ( ~n696 & n3634 ) | ( ~n696 & n7114 ) | ( n3634 & n7114 ) ;
  assign n7818 = ( x125 & ~n1299 ) | ( x125 & n5592 ) | ( ~n1299 & n5592 ) ;
  assign n7819 = ( x51 & n7817 ) | ( x51 & ~n7818 ) | ( n7817 & ~n7818 ) ;
  assign n7820 = n7819 ^ n6429 ^ n992 ;
  assign n7821 = ( n7813 & n7816 ) | ( n7813 & ~n7820 ) | ( n7816 & ~n7820 ) ;
  assign n7822 = ( n7809 & n7811 ) | ( n7809 & n7821 ) | ( n7811 & n7821 ) ;
  assign n7828 = n7827 ^ n7822 ^ n4414 ;
  assign n7836 = n6554 ^ n1243 ^ n129 ;
  assign n7830 = n4576 ^ n2754 ^ n2371 ;
  assign n7831 = n4300 ^ n3834 ^ n931 ;
  assign n7832 = ( ~n4594 & n6576 ) | ( ~n4594 & n7831 ) | ( n6576 & n7831 ) ;
  assign n7833 = ( n1869 & ~n7830 ) | ( n1869 & n7832 ) | ( ~n7830 & n7832 ) ;
  assign n7829 = n2256 ^ n2142 ^ n853 ;
  assign n7834 = n7833 ^ n7829 ^ n3833 ;
  assign n7835 = ( ~n3034 & n4209 ) | ( ~n3034 & n7834 ) | ( n4209 & n7834 ) ;
  assign n7837 = n7836 ^ n7835 ^ n1221 ;
  assign n7842 = ( n1358 & ~n3281 ) | ( n1358 & n6513 ) | ( ~n3281 & n6513 ) ;
  assign n7840 = n4025 ^ n2621 ^ n592 ;
  assign n7841 = ( n472 & n2389 ) | ( n472 & n7840 ) | ( n2389 & n7840 ) ;
  assign n7843 = n7842 ^ n7841 ^ x127 ;
  assign n7838 = n6804 ^ n6515 ^ n401 ;
  assign n7839 = n7838 ^ n6038 ^ n1402 ;
  assign n7844 = n7843 ^ n7839 ^ n7443 ;
  assign n7859 = ( n490 & n3285 ) | ( n490 & ~n3760 ) | ( n3285 & ~n3760 ) ;
  assign n7857 = n2103 ^ n1184 ^ n969 ;
  assign n7854 = ( n1639 & n1978 ) | ( n1639 & ~n2000 ) | ( n1978 & ~n2000 ) ;
  assign n7852 = ( ~n1262 & n2932 ) | ( ~n1262 & n3711 ) | ( n2932 & n3711 ) ;
  assign n7853 = ( n2592 & ~n5477 ) | ( n2592 & n7852 ) | ( ~n5477 & n7852 ) ;
  assign n7855 = n7854 ^ n7853 ^ n6064 ;
  assign n7856 = n7855 ^ n7384 ^ n1420 ;
  assign n7849 = n3388 ^ n586 ^ n373 ;
  assign n7850 = n2736 ^ n1392 ^ n532 ;
  assign n7851 = ( n1214 & n7849 ) | ( n1214 & n7850 ) | ( n7849 & n7850 ) ;
  assign n7858 = n7857 ^ n7856 ^ n7851 ;
  assign n7846 = ( ~n1675 & n2552 ) | ( ~n1675 & n2693 ) | ( n2552 & n2693 ) ;
  assign n7845 = n6076 ^ n5508 ^ n3991 ;
  assign n7847 = n7846 ^ n7845 ^ n1421 ;
  assign n7848 = n7847 ^ n3215 ^ n381 ;
  assign n7860 = n7859 ^ n7858 ^ n7848 ;
  assign n7865 = ( n736 & n3448 ) | ( n736 & n3655 ) | ( n3448 & n3655 ) ;
  assign n7866 = n7865 ^ n4527 ^ n3881 ;
  assign n7867 = ( n3940 & n6932 ) | ( n3940 & n7296 ) | ( n6932 & n7296 ) ;
  assign n7868 = ( n2419 & n7866 ) | ( n2419 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7861 = n4702 ^ n4299 ^ n2487 ;
  assign n7862 = n4822 ^ n3489 ^ n1707 ;
  assign n7863 = n7862 ^ n7436 ^ n6623 ;
  assign n7864 = ( n2469 & n7861 ) | ( n2469 & n7863 ) | ( n7861 & n7863 ) ;
  assign n7869 = n7868 ^ n7864 ^ n460 ;
  assign n7870 = ( ~n1943 & n4781 ) | ( ~n1943 & n7383 ) | ( n4781 & n7383 ) ;
  assign n7871 = ( n164 & ~n7458 ) | ( n164 & n7870 ) | ( ~n7458 & n7870 ) ;
  assign n7872 = ( n5727 & n7869 ) | ( n5727 & ~n7871 ) | ( n7869 & ~n7871 ) ;
  assign n7874 = n7199 ^ n3653 ^ n1694 ;
  assign n7873 = n5549 ^ n2848 ^ n2360 ;
  assign n7875 = n7874 ^ n7873 ^ n7196 ;
  assign n7876 = n7875 ^ n5638 ^ n744 ;
  assign n7877 = n1237 ^ n698 ^ n248 ;
  assign n7878 = n6171 ^ n4402 ^ n1371 ;
  assign n7879 = n7346 ^ n6213 ^ n3618 ;
  assign n7880 = n7879 ^ n3818 ^ n1017 ;
  assign n7881 = ( n7877 & n7878 ) | ( n7877 & n7880 ) | ( n7878 & n7880 ) ;
  assign n7882 = ( n1455 & n4821 ) | ( n1455 & ~n7881 ) | ( n4821 & ~n7881 ) ;
  assign n7883 = ( n4068 & n4077 ) | ( n4068 & ~n7882 ) | ( n4077 & ~n7882 ) ;
  assign n7887 = n7027 ^ n3489 ^ x13 ;
  assign n7884 = n2292 ^ n517 ^ n249 ;
  assign n7885 = ( n1402 & n3071 ) | ( n1402 & ~n7884 ) | ( n3071 & ~n7884 ) ;
  assign n7886 = ( ~n1766 & n4104 ) | ( ~n1766 & n7885 ) | ( n4104 & n7885 ) ;
  assign n7888 = n7887 ^ n7886 ^ n2592 ;
  assign n7889 = ( ~n876 & n3397 ) | ( ~n876 & n5054 ) | ( n3397 & n5054 ) ;
  assign n7890 = ( n2092 & n5080 ) | ( n2092 & n6849 ) | ( n5080 & n6849 ) ;
  assign n7891 = ( n2521 & n3516 ) | ( n2521 & n7890 ) | ( n3516 & n7890 ) ;
  assign n7892 = ( n487 & n7150 ) | ( n487 & ~n7891 ) | ( n7150 & ~n7891 ) ;
  assign n7893 = ( n6393 & ~n7889 ) | ( n6393 & n7892 ) | ( ~n7889 & n7892 ) ;
  assign n7894 = ( n488 & n3667 ) | ( n488 & ~n7893 ) | ( n3667 & ~n7893 ) ;
  assign n7895 = ( ~n2305 & n3052 ) | ( ~n2305 & n4798 ) | ( n3052 & n4798 ) ;
  assign n7896 = ( n900 & ~n2178 ) | ( n900 & n4583 ) | ( ~n2178 & n4583 ) ;
  assign n7897 = ( n1420 & n2138 ) | ( n1420 & ~n7896 ) | ( n2138 & ~n7896 ) ;
  assign n7898 = ( n871 & ~n6633 ) | ( n871 & n7897 ) | ( ~n6633 & n7897 ) ;
  assign n7901 = n5008 ^ n3660 ^ n1883 ;
  assign n7902 = ( n945 & n7759 ) | ( n945 & ~n7901 ) | ( n7759 & ~n7901 ) ;
  assign n7900 = n4559 ^ n4191 ^ n1064 ;
  assign n7899 = ( n1989 & n3297 ) | ( n1989 & ~n3367 ) | ( n3297 & ~n3367 ) ;
  assign n7903 = n7902 ^ n7900 ^ n7899 ;
  assign n7904 = ( n571 & n2735 ) | ( n571 & n3352 ) | ( n2735 & n3352 ) ;
  assign n7905 = ( n6196 & n7903 ) | ( n6196 & ~n7904 ) | ( n7903 & ~n7904 ) ;
  assign n7906 = ( n7895 & n7898 ) | ( n7895 & n7905 ) | ( n7898 & n7905 ) ;
  assign n7910 = n4429 ^ n1266 ^ n674 ;
  assign n7911 = n7910 ^ n2656 ^ n1877 ;
  assign n7908 = ( n1389 & n1539 ) | ( n1389 & ~n2231 ) | ( n1539 & ~n2231 ) ;
  assign n7909 = n7908 ^ n1374 ^ n1303 ;
  assign n7907 = n7510 ^ n635 ^ x4 ;
  assign n7912 = n7911 ^ n7909 ^ n7907 ;
  assign n7913 = ( n1144 & ~n4758 ) | ( n1144 & n4960 ) | ( ~n4758 & n4960 ) ;
  assign n7914 = n7913 ^ n5723 ^ n520 ;
  assign n7915 = n7914 ^ n4176 ^ n2111 ;
  assign n7916 = ( n400 & n7912 ) | ( n400 & n7915 ) | ( n7912 & n7915 ) ;
  assign n7918 = ( n2597 & ~n2916 ) | ( n2597 & n3510 ) | ( ~n2916 & n3510 ) ;
  assign n7919 = n7918 ^ n2773 ^ n1586 ;
  assign n7917 = n6093 ^ n4543 ^ n2978 ;
  assign n7920 = n7919 ^ n7917 ^ n3722 ;
  assign n7921 = ( n3509 & ~n4345 ) | ( n3509 & n7920 ) | ( ~n4345 & n7920 ) ;
  assign n7944 = n4790 ^ n4134 ^ n2369 ;
  assign n7945 = n7944 ^ n2794 ^ n1473 ;
  assign n7939 = n2052 ^ n1338 ^ n1225 ;
  assign n7940 = n7939 ^ n7315 ^ n155 ;
  assign n7941 = ( ~n1422 & n3122 ) | ( ~n1422 & n6056 ) | ( n3122 & n6056 ) ;
  assign n7942 = ( n6814 & n7940 ) | ( n6814 & ~n7941 ) | ( n7940 & ~n7941 ) ;
  assign n7943 = n7942 ^ n5954 ^ n5407 ;
  assign n7946 = n7945 ^ n7943 ^ n2969 ;
  assign n7937 = ( n1764 & n2929 ) | ( n1764 & n6541 ) | ( n2929 & n6541 ) ;
  assign n7938 = ( n1323 & n3652 ) | ( n1323 & n7937 ) | ( n3652 & n7937 ) ;
  assign n7947 = n7946 ^ n7938 ^ n4023 ;
  assign n7925 = ( n389 & n969 ) | ( n389 & ~n4306 ) | ( n969 & ~n4306 ) ;
  assign n7923 = n7896 ^ n2693 ^ n196 ;
  assign n7924 = ( ~n1434 & n4737 ) | ( ~n1434 & n7923 ) | ( n4737 & n7923 ) ;
  assign n7922 = ( n427 & n1539 ) | ( n427 & ~n2620 ) | ( n1539 & ~n2620 ) ;
  assign n7926 = n7925 ^ n7924 ^ n7922 ;
  assign n7927 = ( ~n4229 & n4958 ) | ( ~n4229 & n5403 ) | ( n4958 & n5403 ) ;
  assign n7928 = ( n2183 & ~n5369 ) | ( n2183 & n7927 ) | ( ~n5369 & n7927 ) ;
  assign n7929 = ( n1317 & n7926 ) | ( n1317 & ~n7928 ) | ( n7926 & ~n7928 ) ;
  assign n7930 = n7929 ^ n7074 ^ n1455 ;
  assign n7931 = ( n4687 & ~n4878 ) | ( n4687 & n6357 ) | ( ~n4878 & n6357 ) ;
  assign n7932 = ( ~n849 & n3863 ) | ( ~n849 & n7931 ) | ( n3863 & n7931 ) ;
  assign n7933 = ( ~n1705 & n2194 ) | ( ~n1705 & n7688 ) | ( n2194 & n7688 ) ;
  assign n7934 = ( x94 & n2900 ) | ( x94 & ~n7933 ) | ( n2900 & ~n7933 ) ;
  assign n7935 = ( ~n5636 & n7932 ) | ( ~n5636 & n7934 ) | ( n7932 & n7934 ) ;
  assign n7936 = ( n1933 & ~n7930 ) | ( n1933 & n7935 ) | ( ~n7930 & n7935 ) ;
  assign n7948 = n7947 ^ n7936 ^ n3275 ;
  assign n7958 = ( ~n452 & n1665 ) | ( ~n452 & n2615 ) | ( n1665 & n2615 ) ;
  assign n7959 = n7958 ^ n4113 ^ n2892 ;
  assign n7961 = n7959 ^ n7120 ^ n5551 ;
  assign n7962 = ( ~n5587 & n5862 ) | ( ~n5587 & n7961 ) | ( n5862 & n7961 ) ;
  assign n7953 = ( n1934 & ~n2821 ) | ( n1934 & n5023 ) | ( ~n2821 & n5023 ) ;
  assign n7954 = n7953 ^ n5624 ^ n5273 ;
  assign n7955 = ( n841 & n1210 ) | ( n841 & ~n1788 ) | ( n1210 & ~n1788 ) ;
  assign n7956 = n7955 ^ n4967 ^ n1212 ;
  assign n7957 = ( n4962 & n7954 ) | ( n4962 & n7956 ) | ( n7954 & n7956 ) ;
  assign n7960 = n7959 ^ n7957 ^ n1186 ;
  assign n7951 = n4762 ^ n4644 ^ n2633 ;
  assign n7949 = n1938 ^ n1627 ^ n688 ;
  assign n7950 = ( n1761 & ~n7217 ) | ( n1761 & n7949 ) | ( ~n7217 & n7949 ) ;
  assign n7952 = n7951 ^ n7950 ^ n4683 ;
  assign n7963 = n7962 ^ n7960 ^ n7952 ;
  assign n7966 = ( n2407 & n6609 ) | ( n2407 & n7274 ) | ( n6609 & n7274 ) ;
  assign n7964 = ( ~x107 & n1484 ) | ( ~x107 & n2012 ) | ( n1484 & n2012 ) ;
  assign n7965 = n7964 ^ n3929 ^ n3151 ;
  assign n7967 = n7966 ^ n7965 ^ n4393 ;
  assign n7968 = n7528 ^ n1923 ^ n1843 ;
  assign n7969 = n7968 ^ n7954 ^ n6497 ;
  assign n7970 = n6313 ^ n3237 ^ n2067 ;
  assign n7971 = ( n2174 & ~n4904 ) | ( n2174 & n7970 ) | ( ~n4904 & n7970 ) ;
  assign n7972 = ( n7967 & n7969 ) | ( n7967 & ~n7971 ) | ( n7969 & ~n7971 ) ;
  assign n7973 = ( ~n812 & n7635 ) | ( ~n812 & n7972 ) | ( n7635 & n7972 ) ;
  assign n7976 = ( ~n974 & n6287 ) | ( ~n974 & n6293 ) | ( n6287 & n6293 ) ;
  assign n7974 = n2446 ^ n1805 ^ n1539 ;
  assign n7975 = ( n1073 & n7433 ) | ( n1073 & ~n7974 ) | ( n7433 & ~n7974 ) ;
  assign n7977 = n7976 ^ n7975 ^ n5905 ;
  assign n7978 = n2083 ^ n1626 ^ n1236 ;
  assign n7980 = n3818 ^ n3791 ^ n3225 ;
  assign n7979 = n7809 ^ n1737 ^ n604 ;
  assign n7981 = n7980 ^ n7979 ^ n7322 ;
  assign n7982 = ( n3062 & n3264 ) | ( n3062 & n7981 ) | ( n3264 & n7981 ) ;
  assign n7983 = ( ~n1753 & n7978 ) | ( ~n1753 & n7982 ) | ( n7978 & n7982 ) ;
  assign n7984 = ( n204 & n1386 ) | ( n204 & ~n7983 ) | ( n1386 & ~n7983 ) ;
  assign n7986 = ( n561 & n820 ) | ( n561 & ~n1221 ) | ( n820 & ~n1221 ) ;
  assign n7987 = n2724 ^ n437 ^ n390 ;
  assign n7988 = ( n3613 & n5340 ) | ( n3613 & n7987 ) | ( n5340 & n7987 ) ;
  assign n7989 = ( ~n335 & n7986 ) | ( ~n335 & n7988 ) | ( n7986 & n7988 ) ;
  assign n7985 = ( n303 & n2523 ) | ( n303 & n6995 ) | ( n2523 & n6995 ) ;
  assign n7990 = n7989 ^ n7985 ^ n6803 ;
  assign n7991 = n5690 ^ n3739 ^ n2050 ;
  assign n7996 = ( x114 & n960 ) | ( x114 & ~n2099 ) | ( n960 & ~n2099 ) ;
  assign n7997 = ( n339 & n1257 ) | ( n339 & n7996 ) | ( n1257 & n7996 ) ;
  assign n7998 = ( n2321 & n4061 ) | ( n2321 & n7997 ) | ( n4061 & n7997 ) ;
  assign n7999 = n7998 ^ n5180 ^ n2197 ;
  assign n8000 = ( n2417 & n3494 ) | ( n2417 & ~n7999 ) | ( n3494 & ~n7999 ) ;
  assign n7992 = n4386 ^ n4237 ^ n2628 ;
  assign n7993 = n7992 ^ n6699 ^ n963 ;
  assign n7994 = ( n6312 & n6648 ) | ( n6312 & ~n7993 ) | ( n6648 & ~n7993 ) ;
  assign n7995 = n7994 ^ n6258 ^ n6048 ;
  assign n8001 = n8000 ^ n7995 ^ n3624 ;
  assign n8002 = ( n7990 & n7991 ) | ( n7990 & n8001 ) | ( n7991 & n8001 ) ;
  assign n8003 = ( n954 & n2012 ) | ( n954 & ~n6828 ) | ( n2012 & ~n6828 ) ;
  assign n8004 = ( n1733 & ~n2511 ) | ( n1733 & n8003 ) | ( ~n2511 & n8003 ) ;
  assign n8010 = n5072 ^ n3890 ^ n3254 ;
  assign n8011 = ( n1884 & n2501 ) | ( n1884 & n8010 ) | ( n2501 & n8010 ) ;
  assign n8005 = ( n294 & ~n1161 ) | ( n294 & n1454 ) | ( ~n1161 & n1454 ) ;
  assign n8006 = n8005 ^ n5038 ^ n815 ;
  assign n8007 = n3591 ^ n2555 ^ n557 ;
  assign n8008 = ( ~n2188 & n6820 ) | ( ~n2188 & n8007 ) | ( n6820 & n8007 ) ;
  assign n8009 = ( n6691 & n8006 ) | ( n6691 & ~n8008 ) | ( n8006 & ~n8008 ) ;
  assign n8012 = n8011 ^ n8009 ^ n6225 ;
  assign n8013 = n6545 ^ n2021 ^ x54 ;
  assign n8014 = ( n1474 & n6120 ) | ( n1474 & ~n8013 ) | ( n6120 & ~n8013 ) ;
  assign n8015 = ( n8004 & n8012 ) | ( n8004 & n8014 ) | ( n8012 & n8014 ) ;
  assign n8016 = ( ~n332 & n1598 ) | ( ~n332 & n5037 ) | ( n1598 & n5037 ) ;
  assign n8017 = n2448 ^ n1513 ^ n1206 ;
  assign n8018 = ( n936 & n4104 ) | ( n936 & n7132 ) | ( n4104 & n7132 ) ;
  assign n8019 = ( ~n2586 & n8017 ) | ( ~n2586 & n8018 ) | ( n8017 & n8018 ) ;
  assign n8020 = ( n934 & n6935 ) | ( n934 & n8019 ) | ( n6935 & n8019 ) ;
  assign n8021 = ( ~n7134 & n8016 ) | ( ~n7134 & n8020 ) | ( n8016 & n8020 ) ;
  assign n8022 = n3351 ^ n2595 ^ n558 ;
  assign n8023 = n8022 ^ n6678 ^ n1371 ;
  assign n8024 = ( n2102 & n2224 ) | ( n2102 & ~n2465 ) | ( n2224 & ~n2465 ) ;
  assign n8025 = n1724 ^ n1585 ^ x118 ;
  assign n8026 = ( n2201 & n3688 ) | ( n2201 & ~n5781 ) | ( n3688 & ~n5781 ) ;
  assign n8027 = ( n510 & ~n2885 ) | ( n510 & n3833 ) | ( ~n2885 & n3833 ) ;
  assign n8029 = ( x86 & n1875 ) | ( x86 & ~n6940 ) | ( n1875 & ~n6940 ) ;
  assign n8030 = ( ~n1401 & n4689 ) | ( ~n1401 & n8029 ) | ( n4689 & n8029 ) ;
  assign n8031 = ( ~n2214 & n4477 ) | ( ~n2214 & n8030 ) | ( n4477 & n8030 ) ;
  assign n8028 = n6224 ^ n5208 ^ n3256 ;
  assign n8032 = n8031 ^ n8028 ^ n268 ;
  assign n8033 = ( ~n8026 & n8027 ) | ( ~n8026 & n8032 ) | ( n8027 & n8032 ) ;
  assign n8034 = ( n6825 & n8025 ) | ( n6825 & n8033 ) | ( n8025 & n8033 ) ;
  assign n8035 = n3954 ^ n3160 ^ n569 ;
  assign n8049 = ( n599 & n5244 ) | ( n599 & n6280 ) | ( n5244 & n6280 ) ;
  assign n8054 = ( n672 & n1443 ) | ( n672 & n4180 ) | ( n1443 & n4180 ) ;
  assign n8052 = ( ~n459 & n2317 ) | ( ~n459 & n5079 ) | ( n2317 & n5079 ) ;
  assign n8051 = n7173 ^ n5065 ^ n1450 ;
  assign n8053 = n8052 ^ n8051 ^ n5585 ;
  assign n8050 = ( n1542 & ~n1842 ) | ( n1542 & n4205 ) | ( ~n1842 & n4205 ) ;
  assign n8055 = n8054 ^ n8053 ^ n8050 ;
  assign n8056 = ( ~n1804 & n8049 ) | ( ~n1804 & n8055 ) | ( n8049 & n8055 ) ;
  assign n8047 = n5109 ^ n1633 ^ x47 ;
  assign n8040 = n1386 ^ n766 ^ n691 ;
  assign n8041 = n8040 ^ n2540 ^ n1400 ;
  assign n8042 = n8041 ^ n1210 ^ n1124 ;
  assign n8043 = ( n974 & n3746 ) | ( n974 & n4611 ) | ( n3746 & n4611 ) ;
  assign n8044 = n6491 ^ n6452 ^ n3940 ;
  assign n8045 = ( ~n1565 & n8043 ) | ( ~n1565 & n8044 ) | ( n8043 & n8044 ) ;
  assign n8046 = ( n5797 & n8042 ) | ( n5797 & n8045 ) | ( n8042 & n8045 ) ;
  assign n8036 = n4573 ^ n4045 ^ n3327 ;
  assign n8037 = n8036 ^ n3940 ^ n3513 ;
  assign n8038 = n8037 ^ n4492 ^ n238 ;
  assign n8039 = n8038 ^ n2524 ^ n1421 ;
  assign n8048 = n8047 ^ n8046 ^ n8039 ;
  assign n8057 = n8056 ^ n8048 ^ n6373 ;
  assign n8058 = n6615 ^ n4926 ^ n2803 ;
  assign n8059 = ( n517 & ~n3189 ) | ( n517 & n7964 ) | ( ~n3189 & n7964 ) ;
  assign n8060 = n8059 ^ n2269 ^ n946 ;
  assign n8061 = ( n838 & n8058 ) | ( n838 & ~n8060 ) | ( n8058 & ~n8060 ) ;
  assign n8063 = n3754 ^ n3456 ^ n1514 ;
  assign n8064 = ( n637 & n3101 ) | ( n637 & ~n8063 ) | ( n3101 & ~n8063 ) ;
  assign n8062 = n6412 ^ n4411 ^ n3535 ;
  assign n8065 = n8064 ^ n8062 ^ n354 ;
  assign n8069 = ( n1946 & n4596 ) | ( n1946 & n7759 ) | ( n4596 & n7759 ) ;
  assign n8066 = n2281 ^ n330 ^ x40 ;
  assign n8067 = n8066 ^ n7433 ^ n2498 ;
  assign n8068 = ( n6338 & n7001 ) | ( n6338 & n8067 ) | ( n7001 & n8067 ) ;
  assign n8070 = n8069 ^ n8068 ^ n6411 ;
  assign n8071 = ( n8061 & n8065 ) | ( n8061 & n8070 ) | ( n8065 & n8070 ) ;
  assign n8072 = n2268 ^ n757 ^ x65 ;
  assign n8073 = n8072 ^ n7763 ^ n5712 ;
  assign n8074 = n8073 ^ n7632 ^ n2104 ;
  assign n8075 = n8074 ^ n6263 ^ n1000 ;
  assign n8076 = ( n144 & ~n398 ) | ( n144 & n8075 ) | ( ~n398 & n8075 ) ;
  assign n8077 = n4536 ^ n2421 ^ n1307 ;
  assign n8078 = n8077 ^ n5890 ^ n1292 ;
  assign n8079 = ( n601 & n1052 ) | ( n601 & ~n1991 ) | ( n1052 & ~n1991 ) ;
  assign n8080 = ( n1202 & ~n3985 ) | ( n1202 & n4639 ) | ( ~n3985 & n4639 ) ;
  assign n8081 = ( n7032 & n8079 ) | ( n7032 & ~n8080 ) | ( n8079 & ~n8080 ) ;
  assign n8084 = ( n1454 & ~n3122 ) | ( n1454 & n3504 ) | ( ~n3122 & n3504 ) ;
  assign n8082 = ( ~n3323 & n3703 ) | ( ~n3323 & n4102 ) | ( n3703 & n4102 ) ;
  assign n8083 = ( ~n1396 & n2988 ) | ( ~n1396 & n8082 ) | ( n2988 & n8082 ) ;
  assign n8085 = n8084 ^ n8083 ^ n1345 ;
  assign n8086 = ( n384 & n652 ) | ( n384 & n2943 ) | ( n652 & n2943 ) ;
  assign n8095 = ( n717 & ~n2193 ) | ( n717 & n6208 ) | ( ~n2193 & n6208 ) ;
  assign n8093 = n5339 ^ n3738 ^ n1706 ;
  assign n8090 = ( n2236 & n4192 ) | ( n2236 & n7831 ) | ( n4192 & n7831 ) ;
  assign n8091 = n8090 ^ n1342 ^ n1065 ;
  assign n8092 = n8091 ^ n7016 ^ n2646 ;
  assign n8094 = n8093 ^ n8092 ^ n5336 ;
  assign n8087 = ( ~n3597 & n4576 ) | ( ~n3597 & n6404 ) | ( n4576 & n6404 ) ;
  assign n8088 = n8087 ^ n5993 ^ n3016 ;
  assign n8089 = ( n1870 & n5071 ) | ( n1870 & n8088 ) | ( n5071 & n8088 ) ;
  assign n8096 = n8095 ^ n8094 ^ n8089 ;
  assign n8097 = ( n2081 & n6058 ) | ( n2081 & ~n7410 ) | ( n6058 & ~n7410 ) ;
  assign n8098 = ( n1458 & ~n2792 ) | ( n1458 & n5110 ) | ( ~n2792 & n5110 ) ;
  assign n8099 = n8098 ^ n4588 ^ n2230 ;
  assign n8100 = ( n920 & ~n2465 ) | ( n920 & n7344 ) | ( ~n2465 & n7344 ) ;
  assign n8101 = ( n828 & ~n873 ) | ( n828 & n8100 ) | ( ~n873 & n8100 ) ;
  assign n8102 = ( n1893 & n8099 ) | ( n1893 & n8101 ) | ( n8099 & n8101 ) ;
  assign n8103 = n7239 ^ n4386 ^ n4134 ;
  assign n8104 = ( ~n8097 & n8102 ) | ( ~n8097 & n8103 ) | ( n8102 & n8103 ) ;
  assign n8107 = n6327 ^ n3878 ^ n2581 ;
  assign n8108 = n8107 ^ n3307 ^ n1950 ;
  assign n8109 = n8108 ^ n1100 ^ n320 ;
  assign n8105 = n8077 ^ n7577 ^ n3655 ;
  assign n8106 = n8105 ^ n3633 ^ n637 ;
  assign n8110 = n8109 ^ n8106 ^ n1020 ;
  assign n8111 = n8110 ^ n3836 ^ n980 ;
  assign n8118 = n8054 ^ n4179 ^ n2462 ;
  assign n8112 = n3950 ^ n2454 ^ n1722 ;
  assign n8115 = ( ~n3004 & n3163 ) | ( ~n3004 & n6863 ) | ( n3163 & n6863 ) ;
  assign n8113 = ( ~n980 & n2556 ) | ( ~n980 & n5435 ) | ( n2556 & n5435 ) ;
  assign n8114 = ( n438 & n6065 ) | ( n438 & n8113 ) | ( n6065 & n8113 ) ;
  assign n8116 = n8115 ^ n8114 ^ n764 ;
  assign n8117 = ( n5042 & n8112 ) | ( n5042 & n8116 ) | ( n8112 & n8116 ) ;
  assign n8119 = n8118 ^ n8117 ^ n1714 ;
  assign n8120 = n8119 ^ n3837 ^ n3651 ;
  assign n8122 = n4500 ^ n1146 ^ n653 ;
  assign n8123 = n8122 ^ n2997 ^ n797 ;
  assign n8121 = n2424 ^ n2130 ^ n1652 ;
  assign n8124 = n8123 ^ n8121 ^ n7362 ;
  assign n8133 = n4585 ^ n1314 ^ n544 ;
  assign n8125 = ( n500 & n1534 ) | ( n500 & n2051 ) | ( n1534 & n2051 ) ;
  assign n8126 = ( ~n1419 & n3818 ) | ( ~n1419 & n8125 ) | ( n3818 & n8125 ) ;
  assign n8127 = ( n2170 & n3735 ) | ( n2170 & ~n8126 ) | ( n3735 & ~n8126 ) ;
  assign n8129 = ( ~n630 & n1059 ) | ( ~n630 & n7432 ) | ( n1059 & n7432 ) ;
  assign n8128 = ( n1051 & n1762 ) | ( n1051 & n6816 ) | ( n1762 & n6816 ) ;
  assign n8130 = n8129 ^ n8128 ^ n8088 ;
  assign n8131 = n8130 ^ n2698 ^ n1840 ;
  assign n8132 = ( n3887 & n8127 ) | ( n3887 & n8131 ) | ( n8127 & n8131 ) ;
  assign n8134 = n8133 ^ n8132 ^ n7951 ;
  assign n8136 = n7824 ^ n2441 ^ n1723 ;
  assign n8135 = ( ~n3165 & n6617 ) | ( ~n3165 & n6867 ) | ( n6617 & n6867 ) ;
  assign n8137 = n8136 ^ n8135 ^ n5380 ;
  assign n8138 = ( x125 & n5981 ) | ( x125 & n6014 ) | ( n5981 & n6014 ) ;
  assign n8139 = ( x120 & n2089 ) | ( x120 & ~n8138 ) | ( n2089 & ~n8138 ) ;
  assign n8147 = ( ~n1300 & n1446 ) | ( ~n1300 & n2906 ) | ( n1446 & n2906 ) ;
  assign n8148 = n8147 ^ n6863 ^ n1791 ;
  assign n8145 = n6079 ^ n3539 ^ n966 ;
  assign n8146 = n8145 ^ n4275 ^ n1006 ;
  assign n8140 = ( n2369 & n2621 ) | ( n2369 & ~n2942 ) | ( n2621 & ~n2942 ) ;
  assign n8141 = n8140 ^ n2420 ^ n1381 ;
  assign n8142 = ( ~n2647 & n2894 ) | ( ~n2647 & n8141 ) | ( n2894 & n8141 ) ;
  assign n8143 = n8142 ^ n6278 ^ n912 ;
  assign n8144 = ( ~n1943 & n2982 ) | ( ~n1943 & n8143 ) | ( n2982 & n8143 ) ;
  assign n8149 = n8148 ^ n8146 ^ n8144 ;
  assign n8150 = ( n7840 & ~n8139 ) | ( n7840 & n8149 ) | ( ~n8139 & n8149 ) ;
  assign n8151 = ( ~n5870 & n8137 ) | ( ~n5870 & n8150 ) | ( n8137 & n8150 ) ;
  assign n8152 = ( n915 & n2295 ) | ( n915 & ~n3010 ) | ( n2295 & ~n3010 ) ;
  assign n8153 = n8152 ^ n5411 ^ n522 ;
  assign n8156 = n2502 ^ n995 ^ n462 ;
  assign n8154 = n7057 ^ n5489 ^ n253 ;
  assign n8155 = ( n983 & n7861 ) | ( n983 & ~n8154 ) | ( n7861 & ~n8154 ) ;
  assign n8157 = n8156 ^ n8155 ^ n3135 ;
  assign n8158 = ( n4594 & n8153 ) | ( n4594 & ~n8157 ) | ( n8153 & ~n8157 ) ;
  assign n8173 = n3857 ^ n3608 ^ n1135 ;
  assign n8169 = n2398 ^ n1898 ^ n550 ;
  assign n8170 = ( n1141 & n3637 ) | ( n1141 & ~n8169 ) | ( n3637 & ~n8169 ) ;
  assign n8167 = ( n452 & n2603 ) | ( n452 & n4217 ) | ( n2603 & n4217 ) ;
  assign n8166 = n4501 ^ n3946 ^ n3737 ;
  assign n8168 = n8167 ^ n8166 ^ n2829 ;
  assign n8171 = n8170 ^ n8168 ^ n1895 ;
  assign n8163 = n2607 ^ n2280 ^ n2206 ;
  assign n8164 = ( n2409 & n3659 ) | ( n2409 & n8163 ) | ( n3659 & n8163 ) ;
  assign n8159 = n7265 ^ n5009 ^ n2229 ;
  assign n8160 = n8159 ^ n5089 ^ n1247 ;
  assign n8161 = n8160 ^ n4226 ^ n342 ;
  assign n8162 = ( n546 & n949 ) | ( n546 & ~n8161 ) | ( n949 & ~n8161 ) ;
  assign n8165 = n8164 ^ n8162 ^ n3839 ;
  assign n8172 = n8171 ^ n8165 ^ n4405 ;
  assign n8174 = n8173 ^ n8172 ^ n3348 ;
  assign n8175 = ( ~n1165 & n3773 ) | ( ~n1165 & n5229 ) | ( n3773 & n5229 ) ;
  assign n8176 = ( n2720 & n3271 ) | ( n2720 & n8175 ) | ( n3271 & n8175 ) ;
  assign n8177 = n8176 ^ n5612 ^ n4835 ;
  assign n8178 = ( n3215 & ~n6080 ) | ( n3215 & n7296 ) | ( ~n6080 & n7296 ) ;
  assign n8179 = n8178 ^ n238 ^ x107 ;
  assign n8180 = ( n1761 & ~n2367 ) | ( n1761 & n8179 ) | ( ~n2367 & n8179 ) ;
  assign n8181 = ( n1813 & ~n8177 ) | ( n1813 & n8180 ) | ( ~n8177 & n8180 ) ;
  assign n8182 = n8181 ^ n4323 ^ n1785 ;
  assign n8183 = n8182 ^ n5067 ^ n4504 ;
  assign n8184 = ( n360 & n4683 ) | ( n360 & n8183 ) | ( n4683 & n8183 ) ;
  assign n8185 = n6620 ^ n2738 ^ n398 ;
  assign n8186 = n6825 ^ n5510 ^ n799 ;
  assign n8187 = ( n4053 & n8185 ) | ( n4053 & ~n8186 ) | ( n8185 & ~n8186 ) ;
  assign n8188 = n8187 ^ n6310 ^ n439 ;
  assign n8189 = ( n1209 & n5813 ) | ( n1209 & n7700 ) | ( n5813 & n7700 ) ;
  assign n8190 = ( n3547 & n4945 ) | ( n3547 & ~n8189 ) | ( n4945 & ~n8189 ) ;
  assign n8191 = ( n1261 & n2305 ) | ( n1261 & n5204 ) | ( n2305 & n5204 ) ;
  assign n8192 = n3265 ^ n2808 ^ n1991 ;
  assign n8193 = ( n7270 & ~n8191 ) | ( n7270 & n8192 ) | ( ~n8191 & n8192 ) ;
  assign n8194 = n5804 ^ n4493 ^ n3120 ;
  assign n8195 = ( n2032 & n3585 ) | ( n2032 & n5503 ) | ( n3585 & n5503 ) ;
  assign n8196 = ( n4099 & n7818 ) | ( n4099 & ~n8195 ) | ( n7818 & ~n8195 ) ;
  assign n8197 = ( ~n4511 & n8194 ) | ( ~n4511 & n8196 ) | ( n8194 & n8196 ) ;
  assign n8203 = n4779 ^ n3233 ^ n3198 ;
  assign n8204 = ( n4225 & n4432 ) | ( n4225 & ~n8203 ) | ( n4432 & ~n8203 ) ;
  assign n8200 = n4420 ^ n3606 ^ n850 ;
  assign n8201 = ( n3432 & n6922 ) | ( n3432 & ~n8200 ) | ( n6922 & ~n8200 ) ;
  assign n8198 = n6404 ^ n3241 ^ n902 ;
  assign n8199 = ( ~n319 & n1483 ) | ( ~n319 & n8198 ) | ( n1483 & n8198 ) ;
  assign n8202 = n8201 ^ n8199 ^ n5333 ;
  assign n8205 = n8204 ^ n8202 ^ n5222 ;
  assign n8206 = n7890 ^ n6280 ^ n4887 ;
  assign n8207 = ( n4448 & n4935 ) | ( n4448 & n6773 ) | ( n4935 & n6773 ) ;
  assign n8208 = ( n251 & n3918 ) | ( n251 & ~n5715 ) | ( n3918 & ~n5715 ) ;
  assign n8209 = n3686 ^ n3655 ^ n151 ;
  assign n8210 = ( n7010 & n8208 ) | ( n7010 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8211 = ( n5054 & n8207 ) | ( n5054 & ~n8210 ) | ( n8207 & ~n8210 ) ;
  assign n8212 = ( n6126 & n8206 ) | ( n6126 & ~n8211 ) | ( n8206 & ~n8211 ) ;
  assign n8213 = ( n3039 & ~n8205 ) | ( n3039 & n8212 ) | ( ~n8205 & n8212 ) ;
  assign n8214 = ( n508 & n4461 ) | ( n508 & ~n5724 ) | ( n4461 & ~n5724 ) ;
  assign n8216 = ( n3185 & ~n3490 ) | ( n3185 & n3822 ) | ( ~n3490 & n3822 ) ;
  assign n8215 = ( n1310 & n2819 ) | ( n1310 & n5712 ) | ( n2819 & n5712 ) ;
  assign n8217 = n8216 ^ n8215 ^ n2008 ;
  assign n8218 = ( ~n3867 & n5837 ) | ( ~n3867 & n8217 ) | ( n5837 & n8217 ) ;
  assign n8219 = ( n6819 & ~n8214 ) | ( n6819 & n8218 ) | ( ~n8214 & n8218 ) ;
  assign n8222 = n5879 ^ n1927 ^ n228 ;
  assign n8220 = ( ~x88 & n3688 ) | ( ~x88 & n4264 ) | ( n3688 & n4264 ) ;
  assign n8221 = n8220 ^ n1498 ^ n510 ;
  assign n8223 = n8222 ^ n8221 ^ n6706 ;
  assign n8224 = ( n1273 & n2503 ) | ( n1273 & ~n3182 ) | ( n2503 & ~n3182 ) ;
  assign n8225 = ( ~n2608 & n3529 ) | ( ~n2608 & n7264 ) | ( n3529 & n7264 ) ;
  assign n8226 = ( n162 & n2045 ) | ( n162 & ~n7255 ) | ( n2045 & ~n7255 ) ;
  assign n8227 = n6154 ^ n3690 ^ n3678 ;
  assign n8228 = ( n7832 & n8226 ) | ( n7832 & ~n8227 ) | ( n8226 & ~n8227 ) ;
  assign n8229 = ( ~n6470 & n8225 ) | ( ~n6470 & n8228 ) | ( n8225 & n8228 ) ;
  assign n8230 = n6630 ^ n2187 ^ n808 ;
  assign n8231 = ( ~n5594 & n6393 ) | ( ~n5594 & n8230 ) | ( n6393 & n8230 ) ;
  assign n8232 = ( n6930 & n8229 ) | ( n6930 & n8231 ) | ( n8229 & n8231 ) ;
  assign n8233 = ( n215 & n397 ) | ( n215 & ~n7297 ) | ( n397 & ~n7297 ) ;
  assign n8234 = ( n827 & n1114 ) | ( n827 & n6256 ) | ( n1114 & n6256 ) ;
  assign n8235 = ( n6541 & ~n8233 ) | ( n6541 & n8234 ) | ( ~n8233 & n8234 ) ;
  assign n8236 = n5994 ^ n5101 ^ n2139 ;
  assign n8237 = n6758 ^ n3704 ^ n1319 ;
  assign n8238 = ( ~n2362 & n3772 ) | ( ~n2362 & n8237 ) | ( n3772 & n8237 ) ;
  assign n8239 = ( n1291 & ~n7109 ) | ( n1291 & n8238 ) | ( ~n7109 & n8238 ) ;
  assign n8240 = n8239 ^ n2027 ^ n1520 ;
  assign n8241 = ( ~n1080 & n8236 ) | ( ~n1080 & n8240 ) | ( n8236 & n8240 ) ;
  assign n8253 = ( n2201 & ~n3922 ) | ( n2201 & n7842 ) | ( ~n3922 & n7842 ) ;
  assign n8245 = ( n3238 & ~n3280 ) | ( n3238 & n5582 ) | ( ~n3280 & n5582 ) ;
  assign n8246 = n8245 ^ n5260 ^ n549 ;
  assign n8248 = ( ~n797 & n4002 ) | ( ~n797 & n8108 ) | ( n4002 & n8108 ) ;
  assign n8249 = n8248 ^ n2475 ^ x106 ;
  assign n8247 = ( n2480 & ~n3000 ) | ( n2480 & n3526 ) | ( ~n3000 & n3526 ) ;
  assign n8250 = n8249 ^ n8247 ^ n1799 ;
  assign n8251 = ( n909 & n911 ) | ( n909 & n8250 ) | ( n911 & n8250 ) ;
  assign n8252 = ( ~n7368 & n8246 ) | ( ~n7368 & n8251 ) | ( n8246 & n8251 ) ;
  assign n8254 = n8253 ^ n8252 ^ n5322 ;
  assign n8242 = n3431 ^ n2632 ^ n832 ;
  assign n8243 = ( n4011 & n5369 ) | ( n4011 & ~n8242 ) | ( n5369 & ~n8242 ) ;
  assign n8244 = ( ~n2372 & n7272 ) | ( ~n2372 & n8243 ) | ( n7272 & n8243 ) ;
  assign n8255 = n8254 ^ n8244 ^ n3768 ;
  assign n8256 = ( n1903 & n2571 ) | ( n1903 & n8255 ) | ( n2571 & n8255 ) ;
  assign n8257 = n5579 ^ n2223 ^ n1286 ;
  assign n8258 = ( ~n1216 & n7991 ) | ( ~n1216 & n8257 ) | ( n7991 & n8257 ) ;
  assign n8259 = ( ~n3476 & n7464 ) | ( ~n3476 & n8258 ) | ( n7464 & n8258 ) ;
  assign n8260 = n8259 ^ n6336 ^ n1014 ;
  assign n8261 = ( ~n208 & n5271 ) | ( ~n208 & n8260 ) | ( n5271 & n8260 ) ;
  assign n8262 = ( x92 & n870 ) | ( x92 & n6798 ) | ( n870 & n6798 ) ;
  assign n8263 = n8262 ^ n4991 ^ n1025 ;
  assign n8264 = n8113 ^ n4652 ^ n3000 ;
  assign n8265 = ( n6574 & n8263 ) | ( n6574 & ~n8264 ) | ( n8263 & ~n8264 ) ;
  assign n8272 = ( n427 & ~n2120 ) | ( n427 & n2232 ) | ( ~n2120 & n2232 ) ;
  assign n8266 = ( ~n2435 & n2502 ) | ( ~n2435 & n4794 ) | ( n2502 & n4794 ) ;
  assign n8267 = n4004 ^ n1149 ^ n830 ;
  assign n8268 = ( n1809 & n7007 ) | ( n1809 & n8267 ) | ( n7007 & n8267 ) ;
  assign n8269 = ( n1731 & n2102 ) | ( n1731 & n8268 ) | ( n2102 & n8268 ) ;
  assign n8270 = n8269 ^ n4949 ^ n4124 ;
  assign n8271 = ( n6049 & ~n8266 ) | ( n6049 & n8270 ) | ( ~n8266 & n8270 ) ;
  assign n8273 = n8272 ^ n8271 ^ n4733 ;
  assign n8274 = n2977 ^ n2792 ^ n2285 ;
  assign n8275 = n8274 ^ n1270 ^ n507 ;
  assign n8276 = ( n5125 & ~n7136 ) | ( n5125 & n8275 ) | ( ~n7136 & n8275 ) ;
  assign n8277 = n7251 ^ n5830 ^ n4454 ;
  assign n8278 = ( n1047 & ~n3812 ) | ( n1047 & n8277 ) | ( ~n3812 & n8277 ) ;
  assign n8279 = ( n4649 & ~n8276 ) | ( n4649 & n8278 ) | ( ~n8276 & n8278 ) ;
  assign n8283 = ( n695 & n1164 ) | ( n695 & ~n1241 ) | ( n1164 & ~n1241 ) ;
  assign n8282 = ( ~n3451 & n4432 ) | ( ~n3451 & n4926 ) | ( n4432 & n4926 ) ;
  assign n8280 = n5193 ^ n2058 ^ n572 ;
  assign n8281 = ( n1055 & n6058 ) | ( n1055 & ~n8280 ) | ( n6058 & ~n8280 ) ;
  assign n8284 = n8283 ^ n8282 ^ n8281 ;
  assign n8290 = n2786 ^ n1223 ^ n1110 ;
  assign n8285 = n4674 ^ n2627 ^ n1622 ;
  assign n8286 = ( n1706 & n6321 ) | ( n1706 & n8285 ) | ( n6321 & n8285 ) ;
  assign n8287 = n8286 ^ n8245 ^ n6337 ;
  assign n8288 = n8287 ^ n4235 ^ n2739 ;
  assign n8289 = ( n2567 & n4568 ) | ( n2567 & n8288 ) | ( n4568 & n8288 ) ;
  assign n8291 = n8290 ^ n8289 ^ n4126 ;
  assign n8296 = n3363 ^ n2622 ^ n1369 ;
  assign n8294 = ( ~n719 & n2036 ) | ( ~n719 & n7097 ) | ( n2036 & n7097 ) ;
  assign n8295 = n8294 ^ n5644 ^ n1030 ;
  assign n8292 = ( n285 & n313 ) | ( n285 & ~n873 ) | ( n313 & ~n873 ) ;
  assign n8293 = n8292 ^ n3626 ^ n379 ;
  assign n8297 = n8296 ^ n8295 ^ n8293 ;
  assign n8304 = n4315 ^ n4080 ^ n1692 ;
  assign n8302 = n5356 ^ n729 ^ n278 ;
  assign n8298 = ( x97 & n3654 ) | ( x97 & n7264 ) | ( n3654 & n7264 ) ;
  assign n8299 = n2525 ^ n923 ^ x109 ;
  assign n8300 = n7118 ^ n5124 ^ n3162 ;
  assign n8301 = ( n8298 & n8299 ) | ( n8298 & ~n8300 ) | ( n8299 & ~n8300 ) ;
  assign n8303 = n8302 ^ n8301 ^ n4072 ;
  assign n8305 = n8304 ^ n8303 ^ n2452 ;
  assign n8306 = ( n2667 & ~n3478 ) | ( n2667 & n5039 ) | ( ~n3478 & n5039 ) ;
  assign n8307 = n8306 ^ n7900 ^ n2001 ;
  assign n8310 = n1426 ^ n1166 ^ n711 ;
  assign n8308 = n5059 ^ n2888 ^ n2502 ;
  assign n8309 = ( n4966 & n5483 ) | ( n4966 & n8308 ) | ( n5483 & n8308 ) ;
  assign n8311 = n8310 ^ n8309 ^ n5603 ;
  assign n8312 = ( n402 & ~n1440 ) | ( n402 & n5575 ) | ( ~n1440 & n5575 ) ;
  assign n8313 = n8312 ^ n6013 ^ n4420 ;
  assign n8314 = n4376 ^ n3953 ^ n1703 ;
  assign n8315 = n2628 ^ n853 ^ x72 ;
  assign n8316 = n4175 ^ n3980 ^ n3428 ;
  assign n8317 = ( n1137 & n8315 ) | ( n1137 & n8316 ) | ( n8315 & n8316 ) ;
  assign n8318 = ( n4952 & n5052 ) | ( n4952 & n8317 ) | ( n5052 & n8317 ) ;
  assign n8319 = ( ~n5553 & n8314 ) | ( ~n5553 & n8318 ) | ( n8314 & n8318 ) ;
  assign n8320 = ( n1161 & ~n3044 ) | ( n1161 & n4596 ) | ( ~n3044 & n4596 ) ;
  assign n8321 = ( n5325 & n7935 ) | ( n5325 & ~n8320 ) | ( n7935 & ~n8320 ) ;
  assign n8322 = ( x117 & n571 ) | ( x117 & n4096 ) | ( n571 & n4096 ) ;
  assign n8323 = ( n4829 & ~n7226 ) | ( n4829 & n8322 ) | ( ~n7226 & n8322 ) ;
  assign n8327 = n1151 ^ n1093 ^ n473 ;
  assign n8324 = ( n595 & n642 ) | ( n595 & n1770 ) | ( n642 & n1770 ) ;
  assign n8325 = ( n273 & n641 ) | ( n273 & ~n8324 ) | ( n641 & ~n8324 ) ;
  assign n8326 = n8325 ^ n7473 ^ n703 ;
  assign n8328 = n8327 ^ n8326 ^ n7899 ;
  assign n8329 = ( n694 & n3294 ) | ( n694 & ~n8328 ) | ( n3294 & ~n8328 ) ;
  assign n8341 = n3999 ^ n2327 ^ n1702 ;
  assign n8339 = ( ~n3270 & n4061 ) | ( ~n3270 & n7171 ) | ( n4061 & n7171 ) ;
  assign n8340 = ( n4578 & n6689 ) | ( n4578 & n8339 ) | ( n6689 & n8339 ) ;
  assign n8330 = ( ~n1432 & n6093 ) | ( ~n1432 & n8160 ) | ( n6093 & n8160 ) ;
  assign n8331 = n6638 ^ n1241 ^ n488 ;
  assign n8332 = n2819 ^ n1208 ^ n475 ;
  assign n8333 = ( n641 & n1241 ) | ( n641 & ~n8332 ) | ( n1241 & ~n8332 ) ;
  assign n8334 = ( ~n1828 & n7884 ) | ( ~n1828 & n8333 ) | ( n7884 & n8333 ) ;
  assign n8335 = ( n5180 & n6195 ) | ( n5180 & ~n8334 ) | ( n6195 & ~n8334 ) ;
  assign n8336 = ( n1437 & n5363 ) | ( n1437 & ~n8335 ) | ( n5363 & ~n8335 ) ;
  assign n8337 = ( n579 & n8331 ) | ( n579 & ~n8336 ) | ( n8331 & ~n8336 ) ;
  assign n8338 = ( n3143 & n8330 ) | ( n3143 & ~n8337 ) | ( n8330 & ~n8337 ) ;
  assign n8342 = n8341 ^ n8340 ^ n8338 ;
  assign n8343 = ( n5265 & n8329 ) | ( n5265 & ~n8342 ) | ( n8329 & ~n8342 ) ;
  assign n8345 = n6786 ^ n2780 ^ n1738 ;
  assign n8344 = n5410 ^ n3412 ^ n1959 ;
  assign n8346 = n8345 ^ n8344 ^ n770 ;
  assign n8356 = n6995 ^ n4598 ^ n4193 ;
  assign n8355 = n3131 ^ n2524 ^ n442 ;
  assign n8347 = n2958 ^ n1587 ^ n1235 ;
  assign n8352 = n6861 ^ n3077 ^ n1638 ;
  assign n8351 = n5586 ^ n3050 ^ n2927 ;
  assign n8348 = n6333 ^ n2999 ^ n1334 ;
  assign n8349 = ( n1629 & n3371 ) | ( n1629 & n8348 ) | ( n3371 & n8348 ) ;
  assign n8350 = ( ~n2400 & n3200 ) | ( ~n2400 & n8349 ) | ( n3200 & n8349 ) ;
  assign n8353 = n8352 ^ n8351 ^ n8350 ;
  assign n8354 = ( ~n4318 & n8347 ) | ( ~n4318 & n8353 ) | ( n8347 & n8353 ) ;
  assign n8357 = n8356 ^ n8355 ^ n8354 ;
  assign n8358 = ( n1811 & n2295 ) | ( n1811 & n3049 ) | ( n2295 & n3049 ) ;
  assign n8359 = ( ~n1857 & n3328 ) | ( ~n1857 & n8358 ) | ( n3328 & n8358 ) ;
  assign n8372 = n3837 ^ n3516 ^ n3078 ;
  assign n8369 = ( n2322 & ~n2587 ) | ( n2322 & n7052 ) | ( ~n2587 & n7052 ) ;
  assign n8370 = ( n4090 & ~n8115 ) | ( n4090 & n8369 ) | ( ~n8115 & n8369 ) ;
  assign n8360 = n7760 ^ n735 ^ n239 ;
  assign n8361 = ( x13 & n1905 ) | ( x13 & n4979 ) | ( n1905 & n4979 ) ;
  assign n8362 = ( n4910 & ~n8360 ) | ( n4910 & n8361 ) | ( ~n8360 & n8361 ) ;
  assign n8364 = n5832 ^ n5401 ^ n2628 ;
  assign n8365 = ( ~n1010 & n3326 ) | ( ~n1010 & n5870 ) | ( n3326 & n5870 ) ;
  assign n8366 = ( x55 & n8364 ) | ( x55 & ~n8365 ) | ( n8364 & ~n8365 ) ;
  assign n8363 = ( n289 & n4200 ) | ( n289 & n7500 ) | ( n4200 & n7500 ) ;
  assign n8367 = n8366 ^ n8363 ^ n2795 ;
  assign n8368 = ( n2908 & ~n8362 ) | ( n2908 & n8367 ) | ( ~n8362 & n8367 ) ;
  assign n8371 = n8370 ^ n8368 ^ n2889 ;
  assign n8373 = n8372 ^ n8371 ^ n7429 ;
  assign n8386 = ( n373 & n542 ) | ( n373 & n4146 ) | ( n542 & n4146 ) ;
  assign n8387 = n8386 ^ n7640 ^ n1190 ;
  assign n8383 = ( ~n151 & n3660 ) | ( ~n151 & n4734 ) | ( n3660 & n4734 ) ;
  assign n8384 = ( n3365 & ~n3731 ) | ( n3365 & n8383 ) | ( ~n3731 & n8383 ) ;
  assign n8378 = ( ~n193 & n671 ) | ( ~n193 & n876 ) | ( n671 & n876 ) ;
  assign n8379 = ( ~n592 & n2705 ) | ( ~n592 & n6074 ) | ( n2705 & n6074 ) ;
  assign n8380 = ( ~n260 & n639 ) | ( ~n260 & n8379 ) | ( n639 & n8379 ) ;
  assign n8381 = ( n6973 & n8378 ) | ( n6973 & ~n8380 ) | ( n8378 & ~n8380 ) ;
  assign n8382 = ( n772 & n4650 ) | ( n772 & ~n8381 ) | ( n4650 & ~n8381 ) ;
  assign n8385 = n8384 ^ n8382 ^ n5328 ;
  assign n8374 = ( n847 & n1788 ) | ( n847 & ~n2687 ) | ( n1788 & ~n2687 ) ;
  assign n8375 = n8374 ^ n8169 ^ n5895 ;
  assign n8376 = n8375 ^ n7222 ^ n2477 ;
  assign n8377 = n8376 ^ n7480 ^ n2214 ;
  assign n8388 = n8387 ^ n8385 ^ n8377 ;
  assign n8393 = ( n599 & n766 ) | ( n599 & n1544 ) | ( n766 & n1544 ) ;
  assign n8389 = n1972 ^ n1316 ^ n1272 ;
  assign n8390 = ( n793 & n1921 ) | ( n793 & ~n8389 ) | ( n1921 & ~n8389 ) ;
  assign n8391 = n8390 ^ n4556 ^ n449 ;
  assign n8392 = ( ~n645 & n8093 ) | ( ~n645 & n8391 ) | ( n8093 & n8391 ) ;
  assign n8394 = n8393 ^ n8392 ^ n5675 ;
  assign n8397 = ( n1198 & ~n1893 ) | ( n1198 & n2376 ) | ( ~n1893 & n2376 ) ;
  assign n8395 = n2236 ^ n835 ^ x42 ;
  assign n8396 = n8395 ^ n6209 ^ n2391 ;
  assign n8398 = n8397 ^ n8396 ^ n1783 ;
  assign n8399 = ( n187 & ~n7133 ) | ( n187 & n8398 ) | ( ~n7133 & n8398 ) ;
  assign n8400 = n8399 ^ n6293 ^ n5469 ;
  assign n8414 = ( ~n684 & n1545 ) | ( ~n684 & n7416 ) | ( n1545 & n7416 ) ;
  assign n8410 = n3785 ^ n3066 ^ x18 ;
  assign n8411 = n8410 ^ n4080 ^ n935 ;
  assign n8412 = n8411 ^ n6461 ^ n2538 ;
  assign n8413 = n8412 ^ n4790 ^ n4010 ;
  assign n8415 = n8414 ^ n8413 ^ n1089 ;
  assign n8406 = ( n1174 & n2095 ) | ( n1174 & ~n6726 ) | ( n2095 & ~n6726 ) ;
  assign n8407 = n5383 ^ n3083 ^ n475 ;
  assign n8408 = n8407 ^ n5775 ^ n3462 ;
  assign n8409 = ( n304 & n8406 ) | ( n304 & n8408 ) | ( n8406 & n8408 ) ;
  assign n8401 = ( n2196 & ~n2226 ) | ( n2196 & n6925 ) | ( ~n2226 & n6925 ) ;
  assign n8402 = ( n478 & n600 ) | ( n478 & ~n5216 ) | ( n600 & ~n5216 ) ;
  assign n8403 = ( n597 & ~n1429 ) | ( n597 & n8402 ) | ( ~n1429 & n8402 ) ;
  assign n8404 = ( n3820 & n5748 ) | ( n3820 & n8403 ) | ( n5748 & n8403 ) ;
  assign n8405 = ( n6651 & n8401 ) | ( n6651 & ~n8404 ) | ( n8401 & ~n8404 ) ;
  assign n8416 = n8415 ^ n8409 ^ n8405 ;
  assign n8422 = n3382 ^ n1559 ^ n1435 ;
  assign n8421 = n7136 ^ n2314 ^ n1588 ;
  assign n8419 = ( n1912 & n3026 ) | ( n1912 & n4485 ) | ( n3026 & n4485 ) ;
  assign n8418 = ( n3520 & ~n7865 ) | ( n3520 & n8226 ) | ( ~n7865 & n8226 ) ;
  assign n8417 = n6565 ^ n4835 ^ n1004 ;
  assign n8420 = n8419 ^ n8418 ^ n8417 ;
  assign n8423 = n8422 ^ n8421 ^ n8420 ;
  assign n8424 = ( n3428 & n7278 ) | ( n3428 & n8423 ) | ( n7278 & n8423 ) ;
  assign n8425 = n4326 ^ n2771 ^ n2366 ;
  assign n8426 = ( n686 & ~n6894 ) | ( n686 & n8425 ) | ( ~n6894 & n8425 ) ;
  assign n8429 = ( ~n485 & n1241 ) | ( ~n485 & n6816 ) | ( n1241 & n6816 ) ;
  assign n8427 = ( n6887 & ~n7700 ) | ( n6887 & n7831 ) | ( ~n7700 & n7831 ) ;
  assign n8428 = ( n1718 & n3043 ) | ( n1718 & n8427 ) | ( n3043 & n8427 ) ;
  assign n8430 = n8429 ^ n8428 ^ n845 ;
  assign n8438 = ( x50 & ~n323 ) | ( x50 & n7701 ) | ( ~n323 & n7701 ) ;
  assign n8435 = n5113 ^ n4778 ^ n3728 ;
  assign n8432 = ( n3732 & n3959 ) | ( n3732 & ~n5610 ) | ( n3959 & ~n5610 ) ;
  assign n8431 = ( x115 & ~n7874 ) | ( x115 & n8099 ) | ( ~n7874 & n8099 ) ;
  assign n8433 = n8432 ^ n8431 ^ n8093 ;
  assign n8434 = n8433 ^ n791 ^ n574 ;
  assign n8436 = n8435 ^ n8434 ^ n7088 ;
  assign n8437 = n8436 ^ n1811 ^ n921 ;
  assign n8439 = n8438 ^ n8437 ^ n6156 ;
  assign n8440 = ( ~n7628 & n8430 ) | ( ~n7628 & n8439 ) | ( n8430 & n8439 ) ;
  assign n8453 = n1262 ^ n1166 ^ n377 ;
  assign n8454 = n8453 ^ n3038 ^ n1473 ;
  assign n8445 = ( ~x118 & n2173 ) | ( ~x118 & n3484 ) | ( n2173 & n3484 ) ;
  assign n8446 = ( n2293 & ~n7377 ) | ( n2293 & n8445 ) | ( ~n7377 & n8445 ) ;
  assign n8448 = ( ~n546 & n5178 ) | ( ~n546 & n7759 ) | ( n5178 & n7759 ) ;
  assign n8449 = ( n359 & ~n1751 ) | ( n359 & n8448 ) | ( ~n1751 & n8448 ) ;
  assign n8447 = ( n2039 & n3909 ) | ( n2039 & ~n6291 ) | ( n3909 & ~n6291 ) ;
  assign n8450 = n8449 ^ n8447 ^ n519 ;
  assign n8451 = n8450 ^ n3243 ^ n2329 ;
  assign n8452 = ( n2354 & n8446 ) | ( n2354 & ~n8451 ) | ( n8446 & ~n8451 ) ;
  assign n8441 = n3179 ^ n3150 ^ x36 ;
  assign n8442 = n8441 ^ n8088 ^ n2752 ;
  assign n8443 = ( n775 & ~n5381 ) | ( n775 & n7438 ) | ( ~n5381 & n7438 ) ;
  assign n8444 = ( n5428 & n8442 ) | ( n5428 & ~n8443 ) | ( n8442 & ~n8443 ) ;
  assign n8455 = n8454 ^ n8452 ^ n8444 ;
  assign n8458 = ( ~n1608 & n1676 ) | ( ~n1608 & n6001 ) | ( n1676 & n6001 ) ;
  assign n8459 = ( n2389 & ~n7817 ) | ( n2389 & n8458 ) | ( ~n7817 & n8458 ) ;
  assign n8456 = ( ~n213 & n1865 ) | ( ~n213 & n6014 ) | ( n1865 & n6014 ) ;
  assign n8457 = n8456 ^ n1865 ^ n758 ;
  assign n8460 = n8459 ^ n8457 ^ n7091 ;
  assign n8461 = ( ~n707 & n5939 ) | ( ~n707 & n6537 ) | ( n5939 & n6537 ) ;
  assign n8462 = n8461 ^ n5684 ^ n2669 ;
  assign n8463 = n8225 ^ n2555 ^ n424 ;
  assign n8464 = n3215 ^ n2744 ^ n667 ;
  assign n8465 = n4081 ^ n3734 ^ n2018 ;
  assign n8466 = ( n6935 & n8464 ) | ( n6935 & ~n8465 ) | ( n8464 & ~n8465 ) ;
  assign n8467 = ( n6251 & ~n8463 ) | ( n6251 & n8466 ) | ( ~n8463 & n8466 ) ;
  assign n8468 = ( n7787 & n8462 ) | ( n7787 & ~n8467 ) | ( n8462 & ~n8467 ) ;
  assign n8469 = ( n5095 & ~n8460 ) | ( n5095 & n8468 ) | ( ~n8460 & n8468 ) ;
  assign n8470 = ( n3162 & ~n3745 ) | ( n3162 & n3816 ) | ( ~n3745 & n3816 ) ;
  assign n8471 = ( n1611 & ~n6977 ) | ( n1611 & n8470 ) | ( ~n6977 & n8470 ) ;
  assign n8472 = ( ~n175 & n1347 ) | ( ~n175 & n6590 ) | ( n1347 & n6590 ) ;
  assign n8473 = n4325 ^ n3869 ^ n2597 ;
  assign n8474 = ( n317 & n320 ) | ( n317 & n3252 ) | ( n320 & n3252 ) ;
  assign n8475 = ( n1620 & ~n2708 ) | ( n1620 & n4704 ) | ( ~n2708 & n4704 ) ;
  assign n8476 = ( n4604 & n8474 ) | ( n4604 & ~n8475 ) | ( n8474 & ~n8475 ) ;
  assign n8477 = ( n7121 & ~n8473 ) | ( n7121 & n8476 ) | ( ~n8473 & n8476 ) ;
  assign n8478 = ( n8471 & n8472 ) | ( n8471 & n8477 ) | ( n8472 & n8477 ) ;
  assign n8479 = ( ~n1272 & n1773 ) | ( ~n1272 & n2169 ) | ( n1773 & n2169 ) ;
  assign n8480 = ( ~n5483 & n7964 ) | ( ~n5483 & n8479 ) | ( n7964 & n8479 ) ;
  assign n8481 = ( n5237 & n5903 ) | ( n5237 & ~n8480 ) | ( n5903 & ~n8480 ) ;
  assign n8482 = ( n1612 & n1783 ) | ( n1612 & n8481 ) | ( n1783 & n8481 ) ;
  assign n8483 = ( n676 & n6019 ) | ( n676 & n7316 ) | ( n6019 & n7316 ) ;
  assign n8484 = ( n2849 & n5334 ) | ( n2849 & ~n8483 ) | ( n5334 & ~n8483 ) ;
  assign n8485 = ( n955 & n6148 ) | ( n955 & ~n8484 ) | ( n6148 & ~n8484 ) ;
  assign n8491 = ( ~n185 & n836 ) | ( ~n185 & n1028 ) | ( n836 & n1028 ) ;
  assign n8486 = n2336 ^ n1011 ^ n183 ;
  assign n8487 = ( n1278 & ~n1361 ) | ( n1278 & n8486 ) | ( ~n1361 & n8486 ) ;
  assign n8488 = n7559 ^ n2308 ^ n1071 ;
  assign n8489 = ( n1454 & n8487 ) | ( n1454 & n8488 ) | ( n8487 & n8488 ) ;
  assign n8490 = ( n913 & n1991 ) | ( n913 & ~n8489 ) | ( n1991 & ~n8489 ) ;
  assign n8492 = n8491 ^ n8490 ^ n7170 ;
  assign n8493 = n6825 ^ n5911 ^ n4045 ;
  assign n8494 = ( ~n6440 & n8167 ) | ( ~n6440 & n8493 ) | ( n8167 & n8493 ) ;
  assign n8495 = n8494 ^ n8415 ^ n2279 ;
  assign n8496 = ( n1342 & n2345 ) | ( n1342 & n4536 ) | ( n2345 & n4536 ) ;
  assign n8500 = n1044 ^ n1029 ^ n250 ;
  assign n8501 = ( n208 & n1875 ) | ( n208 & n8500 ) | ( n1875 & n8500 ) ;
  assign n8502 = n5330 ^ n4087 ^ n3810 ;
  assign n8503 = ( n151 & n8501 ) | ( n151 & ~n8502 ) | ( n8501 & ~n8502 ) ;
  assign n8497 = ( n1668 & n1827 ) | ( n1668 & n6424 ) | ( n1827 & n6424 ) ;
  assign n8498 = ( ~n2838 & n8333 ) | ( ~n2838 & n8497 ) | ( n8333 & n8497 ) ;
  assign n8499 = n8498 ^ n7137 ^ n4254 ;
  assign n8504 = n8503 ^ n8499 ^ n2107 ;
  assign n8505 = ( ~n2682 & n8496 ) | ( ~n2682 & n8504 ) | ( n8496 & n8504 ) ;
  assign n8514 = n7246 ^ n5482 ^ n674 ;
  assign n8515 = ( n661 & n1266 ) | ( n661 & ~n2627 ) | ( n1266 & ~n2627 ) ;
  assign n8516 = n8515 ^ n2536 ^ n527 ;
  assign n8517 = ( n3305 & n8514 ) | ( n3305 & n8516 ) | ( n8514 & n8516 ) ;
  assign n8518 = ( n1204 & n7296 ) | ( n1204 & ~n8517 ) | ( n7296 & ~n8517 ) ;
  assign n8511 = ( n1404 & n2536 ) | ( n1404 & n4958 ) | ( n2536 & n4958 ) ;
  assign n8512 = ( n2317 & n2377 ) | ( n2317 & ~n8511 ) | ( n2377 & ~n8511 ) ;
  assign n8513 = ( ~n2730 & n4812 ) | ( ~n2730 & n8512 ) | ( n4812 & n8512 ) ;
  assign n8506 = n7942 ^ n5095 ^ n4046 ;
  assign n8507 = n6046 ^ n3451 ^ x65 ;
  assign n8508 = ( n2190 & n3063 ) | ( n2190 & ~n8507 ) | ( n3063 & ~n8507 ) ;
  assign n8509 = n8508 ^ n2429 ^ n623 ;
  assign n8510 = ( ~n6640 & n8506 ) | ( ~n6640 & n8509 ) | ( n8506 & n8509 ) ;
  assign n8519 = n8518 ^ n8513 ^ n8510 ;
  assign n8520 = n6340 ^ n1107 ^ n926 ;
  assign n8521 = ( n1325 & ~n5609 ) | ( n1325 & n8520 ) | ( ~n5609 & n8520 ) ;
  assign n8524 = n5382 ^ n4088 ^ n492 ;
  assign n8525 = n8524 ^ n4708 ^ n708 ;
  assign n8526 = ( n3340 & ~n4872 ) | ( n3340 & n8525 ) | ( ~n4872 & n8525 ) ;
  assign n8522 = ( ~n770 & n4039 ) | ( ~n770 & n4884 ) | ( n4039 & n4884 ) ;
  assign n8523 = ( n4324 & ~n8101 ) | ( n4324 & n8522 ) | ( ~n8101 & n8522 ) ;
  assign n8527 = n8526 ^ n8523 ^ n7507 ;
  assign n8528 = ( ~n4460 & n8521 ) | ( ~n4460 & n8527 ) | ( n8521 & n8527 ) ;
  assign n8530 = ( n3268 & n5798 ) | ( n3268 & ~n8332 ) | ( n5798 & ~n8332 ) ;
  assign n8529 = n2968 ^ n2912 ^ n240 ;
  assign n8531 = n8530 ^ n8529 ^ n1085 ;
  assign n8532 = n3513 ^ n3016 ^ n1018 ;
  assign n8533 = n5545 ^ n2727 ^ n1971 ;
  assign n8534 = ( n3318 & n5466 ) | ( n3318 & ~n8533 ) | ( n5466 & ~n8533 ) ;
  assign n8535 = ( n4283 & n8532 ) | ( n4283 & n8534 ) | ( n8532 & n8534 ) ;
  assign n8539 = ( n5459 & n6393 ) | ( n5459 & ~n6980 ) | ( n6393 & ~n6980 ) ;
  assign n8536 = n8072 ^ n5264 ^ n4013 ;
  assign n8537 = n8536 ^ n5940 ^ n1500 ;
  assign n8538 = n8537 ^ n5893 ^ n1469 ;
  assign n8540 = n8539 ^ n8538 ^ n1318 ;
  assign n8541 = ( n7056 & ~n8535 ) | ( n7056 & n8540 ) | ( ~n8535 & n8540 ) ;
  assign n8543 = ( n2095 & n4745 ) | ( n2095 & ~n6094 ) | ( n4745 & ~n6094 ) ;
  assign n8544 = n8543 ^ n1059 ^ n650 ;
  assign n8545 = ( ~n6546 & n8476 ) | ( ~n6546 & n8544 ) | ( n8476 & n8544 ) ;
  assign n8546 = n8545 ^ n4124 ^ n694 ;
  assign n8542 = n4131 ^ n3308 ^ n1005 ;
  assign n8547 = n8546 ^ n8542 ^ n5726 ;
  assign n8548 = ( n1175 & n1871 ) | ( n1175 & n3960 ) | ( n1871 & n3960 ) ;
  assign n8549 = n8548 ^ n5359 ^ n2762 ;
  assign n8550 = ( n4763 & n7232 ) | ( n4763 & ~n8549 ) | ( n7232 & ~n8549 ) ;
  assign n8561 = ( n808 & n2225 ) | ( n808 & n4027 ) | ( n2225 & n4027 ) ;
  assign n8559 = n5445 ^ n1534 ^ n1318 ;
  assign n8560 = n8559 ^ n7313 ^ n4206 ;
  assign n8562 = n8561 ^ n8560 ^ n3767 ;
  assign n8563 = n8562 ^ n5329 ^ n4778 ;
  assign n8555 = ( ~n1481 & n5100 ) | ( ~n1481 & n6896 ) | ( n5100 & n6896 ) ;
  assign n8556 = n8555 ^ n3906 ^ n2464 ;
  assign n8557 = n8556 ^ n3524 ^ n1205 ;
  assign n8558 = n8557 ^ n5003 ^ n4587 ;
  assign n8564 = n8563 ^ n8558 ^ n4799 ;
  assign n8565 = ( n4773 & n7280 ) | ( n4773 & ~n8564 ) | ( n7280 & ~n8564 ) ;
  assign n8553 = n7465 ^ n5448 ^ n2170 ;
  assign n8554 = ( n592 & n3535 ) | ( n592 & ~n8553 ) | ( n3535 & ~n8553 ) ;
  assign n8566 = n8565 ^ n8554 ^ n5666 ;
  assign n8551 = ( n4584 & n4929 ) | ( n4584 & n7619 ) | ( n4929 & n7619 ) ;
  assign n8552 = ( n3527 & n6122 ) | ( n3527 & ~n8551 ) | ( n6122 & ~n8551 ) ;
  assign n8567 = n8566 ^ n8552 ^ n2881 ;
  assign n8568 = n4439 ^ n4318 ^ n2854 ;
  assign n8569 = n8568 ^ n1708 ^ n742 ;
  assign n8570 = n8569 ^ n3906 ^ n2925 ;
  assign n8571 = n7930 ^ n3577 ^ n1390 ;
  assign n8572 = ( ~n2928 & n8570 ) | ( ~n2928 & n8571 ) | ( n8570 & n8571 ) ;
  assign n8573 = ( x6 & n1937 ) | ( x6 & n6919 ) | ( n1937 & n6919 ) ;
  assign n8574 = ( n5769 & n8572 ) | ( n5769 & n8573 ) | ( n8572 & n8573 ) ;
  assign n8575 = n4512 ^ n2250 ^ n262 ;
  assign n8576 = ( n1287 & n4426 ) | ( n1287 & ~n4715 ) | ( n4426 & ~n4715 ) ;
  assign n8577 = ( n7325 & n8575 ) | ( n7325 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8578 = ( n8567 & ~n8574 ) | ( n8567 & n8577 ) | ( ~n8574 & n8577 ) ;
  assign n8579 = ( n618 & n771 ) | ( n618 & n8141 ) | ( n771 & n8141 ) ;
  assign n8580 = n7458 ^ n5539 ^ n4680 ;
  assign n8581 = n8580 ^ n1498 ^ n1353 ;
  assign n8591 = ( n3232 & ~n3989 ) | ( n3232 & n5137 ) | ( ~n3989 & n5137 ) ;
  assign n8582 = n3952 ^ n3021 ^ n2609 ;
  assign n8583 = ( n2882 & n4360 ) | ( n2882 & ~n8582 ) | ( n4360 & ~n8582 ) ;
  assign n8584 = n8583 ^ n5317 ^ n3378 ;
  assign n8585 = n6873 ^ n4058 ^ n3667 ;
  assign n8586 = n8585 ^ n5366 ^ n3257 ;
  assign n8587 = n8586 ^ n5336 ^ n2094 ;
  assign n8588 = ( n2607 & n5358 ) | ( n2607 & n7059 ) | ( n5358 & n7059 ) ;
  assign n8589 = ( n7425 & ~n8587 ) | ( n7425 & n8588 ) | ( ~n8587 & n8588 ) ;
  assign n8590 = ( n928 & ~n8584 ) | ( n928 & n8589 ) | ( ~n8584 & n8589 ) ;
  assign n8592 = n8591 ^ n8590 ^ n6880 ;
  assign n8597 = n6069 ^ n1448 ^ n196 ;
  assign n8598 = n8597 ^ n7473 ^ n5450 ;
  assign n8593 = n6940 ^ n2390 ^ n795 ;
  assign n8594 = n4073 ^ n1258 ^ x8 ;
  assign n8595 = ( n1545 & ~n3862 ) | ( n1545 & n8594 ) | ( ~n3862 & n8594 ) ;
  assign n8596 = ( ~n891 & n8593 ) | ( ~n891 & n8595 ) | ( n8593 & n8595 ) ;
  assign n8599 = n8598 ^ n8596 ^ n3254 ;
  assign n8600 = n6251 ^ n5193 ^ n4115 ;
  assign n8601 = ( n1028 & ~n5928 ) | ( n1028 & n8600 ) | ( ~n5928 & n8600 ) ;
  assign n8602 = ( n1821 & n7163 ) | ( n1821 & ~n8601 ) | ( n7163 & ~n8601 ) ;
  assign n8603 = n3108 ^ n1468 ^ n681 ;
  assign n8604 = n8603 ^ n4292 ^ n4186 ;
  assign n8605 = ( n1098 & ~n3046 ) | ( n1098 & n8604 ) | ( ~n3046 & n8604 ) ;
  assign n8606 = ( n1760 & n8251 ) | ( n1760 & n8605 ) | ( n8251 & n8605 ) ;
  assign n8607 = ( n1897 & n3183 ) | ( n1897 & ~n8606 ) | ( n3183 & ~n8606 ) ;
  assign n8608 = n6895 ^ n1516 ^ n1304 ;
  assign n8609 = n6348 ^ n3568 ^ n3473 ;
  assign n8610 = n5695 ^ n2996 ^ n2137 ;
  assign n8611 = ( n8608 & n8609 ) | ( n8608 & n8610 ) | ( n8609 & n8610 ) ;
  assign n8612 = n7071 ^ n3292 ^ n441 ;
  assign n8613 = n8612 ^ n6839 ^ n5289 ;
  assign n8614 = n7007 ^ n2758 ^ n1261 ;
  assign n8615 = ( n2541 & n3991 ) | ( n2541 & ~n8005 ) | ( n3991 & ~n8005 ) ;
  assign n8616 = ( n849 & n8614 ) | ( n849 & n8615 ) | ( n8614 & n8615 ) ;
  assign n8617 = ( n1806 & ~n1902 ) | ( n1806 & n5384 ) | ( ~n1902 & n5384 ) ;
  assign n8618 = ( n2810 & n6145 ) | ( n2810 & n8617 ) | ( n6145 & n8617 ) ;
  assign n8619 = n8618 ^ n3036 ^ n1287 ;
  assign n8620 = n8619 ^ n6043 ^ n4930 ;
  assign n8621 = ( n6314 & n7194 ) | ( n6314 & n8620 ) | ( n7194 & n8620 ) ;
  assign n8622 = ( ~n5287 & n8616 ) | ( ~n5287 & n8621 ) | ( n8616 & n8621 ) ;
  assign n8623 = n8622 ^ n6655 ^ n5556 ;
  assign n8627 = n4147 ^ n1958 ^ n414 ;
  assign n8624 = ( ~n1364 & n5072 ) | ( ~n1364 & n5739 ) | ( n5072 & n5739 ) ;
  assign n8625 = n8624 ^ n4831 ^ n981 ;
  assign n8626 = n8625 ^ n6065 ^ n5763 ;
  assign n8628 = n8627 ^ n8626 ^ n7767 ;
  assign n8629 = ( x115 & n3792 ) | ( x115 & n4894 ) | ( n3792 & n4894 ) ;
  assign n8638 = ( n4437 & ~n5418 ) | ( n4437 & n7051 ) | ( ~n5418 & n7051 ) ;
  assign n8637 = ( n2687 & n7316 ) | ( n2687 & ~n8285 ) | ( n7316 & ~n8285 ) ;
  assign n8634 = ( n913 & n3670 ) | ( n913 & ~n4005 ) | ( n3670 & ~n4005 ) ;
  assign n8632 = ( x120 & n328 ) | ( x120 & n876 ) | ( n328 & n876 ) ;
  assign n8630 = ( n412 & ~n1734 ) | ( n412 & n3441 ) | ( ~n1734 & n3441 ) ;
  assign n8631 = ( n984 & ~n2905 ) | ( n984 & n8630 ) | ( ~n2905 & n8630 ) ;
  assign n8633 = n8632 ^ n8631 ^ n2781 ;
  assign n8635 = n8634 ^ n8633 ^ n1516 ;
  assign n8636 = n8635 ^ n3581 ^ n1673 ;
  assign n8639 = n8638 ^ n8637 ^ n8636 ;
  assign n8640 = ( n6843 & n8629 ) | ( n6843 & n8639 ) | ( n8629 & n8639 ) ;
  assign n8643 = n3810 ^ n1039 ^ n966 ;
  assign n8641 = ( n1996 & n7493 ) | ( n1996 & ~n8632 ) | ( n7493 & ~n8632 ) ;
  assign n8642 = n8641 ^ n3091 ^ n764 ;
  assign n8644 = n8643 ^ n8642 ^ n1871 ;
  assign n8645 = ( ~n198 & n4425 ) | ( ~n198 & n6424 ) | ( n4425 & n6424 ) ;
  assign n8646 = ( n4370 & ~n8496 ) | ( n4370 & n8645 ) | ( ~n8496 & n8645 ) ;
  assign n8653 = n8147 ^ n6817 ^ n2202 ;
  assign n8650 = ( x103 & ~n1866 ) | ( x103 & n6147 ) | ( ~n1866 & n6147 ) ;
  assign n8651 = ( n1755 & n8355 ) | ( n1755 & n8650 ) | ( n8355 & n8650 ) ;
  assign n8652 = ( n2505 & n6024 ) | ( n2505 & n8651 ) | ( n6024 & n8651 ) ;
  assign n8647 = n6441 ^ n3192 ^ n1623 ;
  assign n8648 = n8647 ^ n5724 ^ n2154 ;
  assign n8649 = n8648 ^ n7165 ^ n6169 ;
  assign n8654 = n8653 ^ n8652 ^ n8649 ;
  assign n8655 = n8283 ^ n4124 ^ n294 ;
  assign n8656 = ( n6376 & n8654 ) | ( n6376 & ~n8655 ) | ( n8654 & ~n8655 ) ;
  assign n8658 = n4125 ^ n2419 ^ n1892 ;
  assign n8657 = n5178 ^ n2427 ^ n2321 ;
  assign n8659 = n8658 ^ n8657 ^ n5819 ;
  assign n8660 = n6830 ^ n5301 ^ n2216 ;
  assign n8661 = n8660 ^ n2466 ^ n1097 ;
  assign n8662 = n8661 ^ n4691 ^ x86 ;
  assign n8663 = ( ~n6886 & n7646 ) | ( ~n6886 & n8662 ) | ( n7646 & n8662 ) ;
  assign n8664 = n5400 ^ n4579 ^ n1854 ;
  assign n8665 = ( n1037 & ~n2105 ) | ( n1037 & n8664 ) | ( ~n2105 & n8664 ) ;
  assign n8666 = ( n279 & ~n1720 ) | ( n279 & n2779 ) | ( ~n1720 & n2779 ) ;
  assign n8667 = n8666 ^ n5572 ^ n2220 ;
  assign n8668 = ( ~n483 & n491 ) | ( ~n483 & n5650 ) | ( n491 & n5650 ) ;
  assign n8669 = ( ~n6089 & n7576 ) | ( ~n6089 & n8668 ) | ( n7576 & n8668 ) ;
  assign n8670 = ( ~n1482 & n3557 ) | ( ~n1482 & n8669 ) | ( n3557 & n8669 ) ;
  assign n8671 = ( n6883 & n8667 ) | ( n6883 & ~n8670 ) | ( n8667 & ~n8670 ) ;
  assign n8672 = ( x100 & n8665 ) | ( x100 & n8671 ) | ( n8665 & n8671 ) ;
  assign n8673 = n3331 ^ n1935 ^ n212 ;
  assign n8674 = n8516 ^ n4579 ^ n2627 ;
  assign n8675 = n8553 ^ n1357 ^ n1088 ;
  assign n8676 = ( n8673 & n8674 ) | ( n8673 & n8675 ) | ( n8674 & n8675 ) ;
  assign n8677 = ( n540 & n3294 ) | ( n540 & ~n8630 ) | ( n3294 & ~n8630 ) ;
  assign n8678 = ( n524 & n7190 ) | ( n524 & ~n8677 ) | ( n7190 & ~n8677 ) ;
  assign n8679 = ( n322 & ~n6773 ) | ( n322 & n8678 ) | ( ~n6773 & n8678 ) ;
  assign n8682 = ( n1788 & ~n2998 ) | ( n1788 & n5782 ) | ( ~n2998 & n5782 ) ;
  assign n8680 = ( n892 & n4729 ) | ( n892 & n5528 ) | ( n4729 & n5528 ) ;
  assign n8681 = n8680 ^ n7087 ^ n292 ;
  assign n8683 = n8682 ^ n8681 ^ n614 ;
  assign n8684 = n6142 ^ n5928 ^ n2131 ;
  assign n8685 = n2300 ^ n1213 ^ n818 ;
  assign n8686 = ( n678 & ~n701 ) | ( n678 & n6163 ) | ( ~n701 & n6163 ) ;
  assign n8687 = n8686 ^ n3045 ^ n150 ;
  assign n8688 = ( n294 & n1044 ) | ( n294 & ~n8629 ) | ( n1044 & ~n8629 ) ;
  assign n8689 = n8688 ^ n2802 ^ n906 ;
  assign n8690 = ( n8685 & ~n8687 ) | ( n8685 & n8689 ) | ( ~n8687 & n8689 ) ;
  assign n8691 = ( n1641 & ~n5815 ) | ( n1641 & n8690 ) | ( ~n5815 & n8690 ) ;
  assign n8692 = ( n502 & n660 ) | ( n502 & n8691 ) | ( n660 & n8691 ) ;
  assign n8693 = ( n1066 & n8684 ) | ( n1066 & ~n8692 ) | ( n8684 & ~n8692 ) ;
  assign n8695 = n8680 ^ n8084 ^ n1819 ;
  assign n8694 = n5476 ^ n4611 ^ n1371 ;
  assign n8696 = n8695 ^ n8694 ^ n252 ;
  assign n8697 = n8696 ^ n7862 ^ n1333 ;
  assign n8698 = ( n2412 & n5461 ) | ( n2412 & n8697 ) | ( n5461 & n8697 ) ;
  assign n8699 = n8698 ^ n7756 ^ n4557 ;
  assign n8700 = ( n3935 & n5526 ) | ( n3935 & ~n6162 ) | ( n5526 & ~n6162 ) ;
  assign n8701 = n7332 ^ n3371 ^ n504 ;
  assign n8702 = n2921 ^ n1099 ^ n286 ;
  assign n8703 = ( ~n3773 & n4272 ) | ( ~n3773 & n8702 ) | ( n4272 & n8702 ) ;
  assign n8704 = ( ~n1481 & n3729 ) | ( ~n1481 & n4882 ) | ( n3729 & n4882 ) ;
  assign n8705 = ( n3651 & ~n5042 ) | ( n3651 & n8704 ) | ( ~n5042 & n8704 ) ;
  assign n8706 = ( n3495 & ~n8703 ) | ( n3495 & n8705 ) | ( ~n8703 & n8705 ) ;
  assign n8707 = ( n2459 & ~n6257 ) | ( n2459 & n6945 ) | ( ~n6257 & n6945 ) ;
  assign n8708 = ( n499 & ~n1947 ) | ( n499 & n4299 ) | ( ~n1947 & n4299 ) ;
  assign n8709 = n8708 ^ n5118 ^ n4429 ;
  assign n8710 = n8626 ^ n6534 ^ n5590 ;
  assign n8713 = ( n317 & n548 ) | ( n317 & n3392 ) | ( n548 & n3392 ) ;
  assign n8714 = ( n1002 & n1187 ) | ( n1002 & ~n8713 ) | ( n1187 & ~n8713 ) ;
  assign n8711 = n7713 ^ n4563 ^ n496 ;
  assign n8712 = ( n2836 & n7798 ) | ( n2836 & ~n8711 ) | ( n7798 & ~n8711 ) ;
  assign n8715 = n8714 ^ n8712 ^ n501 ;
  assign n8716 = n2996 ^ n428 ^ n364 ;
  assign n8717 = ( n1506 & n2224 ) | ( n1506 & n8716 ) | ( n2224 & n8716 ) ;
  assign n8718 = n8717 ^ n2767 ^ n965 ;
  assign n8719 = n8718 ^ n3600 ^ n781 ;
  assign n8720 = n8719 ^ n7776 ^ n2908 ;
  assign n8721 = n8367 ^ n5911 ^ n1184 ;
  assign n8722 = ( n626 & n2704 ) | ( n626 & n2826 ) | ( n2704 & n2826 ) ;
  assign n8723 = n8722 ^ n3433 ^ n1633 ;
  assign n8724 = ( n1143 & n1503 ) | ( n1143 & n5466 ) | ( n1503 & n5466 ) ;
  assign n8725 = ( n6217 & n6817 ) | ( n6217 & n7649 ) | ( n6817 & n7649 ) ;
  assign n8726 = ( ~n8723 & n8724 ) | ( ~n8723 & n8725 ) | ( n8724 & n8725 ) ;
  assign n8728 = ( ~n1005 & n1437 ) | ( ~n1005 & n1714 ) | ( n1437 & n1714 ) ;
  assign n8727 = ( n3202 & ~n3927 ) | ( n3202 & n5968 ) | ( ~n3927 & n5968 ) ;
  assign n8729 = n8728 ^ n8727 ^ n8077 ;
  assign n8730 = ( n5538 & n8466 ) | ( n5538 & ~n8729 ) | ( n8466 & ~n8729 ) ;
  assign n8731 = ( ~n7071 & n7162 ) | ( ~n7071 & n8730 ) | ( n7162 & n8730 ) ;
  assign n8741 = n7150 ^ n2109 ^ n795 ;
  assign n8742 = n8741 ^ n2409 ^ n1327 ;
  assign n8743 = n8742 ^ n4970 ^ n310 ;
  assign n8738 = ( ~n740 & n4029 ) | ( ~n740 & n4172 ) | ( n4029 & n4172 ) ;
  assign n8739 = n8738 ^ n7956 ^ n4112 ;
  assign n8734 = ( n657 & n844 ) | ( n657 & ~n1832 ) | ( n844 & ~n1832 ) ;
  assign n8735 = ( ~n4572 & n5432 ) | ( ~n4572 & n6097 ) | ( n5432 & n6097 ) ;
  assign n8736 = ( n386 & n8734 ) | ( n386 & n8735 ) | ( n8734 & n8735 ) ;
  assign n8737 = n8736 ^ n4384 ^ n2311 ;
  assign n8740 = n8739 ^ n8737 ^ n2696 ;
  assign n8732 = n6667 ^ n4480 ^ n3059 ;
  assign n8733 = ( n1715 & n3603 ) | ( n1715 & ~n8732 ) | ( n3603 & ~n8732 ) ;
  assign n8744 = n8743 ^ n8740 ^ n8733 ;
  assign n8745 = ( n2234 & n2902 ) | ( n2234 & ~n2975 ) | ( n2902 & ~n2975 ) ;
  assign n8746 = ( n952 & n2001 ) | ( n952 & n4810 ) | ( n2001 & n4810 ) ;
  assign n8747 = ( n1766 & n1819 ) | ( n1766 & ~n2411 ) | ( n1819 & ~n2411 ) ;
  assign n8748 = ( n2555 & n7083 ) | ( n2555 & n8747 ) | ( n7083 & n8747 ) ;
  assign n8749 = ( n3936 & ~n8746 ) | ( n3936 & n8748 ) | ( ~n8746 & n8748 ) ;
  assign n8750 = n8749 ^ n7512 ^ n5903 ;
  assign n8751 = ( n642 & n8745 ) | ( n642 & n8750 ) | ( n8745 & n8750 ) ;
  assign n8752 = ( n2910 & n3243 ) | ( n2910 & ~n6502 ) | ( n3243 & ~n6502 ) ;
  assign n8753 = n5054 ^ n1290 ^ x9 ;
  assign n8754 = n2037 ^ n1439 ^ n613 ;
  assign n8755 = ( ~n3132 & n4364 ) | ( ~n3132 & n8754 ) | ( n4364 & n8754 ) ;
  assign n8756 = n8755 ^ n4300 ^ n807 ;
  assign n8757 = n8756 ^ n5741 ^ n5051 ;
  assign n8758 = n2764 ^ n2252 ^ n850 ;
  assign n8759 = ( ~n1323 & n4686 ) | ( ~n1323 & n8758 ) | ( n4686 & n8758 ) ;
  assign n8760 = ( ~n8753 & n8757 ) | ( ~n8753 & n8759 ) | ( n8757 & n8759 ) ;
  assign n8761 = n8597 ^ n3997 ^ n2323 ;
  assign n8762 = ( n416 & n8760 ) | ( n416 & n8761 ) | ( n8760 & n8761 ) ;
  assign n8763 = ( n1699 & n6463 ) | ( n1699 & n8762 ) | ( n6463 & n8762 ) ;
  assign n8764 = ( n1218 & ~n1287 ) | ( n1218 & n8763 ) | ( ~n1287 & n8763 ) ;
  assign n8775 = ( n2543 & ~n5256 ) | ( n2543 & n5408 ) | ( ~n5256 & n5408 ) ;
  assign n8765 = ( n1501 & ~n1734 ) | ( n1501 & n2880 ) | ( ~n1734 & n2880 ) ;
  assign n8766 = ( n2829 & n2934 ) | ( n2829 & n4364 ) | ( n2934 & n4364 ) ;
  assign n8767 = ( n2218 & ~n8765 ) | ( n2218 & n8766 ) | ( ~n8765 & n8766 ) ;
  assign n8768 = n8767 ^ n4954 ^ n1369 ;
  assign n8769 = n2330 ^ n2014 ^ n1603 ;
  assign n8770 = ( n268 & ~n3192 ) | ( n268 & n8769 ) | ( ~n3192 & n8769 ) ;
  assign n8771 = ( n388 & ~n815 ) | ( n388 & n4122 ) | ( ~n815 & n4122 ) ;
  assign n8772 = n8771 ^ n6292 ^ n2908 ;
  assign n8773 = ( n1872 & ~n8770 ) | ( n1872 & n8772 ) | ( ~n8770 & n8772 ) ;
  assign n8774 = ( ~n6616 & n8768 ) | ( ~n6616 & n8773 ) | ( n8768 & n8773 ) ;
  assign n8776 = n8775 ^ n8774 ^ n5426 ;
  assign n8782 = ( x123 & n3812 ) | ( x123 & ~n5859 ) | ( n3812 & ~n5859 ) ;
  assign n8783 = n8782 ^ n7890 ^ n222 ;
  assign n8778 = ( ~n1168 & n1246 ) | ( ~n1168 & n4052 ) | ( n1246 & n4052 ) ;
  assign n8779 = n8778 ^ n2259 ^ n1546 ;
  assign n8777 = n2834 ^ n2324 ^ n1280 ;
  assign n8780 = n8779 ^ n8777 ^ x8 ;
  assign n8781 = n8780 ^ n8472 ^ n823 ;
  assign n8784 = n8783 ^ n8781 ^ n242 ;
  assign n8786 = ( n1685 & ~n3429 ) | ( n1685 & n3804 ) | ( ~n3429 & n3804 ) ;
  assign n8785 = ( n594 & n1260 ) | ( n594 & ~n2449 ) | ( n1260 & ~n2449 ) ;
  assign n8787 = n8786 ^ n8785 ^ n2957 ;
  assign n8788 = n4566 ^ n2286 ^ n1953 ;
  assign n8789 = n5624 ^ n3001 ^ n2077 ;
  assign n8790 = ( n1873 & ~n4359 ) | ( n1873 & n8789 ) | ( ~n4359 & n8789 ) ;
  assign n8791 = ( n1994 & ~n5451 ) | ( n1994 & n8790 ) | ( ~n5451 & n8790 ) ;
  assign n8792 = ( n4471 & ~n8788 ) | ( n4471 & n8791 ) | ( ~n8788 & n8791 ) ;
  assign n8793 = ( ~n2287 & n4228 ) | ( ~n2287 & n8792 ) | ( n4228 & n8792 ) ;
  assign n8794 = ( ~n3206 & n3522 ) | ( ~n3206 & n5263 ) | ( n3522 & n5263 ) ;
  assign n8795 = n8794 ^ n5040 ^ n928 ;
  assign n8796 = ( n172 & n206 ) | ( n172 & n8795 ) | ( n206 & n8795 ) ;
  assign n8797 = ( n2211 & n2325 ) | ( n2211 & ~n8060 ) | ( n2325 & ~n8060 ) ;
  assign n8798 = n8797 ^ n6189 ^ n1485 ;
  assign n8799 = n8798 ^ n4733 ^ n2891 ;
  assign n8807 = n4444 ^ n842 ^ n373 ;
  assign n8804 = n973 ^ n482 ^ n462 ;
  assign n8805 = n8804 ^ n8630 ^ n5428 ;
  assign n8806 = ( n5007 & n6690 ) | ( n5007 & ~n8805 ) | ( n6690 & ~n8805 ) ;
  assign n8800 = n5709 ^ n2657 ^ n1082 ;
  assign n8801 = n8800 ^ n5983 ^ n2054 ;
  assign n8802 = n8801 ^ n4507 ^ n3603 ;
  assign n8803 = n8802 ^ n4085 ^ n1598 ;
  assign n8808 = n8807 ^ n8806 ^ n8803 ;
  assign n8809 = ( ~n8796 & n8799 ) | ( ~n8796 & n8808 ) | ( n8799 & n8808 ) ;
  assign n8810 = ( ~x24 & n3035 ) | ( ~x24 & n6483 ) | ( n3035 & n6483 ) ;
  assign n8811 = n8810 ^ n6301 ^ n2899 ;
  assign n8812 = n8811 ^ n5155 ^ n5125 ;
  assign n8814 = ( ~n2699 & n4616 ) | ( ~n2699 & n6085 ) | ( n4616 & n6085 ) ;
  assign n8813 = ( ~n484 & n1961 ) | ( ~n484 & n2084 ) | ( n1961 & n2084 ) ;
  assign n8815 = n8814 ^ n8813 ^ n2784 ;
  assign n8816 = ( n376 & n3096 ) | ( n376 & ~n8815 ) | ( n3096 & ~n8815 ) ;
  assign n8817 = ( n2377 & ~n4642 ) | ( n2377 & n6643 ) | ( ~n4642 & n6643 ) ;
  assign n8818 = n3960 ^ n871 ^ n715 ;
  assign n8819 = ( n877 & ~n8817 ) | ( n877 & n8818 ) | ( ~n8817 & n8818 ) ;
  assign n8825 = ( n1256 & ~n1715 ) | ( n1256 & n6356 ) | ( ~n1715 & n6356 ) ;
  assign n8824 = n1352 ^ n1228 ^ n838 ;
  assign n8820 = ( n1190 & n1577 ) | ( n1190 & ~n2145 ) | ( n1577 & ~n2145 ) ;
  assign n8821 = n4158 ^ n3544 ^ n1451 ;
  assign n8822 = ( n707 & n5857 ) | ( n707 & n8821 ) | ( n5857 & n8821 ) ;
  assign n8823 = ( n7830 & n8820 ) | ( n7830 & ~n8822 ) | ( n8820 & ~n8822 ) ;
  assign n8826 = n8825 ^ n8824 ^ n8823 ;
  assign n8831 = n4434 ^ n2095 ^ n508 ;
  assign n8827 = ( n1459 & ~n1568 ) | ( n1459 & n3528 ) | ( ~n1568 & n3528 ) ;
  assign n8828 = ( n146 & n3399 ) | ( n146 & n5953 ) | ( n3399 & n5953 ) ;
  assign n8829 = n8828 ^ n4816 ^ n1404 ;
  assign n8830 = ( ~n8383 & n8827 ) | ( ~n8383 & n8829 ) | ( n8827 & n8829 ) ;
  assign n8832 = n8831 ^ n8830 ^ n5978 ;
  assign n8833 = n7864 ^ n5666 ^ n1983 ;
  assign n8834 = n2062 ^ n1732 ^ n146 ;
  assign n8836 = n2189 ^ n1628 ^ n671 ;
  assign n8837 = ( ~n540 & n2452 ) | ( ~n540 & n8836 ) | ( n2452 & n8836 ) ;
  assign n8838 = n8837 ^ n3864 ^ n3199 ;
  assign n8835 = n6425 ^ n6222 ^ n2288 ;
  assign n8839 = n8838 ^ n8835 ^ n3071 ;
  assign n8840 = ( n3525 & ~n8834 ) | ( n3525 & n8839 ) | ( ~n8834 & n8839 ) ;
  assign n8841 = ( n4263 & ~n8833 ) | ( n4263 & n8840 ) | ( ~n8833 & n8840 ) ;
  assign n8842 = ( ~n2788 & n2840 ) | ( ~n2788 & n3212 ) | ( n2840 & n3212 ) ;
  assign n8843 = ( n2359 & n2606 ) | ( n2359 & ~n5871 ) | ( n2606 & ~n5871 ) ;
  assign n8844 = ( n892 & n3827 ) | ( n892 & ~n8843 ) | ( n3827 & ~n8843 ) ;
  assign n8845 = ( n5295 & n8842 ) | ( n5295 & n8844 ) | ( n8842 & n8844 ) ;
  assign n8846 = ( n2133 & ~n3466 ) | ( n2133 & n8845 ) | ( ~n3466 & n8845 ) ;
  assign n8847 = ( n5724 & n6795 ) | ( n5724 & ~n8846 ) | ( n6795 & ~n8846 ) ;
  assign n8848 = ( n2148 & n2790 ) | ( n2148 & n3736 ) | ( n2790 & n3736 ) ;
  assign n8849 = n8848 ^ n4881 ^ n2649 ;
  assign n8850 = n8849 ^ n7665 ^ n4416 ;
  assign n8851 = n3624 ^ n2928 ^ n1830 ;
  assign n8852 = n4537 ^ n1662 ^ n235 ;
  assign n8853 = ( n1237 & ~n4157 ) | ( n1237 & n8852 ) | ( ~n4157 & n8852 ) ;
  assign n8854 = ( n3950 & n4250 ) | ( n3950 & n8853 ) | ( n4250 & n8853 ) ;
  assign n8855 = ( ~x106 & n4207 ) | ( ~x106 & n4869 ) | ( n4207 & n4869 ) ;
  assign n8856 = ( n1494 & n7238 ) | ( n1494 & n8855 ) | ( n7238 & n8855 ) ;
  assign n8857 = ( n1087 & n7671 ) | ( n1087 & ~n8856 ) | ( n7671 & ~n8856 ) ;
  assign n8858 = ( ~n2690 & n2701 ) | ( ~n2690 & n8857 ) | ( n2701 & n8857 ) ;
  assign n8859 = ( n1076 & ~n2943 ) | ( n1076 & n3100 ) | ( ~n2943 & n3100 ) ;
  assign n8860 = ( ~n5621 & n8858 ) | ( ~n5621 & n8859 ) | ( n8858 & n8859 ) ;
  assign n8861 = ( n5386 & n8854 ) | ( n5386 & n8860 ) | ( n8854 & n8860 ) ;
  assign n8862 = ( n1694 & n8851 ) | ( n1694 & n8861 ) | ( n8851 & n8861 ) ;
  assign n8863 = n8657 ^ n2731 ^ x118 ;
  assign n8864 = ( ~n1120 & n2095 ) | ( ~n1120 & n2872 ) | ( n2095 & n2872 ) ;
  assign n8865 = n2855 ^ n1587 ^ n298 ;
  assign n8866 = ( ~n2007 & n3254 ) | ( ~n2007 & n8865 ) | ( n3254 & n8865 ) ;
  assign n8867 = ( n2313 & n4285 ) | ( n2313 & n6055 ) | ( n4285 & n6055 ) ;
  assign n8868 = n8059 ^ n5521 ^ n2526 ;
  assign n8869 = ( n6787 & ~n8867 ) | ( n6787 & n8868 ) | ( ~n8867 & n8868 ) ;
  assign n8870 = ( n4005 & ~n8866 ) | ( n4005 & n8869 ) | ( ~n8866 & n8869 ) ;
  assign n8871 = n8870 ^ n8716 ^ n4849 ;
  assign n8872 = ( n8863 & ~n8864 ) | ( n8863 & n8871 ) | ( ~n8864 & n8871 ) ;
  assign n8873 = ( ~n2566 & n2661 ) | ( ~n2566 & n5120 ) | ( n2661 & n5120 ) ;
  assign n8874 = n8873 ^ n6404 ^ n2759 ;
  assign n8875 = n4210 ^ n2108 ^ n273 ;
  assign n8877 = ( n7470 & n7700 ) | ( n7470 & ~n8741 ) | ( n7700 & ~n8741 ) ;
  assign n8876 = ( ~n1749 & n4484 ) | ( ~n1749 & n6603 ) | ( n4484 & n6603 ) ;
  assign n8878 = n8877 ^ n8876 ^ n1128 ;
  assign n8885 = n7162 ^ n6210 ^ n1412 ;
  assign n8879 = ( n2560 & ~n2942 ) | ( n2560 & n3937 ) | ( ~n2942 & n3937 ) ;
  assign n8880 = n3458 ^ n1080 ^ n1018 ;
  assign n8881 = n8880 ^ n706 ^ n552 ;
  assign n8882 = n5567 ^ n5360 ^ n3138 ;
  assign n8883 = ( n6188 & n8881 ) | ( n6188 & n8882 ) | ( n8881 & n8882 ) ;
  assign n8884 = ( n5945 & n8879 ) | ( n5945 & ~n8883 ) | ( n8879 & ~n8883 ) ;
  assign n8886 = n8885 ^ n8884 ^ n3645 ;
  assign n8887 = ( n8875 & n8878 ) | ( n8875 & ~n8886 ) | ( n8878 & ~n8886 ) ;
  assign n8888 = ( n2160 & n3884 ) | ( n2160 & n5797 ) | ( n3884 & n5797 ) ;
  assign n8890 = n3108 ^ n2245 ^ x47 ;
  assign n8891 = ( ~n6206 & n6882 ) | ( ~n6206 & n8890 ) | ( n6882 & n8890 ) ;
  assign n8889 = ( n701 & ~n3730 ) | ( n701 & n5949 ) | ( ~n3730 & n5949 ) ;
  assign n8892 = n8891 ^ n8889 ^ n8161 ;
  assign n8893 = n8892 ^ n7713 ^ n2351 ;
  assign n8894 = ( ~n1064 & n3236 ) | ( ~n1064 & n4852 ) | ( n3236 & n4852 ) ;
  assign n8895 = ( n1761 & n2292 ) | ( n1761 & n5251 ) | ( n2292 & n5251 ) ;
  assign n8896 = n8895 ^ n6366 ^ n790 ;
  assign n8897 = ( n1914 & n8724 ) | ( n1914 & ~n8896 ) | ( n8724 & ~n8896 ) ;
  assign n8905 = ( n1060 & ~n2746 ) | ( n1060 & n4641 ) | ( ~n2746 & n4641 ) ;
  assign n8906 = n8905 ^ n7277 ^ n2872 ;
  assign n8907 = ( ~n443 & n3830 ) | ( ~n443 & n8749 ) | ( n3830 & n8749 ) ;
  assign n8908 = ( n8210 & ~n8906 ) | ( n8210 & n8907 ) | ( ~n8906 & n8907 ) ;
  assign n8898 = n4459 ^ n1438 ^ n1280 ;
  assign n8899 = ( n826 & ~n4167 ) | ( n826 & n8898 ) | ( ~n4167 & n8898 ) ;
  assign n8900 = n8899 ^ n2757 ^ n1989 ;
  assign n8901 = n7788 ^ n3388 ^ n2920 ;
  assign n8902 = ( n460 & ~n4992 ) | ( n460 & n8901 ) | ( ~n4992 & n8901 ) ;
  assign n8903 = ( n2664 & ~n7970 ) | ( n2664 & n8902 ) | ( ~n7970 & n8902 ) ;
  assign n8904 = ( n1062 & ~n8900 ) | ( n1062 & n8903 ) | ( ~n8900 & n8903 ) ;
  assign n8909 = n8908 ^ n8904 ^ n4864 ;
  assign n8911 = ( n2179 & ~n3427 ) | ( n2179 & n5196 ) | ( ~n3427 & n5196 ) ;
  assign n8912 = n4687 ^ n2820 ^ x2 ;
  assign n8913 = ( n491 & n1327 ) | ( n491 & n8912 ) | ( n1327 & n8912 ) ;
  assign n8914 = n8913 ^ n7475 ^ n2984 ;
  assign n8915 = ( n1271 & n8911 ) | ( n1271 & n8914 ) | ( n8911 & n8914 ) ;
  assign n8910 = ( ~n3201 & n3897 ) | ( ~n3201 & n6143 ) | ( n3897 & n6143 ) ;
  assign n8916 = n8915 ^ n8910 ^ n1928 ;
  assign n8926 = ( n3687 & ~n5309 ) | ( n3687 & n6936 ) | ( ~n5309 & n6936 ) ;
  assign n8917 = n7582 ^ n5472 ^ n4939 ;
  assign n8918 = n3959 ^ n551 ^ n359 ;
  assign n8919 = n8918 ^ n949 ^ n488 ;
  assign n8920 = n8919 ^ n879 ^ n732 ;
  assign n8921 = n5178 ^ n1623 ^ n238 ;
  assign n8922 = n8921 ^ n6995 ^ n4689 ;
  assign n8923 = ( n3676 & n8920 ) | ( n3676 & n8922 ) | ( n8920 & n8922 ) ;
  assign n8924 = ( n3205 & ~n3874 ) | ( n3205 & n4506 ) | ( ~n3874 & n4506 ) ;
  assign n8925 = ( n8917 & ~n8923 ) | ( n8917 & n8924 ) | ( ~n8923 & n8924 ) ;
  assign n8927 = n8926 ^ n8925 ^ n881 ;
  assign n8934 = n6015 ^ n3665 ^ n2225 ;
  assign n8935 = n8934 ^ n8390 ^ n5401 ;
  assign n8936 = n8935 ^ n3134 ^ n2305 ;
  assign n8928 = n4498 ^ n900 ^ n479 ;
  assign n8929 = ( n6019 & n8515 ) | ( n6019 & ~n8928 ) | ( n8515 & ~n8928 ) ;
  assign n8930 = n8929 ^ n1562 ^ n464 ;
  assign n8931 = n6439 ^ n585 ^ n333 ;
  assign n8932 = n8931 ^ n5153 ^ n2550 ;
  assign n8933 = ( n5616 & ~n8930 ) | ( n5616 & n8932 ) | ( ~n8930 & n8932 ) ;
  assign n8937 = n8936 ^ n8933 ^ n3036 ;
  assign n8960 = n7987 ^ n5040 ^ n454 ;
  assign n8949 = ( n3281 & ~n5073 ) | ( n3281 & n8283 ) | ( ~n5073 & n8283 ) ;
  assign n8950 = n8949 ^ n5627 ^ n881 ;
  assign n8951 = ( n1294 & ~n4647 ) | ( n1294 & n4686 ) | ( ~n4647 & n4686 ) ;
  assign n8952 = n1669 ^ n715 ^ n430 ;
  assign n8953 = n8952 ^ n4856 ^ x5 ;
  assign n8954 = n8128 ^ n7520 ^ n5007 ;
  assign n8955 = ( n3114 & n8133 ) | ( n3114 & n8954 ) | ( n8133 & n8954 ) ;
  assign n8956 = ( ~n2889 & n8953 ) | ( ~n2889 & n8955 ) | ( n8953 & n8955 ) ;
  assign n8957 = ( n7627 & n8951 ) | ( n7627 & ~n8956 ) | ( n8951 & ~n8956 ) ;
  assign n8958 = ( n2239 & n8906 ) | ( n2239 & n8957 ) | ( n8906 & n8957 ) ;
  assign n8959 = ( n1977 & n8950 ) | ( n1977 & ~n8958 ) | ( n8950 & ~n8958 ) ;
  assign n8938 = n4166 ^ n3283 ^ n2892 ;
  assign n8939 = ( n3150 & n7577 ) | ( n3150 & ~n8938 ) | ( n7577 & ~n8938 ) ;
  assign n8943 = n3968 ^ n3726 ^ n776 ;
  assign n8940 = ( n1016 & n1080 ) | ( n1016 & n1828 ) | ( n1080 & n1828 ) ;
  assign n8941 = ( n198 & n3986 ) | ( n198 & n7310 ) | ( n3986 & n7310 ) ;
  assign n8942 = ( ~n375 & n8940 ) | ( ~n375 & n8941 ) | ( n8940 & n8941 ) ;
  assign n8944 = n8943 ^ n8942 ^ n4170 ;
  assign n8945 = ( n5150 & n8939 ) | ( n5150 & n8944 ) | ( n8939 & n8944 ) ;
  assign n8946 = n7954 ^ n6793 ^ n1875 ;
  assign n8947 = n8946 ^ n3822 ^ n771 ;
  assign n8948 = ( n7858 & ~n8945 ) | ( n7858 & n8947 ) | ( ~n8945 & n8947 ) ;
  assign n8961 = n8960 ^ n8959 ^ n8948 ;
  assign n8963 = ( n489 & ~n539 ) | ( n489 & n1760 ) | ( ~n539 & n1760 ) ;
  assign n8962 = ( n2927 & n7459 ) | ( n2927 & ~n7746 ) | ( n7459 & ~n7746 ) ;
  assign n8964 = n8963 ^ n8962 ^ n7688 ;
  assign n8967 = n7762 ^ n3554 ^ n1792 ;
  assign n8968 = ( n2318 & n2375 ) | ( n2318 & n8967 ) | ( n2375 & n8967 ) ;
  assign n8969 = ( ~n3972 & n4405 ) | ( ~n3972 & n8512 ) | ( n4405 & n8512 ) ;
  assign n8970 = ( n2606 & n8968 ) | ( n2606 & ~n8969 ) | ( n8968 & ~n8969 ) ;
  assign n8965 = ( n1233 & n6733 ) | ( n1233 & n8637 ) | ( n6733 & n8637 ) ;
  assign n8966 = ( n925 & n5251 ) | ( n925 & n8965 ) | ( n5251 & n8965 ) ;
  assign n8971 = n8970 ^ n8966 ^ n7767 ;
  assign n8972 = ( x112 & n6460 ) | ( x112 & ~n7093 ) | ( n6460 & ~n7093 ) ;
  assign n8973 = n8972 ^ n3976 ^ n1238 ;
  assign n8974 = ( n2703 & n4997 ) | ( n2703 & n6358 ) | ( n4997 & n6358 ) ;
  assign n8975 = ( n491 & ~n3078 ) | ( n491 & n8974 ) | ( ~n3078 & n8974 ) ;
  assign n8976 = ( n748 & n1999 ) | ( n748 & ~n8975 ) | ( n1999 & ~n8975 ) ;
  assign n8977 = ( n846 & ~n1049 ) | ( n846 & n7679 ) | ( ~n1049 & n7679 ) ;
  assign n8978 = ( ~n8309 & n8939 ) | ( ~n8309 & n8977 ) | ( n8939 & n8977 ) ;
  assign n8979 = n8480 ^ n3489 ^ n2362 ;
  assign n8980 = ( n1771 & n5680 ) | ( n1771 & ~n6760 ) | ( n5680 & ~n6760 ) ;
  assign n8981 = n6669 ^ n5763 ^ n1975 ;
  assign n8982 = n8981 ^ n2602 ^ n288 ;
  assign n8983 = n8982 ^ n7755 ^ n2991 ;
  assign n8986 = n2061 ^ n1053 ^ x88 ;
  assign n8984 = n8310 ^ n2496 ^ n2423 ;
  assign n8985 = ( n3069 & n4926 ) | ( n3069 & ~n8984 ) | ( n4926 & ~n8984 ) ;
  assign n8987 = n8986 ^ n8985 ^ n4743 ;
  assign n8988 = ( ~n475 & n7558 ) | ( ~n475 & n8987 ) | ( n7558 & n8987 ) ;
  assign n8989 = ( n2920 & n3380 ) | ( n2920 & ~n8988 ) | ( n3380 & ~n8988 ) ;
  assign n8990 = n8989 ^ n8675 ^ n8436 ;
  assign n8991 = ( n8980 & n8983 ) | ( n8980 & n8990 ) | ( n8983 & n8990 ) ;
  assign n8992 = ( ~n639 & n4855 ) | ( ~n639 & n8837 ) | ( n4855 & n8837 ) ;
  assign n8993 = ( n465 & n5563 ) | ( n465 & ~n8992 ) | ( n5563 & ~n8992 ) ;
  assign n8994 = ( n2224 & n7085 ) | ( n2224 & ~n8717 ) | ( n7085 & ~n8717 ) ;
  assign n8995 = n8994 ^ n8189 ^ n7383 ;
  assign n8996 = ( n390 & ~n6262 ) | ( n390 & n6263 ) | ( ~n6262 & n6263 ) ;
  assign n8997 = n8996 ^ n7114 ^ n1971 ;
  assign n8998 = n8997 ^ n6684 ^ n5581 ;
  assign n8999 = n8998 ^ n5142 ^ n2794 ;
  assign n9000 = n6734 ^ n5315 ^ n3875 ;
  assign n9001 = n9000 ^ n6163 ^ n1854 ;
  assign n9002 = ( n3046 & ~n4126 ) | ( n3046 & n9001 ) | ( ~n4126 & n9001 ) ;
  assign n9003 = n5237 ^ n4315 ^ n3436 ;
  assign n9004 = ( ~n4823 & n5315 ) | ( ~n4823 & n9003 ) | ( n5315 & n9003 ) ;
  assign n9005 = n6736 ^ n5708 ^ n4238 ;
  assign n9006 = ( ~n363 & n1955 ) | ( ~n363 & n4150 ) | ( n1955 & n4150 ) ;
  assign n9007 = n9006 ^ n3243 ^ n1145 ;
  assign n9013 = ( x43 & ~n2057 ) | ( x43 & n3175 ) | ( ~n2057 & n3175 ) ;
  assign n9014 = ( n540 & n5798 ) | ( n540 & n9013 ) | ( n5798 & n9013 ) ;
  assign n9008 = ( ~n434 & n2473 ) | ( ~n434 & n3433 ) | ( n2473 & n3433 ) ;
  assign n9009 = n9008 ^ n1571 ^ n656 ;
  assign n9010 = ( n480 & n1672 ) | ( n480 & n4351 ) | ( n1672 & n4351 ) ;
  assign n9011 = n9010 ^ n7490 ^ n5698 ;
  assign n9012 = ( ~n4640 & n9009 ) | ( ~n4640 & n9011 ) | ( n9009 & n9011 ) ;
  assign n9015 = n9014 ^ n9012 ^ n4527 ;
  assign n9016 = ( ~n3544 & n9007 ) | ( ~n3544 & n9015 ) | ( n9007 & n9015 ) ;
  assign n9017 = ( ~n386 & n9005 ) | ( ~n386 & n9016 ) | ( n9005 & n9016 ) ;
  assign n9018 = ( n2867 & ~n9004 ) | ( n2867 & n9017 ) | ( ~n9004 & n9017 ) ;
  assign n9019 = ( n328 & n1529 ) | ( n328 & ~n4370 ) | ( n1529 & ~n4370 ) ;
  assign n9020 = n8759 ^ n4731 ^ n2386 ;
  assign n9021 = n9020 ^ n8127 ^ n5097 ;
  assign n9022 = ( n2673 & n5176 ) | ( n2673 & n8918 ) | ( n5176 & n8918 ) ;
  assign n9023 = ( n9019 & ~n9021 ) | ( n9019 & n9022 ) | ( ~n9021 & n9022 ) ;
  assign n9025 = ( ~n388 & n1684 ) | ( ~n388 & n2475 ) | ( n1684 & n2475 ) ;
  assign n9024 = n3962 ^ n1570 ^ n1453 ;
  assign n9026 = n9025 ^ n9024 ^ n2228 ;
  assign n9027 = ( n3244 & n7709 ) | ( n3244 & ~n9026 ) | ( n7709 & ~n9026 ) ;
  assign n9029 = ( n170 & ~n2216 ) | ( n170 & n7007 ) | ( ~n2216 & n7007 ) ;
  assign n9028 = n8666 ^ n1977 ^ n1341 ;
  assign n9030 = n9029 ^ n9028 ^ n8300 ;
  assign n9031 = ( ~n2293 & n7272 ) | ( ~n2293 & n8507 ) | ( n7272 & n8507 ) ;
  assign n9032 = ( n1734 & n2868 ) | ( n1734 & ~n8912 ) | ( n2868 & ~n8912 ) ;
  assign n9033 = ( ~n1766 & n5841 ) | ( ~n1766 & n9032 ) | ( n5841 & n9032 ) ;
  assign n9034 = ( n3310 & ~n3557 ) | ( n3310 & n9033 ) | ( ~n3557 & n9033 ) ;
  assign n9035 = ( n3221 & n5968 ) | ( n3221 & n9034 ) | ( n5968 & n9034 ) ;
  assign n9036 = ( ~n6949 & n9031 ) | ( ~n6949 & n9035 ) | ( n9031 & n9035 ) ;
  assign n9037 = n8238 ^ n6155 ^ n4028 ;
  assign n9038 = n5214 ^ n3744 ^ n1539 ;
  assign n9039 = ( ~n2060 & n2632 ) | ( ~n2060 & n9038 ) | ( n2632 & n9038 ) ;
  assign n9040 = n9039 ^ n3927 ^ n1473 ;
  assign n9041 = ( n2237 & n8163 ) | ( n2237 & ~n9040 ) | ( n8163 & ~n9040 ) ;
  assign n9042 = n9041 ^ n5879 ^ n5090 ;
  assign n9045 = n3808 ^ n2258 ^ x93 ;
  assign n9046 = n9045 ^ n2148 ^ n716 ;
  assign n9047 = ( n1418 & n3790 ) | ( n1418 & n9046 ) | ( n3790 & n9046 ) ;
  assign n9043 = ( n1029 & ~n2706 ) | ( n1029 & n5318 ) | ( ~n2706 & n5318 ) ;
  assign n9044 = n9043 ^ n2678 ^ n1504 ;
  assign n9048 = n9047 ^ n9044 ^ n3218 ;
  assign n9049 = n9048 ^ n7670 ^ n6240 ;
  assign n9058 = n5497 ^ n3831 ^ n2051 ;
  assign n9059 = n9058 ^ n6513 ^ n716 ;
  assign n9060 = ( n4631 & n5176 ) | ( n4631 & ~n9059 ) | ( n5176 & ~n9059 ) ;
  assign n9050 = n1972 ^ n1767 ^ n496 ;
  assign n9051 = ( ~n705 & n4512 ) | ( ~n705 & n9050 ) | ( n4512 & n9050 ) ;
  assign n9052 = ( n3699 & n7548 ) | ( n3699 & n9051 ) | ( n7548 & n9051 ) ;
  assign n9055 = n7902 ^ n5313 ^ n3168 ;
  assign n9053 = n3984 ^ n1812 ^ n295 ;
  assign n9054 = ( ~n1403 & n4210 ) | ( ~n1403 & n9053 ) | ( n4210 & n9053 ) ;
  assign n9056 = n9055 ^ n9054 ^ n7484 ;
  assign n9057 = ( ~n7595 & n9052 ) | ( ~n7595 & n9056 ) | ( n9052 & n9056 ) ;
  assign n9061 = n9060 ^ n9057 ^ n3775 ;
  assign n9062 = ( n1985 & n2024 ) | ( n1985 & ~n8734 ) | ( n2024 & ~n8734 ) ;
  assign n9063 = ( ~x48 & n465 ) | ( ~x48 & n1752 ) | ( n465 & n1752 ) ;
  assign n9064 = n9063 ^ n4383 ^ n3793 ;
  assign n9065 = ( n5895 & n9062 ) | ( n5895 & n9064 ) | ( n9062 & n9064 ) ;
  assign n9066 = n6600 ^ n1320 ^ n504 ;
  assign n9067 = n9066 ^ n4885 ^ n3068 ;
  assign n9068 = ( n4626 & n5855 ) | ( n4626 & ~n9067 ) | ( n5855 & ~n9067 ) ;
  assign n9069 = n8686 ^ n2294 ^ n1280 ;
  assign n9070 = n9069 ^ n876 ^ n396 ;
  assign n9071 = ( n9065 & n9068 ) | ( n9065 & n9070 ) | ( n9068 & n9070 ) ;
  assign n9081 = n5476 ^ n5175 ^ n795 ;
  assign n9082 = ( ~n1197 & n6382 ) | ( ~n1197 & n9081 ) | ( n6382 & n9081 ) ;
  assign n9072 = n1829 ^ n1780 ^ n1749 ;
  assign n9073 = ( n1948 & n5702 ) | ( n1948 & n8107 ) | ( n5702 & n8107 ) ;
  assign n9074 = ( n2206 & n4251 ) | ( n2206 & n9073 ) | ( n4251 & n9073 ) ;
  assign n9075 = ( n6859 & n9072 ) | ( n6859 & ~n9074 ) | ( n9072 & ~n9074 ) ;
  assign n9078 = n8920 ^ n8169 ^ n3900 ;
  assign n9076 = n8852 ^ n4853 ^ n3333 ;
  assign n9077 = ( n6154 & n7838 ) | ( n6154 & n9076 ) | ( n7838 & n9076 ) ;
  assign n9079 = n9078 ^ n9077 ^ n5244 ;
  assign n9080 = ( n1748 & n9075 ) | ( n1748 & ~n9079 ) | ( n9075 & ~n9079 ) ;
  assign n9083 = n9082 ^ n9080 ^ n7869 ;
  assign n9084 = n6031 ^ n1853 ^ x51 ;
  assign n9085 = ( n1055 & n7642 ) | ( n1055 & ~n8471 ) | ( n7642 & ~n8471 ) ;
  assign n9086 = n9085 ^ n6038 ^ n523 ;
  assign n9087 = ( ~n451 & n1686 ) | ( ~n451 & n3606 ) | ( n1686 & n3606 ) ;
  assign n9088 = n9087 ^ n6281 ^ n4065 ;
  assign n9089 = n2353 ^ n2106 ^ n207 ;
  assign n9090 = ( n164 & n1348 ) | ( n164 & n9089 ) | ( n1348 & n9089 ) ;
  assign n9091 = n9090 ^ n6237 ^ n1409 ;
  assign n9092 = ( ~n191 & n388 ) | ( ~n191 & n1124 ) | ( n388 & n1124 ) ;
  assign n9093 = n9092 ^ n2309 ^ n2209 ;
  assign n9094 = n9093 ^ n7160 ^ n3557 ;
  assign n9095 = ( n3501 & ~n4914 ) | ( n3501 & n9094 ) | ( ~n4914 & n9094 ) ;
  assign n9096 = n9095 ^ n7253 ^ n3812 ;
  assign n9097 = ( ~n1368 & n6215 ) | ( ~n1368 & n6525 ) | ( n6215 & n6525 ) ;
  assign n9098 = ( n3539 & n7371 ) | ( n3539 & ~n9097 ) | ( n7371 & ~n9097 ) ;
  assign n9099 = n2993 ^ n707 ^ x17 ;
  assign n9100 = n6576 ^ n5969 ^ n4374 ;
  assign n9101 = ( n6972 & ~n9099 ) | ( n6972 & n9100 ) | ( ~n9099 & n9100 ) ;
  assign n9102 = ( n3701 & n7899 ) | ( n3701 & ~n9101 ) | ( n7899 & ~n9101 ) ;
  assign n9103 = n8741 ^ n772 ^ n259 ;
  assign n9104 = ( n2033 & n2487 ) | ( n2033 & ~n9103 ) | ( n2487 & ~n9103 ) ;
  assign n9105 = n9104 ^ n3095 ^ n1919 ;
  assign n9106 = ( n1915 & n9102 ) | ( n1915 & n9105 ) | ( n9102 & n9105 ) ;
  assign n9107 = n5544 ^ n5463 ^ n2311 ;
  assign n9108 = ( ~n216 & n2579 ) | ( ~n216 & n9107 ) | ( n2579 & n9107 ) ;
  assign n9109 = ( ~n7877 & n9106 ) | ( ~n7877 & n9108 ) | ( n9106 & n9108 ) ;
  assign n9110 = ( n2374 & n9098 ) | ( n2374 & ~n9109 ) | ( n9098 & ~n9109 ) ;
  assign n9111 = ( n9091 & ~n9096 ) | ( n9091 & n9110 ) | ( ~n9096 & n9110 ) ;
  assign n9116 = n2927 ^ n1643 ^ n752 ;
  assign n9117 = ( ~n1167 & n3657 ) | ( ~n1167 & n9116 ) | ( n3657 & n9116 ) ;
  assign n9112 = ( n2383 & ~n5639 ) | ( n2383 & n8040 ) | ( ~n5639 & n8040 ) ;
  assign n9113 = n9112 ^ n4492 ^ n752 ;
  assign n9114 = n9113 ^ n7177 ^ n1778 ;
  assign n9115 = n9114 ^ n6143 ^ n1755 ;
  assign n9118 = n9117 ^ n9115 ^ n8274 ;
  assign n9120 = n2354 ^ n2046 ^ n405 ;
  assign n9119 = n6887 ^ n3605 ^ n2897 ;
  assign n9121 = n9120 ^ n9119 ^ n2835 ;
  assign n9122 = n9121 ^ n3609 ^ n2292 ;
  assign n9123 = ( n3773 & ~n6188 ) | ( n3773 & n9122 ) | ( ~n6188 & n9122 ) ;
  assign n9133 = n2427 ^ n1730 ^ n1407 ;
  assign n9134 = ( n450 & n6910 ) | ( n450 & n9133 ) | ( n6910 & n9133 ) ;
  assign n9136 = n4055 ^ n3193 ^ n1400 ;
  assign n9137 = ( n1137 & ~n1303 ) | ( n1137 & n9136 ) | ( ~n1303 & n9136 ) ;
  assign n9135 = ( n2820 & n4706 ) | ( n2820 & n5719 ) | ( n4706 & n5719 ) ;
  assign n9138 = n9137 ^ n9135 ^ n3467 ;
  assign n9139 = ( ~n7953 & n9134 ) | ( ~n7953 & n9138 ) | ( n9134 & n9138 ) ;
  assign n9130 = n5407 ^ n1997 ^ n1189 ;
  assign n9131 = ( n1173 & n4357 ) | ( n1173 & n9130 ) | ( n4357 & n9130 ) ;
  assign n9132 = ( n971 & n7530 ) | ( n971 & n9131 ) | ( n7530 & n9131 ) ;
  assign n9124 = ( n418 & ~n977 ) | ( n418 & n2329 ) | ( ~n977 & n2329 ) ;
  assign n9125 = n9124 ^ n1426 ^ n586 ;
  assign n9126 = ( ~x22 & n4369 ) | ( ~x22 & n9125 ) | ( n4369 & n9125 ) ;
  assign n9127 = n9126 ^ n1229 ^ n1028 ;
  assign n9128 = ( n2409 & n2584 ) | ( n2409 & n9127 ) | ( n2584 & n9127 ) ;
  assign n9129 = n9128 ^ n5729 ^ n2916 ;
  assign n9140 = n9139 ^ n9132 ^ n9129 ;
  assign n9141 = n5684 ^ n2938 ^ n1832 ;
  assign n9142 = n9141 ^ n6341 ^ n339 ;
  assign n9143 = n7070 ^ n5715 ^ n4146 ;
  assign n9144 = ( n787 & ~n1981 ) | ( n787 & n3581 ) | ( ~n1981 & n3581 ) ;
  assign n9145 = ( n307 & n1010 ) | ( n307 & ~n9144 ) | ( n1010 & ~n9144 ) ;
  assign n9146 = ( n2143 & n2665 ) | ( n2143 & n9145 ) | ( n2665 & n9145 ) ;
  assign n9147 = ( ~n7228 & n9143 ) | ( ~n7228 & n9146 ) | ( n9143 & n9146 ) ;
  assign n9148 = ( n1218 & n4322 ) | ( n1218 & n6751 ) | ( n4322 & n6751 ) ;
  assign n9149 = ( n701 & n1432 ) | ( n701 & ~n3206 ) | ( n1432 & ~n3206 ) ;
  assign n9150 = n9149 ^ n4559 ^ n2191 ;
  assign n9151 = n9150 ^ n960 ^ n162 ;
  assign n9152 = ( n6534 & ~n9148 ) | ( n6534 & n9151 ) | ( ~n9148 & n9151 ) ;
  assign n9153 = ( n1125 & n2425 ) | ( n1125 & n3905 ) | ( n2425 & n3905 ) ;
  assign n9154 = ( n1955 & n9152 ) | ( n1955 & n9153 ) | ( n9152 & n9153 ) ;
  assign n9155 = ( n2693 & n6281 ) | ( n2693 & ~n7099 ) | ( n6281 & ~n7099 ) ;
  assign n9156 = n3682 ^ n2008 ^ x5 ;
  assign n9157 = ( ~n5826 & n9155 ) | ( ~n5826 & n9156 ) | ( n9155 & n9156 ) ;
  assign n9158 = n9157 ^ n8347 ^ n5141 ;
  assign n9159 = ( n4537 & ~n4895 ) | ( n4537 & n9158 ) | ( ~n4895 & n9158 ) ;
  assign n9166 = ( n288 & n1414 ) | ( n288 & ~n7840 ) | ( n1414 & ~n7840 ) ;
  assign n9164 = ( n1862 & ~n4686 ) | ( n1862 & n8058 ) | ( ~n4686 & n8058 ) ;
  assign n9165 = ( ~n2182 & n7359 ) | ( ~n2182 & n9164 ) | ( n7359 & n9164 ) ;
  assign n9161 = ( n560 & ~n1821 ) | ( n560 & n2688 ) | ( ~n1821 & n2688 ) ;
  assign n9160 = n6579 ^ n4733 ^ n2247 ;
  assign n9162 = n9161 ^ n9160 ^ n3349 ;
  assign n9163 = ( n1942 & ~n3587 ) | ( n1942 & n9162 ) | ( ~n3587 & n9162 ) ;
  assign n9167 = n9166 ^ n9165 ^ n9163 ;
  assign n9168 = ( ~n3713 & n3943 ) | ( ~n3713 & n6714 ) | ( n3943 & n6714 ) ;
  assign n9169 = n2279 ^ n1783 ^ n1730 ;
  assign n9170 = n9169 ^ n3428 ^ n495 ;
  assign n9171 = ( n573 & ~n9168 ) | ( n573 & n9170 ) | ( ~n9168 & n9170 ) ;
  assign n9196 = ( ~x22 & n2203 ) | ( ~x22 & n6126 ) | ( n2203 & n6126 ) ;
  assign n9190 = ( n595 & n1133 ) | ( n595 & n1570 ) | ( n1133 & n1570 ) ;
  assign n9191 = ( ~n4715 & n8790 ) | ( ~n4715 & n9190 ) | ( n8790 & n9190 ) ;
  assign n9192 = ( x104 & ~n326 ) | ( x104 & n882 ) | ( ~n326 & n882 ) ;
  assign n9193 = ( ~n4572 & n8099 ) | ( ~n4572 & n9192 ) | ( n8099 & n9192 ) ;
  assign n9194 = ( n2516 & n2984 ) | ( n2516 & ~n9193 ) | ( n2984 & ~n9193 ) ;
  assign n9195 = ( n1993 & ~n9191 ) | ( n1993 & n9194 ) | ( ~n9191 & n9194 ) ;
  assign n9185 = n5372 ^ n3247 ^ n2464 ;
  assign n9186 = n9185 ^ n4567 ^ n4470 ;
  assign n9187 = ( n2320 & n4519 ) | ( n2320 & n9186 ) | ( n4519 & n9186 ) ;
  assign n9188 = n9187 ^ n8017 ^ n1759 ;
  assign n9182 = ( n1863 & n4585 ) | ( n1863 & n4848 ) | ( n4585 & n4848 ) ;
  assign n9183 = n9182 ^ n2040 ^ n1915 ;
  assign n9180 = n8865 ^ n3297 ^ n518 ;
  assign n9181 = ( n2623 & n6072 ) | ( n2623 & ~n9180 ) | ( n6072 & ~n9180 ) ;
  assign n9178 = n8931 ^ n6658 ^ x82 ;
  assign n9174 = ( n1629 & n2288 ) | ( n1629 & ~n2536 ) | ( n2288 & ~n2536 ) ;
  assign n9173 = n8011 ^ n3971 ^ n3199 ;
  assign n9175 = n9174 ^ n9173 ^ n6071 ;
  assign n9176 = ( n898 & ~n3360 ) | ( n898 & n9175 ) | ( ~n3360 & n9175 ) ;
  assign n9177 = n9176 ^ n6235 ^ n1328 ;
  assign n9172 = ( n1292 & n4132 ) | ( n1292 & ~n6239 ) | ( n4132 & ~n6239 ) ;
  assign n9179 = n9178 ^ n9177 ^ n9172 ;
  assign n9184 = n9183 ^ n9181 ^ n9179 ;
  assign n9189 = n9188 ^ n9184 ^ n7196 ;
  assign n9197 = n9196 ^ n9195 ^ n9189 ;
  assign n9199 = n3116 ^ n2150 ^ n1147 ;
  assign n9200 = ( n3678 & n4537 ) | ( n3678 & ~n9199 ) | ( n4537 & ~n9199 ) ;
  assign n9201 = n9200 ^ n7760 ^ n6578 ;
  assign n9198 = ( n301 & n1967 ) | ( n301 & ~n3714 ) | ( n1967 & ~n3714 ) ;
  assign n9202 = n9201 ^ n9198 ^ n1495 ;
  assign n9209 = ( ~n381 & n7852 ) | ( ~n381 & n8380 ) | ( n7852 & n8380 ) ;
  assign n9208 = n6498 ^ n6452 ^ n2517 ;
  assign n9203 = ( n530 & n2256 ) | ( n530 & n5885 ) | ( n2256 & n5885 ) ;
  assign n9204 = ( n6554 & n7694 ) | ( n6554 & ~n8516 ) | ( n7694 & ~n8516 ) ;
  assign n9205 = n9204 ^ n5956 ^ n2096 ;
  assign n9206 = ( n2279 & n5152 ) | ( n2279 & ~n9205 ) | ( n5152 & ~n9205 ) ;
  assign n9207 = ( ~n2863 & n9203 ) | ( ~n2863 & n9206 ) | ( n9203 & n9206 ) ;
  assign n9210 = n9209 ^ n9208 ^ n9207 ;
  assign n9213 = ( n1524 & ~n2112 ) | ( n1524 & n7753 ) | ( ~n2112 & n7753 ) ;
  assign n9211 = ( n2178 & n2181 ) | ( n2178 & n5509 ) | ( n2181 & n5509 ) ;
  assign n9212 = ( n2965 & n8712 ) | ( n2965 & ~n9211 ) | ( n8712 & ~n9211 ) ;
  assign n9214 = n9213 ^ n9212 ^ n5824 ;
  assign n9219 = ( ~n1565 & n3738 ) | ( ~n1565 & n5451 ) | ( n3738 & n5451 ) ;
  assign n9218 = n3644 ^ n3438 ^ n2419 ;
  assign n9220 = n9219 ^ n9218 ^ n3033 ;
  assign n9221 = ( ~n3973 & n5639 ) | ( ~n3973 & n8821 ) | ( n5639 & n8821 ) ;
  assign n9222 = ( n1546 & n3990 ) | ( n1546 & ~n9221 ) | ( n3990 & ~n9221 ) ;
  assign n9223 = ( ~n952 & n2757 ) | ( ~n952 & n6770 ) | ( n2757 & n6770 ) ;
  assign n9224 = ( n7988 & n9222 ) | ( n7988 & ~n9223 ) | ( n9222 & ~n9223 ) ;
  assign n9225 = n9224 ^ n6427 ^ x67 ;
  assign n9226 = ( n7538 & n9220 ) | ( n7538 & n9225 ) | ( n9220 & n9225 ) ;
  assign n9215 = ( n391 & n769 ) | ( n391 & n5049 ) | ( n769 & n5049 ) ;
  assign n9216 = ( n2824 & n6953 ) | ( n2824 & n9215 ) | ( n6953 & n9215 ) ;
  assign n9217 = ( n1117 & n4922 ) | ( n1117 & ~n9216 ) | ( n4922 & ~n9216 ) ;
  assign n9227 = n9226 ^ n9217 ^ n1895 ;
  assign n9228 = ( n2154 & n3473 ) | ( n2154 & n9099 ) | ( n3473 & n9099 ) ;
  assign n9229 = n9228 ^ n6319 ^ n494 ;
  assign n9230 = ( n407 & ~n9143 ) | ( n407 & n9229 ) | ( ~n9143 & n9229 ) ;
  assign n9231 = ( n721 & n9227 ) | ( n721 & ~n9230 ) | ( n9227 & ~n9230 ) ;
  assign n9232 = n3645 ^ n2712 ^ n1760 ;
  assign n9233 = n9232 ^ n8330 ^ n2045 ;
  assign n9237 = ( ~n1516 & n1812 ) | ( ~n1516 & n4256 ) | ( n1812 & n4256 ) ;
  assign n9238 = n9237 ^ n4711 ^ n4493 ;
  assign n9239 = n9238 ^ n1595 ^ n186 ;
  assign n9234 = ( n4475 & n4577 ) | ( n4475 & n4944 ) | ( n4577 & n4944 ) ;
  assign n9235 = n9234 ^ n6340 ^ n135 ;
  assign n9236 = n9235 ^ n6816 ^ n1642 ;
  assign n9240 = n9239 ^ n9236 ^ n6894 ;
  assign n9242 = ( ~n757 & n4275 ) | ( ~n757 & n6163 ) | ( n4275 & n6163 ) ;
  assign n9243 = ( n452 & n1530 ) | ( n452 & ~n9242 ) | ( n1530 & ~n9242 ) ;
  assign n9244 = n9243 ^ n4221 ^ n572 ;
  assign n9241 = n8366 ^ n7406 ^ n1841 ;
  assign n9245 = n9244 ^ n9241 ^ n485 ;
  assign n9246 = ( n6055 & n6645 ) | ( n6055 & ~n9245 ) | ( n6645 & ~n9245 ) ;
  assign n9247 = ( n5585 & n5849 ) | ( n5585 & n6806 ) | ( n5849 & n6806 ) ;
  assign n9248 = ( ~n1808 & n1861 ) | ( ~n1808 & n3479 ) | ( n1861 & n3479 ) ;
  assign n9249 = n9248 ^ n4883 ^ n3483 ;
  assign n9250 = n9249 ^ n3419 ^ n1758 ;
  assign n9253 = ( n1066 & ~n6323 ) | ( n1066 & n6486 ) | ( ~n6323 & n6486 ) ;
  assign n9251 = n4005 ^ n810 ^ n255 ;
  assign n9252 = ( n3165 & n6928 ) | ( n3165 & ~n9251 ) | ( n6928 & ~n9251 ) ;
  assign n9254 = n9253 ^ n9252 ^ n7760 ;
  assign n9255 = ( ~n832 & n1480 ) | ( ~n832 & n3970 ) | ( n1480 & n3970 ) ;
  assign n9256 = ( ~n3204 & n6320 ) | ( ~n3204 & n9255 ) | ( n6320 & n9255 ) ;
  assign n9257 = ( n4065 & ~n5946 ) | ( n4065 & n7472 ) | ( ~n5946 & n7472 ) ;
  assign n9258 = ( n471 & n9256 ) | ( n471 & ~n9257 ) | ( n9256 & ~n9257 ) ;
  assign n9259 = n852 ^ n851 ^ x96 ;
  assign n9260 = n9259 ^ n997 ^ n848 ;
  assign n9264 = ( n534 & n3449 ) | ( n534 & n6443 ) | ( n3449 & n6443 ) ;
  assign n9265 = ( n2701 & n3966 ) | ( n2701 & ~n9264 ) | ( n3966 & ~n9264 ) ;
  assign n9266 = ( n6048 & n6101 ) | ( n6048 & ~n9265 ) | ( n6101 & ~n9265 ) ;
  assign n9267 = n1851 ^ n1635 ^ n1412 ;
  assign n9268 = ( x92 & ~n268 ) | ( x92 & n3757 ) | ( ~n268 & n3757 ) ;
  assign n9269 = ( n2076 & n3062 ) | ( n2076 & ~n9268 ) | ( n3062 & ~n9268 ) ;
  assign n9270 = ( n2360 & ~n6944 ) | ( n2360 & n9269 ) | ( ~n6944 & n9269 ) ;
  assign n9271 = ( ~n9266 & n9267 ) | ( ~n9266 & n9270 ) | ( n9267 & n9270 ) ;
  assign n9261 = ( n176 & n4714 ) | ( n176 & n6849 ) | ( n4714 & n6849 ) ;
  assign n9262 = ( n5544 & n8271 ) | ( n5544 & ~n9261 ) | ( n8271 & ~n9261 ) ;
  assign n9263 = ( n1525 & n8617 ) | ( n1525 & n9262 ) | ( n8617 & n9262 ) ;
  assign n9272 = n9271 ^ n9263 ^ n7874 ;
  assign n9273 = ( ~n2203 & n3133 ) | ( ~n2203 & n3427 ) | ( n3133 & n3427 ) ;
  assign n9274 = ( n476 & n2184 ) | ( n476 & ~n9273 ) | ( n2184 & ~n9273 ) ;
  assign n9275 = n9274 ^ n4460 ^ n548 ;
  assign n9276 = ( x6 & ~n459 ) | ( x6 & n9275 ) | ( ~n459 & n9275 ) ;
  assign n9278 = ( n1946 & n4285 ) | ( n1946 & n4821 ) | ( n4285 & n4821 ) ;
  assign n9277 = n8274 ^ n7964 ^ n3836 ;
  assign n9279 = n9278 ^ n9277 ^ n7402 ;
  assign n9280 = ( n787 & ~n6979 ) | ( n787 & n7991 ) | ( ~n6979 & n7991 ) ;
  assign n9281 = n8060 ^ n5445 ^ n5356 ;
  assign n9282 = n9281 ^ n7497 ^ n5781 ;
  assign n9283 = n9282 ^ n3383 ^ n1719 ;
  assign n9284 = ( n5031 & n9280 ) | ( n5031 & ~n9283 ) | ( n9280 & ~n9283 ) ;
  assign n9285 = ( ~n4321 & n4540 ) | ( ~n4321 & n7457 ) | ( n4540 & n7457 ) ;
  assign n9286 = n9285 ^ n8734 ^ n1052 ;
  assign n9287 = ( x48 & n945 ) | ( x48 & ~n2209 ) | ( n945 & ~n2209 ) ;
  assign n9288 = n2410 ^ n1557 ^ n1472 ;
  assign n9289 = ( n3213 & n9287 ) | ( n3213 & ~n9288 ) | ( n9287 & ~n9288 ) ;
  assign n9290 = n9289 ^ n5721 ^ n5119 ;
  assign n9291 = n9169 ^ n2457 ^ n376 ;
  assign n9292 = n5541 ^ n2733 ^ n2581 ;
  assign n9294 = ( ~x41 & n917 ) | ( ~x41 & n4827 ) | ( n917 & n4827 ) ;
  assign n9293 = n6688 ^ n6656 ^ n582 ;
  assign n9295 = n9294 ^ n9293 ^ n3030 ;
  assign n9296 = ( n9291 & ~n9292 ) | ( n9291 & n9295 ) | ( ~n9292 & n9295 ) ;
  assign n9297 = ( n1665 & n3687 ) | ( n1665 & n8556 ) | ( n3687 & n8556 ) ;
  assign n9298 = ( n2073 & ~n7991 ) | ( n2073 & n9297 ) | ( ~n7991 & n9297 ) ;
  assign n9301 = n8713 ^ n3520 ^ n1410 ;
  assign n9302 = ( n529 & n2827 ) | ( n529 & n9301 ) | ( n2827 & n9301 ) ;
  assign n9303 = n9302 ^ n4386 ^ n3735 ;
  assign n9299 = ( ~n257 & n3370 ) | ( ~n257 & n8327 ) | ( n3370 & n8327 ) ;
  assign n9300 = n9299 ^ n8521 ^ n1876 ;
  assign n9304 = n9303 ^ n9300 ^ n5286 ;
  assign n9305 = ( ~n1782 & n9298 ) | ( ~n1782 & n9304 ) | ( n9298 & n9304 ) ;
  assign n9306 = n8994 ^ n5649 ^ n3019 ;
  assign n9307 = ( ~n4834 & n6029 ) | ( ~n4834 & n9306 ) | ( n6029 & n9306 ) ;
  assign n9308 = n9307 ^ n8806 ^ n541 ;
  assign n9309 = ( ~n433 & n8545 ) | ( ~n433 & n9308 ) | ( n8545 & n9308 ) ;
  assign n9310 = ( ~x43 & x44 ) | ( ~x43 & n323 ) | ( x44 & n323 ) ;
  assign n9311 = n9310 ^ n4344 ^ n1927 ;
  assign n9312 = n6574 ^ n5456 ^ n4308 ;
  assign n9313 = n9312 ^ n8562 ^ n2834 ;
  assign n9314 = n3081 ^ n1478 ^ n668 ;
  assign n9315 = ( n3499 & n4407 ) | ( n3499 & n6638 ) | ( n4407 & n6638 ) ;
  assign n9316 = ( x110 & n9314 ) | ( x110 & ~n9315 ) | ( n9314 & ~n9315 ) ;
  assign n9317 = n9316 ^ n3550 ^ n2001 ;
  assign n9319 = ( n656 & n3006 ) | ( n656 & n6814 ) | ( n3006 & n6814 ) ;
  assign n9318 = ( n392 & ~n2751 ) | ( n392 & n8905 ) | ( ~n2751 & n8905 ) ;
  assign n9320 = n9319 ^ n9318 ^ n7490 ;
  assign n9321 = ( ~n1662 & n4585 ) | ( ~n1662 & n5138 ) | ( n4585 & n5138 ) ;
  assign n9322 = ( n3514 & ~n5233 ) | ( n3514 & n9321 ) | ( ~n5233 & n9321 ) ;
  assign n9323 = n9322 ^ n7542 ^ n5420 ;
  assign n9325 = ( n1333 & ~n1884 ) | ( n1333 & n2542 ) | ( ~n1884 & n2542 ) ;
  assign n9324 = ( n2436 & ~n2706 ) | ( n2436 & n3744 ) | ( ~n2706 & n3744 ) ;
  assign n9326 = n9325 ^ n9324 ^ n6963 ;
  assign n9327 = ( n1842 & ~n9323 ) | ( n1842 & n9326 ) | ( ~n9323 & n9326 ) ;
  assign n9329 = n6666 ^ n3962 ^ n3539 ;
  assign n9328 = n8395 ^ n4789 ^ n3798 ;
  assign n9330 = n9329 ^ n9328 ^ n4734 ;
  assign n9331 = n9330 ^ n5668 ^ n4040 ;
  assign n9333 = n6120 ^ n4271 ^ n3674 ;
  assign n9334 = ( n451 & n3385 ) | ( n451 & n9333 ) | ( n3385 & n9333 ) ;
  assign n9335 = n9334 ^ n3433 ^ n2352 ;
  assign n9336 = n9335 ^ n7850 ^ n3325 ;
  assign n9332 = ( ~n3118 & n3209 ) | ( ~n3118 & n3301 ) | ( n3209 & n3301 ) ;
  assign n9337 = n9336 ^ n9332 ^ n8739 ;
  assign n9338 = n4158 ^ n3666 ^ n3566 ;
  assign n9341 = n3202 ^ n2620 ^ n1833 ;
  assign n9340 = n8773 ^ n4546 ^ n3636 ;
  assign n9339 = ( ~n2762 & n3839 ) | ( ~n2762 & n6964 ) | ( n3839 & n6964 ) ;
  assign n9342 = n9341 ^ n9340 ^ n9339 ;
  assign n9348 = ( x66 & n933 ) | ( x66 & n3887 ) | ( n933 & n3887 ) ;
  assign n9347 = n9058 ^ n8356 ^ n4812 ;
  assign n9349 = n9348 ^ n9347 ^ n6458 ;
  assign n9345 = n5863 ^ n5155 ^ n4042 ;
  assign n9343 = ( n2514 & n2557 ) | ( n2514 & ~n4440 ) | ( n2557 & ~n4440 ) ;
  assign n9344 = ( n2161 & n6876 ) | ( n2161 & n9343 ) | ( n6876 & n9343 ) ;
  assign n9346 = n9345 ^ n9344 ^ n3686 ;
  assign n9350 = n9349 ^ n9346 ^ n3600 ;
  assign n9353 = n3928 ^ n2126 ^ n1779 ;
  assign n9351 = ( n1982 & n2273 ) | ( n1982 & n7159 ) | ( n2273 & n7159 ) ;
  assign n9352 = ( ~n4237 & n4679 ) | ( ~n4237 & n9351 ) | ( n4679 & n9351 ) ;
  assign n9354 = n9353 ^ n9352 ^ n1352 ;
  assign n9355 = n9354 ^ n7917 ^ n5438 ;
  assign n9356 = ( n2240 & n3084 ) | ( n2240 & ~n7867 ) | ( n3084 & ~n7867 ) ;
  assign n9357 = ( n4418 & n7588 ) | ( n4418 & n9222 ) | ( n7588 & n9222 ) ;
  assign n9358 = n6660 ^ n4697 ^ n455 ;
  assign n9359 = ( n2502 & ~n9357 ) | ( n2502 & n9358 ) | ( ~n9357 & n9358 ) ;
  assign n9360 = ( n4285 & n6948 ) | ( n4285 & ~n9359 ) | ( n6948 & ~n9359 ) ;
  assign n9361 = ( ~n9355 & n9356 ) | ( ~n9355 & n9360 ) | ( n9356 & n9360 ) ;
  assign n9362 = ( ~n1159 & n1187 ) | ( ~n1159 & n5428 ) | ( n1187 & n5428 ) ;
  assign n9363 = n9362 ^ n6254 ^ n5229 ;
  assign n9370 = ( n3664 & n9058 ) | ( n3664 & n9101 ) | ( n9058 & n9101 ) ;
  assign n9366 = n6618 ^ n2110 ^ n832 ;
  assign n9367 = ( n1196 & n2361 ) | ( n1196 & ~n9366 ) | ( n2361 & ~n9366 ) ;
  assign n9368 = ( n2032 & n4360 ) | ( n2032 & n8115 ) | ( n4360 & n8115 ) ;
  assign n9369 = ( n3730 & ~n9367 ) | ( n3730 & n9368 ) | ( ~n9367 & n9368 ) ;
  assign n9364 = n7511 ^ n5769 ^ n584 ;
  assign n9365 = ( n3634 & n7776 ) | ( n3634 & n9364 ) | ( n7776 & n9364 ) ;
  assign n9371 = n9370 ^ n9369 ^ n9365 ;
  assign n9372 = ( n6369 & n9363 ) | ( n6369 & ~n9371 ) | ( n9363 & ~n9371 ) ;
  assign n9373 = n8411 ^ n1679 ^ n621 ;
  assign n9374 = n9373 ^ n7606 ^ n2623 ;
  assign n9375 = ( n6539 & n9307 ) | ( n6539 & n9374 ) | ( n9307 & n9374 ) ;
  assign n9377 = ( n431 & n1631 ) | ( n431 & n3651 ) | ( n1631 & n3651 ) ;
  assign n9376 = ( n4484 & n4550 ) | ( n4484 & n5184 ) | ( n4550 & n5184 ) ;
  assign n9378 = n9377 ^ n9376 ^ n8539 ;
  assign n9379 = n8595 ^ n3413 ^ n3348 ;
  assign n9380 = n5457 ^ n4479 ^ n3205 ;
  assign n9381 = n9380 ^ n5204 ^ n2810 ;
  assign n9382 = n9381 ^ n4898 ^ n563 ;
  assign n9384 = ( ~n3810 & n5345 ) | ( ~n3810 & n5745 ) | ( n5345 & n5745 ) ;
  assign n9383 = n6132 ^ n3816 ^ n1195 ;
  assign n9385 = n9384 ^ n9383 ^ n3513 ;
  assign n9388 = ( ~n2671 & n3506 ) | ( ~n2671 & n5237 ) | ( n3506 & n5237 ) ;
  assign n9389 = n9388 ^ n7098 ^ n4789 ;
  assign n9386 = n4287 ^ n2455 ^ n2175 ;
  assign n9387 = n9386 ^ n9349 ^ n604 ;
  assign n9390 = n9389 ^ n9387 ^ n640 ;
  assign n9394 = n4764 ^ n2818 ^ n1763 ;
  assign n9391 = n4714 ^ n2866 ^ n442 ;
  assign n9392 = ( n1048 & n3322 ) | ( n1048 & ~n9391 ) | ( n3322 & ~n9391 ) ;
  assign n9393 = n9392 ^ n7999 ^ n5172 ;
  assign n9395 = n9394 ^ n9393 ^ n7934 ;
  assign n9405 = n2626 ^ n1811 ^ n1502 ;
  assign n9406 = ( x63 & n3530 ) | ( x63 & ~n4902 ) | ( n3530 & ~n4902 ) ;
  assign n9407 = ( n1156 & n9405 ) | ( n1156 & ~n9406 ) | ( n9405 & ~n9406 ) ;
  assign n9402 = ( n3724 & n4653 ) | ( n3724 & ~n9125 ) | ( n4653 & ~n9125 ) ;
  assign n9401 = n8516 ^ n3117 ^ n3111 ;
  assign n9399 = n8166 ^ n5411 ^ n139 ;
  assign n9400 = ( n5823 & n6913 ) | ( n5823 & n9399 ) | ( n6913 & n9399 ) ;
  assign n9403 = n9402 ^ n9401 ^ n9400 ;
  assign n9396 = n7964 ^ n5876 ^ n1012 ;
  assign n9397 = n9396 ^ n4442 ^ n1391 ;
  assign n9398 = ( ~n3963 & n6187 ) | ( ~n3963 & n9397 ) | ( n6187 & n9397 ) ;
  assign n9404 = n9403 ^ n9398 ^ n1598 ;
  assign n9408 = n9407 ^ n9404 ^ n7629 ;
  assign n9409 = ( n2357 & n4269 ) | ( n2357 & n9408 ) | ( n4269 & n9408 ) ;
  assign n9410 = n4259 ^ n1502 ^ n1198 ;
  assign n9413 = n7498 ^ n671 ^ n654 ;
  assign n9411 = ( ~n2492 & n2948 ) | ( ~n2492 & n4191 ) | ( n2948 & n4191 ) ;
  assign n9412 = ( n1006 & n2386 ) | ( n1006 & n9411 ) | ( n2386 & n9411 ) ;
  assign n9414 = n9413 ^ n9412 ^ n1790 ;
  assign n9415 = ( ~n3067 & n9410 ) | ( ~n3067 & n9414 ) | ( n9410 & n9414 ) ;
  assign n9416 = ( n1018 & ~n8427 ) | ( n1018 & n9415 ) | ( ~n8427 & n9415 ) ;
  assign n9417 = ( n2072 & n3104 ) | ( n2072 & ~n9416 ) | ( n3104 & ~n9416 ) ;
  assign n9423 = ( ~x79 & n1831 ) | ( ~x79 & n3835 ) | ( n1831 & n3835 ) ;
  assign n9424 = n9423 ^ n9325 ^ n4091 ;
  assign n9425 = n9424 ^ n2381 ^ n908 ;
  assign n9422 = n5798 ^ n5336 ^ n3855 ;
  assign n9418 = n4431 ^ n2688 ^ n1377 ;
  assign n9419 = ( n1880 & ~n2388 ) | ( n1880 & n9418 ) | ( ~n2388 & n9418 ) ;
  assign n9420 = ( ~n6343 & n8129 ) | ( ~n6343 & n9419 ) | ( n8129 & n9419 ) ;
  assign n9421 = ( ~n4984 & n8827 ) | ( ~n4984 & n9420 ) | ( n8827 & n9420 ) ;
  assign n9426 = n9425 ^ n9422 ^ n9421 ;
  assign n9427 = n9426 ^ n3961 ^ n905 ;
  assign n9428 = ( n1951 & ~n4901 ) | ( n1951 & n4949 ) | ( ~n4901 & n4949 ) ;
  assign n9429 = ( n2161 & ~n6218 ) | ( n2161 & n9428 ) | ( ~n6218 & n9428 ) ;
  assign n9430 = n3699 ^ n1051 ^ n434 ;
  assign n9431 = ( ~n9165 & n9370 ) | ( ~n9165 & n9430 ) | ( n9370 & n9430 ) ;
  assign n9432 = n9431 ^ n4921 ^ n890 ;
  assign n9444 = n5180 ^ n1845 ^ n1268 ;
  assign n9445 = n9444 ^ n5070 ^ n4274 ;
  assign n9435 = ( n938 & n5078 ) | ( n938 & ~n5956 ) | ( n5078 & ~n5956 ) ;
  assign n9436 = ( n778 & n1714 ) | ( n778 & ~n4911 ) | ( n1714 & ~n4911 ) ;
  assign n9437 = n9436 ^ n6708 ^ n3299 ;
  assign n9438 = ( n429 & n3157 ) | ( n429 & ~n8759 ) | ( n3157 & ~n8759 ) ;
  assign n9439 = n2607 ^ n1111 ^ n517 ;
  assign n9440 = n9043 ^ n3452 ^ n1496 ;
  assign n9441 = ( ~n494 & n9439 ) | ( ~n494 & n9440 ) | ( n9439 & n9440 ) ;
  assign n9442 = ( ~n397 & n9438 ) | ( ~n397 & n9441 ) | ( n9438 & n9441 ) ;
  assign n9443 = ( ~n9435 & n9437 ) | ( ~n9435 & n9442 ) | ( n9437 & n9442 ) ;
  assign n9433 = ( n1891 & n2006 ) | ( n1891 & n6486 ) | ( n2006 & n6486 ) ;
  assign n9434 = n9433 ^ n7561 ^ n1507 ;
  assign n9446 = n9445 ^ n9443 ^ n9434 ;
  assign n9447 = ( ~n1418 & n6397 ) | ( ~n1418 & n9446 ) | ( n6397 & n9446 ) ;
  assign n9448 = ( n3795 & n9432 ) | ( n3795 & ~n9447 ) | ( n9432 & ~n9447 ) ;
  assign n9449 = n2116 ^ n496 ^ n213 ;
  assign n9450 = ( n1752 & n7805 ) | ( n1752 & ~n9449 ) | ( n7805 & ~n9449 ) ;
  assign n9451 = n3531 ^ n2283 ^ n1049 ;
  assign n9453 = ( ~n6296 & n8694 ) | ( ~n6296 & n8844 ) | ( n8694 & n8844 ) ;
  assign n9452 = n8306 ^ n5311 ^ n4727 ;
  assign n9454 = n9453 ^ n9452 ^ n2171 ;
  assign n9455 = n5448 ^ n3737 ^ n566 ;
  assign n9456 = ( n9451 & n9454 ) | ( n9451 & n9455 ) | ( n9454 & n9455 ) ;
  assign n9457 = ( n1870 & n6129 ) | ( n1870 & n9456 ) | ( n6129 & n9456 ) ;
  assign n9467 = n5058 ^ n3606 ^ n3372 ;
  assign n9458 = n6094 ^ n3966 ^ n1847 ;
  assign n9459 = ( n145 & n1134 ) | ( n145 & n9458 ) | ( n1134 & n9458 ) ;
  assign n9462 = ( n2884 & n6524 ) | ( n2884 & n7790 ) | ( n6524 & n7790 ) ;
  assign n9460 = ( ~n1090 & n1898 ) | ( ~n1090 & n7030 ) | ( n1898 & n7030 ) ;
  assign n9461 = ( n947 & ~n5436 ) | ( n947 & n9460 ) | ( ~n5436 & n9460 ) ;
  assign n9463 = n9462 ^ n9461 ^ n353 ;
  assign n9464 = ( ~n2239 & n9459 ) | ( ~n2239 & n9463 ) | ( n9459 & n9463 ) ;
  assign n9465 = n1816 ^ n876 ^ n614 ;
  assign n9466 = ( ~n6497 & n9464 ) | ( ~n6497 & n9465 ) | ( n9464 & n9465 ) ;
  assign n9468 = n9467 ^ n9466 ^ n6975 ;
  assign n9476 = n2972 ^ n1366 ^ n1156 ;
  assign n9477 = ( ~n1259 & n3736 ) | ( ~n1259 & n9476 ) | ( n3736 & n9476 ) ;
  assign n9478 = n9477 ^ n4034 ^ n2944 ;
  assign n9479 = ( ~n812 & n3814 ) | ( ~n812 & n9478 ) | ( n3814 & n9478 ) ;
  assign n9475 = n8350 ^ n8253 ^ n2319 ;
  assign n9480 = n9479 ^ n9475 ^ n7087 ;
  assign n9471 = n7200 ^ n2887 ^ n2034 ;
  assign n9472 = n4572 ^ n3034 ^ n1395 ;
  assign n9473 = ( n4465 & ~n5483 ) | ( n4465 & n9472 ) | ( ~n5483 & n9472 ) ;
  assign n9474 = ( n3549 & n9471 ) | ( n3549 & n9473 ) | ( n9471 & n9473 ) ;
  assign n9469 = n8665 ^ n6222 ^ n3104 ;
  assign n9470 = ( ~n7890 & n8873 ) | ( ~n7890 & n9469 ) | ( n8873 & n9469 ) ;
  assign n9481 = n9480 ^ n9474 ^ n9470 ;
  assign n9482 = n1090 ^ n854 ^ n640 ;
  assign n9483 = ( ~n4908 & n6568 ) | ( ~n4908 & n9482 ) | ( n6568 & n9482 ) ;
  assign n9484 = n8403 ^ n3126 ^ n2799 ;
  assign n9485 = ( n7829 & n9483 ) | ( n7829 & n9484 ) | ( n9483 & n9484 ) ;
  assign n9486 = n9485 ^ n7949 ^ n1318 ;
  assign n9487 = n9221 ^ n5225 ^ n4293 ;
  assign n9488 = ( ~n2338 & n7165 ) | ( ~n2338 & n9487 ) | ( n7165 & n9487 ) ;
  assign n9489 = n3371 ^ n1426 ^ n988 ;
  assign n9490 = n9489 ^ n3102 ^ n2043 ;
  assign n9491 = ( n345 & n3208 ) | ( n345 & ~n8559 ) | ( n3208 & ~n8559 ) ;
  assign n9492 = n9491 ^ n4641 ^ n2774 ;
  assign n9493 = n9492 ^ n3204 ^ n3008 ;
  assign n9494 = ( x79 & n9490 ) | ( x79 & n9493 ) | ( n9490 & n9493 ) ;
  assign n9495 = ( n450 & n9488 ) | ( n450 & n9494 ) | ( n9488 & n9494 ) ;
  assign n9497 = ( x57 & n1213 ) | ( x57 & n2854 ) | ( n1213 & n2854 ) ;
  assign n9496 = ( n309 & ~n4855 ) | ( n309 & n5440 ) | ( ~n4855 & n5440 ) ;
  assign n9498 = n9497 ^ n9496 ^ n8632 ;
  assign n9502 = ( n522 & n6515 ) | ( n522 & ~n8792 ) | ( n6515 & ~n8792 ) ;
  assign n9501 = n7874 ^ n6421 ^ n2687 ;
  assign n9499 = ( n4703 & n8107 ) | ( n4703 & ~n8789 ) | ( n8107 & ~n8789 ) ;
  assign n9500 = ( ~n209 & n7658 ) | ( ~n209 & n9499 ) | ( n7658 & n9499 ) ;
  assign n9503 = n9502 ^ n9501 ^ n9500 ;
  assign n9504 = ( n1419 & n9498 ) | ( n1419 & n9503 ) | ( n9498 & n9503 ) ;
  assign n9505 = ( n3990 & n6434 ) | ( n3990 & ~n9504 ) | ( n6434 & ~n9504 ) ;
  assign n9506 = ( x14 & n6420 ) | ( x14 & n8180 ) | ( n6420 & n8180 ) ;
  assign n9507 = n9506 ^ n9255 ^ n5454 ;
  assign n9508 = ( n3897 & ~n5015 ) | ( n3897 & n6023 ) | ( ~n5015 & n6023 ) ;
  assign n9509 = ( n2054 & n2742 ) | ( n2054 & ~n3669 ) | ( n2742 & ~n3669 ) ;
  assign n9510 = n9509 ^ n8109 ^ n3185 ;
  assign n9511 = ( n3514 & n5041 ) | ( n3514 & ~n8685 ) | ( n5041 & ~n8685 ) ;
  assign n9512 = ( n9508 & n9510 ) | ( n9508 & ~n9511 ) | ( n9510 & ~n9511 ) ;
  assign n9513 = n9512 ^ n3729 ^ n3485 ;
  assign n9514 = ( n5097 & n9507 ) | ( n5097 & ~n9513 ) | ( n9507 & ~n9513 ) ;
  assign n9515 = ( n6083 & n7189 ) | ( n6083 & n9514 ) | ( n7189 & n9514 ) ;
  assign n9519 = n6802 ^ n2238 ^ n964 ;
  assign n9520 = n6532 ^ n2248 ^ n1108 ;
  assign n9521 = n9520 ^ n1881 ^ n1615 ;
  assign n9522 = ( n2394 & n5721 ) | ( n2394 & n8660 ) | ( n5721 & n8660 ) ;
  assign n9523 = ( n9519 & n9521 ) | ( n9519 & ~n9522 ) | ( n9521 & ~n9522 ) ;
  assign n9516 = ( n1689 & n2689 ) | ( n1689 & ~n2710 ) | ( n2689 & ~n2710 ) ;
  assign n9517 = ( n1148 & n2203 ) | ( n1148 & ~n9516 ) | ( n2203 & ~n9516 ) ;
  assign n9518 = ( n1603 & ~n7335 ) | ( n1603 & n9517 ) | ( ~n7335 & n9517 ) ;
  assign n9524 = n9523 ^ n9518 ^ n5946 ;
  assign n9527 = n9440 ^ n3863 ^ n610 ;
  assign n9525 = n823 ^ x108 ^ x82 ;
  assign n9526 = n9525 ^ n5674 ^ n4495 ;
  assign n9528 = n9527 ^ n9526 ^ n7161 ;
  assign n9529 = ( n5999 & n9524 ) | ( n5999 & ~n9528 ) | ( n9524 & ~n9528 ) ;
  assign n9530 = ( n864 & ~n934 ) | ( n864 & n1881 ) | ( ~n934 & n1881 ) ;
  assign n9531 = ( n6019 & ~n6082 ) | ( n6019 & n7382 ) | ( ~n6082 & n7382 ) ;
  assign n9532 = ( n3630 & ~n4374 ) | ( n3630 & n9531 ) | ( ~n4374 & n9531 ) ;
  assign n9533 = ( n4570 & ~n9530 ) | ( n4570 & n9532 ) | ( ~n9530 & n9532 ) ;
  assign n9534 = ( ~n638 & n5267 ) | ( ~n638 & n8490 ) | ( n5267 & n8490 ) ;
  assign n9535 = ( ~n3971 & n4289 ) | ( ~n3971 & n6870 ) | ( n4289 & n6870 ) ;
  assign n9536 = ( ~n1626 & n1650 ) | ( ~n1626 & n4471 ) | ( n1650 & n4471 ) ;
  assign n9537 = n9536 ^ n5893 ^ n2486 ;
  assign n9538 = n7097 ^ n4660 ^ n3315 ;
  assign n9539 = ( n5509 & n6053 ) | ( n5509 & ~n9538 ) | ( n6053 & ~n9538 ) ;
  assign n9540 = n4420 ^ n3842 ^ n3196 ;
  assign n9541 = ( ~n3518 & n7835 ) | ( ~n3518 & n9540 ) | ( n7835 & n9540 ) ;
  assign n9545 = n2367 ^ n1810 ^ n1473 ;
  assign n9542 = n5922 ^ n3947 ^ n1944 ;
  assign n9543 = n9542 ^ n6326 ^ n1551 ;
  assign n9544 = n9543 ^ n8742 ^ n7239 ;
  assign n9546 = n9545 ^ n9544 ^ n5631 ;
  assign n9547 = ( n9539 & ~n9541 ) | ( n9539 & n9546 ) | ( ~n9541 & n9546 ) ;
  assign n9556 = n8604 ^ n7873 ^ n2221 ;
  assign n9554 = n2607 ^ n1124 ^ n650 ;
  assign n9555 = n9554 ^ n5954 ^ n1118 ;
  assign n9552 = n4059 ^ n2952 ^ n2462 ;
  assign n9548 = n2562 ^ n1702 ^ n859 ;
  assign n9549 = ( ~x52 & n1621 ) | ( ~x52 & n5280 ) | ( n1621 & n5280 ) ;
  assign n9550 = n9549 ^ n7266 ^ n2028 ;
  assign n9551 = ( n8743 & n9548 ) | ( n8743 & n9550 ) | ( n9548 & n9550 ) ;
  assign n9553 = n9552 ^ n9551 ^ n5168 ;
  assign n9557 = n9556 ^ n9555 ^ n9553 ;
  assign n9558 = ( n198 & n2759 ) | ( n198 & n4119 ) | ( n2759 & n4119 ) ;
  assign n9559 = ( n5363 & n8740 ) | ( n5363 & ~n9558 ) | ( n8740 & ~n9558 ) ;
  assign n9560 = ( n8083 & n9557 ) | ( n8083 & ~n9559 ) | ( n9557 & ~n9559 ) ;
  assign n9561 = ( n1605 & n2835 ) | ( n1605 & n3434 ) | ( n2835 & n3434 ) ;
  assign n9562 = ( n1355 & ~n8496 ) | ( n1355 & n9561 ) | ( ~n8496 & n9561 ) ;
  assign n9563 = n4550 ^ n4026 ^ n2413 ;
  assign n9564 = ( n8009 & n9562 ) | ( n8009 & ~n9563 ) | ( n9562 & ~n9563 ) ;
  assign n9565 = n9564 ^ n1486 ^ n797 ;
  assign n9566 = n9565 ^ n7494 ^ n7011 ;
  assign n9570 = ( ~n1203 & n1544 ) | ( ~n1203 & n4091 ) | ( n1544 & n4091 ) ;
  assign n9567 = ( n178 & ~n609 ) | ( n178 & n3947 ) | ( ~n609 & n3947 ) ;
  assign n9568 = n9567 ^ n4293 ^ n3217 ;
  assign n9569 = n9568 ^ n2206 ^ n962 ;
  assign n9571 = n9570 ^ n9569 ^ n655 ;
  assign n9573 = n5356 ^ n3044 ^ n585 ;
  assign n9574 = ( n683 & n2703 ) | ( n683 & n9573 ) | ( n2703 & n9573 ) ;
  assign n9572 = n9469 ^ n8997 ^ n6823 ;
  assign n9575 = n9574 ^ n9572 ^ n413 ;
  assign n9576 = n9575 ^ n4891 ^ n2924 ;
  assign n9577 = n9576 ^ n5487 ^ n2253 ;
  assign n9578 = ( ~n3156 & n5434 ) | ( ~n3156 & n7530 ) | ( n5434 & n7530 ) ;
  assign n9579 = n9578 ^ n5897 ^ n4369 ;
  assign n9580 = n9579 ^ n3785 ^ n3726 ;
  assign n9582 = ( n909 & n1491 ) | ( n909 & n1959 ) | ( n1491 & n1959 ) ;
  assign n9583 = n9582 ^ n7704 ^ n3923 ;
  assign n9581 = ( n4499 & ~n6881 ) | ( n4499 & n9039 ) | ( ~n6881 & n9039 ) ;
  assign n9584 = n9583 ^ n9581 ^ n8780 ;
  assign n9585 = n9584 ^ n3866 ^ n370 ;
  assign n9589 = ( n1576 & n1635 ) | ( n1576 & n4293 ) | ( n1635 & n4293 ) ;
  assign n9587 = ( n2558 & n2995 ) | ( n2558 & ~n6202 ) | ( n2995 & ~n6202 ) ;
  assign n9586 = n8943 ^ n8316 ^ n2315 ;
  assign n9588 = n9587 ^ n9586 ^ n4297 ;
  assign n9590 = n9589 ^ n9588 ^ n1094 ;
  assign n9591 = ( n2733 & n6260 ) | ( n2733 & ~n8005 ) | ( n6260 & ~n8005 ) ;
  assign n9599 = n2687 ^ n2512 ^ n2223 ;
  assign n9600 = ( n2724 & n4548 ) | ( n2724 & n9599 ) | ( n4548 & n9599 ) ;
  assign n9598 = ( n6470 & n7945 ) | ( n6470 & ~n8586 ) | ( n7945 & ~n8586 ) ;
  assign n9601 = n9600 ^ n9598 ^ n3978 ;
  assign n9592 = ( n403 & n3421 ) | ( n403 & ~n6350 ) | ( n3421 & ~n6350 ) ;
  assign n9593 = ( n4446 & ~n4766 ) | ( n4446 & n6012 ) | ( ~n4766 & n6012 ) ;
  assign n9594 = ( ~n1191 & n4789 ) | ( ~n1191 & n6175 ) | ( n4789 & n6175 ) ;
  assign n9595 = n9594 ^ n5939 ^ n1914 ;
  assign n9596 = ( n9592 & ~n9593 ) | ( n9592 & n9595 ) | ( ~n9593 & n9595 ) ;
  assign n9597 = ( ~n3087 & n3603 ) | ( ~n3087 & n9596 ) | ( n3603 & n9596 ) ;
  assign n9602 = n9601 ^ n9597 ^ n6146 ;
  assign n9603 = ( n1430 & n9591 ) | ( n1430 & n9602 ) | ( n9591 & n9602 ) ;
  assign n9604 = n4218 ^ n4158 ^ n3106 ;
  assign n9605 = n4908 ^ n1680 ^ n452 ;
  assign n9606 = n9605 ^ n7705 ^ n1818 ;
  assign n9607 = n6524 ^ n2734 ^ n1143 ;
  assign n9608 = ( n7390 & n9606 ) | ( n7390 & n9607 ) | ( n9606 & n9607 ) ;
  assign n9609 = ( n3908 & n4658 ) | ( n3908 & ~n8620 ) | ( n4658 & ~n8620 ) ;
  assign n9610 = ( n3421 & ~n5691 ) | ( n3421 & n7734 ) | ( ~n5691 & n7734 ) ;
  assign n9611 = n9610 ^ n7207 ^ n4149 ;
  assign n9612 = n9611 ^ n3894 ^ n1600 ;
  assign n9613 = ( n1353 & n4790 ) | ( n1353 & n9612 ) | ( n4790 & n9612 ) ;
  assign n9614 = ( ~n4146 & n4516 ) | ( ~n4146 & n7458 ) | ( n4516 & n7458 ) ;
  assign n9615 = n9477 ^ n8143 ^ n6102 ;
  assign n9616 = ( ~n1152 & n4137 ) | ( ~n1152 & n9615 ) | ( n4137 & n9615 ) ;
  assign n9621 = ( n1000 & n1506 ) | ( n1000 & ~n5135 ) | ( n1506 & ~n5135 ) ;
  assign n9622 = ( x115 & ~n933 ) | ( x115 & n1354 ) | ( ~n933 & n1354 ) ;
  assign n9623 = ( n1007 & ~n9621 ) | ( n1007 & n9622 ) | ( ~n9621 & n9622 ) ;
  assign n9619 = n7019 ^ n1869 ^ n232 ;
  assign n9620 = ( ~n1447 & n8383 ) | ( ~n1447 & n9619 ) | ( n8383 & n9619 ) ;
  assign n9617 = ( ~n3056 & n3430 ) | ( ~n3056 & n8479 ) | ( n3430 & n8479 ) ;
  assign n9618 = n9617 ^ n4136 ^ n1007 ;
  assign n9624 = n9623 ^ n9620 ^ n9618 ;
  assign n9625 = n9624 ^ n9289 ^ n5340 ;
  assign n9630 = ( n2354 & n3036 ) | ( n2354 & n7406 ) | ( n3036 & n7406 ) ;
  assign n9629 = ( n867 & n2363 ) | ( n867 & ~n3291 ) | ( n2363 & ~n3291 ) ;
  assign n9626 = ( n2999 & n3559 ) | ( n2999 & ~n5356 ) | ( n3559 & ~n5356 ) ;
  assign n9627 = n8496 ^ n3644 ^ n234 ;
  assign n9628 = ( n1022 & ~n9626 ) | ( n1022 & n9627 ) | ( ~n9626 & n9627 ) ;
  assign n9631 = n9630 ^ n9629 ^ n9628 ;
  assign n9632 = ( ~n1619 & n3906 ) | ( ~n1619 & n9631 ) | ( n3906 & n9631 ) ;
  assign n9633 = n3973 ^ n3515 ^ n1127 ;
  assign n9634 = ( n1571 & ~n5549 ) | ( n1571 & n9633 ) | ( ~n5549 & n9633 ) ;
  assign n9635 = ( ~n1820 & n7647 ) | ( ~n1820 & n9634 ) | ( n7647 & n9634 ) ;
  assign n9640 = ( n1686 & ~n5407 ) | ( n1686 & n9633 ) | ( ~n5407 & n9633 ) ;
  assign n9636 = ( n1855 & n1904 ) | ( n1855 & n7788 ) | ( n1904 & n7788 ) ;
  assign n9637 = n4721 ^ n4172 ^ n3068 ;
  assign n9638 = ( n9462 & n9636 ) | ( n9462 & n9637 ) | ( n9636 & n9637 ) ;
  assign n9639 = n9638 ^ n8108 ^ n5838 ;
  assign n9641 = n9640 ^ n9639 ^ n2809 ;
  assign n9645 = ( n4396 & ~n4689 ) | ( n4396 & n7703 ) | ( ~n4689 & n7703 ) ;
  assign n9646 = ( ~n3667 & n4708 ) | ( ~n3667 & n9645 ) | ( n4708 & n9645 ) ;
  assign n9642 = n4432 ^ n1668 ^ n1587 ;
  assign n9643 = ( n6189 & n6955 ) | ( n6189 & ~n9642 ) | ( n6955 & ~n9642 ) ;
  assign n9644 = ( n3141 & n8856 ) | ( n3141 & n9643 ) | ( n8856 & n9643 ) ;
  assign n9647 = n9646 ^ n9644 ^ n7190 ;
  assign n9648 = ( n1034 & ~n5892 ) | ( n1034 & n9647 ) | ( ~n5892 & n9647 ) ;
  assign n9652 = ( n1343 & ~n2054 ) | ( n1343 & n5446 ) | ( ~n2054 & n5446 ) ;
  assign n9650 = n7850 ^ n6959 ^ n6461 ;
  assign n9649 = ( ~n5382 & n8247 ) | ( ~n5382 & n9507 ) | ( n8247 & n9507 ) ;
  assign n9651 = n9650 ^ n9649 ^ n2679 ;
  assign n9653 = n9652 ^ n9651 ^ n9033 ;
  assign n9654 = n4035 ^ n2772 ^ n1088 ;
  assign n9655 = ( n3672 & n4543 ) | ( n3672 & n9212 ) | ( n4543 & n9212 ) ;
  assign n9656 = ( n2011 & n9654 ) | ( n2011 & n9655 ) | ( n9654 & n9655 ) ;
  assign n9657 = ( n1904 & n8593 ) | ( n1904 & n9656 ) | ( n8593 & n9656 ) ;
  assign n9658 = n4858 ^ n1593 ^ n1252 ;
  assign n9659 = ( n304 & n895 ) | ( n304 & ~n8298 ) | ( n895 & ~n8298 ) ;
  assign n9660 = ( n5773 & n9658 ) | ( n5773 & ~n9659 ) | ( n9658 & ~n9659 ) ;
  assign n9661 = n9660 ^ n4241 ^ n1258 ;
  assign n9662 = n5726 ^ n4583 ^ n2421 ;
  assign n9663 = ( n3923 & n8302 ) | ( n3923 & ~n9662 ) | ( n8302 & ~n9662 ) ;
  assign n9664 = n9662 ^ n7345 ^ n3753 ;
  assign n9665 = ( x106 & n1396 ) | ( x106 & n2946 ) | ( n1396 & n2946 ) ;
  assign n9666 = ( n2259 & n2404 ) | ( n2259 & n4055 ) | ( n2404 & n4055 ) ;
  assign n9667 = n9666 ^ n5048 ^ n4278 ;
  assign n9668 = n9667 ^ n6160 ^ n3345 ;
  assign n9669 = n9668 ^ n7794 ^ n1713 ;
  assign n9670 = ( ~n816 & n9665 ) | ( ~n816 & n9669 ) | ( n9665 & n9669 ) ;
  assign n9671 = n9670 ^ n4993 ^ n4708 ;
  assign n9672 = ( ~n5053 & n5600 ) | ( ~n5053 & n8871 ) | ( n5600 & n8871 ) ;
  assign n9676 = n6042 ^ n2204 ^ n269 ;
  assign n9677 = n9676 ^ n7704 ^ n1694 ;
  assign n9678 = ( n2181 & n4192 ) | ( n2181 & ~n6736 ) | ( n4192 & ~n6736 ) ;
  assign n9679 = n9678 ^ n9136 ^ n5581 ;
  assign n9680 = ( n1177 & n2793 ) | ( n1177 & n9679 ) | ( n2793 & n9679 ) ;
  assign n9681 = ( n5639 & n9677 ) | ( n5639 & ~n9680 ) | ( n9677 & ~n9680 ) ;
  assign n9673 = ( ~n142 & n2075 ) | ( ~n142 & n2718 ) | ( n2075 & n2718 ) ;
  assign n9674 = ( n620 & n5283 ) | ( n620 & ~n9673 ) | ( n5283 & ~n9673 ) ;
  assign n9675 = ( n3167 & n4596 ) | ( n3167 & n9674 ) | ( n4596 & n9674 ) ;
  assign n9682 = n9681 ^ n9675 ^ n1273 ;
  assign n9683 = n2762 ^ n1685 ^ n644 ;
  assign n9684 = n9683 ^ n3286 ^ n875 ;
  assign n9685 = ( n2237 & ~n4636 ) | ( n2237 & n6005 ) | ( ~n4636 & n6005 ) ;
  assign n9686 = ( n1648 & n5655 ) | ( n1648 & n9677 ) | ( n5655 & n9677 ) ;
  assign n9687 = ( x78 & n394 ) | ( x78 & n2346 ) | ( n394 & n2346 ) ;
  assign n9688 = n9687 ^ n1572 ^ n627 ;
  assign n9689 = ( n854 & ~n2075 ) | ( n854 & n5416 ) | ( ~n2075 & n5416 ) ;
  assign n9690 = ( n2329 & ~n9688 ) | ( n2329 & n9689 ) | ( ~n9688 & n9689 ) ;
  assign n9691 = ( n5084 & ~n9686 ) | ( n5084 & n9690 ) | ( ~n9686 & n9690 ) ;
  assign n9692 = ( ~n9684 & n9685 ) | ( ~n9684 & n9691 ) | ( n9685 & n9691 ) ;
  assign n9693 = ( ~n2191 & n4804 ) | ( ~n2191 & n9692 ) | ( n4804 & n9692 ) ;
  assign n9694 = ( ~n5380 & n6241 ) | ( ~n5380 & n9693 ) | ( n6241 & n9693 ) ;
  assign n9695 = n3248 ^ n3025 ^ n2133 ;
  assign n9696 = ( n2661 & n4235 ) | ( n2661 & ~n6085 ) | ( n4235 & ~n6085 ) ;
  assign n9697 = ( n2568 & n9261 ) | ( n2568 & n9696 ) | ( n9261 & n9696 ) ;
  assign n9701 = ( n5218 & ~n5340 ) | ( n5218 & n6904 ) | ( ~n5340 & n6904 ) ;
  assign n9698 = n4439 ^ n479 ^ x72 ;
  assign n9699 = n4881 ^ n3001 ^ n1298 ;
  assign n9700 = ( n4019 & n9698 ) | ( n4019 & n9699 ) | ( n9698 & n9699 ) ;
  assign n9702 = n9701 ^ n9700 ^ n1633 ;
  assign n9703 = n9702 ^ n5763 ^ n4597 ;
  assign n9704 = n3282 ^ n1342 ^ n173 ;
  assign n9705 = ( ~n5138 & n6158 ) | ( ~n5138 & n9704 ) | ( n6158 & n9704 ) ;
  assign n9706 = ( n4251 & ~n5122 ) | ( n4251 & n9650 ) | ( ~n5122 & n9650 ) ;
  assign n9707 = n8412 ^ n6892 ^ n5757 ;
  assign n9708 = n9707 ^ n7158 ^ n3534 ;
  assign n9709 = ( n217 & n3213 ) | ( n217 & ~n8170 ) | ( n3213 & ~n8170 ) ;
  assign n9716 = ( n819 & n2809 ) | ( n819 & n4438 ) | ( n2809 & n4438 ) ;
  assign n9717 = n9716 ^ n5928 ^ n754 ;
  assign n9710 = ( x76 & n1236 ) | ( x76 & ~n4660 ) | ( n1236 & ~n4660 ) ;
  assign n9711 = ( ~n880 & n3094 ) | ( ~n880 & n6660 ) | ( n3094 & n6660 ) ;
  assign n9712 = ( n3725 & n4660 ) | ( n3725 & ~n9711 ) | ( n4660 & ~n9711 ) ;
  assign n9713 = ( n2247 & ~n9710 ) | ( n2247 & n9712 ) | ( ~n9710 & n9712 ) ;
  assign n9714 = n9713 ^ n2952 ^ n1914 ;
  assign n9715 = n9714 ^ n5601 ^ n4513 ;
  assign n9718 = n9717 ^ n9715 ^ n7173 ;
  assign n9719 = ( ~n1377 & n9709 ) | ( ~n1377 & n9718 ) | ( n9709 & n9718 ) ;
  assign n9720 = ( ~n3624 & n3732 ) | ( ~n3624 & n4525 ) | ( n3732 & n4525 ) ;
  assign n9721 = n9720 ^ n8358 ^ n7412 ;
  assign n9722 = ( n2633 & n3334 ) | ( n2633 & ~n5155 ) | ( n3334 & ~n5155 ) ;
  assign n9723 = ( ~n692 & n4055 ) | ( ~n692 & n4842 ) | ( n4055 & n4842 ) ;
  assign n9724 = ( n4064 & ~n8879 ) | ( n4064 & n9723 ) | ( ~n8879 & n9723 ) ;
  assign n9725 = n7296 ^ n1029 ^ n650 ;
  assign n9726 = ( n379 & n5510 ) | ( n379 & ~n9725 ) | ( n5510 & ~n9725 ) ;
  assign n9727 = ( n563 & n2154 ) | ( n563 & n5367 ) | ( n2154 & n5367 ) ;
  assign n9728 = n2870 ^ n1292 ^ n508 ;
  assign n9729 = ( n350 & n9727 ) | ( n350 & ~n9728 ) | ( n9727 & ~n9728 ) ;
  assign n9730 = ( n2299 & n7955 ) | ( n2299 & n9729 ) | ( n7955 & n9729 ) ;
  assign n9731 = ( n9724 & n9726 ) | ( n9724 & ~n9730 ) | ( n9726 & ~n9730 ) ;
  assign n9732 = n9731 ^ n7646 ^ n256 ;
  assign n9735 = ( ~n679 & n1073 ) | ( ~n679 & n3859 ) | ( n1073 & n3859 ) ;
  assign n9733 = ( n2270 & ~n3698 ) | ( n2270 & n8758 ) | ( ~n3698 & n8758 ) ;
  assign n9734 = n9733 ^ n8050 ^ n2465 ;
  assign n9736 = n9735 ^ n9734 ^ n1944 ;
  assign n9740 = n3326 ^ n3128 ^ n193 ;
  assign n9741 = ( n3047 & ~n3170 ) | ( n3047 & n9740 ) | ( ~n3170 & n9740 ) ;
  assign n9742 = n9741 ^ n8464 ^ n2354 ;
  assign n9737 = n4429 ^ n1349 ^ n1192 ;
  assign n9738 = n9737 ^ n2917 ^ n1839 ;
  assign n9739 = ( n708 & n2533 ) | ( n708 & ~n9738 ) | ( n2533 & ~n9738 ) ;
  assign n9743 = n9742 ^ n9739 ^ n6987 ;
  assign n9744 = ( ~n1147 & n2390 ) | ( ~n1147 & n6333 ) | ( n2390 & n6333 ) ;
  assign n9745 = ( ~n4705 & n7294 ) | ( ~n4705 & n9744 ) | ( n7294 & n9744 ) ;
  assign n9747 = ( n1780 & n4090 ) | ( n1780 & ~n5121 ) | ( n4090 & ~n5121 ) ;
  assign n9746 = ( n362 & ~n5725 ) | ( n362 & n7753 ) | ( ~n5725 & n7753 ) ;
  assign n9748 = n9747 ^ n9746 ^ n1277 ;
  assign n9749 = ( ~n2012 & n9745 ) | ( ~n2012 & n9748 ) | ( n9745 & n9748 ) ;
  assign n9750 = ( n1193 & ~n1363 ) | ( n1193 & n5434 ) | ( ~n1363 & n5434 ) ;
  assign n9751 = n9750 ^ n5811 ^ n440 ;
  assign n9752 = n9751 ^ n7901 ^ n3321 ;
  assign n9753 = n9752 ^ n3515 ^ n362 ;
  assign n9758 = n6898 ^ n3592 ^ n753 ;
  assign n9756 = ( n4717 & ~n6315 ) | ( n4717 & n9242 ) | ( ~n6315 & n9242 ) ;
  assign n9754 = n6952 ^ n2687 ^ n1646 ;
  assign n9755 = n9754 ^ n3323 ^ x33 ;
  assign n9757 = n9756 ^ n9755 ^ n7395 ;
  assign n9759 = n9758 ^ n9757 ^ n2525 ;
  assign n9760 = ( n494 & n2736 ) | ( n494 & n8854 ) | ( n2736 & n8854 ) ;
  assign n9761 = ( ~n418 & n951 ) | ( ~n418 & n4411 ) | ( n951 & n4411 ) ;
  assign n9762 = n9761 ^ n2665 ^ n1871 ;
  assign n9763 = n9762 ^ n3798 ^ n1693 ;
  assign n9764 = n3699 ^ n3512 ^ n1998 ;
  assign n9765 = n9764 ^ n5983 ^ n240 ;
  assign n9766 = n6443 ^ n5577 ^ n608 ;
  assign n9767 = ( n6077 & ~n9765 ) | ( n6077 & n9766 ) | ( ~n9765 & n9766 ) ;
  assign n9768 = n3663 ^ n3629 ^ n419 ;
  assign n9769 = ( ~n6615 & n8058 ) | ( ~n6615 & n9768 ) | ( n8058 & n9768 ) ;
  assign n9772 = n4445 ^ n2414 ^ x105 ;
  assign n9771 = ( ~n2106 & n4879 ) | ( ~n2106 & n5179 ) | ( n4879 & n5179 ) ;
  assign n9773 = n9772 ^ n9771 ^ n2026 ;
  assign n9777 = n8918 ^ n4274 ^ n2307 ;
  assign n9778 = ( ~n1878 & n6765 ) | ( ~n1878 & n9777 ) | ( n6765 & n9777 ) ;
  assign n9779 = ( ~n1223 & n1739 ) | ( ~n1223 & n9778 ) | ( n1739 & n9778 ) ;
  assign n9780 = n9779 ^ n8662 ^ n411 ;
  assign n9774 = n6219 ^ n3213 ^ n1650 ;
  assign n9775 = n9774 ^ n7745 ^ n920 ;
  assign n9776 = ( n2600 & n4085 ) | ( n2600 & n9775 ) | ( n4085 & n9775 ) ;
  assign n9781 = n9780 ^ n9776 ^ n8325 ;
  assign n9782 = ( ~n5705 & n9773 ) | ( ~n5705 & n9781 ) | ( n9773 & n9781 ) ;
  assign n9783 = ( ~n5518 & n6460 ) | ( ~n5518 & n9782 ) | ( n6460 & n9782 ) ;
  assign n9770 = n9742 ^ n8047 ^ n4770 ;
  assign n9784 = n9783 ^ n9770 ^ n7899 ;
  assign n9785 = ( n3469 & n8483 ) | ( n3469 & ~n8725 ) | ( n8483 & ~n8725 ) ;
  assign n9790 = ( n1033 & n1218 ) | ( n1033 & ~n4214 ) | ( n1218 & ~n4214 ) ;
  assign n9791 = n9790 ^ n4608 ^ n3247 ;
  assign n9789 = n4010 ^ n3765 ^ n790 ;
  assign n9792 = n9791 ^ n9789 ^ n4485 ;
  assign n9794 = ( n472 & ~n849 ) | ( n472 & n946 ) | ( ~n849 & n946 ) ;
  assign n9793 = n5482 ^ n1902 ^ n491 ;
  assign n9795 = n9794 ^ n9793 ^ n626 ;
  assign n9796 = ( n2013 & n7933 ) | ( n2013 & n9795 ) | ( n7933 & n9795 ) ;
  assign n9797 = ( n4950 & ~n9792 ) | ( n4950 & n9796 ) | ( ~n9792 & n9796 ) ;
  assign n9786 = ( n608 & n7685 ) | ( n608 & n8769 ) | ( n7685 & n8769 ) ;
  assign n9787 = ( ~n6562 & n7940 ) | ( ~n6562 & n9786 ) | ( n7940 & n9786 ) ;
  assign n9788 = ( n882 & ~n5329 ) | ( n882 & n9787 ) | ( ~n5329 & n9787 ) ;
  assign n9798 = n9797 ^ n9788 ^ n3779 ;
  assign n9799 = ( n1878 & n9785 ) | ( n1878 & n9798 ) | ( n9785 & n9798 ) ;
  assign n9806 = n2356 ^ n729 ^ n308 ;
  assign n9802 = ( n1562 & n2707 ) | ( n1562 & n5402 ) | ( n2707 & n5402 ) ;
  assign n9803 = ( ~n1031 & n6702 ) | ( ~n1031 & n9802 ) | ( n6702 & n9802 ) ;
  assign n9804 = n9803 ^ n7901 ^ n2074 ;
  assign n9805 = ( n2431 & n7181 ) | ( n2431 & ~n9804 ) | ( n7181 & ~n9804 ) ;
  assign n9807 = n9806 ^ n9805 ^ n1133 ;
  assign n9800 = n5720 ^ n2519 ^ n2195 ;
  assign n9801 = n9800 ^ n2177 ^ n882 ;
  assign n9808 = n9807 ^ n9801 ^ n6337 ;
  assign n9809 = ( n258 & n4740 ) | ( n258 & n9808 ) | ( n4740 & n9808 ) ;
  assign n9810 = ( x80 & n2458 ) | ( x80 & n3331 ) | ( n2458 & n3331 ) ;
  assign n9811 = ( ~n3120 & n8163 ) | ( ~n3120 & n9810 ) | ( n8163 & n9810 ) ;
  assign n9812 = ( n3344 & ~n5668 ) | ( n3344 & n9811 ) | ( ~n5668 & n9811 ) ;
  assign n9813 = n9399 ^ n6507 ^ n895 ;
  assign n9814 = ( n630 & n4922 ) | ( n630 & ~n9813 ) | ( n4922 & ~n9813 ) ;
  assign n9815 = ( n2139 & ~n7016 ) | ( n2139 & n8791 ) | ( ~n7016 & n8791 ) ;
  assign n9816 = ( ~x33 & n1684 ) | ( ~x33 & n2880 ) | ( n1684 & n2880 ) ;
  assign n9817 = ( n5178 & ~n9815 ) | ( n5178 & n9816 ) | ( ~n9815 & n9816 ) ;
  assign n9818 = n5683 ^ n4816 ^ n736 ;
  assign n9819 = n9187 ^ n7988 ^ n4536 ;
  assign n9820 = ( n2550 & n9818 ) | ( n2550 & ~n9819 ) | ( n9818 & ~n9819 ) ;
  assign n9821 = ( n5940 & n8091 ) | ( n5940 & ~n9820 ) | ( n8091 & ~n9820 ) ;
  assign n9822 = n5858 ^ n4872 ^ n1030 ;
  assign n9823 = ( n233 & n6609 ) | ( n233 & ~n8583 ) | ( n6609 & ~n8583 ) ;
  assign n9824 = ( n749 & ~n5723 ) | ( n749 & n6443 ) | ( ~n5723 & n6443 ) ;
  assign n9825 = n9824 ^ n9079 ^ n5926 ;
  assign n9826 = n2076 ^ n1563 ^ n281 ;
  assign n9828 = n1095 ^ n967 ^ n782 ;
  assign n9827 = ( n1978 & ~n7874 ) | ( n1978 & n8036 ) | ( ~n7874 & n8036 ) ;
  assign n9829 = n9828 ^ n9827 ^ n1513 ;
  assign n9830 = ( n5575 & n9060 ) | ( n5575 & n9829 ) | ( n9060 & n9829 ) ;
  assign n9831 = ( n6039 & n9826 ) | ( n6039 & ~n9830 ) | ( n9826 & ~n9830 ) ;
  assign n9832 = ( n4300 & ~n8370 ) | ( n4300 & n9831 ) | ( ~n8370 & n9831 ) ;
  assign n9833 = ( x29 & n8003 ) | ( x29 & n8548 ) | ( n8003 & n8548 ) ;
  assign n9834 = ( n4962 & ~n5701 ) | ( n4962 & n9833 ) | ( ~n5701 & n9833 ) ;
  assign n9835 = ( n1578 & n1725 ) | ( n1578 & n9834 ) | ( n1725 & n9834 ) ;
  assign n9836 = ( ~n1046 & n2413 ) | ( ~n1046 & n2720 ) | ( n2413 & n2720 ) ;
  assign n9837 = ( n3547 & ~n8227 ) | ( n3547 & n9836 ) | ( ~n8227 & n9836 ) ;
  assign n9838 = n4397 ^ n1588 ^ x104 ;
  assign n9839 = n2867 ^ n1010 ^ n412 ;
  assign n9840 = ( n241 & ~n9838 ) | ( n241 & n9839 ) | ( ~n9838 & n9839 ) ;
  assign n9841 = n9840 ^ n5054 ^ n3618 ;
  assign n9842 = ( n1514 & n7025 ) | ( n1514 & n9841 ) | ( n7025 & n9841 ) ;
  assign n9843 = n6674 ^ n3723 ^ n1355 ;
  assign n9844 = n9843 ^ n4613 ^ n508 ;
  assign n9845 = n7689 ^ n7084 ^ n639 ;
  assign n9846 = n5836 ^ n1116 ^ n289 ;
  assign n9847 = ( n3735 & n5897 ) | ( n3735 & n9846 ) | ( n5897 & n9846 ) ;
  assign n9848 = n9847 ^ n7554 ^ n4267 ;
  assign n9858 = ( n635 & ~n1167 ) | ( n635 & n6594 ) | ( ~n1167 & n6594 ) ;
  assign n9857 = n9741 ^ n6989 ^ n2139 ;
  assign n9853 = n3918 ^ n3315 ^ n2156 ;
  assign n9854 = n9853 ^ n1423 ^ n1300 ;
  assign n9851 = ( n597 & n1152 ) | ( n597 & ~n5608 ) | ( n1152 & ~n5608 ) ;
  assign n9852 = n9851 ^ n9397 ^ n7229 ;
  assign n9855 = n9854 ^ n9852 ^ n2235 ;
  assign n9849 = ( x107 & n3608 ) | ( x107 & ~n3978 ) | ( n3608 & ~n3978 ) ;
  assign n9850 = ( n6507 & n9224 ) | ( n6507 & ~n9849 ) | ( n9224 & ~n9849 ) ;
  assign n9856 = n9855 ^ n9850 ^ n3039 ;
  assign n9859 = n9858 ^ n9857 ^ n9856 ;
  assign n9861 = ( n313 & n1798 ) | ( n313 & ~n6685 ) | ( n1798 & ~n6685 ) ;
  assign n9862 = n9861 ^ n6317 ^ n4331 ;
  assign n9863 = n9862 ^ n3802 ^ n2403 ;
  assign n9860 = ( n297 & n5731 ) | ( n297 & n7426 ) | ( n5731 & n7426 ) ;
  assign n9864 = n9863 ^ n9860 ^ n5806 ;
  assign n9865 = n8806 ^ n4881 ^ n1014 ;
  assign n9866 = n9865 ^ n5762 ^ n1695 ;
  assign n9867 = n8666 ^ n8555 ^ n5586 ;
  assign n9868 = n9867 ^ n6925 ^ n2986 ;
  assign n9869 = ( ~n227 & n2257 ) | ( ~n227 & n4704 ) | ( n2257 & n4704 ) ;
  assign n9870 = ( n7511 & n9868 ) | ( n7511 & n9869 ) | ( n9868 & n9869 ) ;
  assign n9871 = ( n545 & n1471 ) | ( n545 & ~n3830 ) | ( n1471 & ~n3830 ) ;
  assign n9872 = n6302 ^ n3865 ^ n1803 ;
  assign n9873 = ( n4933 & ~n5028 ) | ( n4933 & n9872 ) | ( ~n5028 & n9872 ) ;
  assign n9874 = ( n4596 & n9871 ) | ( n4596 & ~n9873 ) | ( n9871 & ~n9873 ) ;
  assign n9876 = n5953 ^ n2688 ^ n2159 ;
  assign n9877 = ( n1894 & n5351 ) | ( n1894 & ~n9876 ) | ( n5351 & ~n9876 ) ;
  assign n9875 = ( n3354 & n3871 ) | ( n3354 & n8906 ) | ( n3871 & n8906 ) ;
  assign n9878 = n9877 ^ n9875 ^ n990 ;
  assign n9881 = ( n1401 & n2504 ) | ( n1401 & n8410 ) | ( n2504 & n8410 ) ;
  assign n9882 = n9881 ^ n8866 ^ n5220 ;
  assign n9883 = ( n443 & n4585 ) | ( n443 & n5116 ) | ( n4585 & n5116 ) ;
  assign n9884 = ( n1891 & n9882 ) | ( n1891 & n9883 ) | ( n9882 & n9883 ) ;
  assign n9879 = n6210 ^ n5742 ^ n1880 ;
  assign n9880 = n9879 ^ n6435 ^ n2178 ;
  assign n9885 = n9884 ^ n9880 ^ n1109 ;
  assign n9895 = n6498 ^ n3144 ^ n2390 ;
  assign n9896 = n9895 ^ n3774 ^ n1593 ;
  assign n9889 = ( x82 & n291 ) | ( x82 & ~n4275 ) | ( n291 & ~n4275 ) ;
  assign n9892 = ( n857 & ~n2810 ) | ( n857 & n5847 ) | ( ~n2810 & n5847 ) ;
  assign n9890 = n4711 ^ n3932 ^ n3257 ;
  assign n9891 = ( n5057 & n6037 ) | ( n5057 & n9890 ) | ( n6037 & n9890 ) ;
  assign n9893 = n9892 ^ n9891 ^ n3696 ;
  assign n9894 = ( n6651 & n9889 ) | ( n6651 & ~n9893 ) | ( n9889 & ~n9893 ) ;
  assign n9897 = n9896 ^ n9894 ^ n1939 ;
  assign n9886 = n8940 ^ n6765 ^ n2701 ;
  assign n9887 = n9886 ^ n1923 ^ n1569 ;
  assign n9888 = n9887 ^ n9709 ^ n3343 ;
  assign n9898 = n9897 ^ n9888 ^ x32 ;
  assign n9899 = ( n9878 & ~n9885 ) | ( n9878 & n9898 ) | ( ~n9885 & n9898 ) ;
  assign n9900 = ( n3387 & n7092 ) | ( n3387 & ~n8516 ) | ( n7092 & ~n8516 ) ;
  assign n9901 = ( n2769 & ~n3798 ) | ( n2769 & n9900 ) | ( ~n3798 & n9900 ) ;
  assign n9902 = n7688 ^ n7564 ^ n3530 ;
  assign n9903 = ( ~n1549 & n4420 ) | ( ~n1549 & n9007 ) | ( n4420 & n9007 ) ;
  assign n9904 = ( n425 & ~n8285 ) | ( n425 & n9903 ) | ( ~n8285 & n9903 ) ;
  assign n9905 = n6553 ^ n3476 ^ n710 ;
  assign n9906 = n9905 ^ n4908 ^ n4623 ;
  assign n9907 = n8475 ^ n4265 ^ n1529 ;
  assign n9910 = n6765 ^ n6008 ^ n751 ;
  assign n9911 = n9910 ^ n8310 ^ n182 ;
  assign n9908 = n8643 ^ n5966 ^ n509 ;
  assign n9909 = ( n520 & n6011 ) | ( n520 & n9908 ) | ( n6011 & n9908 ) ;
  assign n9912 = n9911 ^ n9909 ^ n3836 ;
  assign n9913 = ( n4774 & n9907 ) | ( n4774 & n9912 ) | ( n9907 & n9912 ) ;
  assign n9914 = n6638 ^ n5969 ^ n5631 ;
  assign n9915 = n9914 ^ n2479 ^ n1763 ;
  assign n9916 = ( n2327 & ~n4121 ) | ( n2327 & n9915 ) | ( ~n4121 & n9915 ) ;
  assign n9921 = ( ~n1006 & n2742 ) | ( ~n1006 & n6153 ) | ( n2742 & n6153 ) ;
  assign n9922 = n9921 ^ n9064 ^ n4924 ;
  assign n9923 = ( n2881 & n3857 ) | ( n2881 & n4353 ) | ( n3857 & n4353 ) ;
  assign n9924 = ( n5577 & n6469 ) | ( n5577 & ~n9923 ) | ( n6469 & ~n9923 ) ;
  assign n9925 = ( n3025 & n3299 ) | ( n3025 & ~n9924 ) | ( n3299 & ~n9924 ) ;
  assign n9926 = ( n7907 & ~n9922 ) | ( n7907 & n9925 ) | ( ~n9922 & n9925 ) ;
  assign n9919 = ( n931 & n4265 ) | ( n931 & ~n6063 ) | ( n4265 & ~n6063 ) ;
  assign n9917 = ( n658 & n3636 ) | ( n658 & ~n5346 ) | ( n3636 & ~n5346 ) ;
  assign n9918 = ( n733 & n1365 ) | ( n733 & n9917 ) | ( n1365 & n9917 ) ;
  assign n9920 = n9919 ^ n9918 ^ n3684 ;
  assign n9927 = n9926 ^ n9920 ^ n2046 ;
  assign n9928 = ( n558 & ~n2158 ) | ( n558 & n3164 ) | ( ~n2158 & n3164 ) ;
  assign n9929 = n6147 ^ n4759 ^ n3929 ;
  assign n9930 = ( n2462 & ~n3909 ) | ( n2462 & n9929 ) | ( ~n3909 & n9929 ) ;
  assign n9931 = n9930 ^ n8524 ^ n1999 ;
  assign n9932 = n9931 ^ n7808 ^ n2650 ;
  assign n9933 = n9932 ^ n2052 ^ n694 ;
  assign n9934 = ( n8518 & n9928 ) | ( n8518 & ~n9933 ) | ( n9928 & ~n9933 ) ;
  assign n9935 = ( n2507 & n3434 ) | ( n2507 & n8525 ) | ( n3434 & n8525 ) ;
  assign n9938 = ( n732 & ~n1081 ) | ( n732 & n3385 ) | ( ~n1081 & n3385 ) ;
  assign n9936 = n7170 ^ n1612 ^ n738 ;
  assign n9937 = n9936 ^ n5296 ^ n898 ;
  assign n9939 = n9938 ^ n9937 ^ n653 ;
  assign n9940 = n6988 ^ n4796 ^ n2983 ;
  assign n9941 = ( ~n2684 & n7811 ) | ( ~n2684 & n9940 ) | ( n7811 & n9940 ) ;
  assign n9942 = ( n2619 & ~n6593 ) | ( n2619 & n8322 ) | ( ~n6593 & n8322 ) ;
  assign n9943 = n7248 ^ n3862 ^ n177 ;
  assign n9944 = ( ~n5819 & n9942 ) | ( ~n5819 & n9943 ) | ( n9942 & n9943 ) ;
  assign n9947 = n5302 ^ n4910 ^ n561 ;
  assign n9945 = ( ~x26 & n3096 ) | ( ~x26 & n5228 ) | ( n3096 & n5228 ) ;
  assign n9946 = ( n646 & n9830 ) | ( n646 & ~n9945 ) | ( n9830 & ~n9945 ) ;
  assign n9948 = n9947 ^ n9946 ^ n967 ;
  assign n9949 = ( n3811 & n9944 ) | ( n3811 & n9948 ) | ( n9944 & n9948 ) ;
  assign n9950 = ( ~n411 & n3845 ) | ( ~n411 & n6288 ) | ( n3845 & n6288 ) ;
  assign n9951 = n9950 ^ n6293 ^ n3856 ;
  assign n9952 = ( n819 & ~n2907 ) | ( n819 & n9518 ) | ( ~n2907 & n9518 ) ;
  assign n9953 = ( ~n3760 & n5456 ) | ( ~n3760 & n9952 ) | ( n5456 & n9952 ) ;
  assign n9963 = n5604 ^ n1523 ^ n978 ;
  assign n9962 = ( ~n1230 & n2592 ) | ( ~n1230 & n9538 ) | ( n2592 & n9538 ) ;
  assign n9954 = n4884 ^ n2661 ^ n807 ;
  assign n9955 = ( n1758 & n4321 ) | ( n1758 & ~n7658 ) | ( n4321 & ~n7658 ) ;
  assign n9956 = ( x91 & n7218 ) | ( x91 & n9955 ) | ( n7218 & n9955 ) ;
  assign n9957 = ( n3248 & n9733 ) | ( n3248 & n9956 ) | ( n9733 & n9956 ) ;
  assign n9958 = ( n328 & ~n1233 ) | ( n328 & n1267 ) | ( ~n1233 & n1267 ) ;
  assign n9959 = ( n4387 & ~n5810 ) | ( n4387 & n9958 ) | ( ~n5810 & n9958 ) ;
  assign n9960 = ( n9954 & n9957 ) | ( n9954 & ~n9959 ) | ( n9957 & ~n9959 ) ;
  assign n9961 = ( ~n2856 & n6126 ) | ( ~n2856 & n9960 ) | ( n6126 & n9960 ) ;
  assign n9964 = n9963 ^ n9962 ^ n9961 ;
  assign n9965 = n1685 ^ n1268 ^ n320 ;
  assign n9966 = n7296 ^ n2353 ^ n306 ;
  assign n9967 = ( n1630 & n2337 ) | ( n1630 & ~n7410 ) | ( n2337 & ~n7410 ) ;
  assign n9968 = ( ~n2901 & n9966 ) | ( ~n2901 & n9967 ) | ( n9966 & n9967 ) ;
  assign n9969 = ( n8165 & n9965 ) | ( n8165 & n9968 ) | ( n9965 & n9968 ) ;
  assign n9970 = n9039 ^ n5202 ^ n2747 ;
  assign n9971 = ( n4340 & ~n5052 ) | ( n4340 & n9970 ) | ( ~n5052 & n9970 ) ;
  assign n9972 = n8360 ^ n2710 ^ n2644 ;
  assign n9973 = n9972 ^ n8041 ^ n5327 ;
  assign n9974 = n5609 ^ n2120 ^ n1388 ;
  assign n9975 = n9974 ^ n7056 ^ n6029 ;
  assign n9976 = ( ~n2075 & n2396 ) | ( ~n2075 & n9975 ) | ( n2396 & n9975 ) ;
  assign n9977 = n9976 ^ n3783 ^ n2429 ;
  assign n9978 = ( ~n1944 & n5234 ) | ( ~n1944 & n9574 ) | ( n5234 & n9574 ) ;
  assign n9979 = n9978 ^ n7217 ^ n7129 ;
  assign n9980 = ( n8292 & n8732 ) | ( n8292 & ~n9256 ) | ( n8732 & ~n9256 ) ;
  assign n9981 = ( ~n1032 & n7938 ) | ( ~n1032 & n9980 ) | ( n7938 & n9980 ) ;
  assign n9992 = n6156 ^ n1790 ^ n1054 ;
  assign n9991 = ( ~x89 & n668 ) | ( ~x89 & n7384 ) | ( n668 & n7384 ) ;
  assign n9993 = n9992 ^ n9991 ^ n7651 ;
  assign n9982 = ( n2342 & ~n5807 ) | ( n2342 & n7801 ) | ( ~n5807 & n7801 ) ;
  assign n9985 = ( ~n1262 & n1422 ) | ( ~n1262 & n2034 ) | ( n1422 & n2034 ) ;
  assign n9983 = ( ~n1329 & n1787 ) | ( ~n1329 & n4272 ) | ( n1787 & n4272 ) ;
  assign n9984 = ( n913 & n4101 ) | ( n913 & n9983 ) | ( n4101 & n9983 ) ;
  assign n9986 = n9985 ^ n9984 ^ n4956 ;
  assign n9987 = ( ~x87 & n9982 ) | ( ~x87 & n9986 ) | ( n9982 & n9986 ) ;
  assign n9988 = n7570 ^ n4804 ^ n4539 ;
  assign n9989 = ( n4939 & n8797 ) | ( n4939 & ~n9988 ) | ( n8797 & ~n9988 ) ;
  assign n9990 = ( ~n6806 & n9987 ) | ( ~n6806 & n9989 ) | ( n9987 & n9989 ) ;
  assign n9994 = n9993 ^ n9990 ^ n9158 ;
  assign n9995 = n3695 ^ n2683 ^ n458 ;
  assign n9996 = ( ~n6292 & n7533 ) | ( ~n6292 & n9995 ) | ( n7533 & n9995 ) ;
  assign n9997 = ( n2206 & ~n6611 ) | ( n2206 & n7245 ) | ( ~n6611 & n7245 ) ;
  assign n9998 = ( n3235 & n9996 ) | ( n3235 & ~n9997 ) | ( n9996 & ~n9997 ) ;
  assign n10002 = ( n2019 & ~n5795 ) | ( n2019 & n8555 ) | ( ~n5795 & n8555 ) ;
  assign n10003 = n10002 ^ n3332 ^ n3217 ;
  assign n10004 = n10003 ^ n9281 ^ n6238 ;
  assign n9999 = n3506 ^ n2943 ^ n1309 ;
  assign n10000 = ( n4464 & n5077 ) | ( n4464 & n9999 ) | ( n5077 & n9999 ) ;
  assign n10001 = ( n2147 & n3917 ) | ( n2147 & n10000 ) | ( n3917 & n10000 ) ;
  assign n10005 = n10004 ^ n10001 ^ n2240 ;
  assign n10006 = n3009 ^ n1935 ^ n389 ;
  assign n10007 = n5646 ^ n5202 ^ n2094 ;
  assign n10008 = ( n9917 & ~n10006 ) | ( n9917 & n10007 ) | ( ~n10006 & n10007 ) ;
  assign n10013 = ( n2656 & n3203 ) | ( n2656 & n8449 ) | ( n3203 & n8449 ) ;
  assign n10014 = n10013 ^ n7265 ^ n3950 ;
  assign n10015 = n10014 ^ n6308 ^ n562 ;
  assign n10009 = n7910 ^ n7085 ^ n4519 ;
  assign n10010 = ( n900 & n1755 ) | ( n900 & n4747 ) | ( n1755 & n4747 ) ;
  assign n10011 = ( n2636 & n10009 ) | ( n2636 & ~n10010 ) | ( n10009 & ~n10010 ) ;
  assign n10012 = n10011 ^ n6836 ^ n6301 ;
  assign n10016 = n10015 ^ n10012 ^ n3873 ;
  assign n10022 = n5432 ^ n3971 ^ n2856 ;
  assign n10019 = n5904 ^ n1154 ^ n751 ;
  assign n10020 = ( ~n2631 & n3249 ) | ( ~n2631 & n10019 ) | ( n3249 & n10019 ) ;
  assign n10017 = ( n2850 & n3942 ) | ( n2850 & n4878 ) | ( n3942 & n4878 ) ;
  assign n10018 = n10017 ^ n5759 ^ n4539 ;
  assign n10021 = n10020 ^ n10018 ^ n8145 ;
  assign n10023 = n10022 ^ n10021 ^ n8442 ;
  assign n10024 = ( ~n5570 & n6996 ) | ( ~n5570 & n10023 ) | ( n6996 & n10023 ) ;
  assign n10025 = n6862 ^ n3126 ^ n1445 ;
  assign n10026 = n10025 ^ n2519 ^ n1586 ;
  assign n10027 = n10026 ^ n3395 ^ n1137 ;
  assign n10028 = ( ~n815 & n5275 ) | ( ~n815 & n9626 ) | ( n5275 & n9626 ) ;
  assign n10029 = n8802 ^ n5435 ^ n1108 ;
  assign n10030 = ( n10027 & ~n10028 ) | ( n10027 & n10029 ) | ( ~n10028 & n10029 ) ;
  assign n10031 = ( n191 & n8817 ) | ( n191 & n9043 ) | ( n8817 & n9043 ) ;
  assign n10032 = n10031 ^ n3559 ^ n2423 ;
  assign n10033 = ( n2894 & n5043 ) | ( n2894 & ~n10032 ) | ( n5043 & ~n10032 ) ;
  assign n10034 = ( n6928 & ~n8368 ) | ( n6928 & n10033 ) | ( ~n8368 & n10033 ) ;
  assign n10035 = n2043 ^ n1977 ^ n1188 ;
  assign n10036 = n10035 ^ n9867 ^ n2353 ;
  assign n10037 = ( n3586 & ~n7256 ) | ( n3586 & n10036 ) | ( ~n7256 & n10036 ) ;
  assign n10039 = n2952 ^ n2457 ^ n1368 ;
  assign n10040 = n10039 ^ n5938 ^ n5885 ;
  assign n10038 = n9256 ^ n7831 ^ n3365 ;
  assign n10041 = n10040 ^ n10038 ^ n6889 ;
  assign n10042 = n3184 ^ n2440 ^ n980 ;
  assign n10043 = n10042 ^ n6095 ^ n2735 ;
  assign n10044 = ( ~x12 & n2746 ) | ( ~x12 & n3946 ) | ( n2746 & n3946 ) ;
  assign n10045 = ( n6044 & n9221 ) | ( n6044 & n10044 ) | ( n9221 & n10044 ) ;
  assign n10046 = ( n4327 & n10043 ) | ( n4327 & ~n10045 ) | ( n10043 & ~n10045 ) ;
  assign n10048 = n4384 ^ n3837 ^ x76 ;
  assign n10047 = n6776 ^ n5211 ^ n3385 ;
  assign n10049 = n10048 ^ n10047 ^ n237 ;
  assign n10050 = n10049 ^ n2840 ^ n207 ;
  assign n10051 = n10050 ^ n10048 ^ n568 ;
  assign n10052 = ( ~n4587 & n7942 ) | ( ~n4587 & n10051 ) | ( n7942 & n10051 ) ;
  assign n10053 = ( n1213 & ~n2984 ) | ( n1213 & n3961 ) | ( ~n2984 & n3961 ) ;
  assign n10054 = ( n915 & ~n5659 ) | ( n915 & n10053 ) | ( ~n5659 & n10053 ) ;
  assign n10055 = n10054 ^ n7858 ^ n4962 ;
  assign n10056 = n7544 ^ n4111 ^ n1738 ;
  assign n10057 = ( x62 & ~n487 ) | ( x62 & n3160 ) | ( ~n487 & n3160 ) ;
  assign n10058 = ( n3691 & n4473 ) | ( n3691 & n10057 ) | ( n4473 & n10057 ) ;
  assign n10059 = ( ~n163 & n8107 ) | ( ~n163 & n8299 ) | ( n8107 & n8299 ) ;
  assign n10060 = ( n540 & n4409 ) | ( n540 & n10059 ) | ( n4409 & n10059 ) ;
  assign n10061 = ( n3812 & ~n10058 ) | ( n3812 & n10060 ) | ( ~n10058 & n10060 ) ;
  assign n10062 = n5600 ^ n5232 ^ n565 ;
  assign n10063 = ( n4123 & n5710 ) | ( n4123 & n10062 ) | ( n5710 & n10062 ) ;
  assign n10064 = ( n10056 & n10061 ) | ( n10056 & ~n10063 ) | ( n10061 & ~n10063 ) ;
  assign n10067 = n9967 ^ n5887 ^ n5133 ;
  assign n10065 = n8657 ^ n3582 ^ n782 ;
  assign n10066 = n10065 ^ n7043 ^ n242 ;
  assign n10068 = n10067 ^ n10066 ^ n6274 ;
  assign n10069 = n10068 ^ n5174 ^ n490 ;
  assign n10070 = ( n1987 & n5010 ) | ( n1987 & ~n5735 ) | ( n5010 & ~n5735 ) ;
  assign n10074 = ( x69 & ~n4894 ) | ( x69 & n5351 ) | ( ~n4894 & n5351 ) ;
  assign n10071 = n1610 ^ n456 ^ x60 ;
  assign n10072 = ( n1283 & n5791 ) | ( n1283 & ~n10071 ) | ( n5791 & ~n10071 ) ;
  assign n10073 = ( n1654 & n10019 ) | ( n1654 & n10072 ) | ( n10019 & n10072 ) ;
  assign n10075 = n10074 ^ n10073 ^ n1566 ;
  assign n10076 = ( ~n2066 & n5077 ) | ( ~n2066 & n10075 ) | ( n5077 & n10075 ) ;
  assign n10077 = ( n1244 & n1474 ) | ( n1244 & n5439 ) | ( n1474 & n5439 ) ;
  assign n10078 = ( n1978 & n6024 ) | ( n1978 & n10077 ) | ( n6024 & n10077 ) ;
  assign n10079 = n10078 ^ n6257 ^ n652 ;
  assign n10080 = ( n723 & n4412 ) | ( n723 & n6117 ) | ( n4412 & n6117 ) ;
  assign n10081 = ( n449 & n663 ) | ( n449 & n10080 ) | ( n663 & n10080 ) ;
  assign n10085 = ( n6550 & n7760 ) | ( n6550 & n7939 ) | ( n7760 & n7939 ) ;
  assign n10082 = ( n3837 & n5120 ) | ( n3837 & ~n5282 ) | ( n5120 & ~n5282 ) ;
  assign n10083 = ( n196 & n4639 ) | ( n196 & ~n10082 ) | ( n4639 & ~n10082 ) ;
  assign n10084 = ( ~n5796 & n9905 ) | ( ~n5796 & n10083 ) | ( n9905 & n10083 ) ;
  assign n10086 = n10085 ^ n10084 ^ n3875 ;
  assign n10096 = ( n2152 & n3015 ) | ( n2152 & ~n3127 ) | ( n3015 & ~n3127 ) ;
  assign n10094 = n8067 ^ n7252 ^ n3339 ;
  assign n10095 = n10094 ^ n7475 ^ n824 ;
  assign n10092 = ( ~n3888 & n5485 ) | ( ~n3888 & n8836 ) | ( n5485 & n8836 ) ;
  assign n10091 = n2413 ^ n1062 ^ n752 ;
  assign n10087 = n3686 ^ n3670 ^ n2848 ;
  assign n10088 = ( n3485 & ~n3799 ) | ( n3485 & n10087 ) | ( ~n3799 & n10087 ) ;
  assign n10089 = ( n652 & ~n1883 ) | ( n652 & n10088 ) | ( ~n1883 & n10088 ) ;
  assign n10090 = ( n1639 & n7931 ) | ( n1639 & n10089 ) | ( n7931 & n10089 ) ;
  assign n10093 = n10092 ^ n10091 ^ n10090 ;
  assign n10097 = n10096 ^ n10095 ^ n10093 ;
  assign n10098 = ( n2926 & ~n7271 ) | ( n2926 & n8365 ) | ( ~n7271 & n8365 ) ;
  assign n10099 = ( ~n3740 & n6943 ) | ( ~n3740 & n7316 ) | ( n6943 & n7316 ) ;
  assign n10100 = n10099 ^ n6537 ^ n5052 ;
  assign n10101 = ( n3747 & n10098 ) | ( n3747 & ~n10100 ) | ( n10098 & ~n10100 ) ;
  assign n10102 = ( ~n737 & n2888 ) | ( ~n737 & n5621 ) | ( n2888 & n5621 ) ;
  assign n10103 = n9455 ^ n6496 ^ n4129 ;
  assign n10104 = ( n981 & n5554 ) | ( n981 & n10103 ) | ( n5554 & n10103 ) ;
  assign n10105 = n7483 ^ n2731 ^ n215 ;
  assign n10106 = n3637 ^ n1305 ^ n310 ;
  assign n10107 = n10106 ^ n5784 ^ n4750 ;
  assign n10108 = n10107 ^ n7985 ^ n330 ;
  assign n10109 = n10108 ^ n7145 ^ n2309 ;
  assign n10110 = ( n1479 & n6922 ) | ( n1479 & n7435 ) | ( n6922 & n7435 ) ;
  assign n10111 = ( ~n3311 & n9161 ) | ( ~n3311 & n10110 ) | ( n9161 & n10110 ) ;
  assign n10112 = ( n4407 & n7009 ) | ( n4407 & n10111 ) | ( n7009 & n10111 ) ;
  assign n10113 = ( ~n4769 & n10109 ) | ( ~n4769 & n10112 ) | ( n10109 & n10112 ) ;
  assign n10114 = n2994 ^ n2635 ^ n2041 ;
  assign n10115 = ( n2115 & n6325 ) | ( n2115 & n8593 ) | ( n6325 & n8593 ) ;
  assign n10116 = ( n2395 & ~n6470 ) | ( n2395 & n10115 ) | ( ~n6470 & n10115 ) ;
  assign n10117 = ( n3020 & n10114 ) | ( n3020 & ~n10116 ) | ( n10114 & ~n10116 ) ;
  assign n10118 = ( n3741 & n5169 ) | ( n3741 & ~n10117 ) | ( n5169 & ~n10117 ) ;
  assign n10121 = ( ~n2754 & n4640 ) | ( ~n2754 & n8026 ) | ( n4640 & n8026 ) ;
  assign n10119 = ( ~n5037 & n5721 ) | ( ~n5037 & n7368 ) | ( n5721 & n7368 ) ;
  assign n10120 = ( n7852 & ~n9846 ) | ( n7852 & n10119 ) | ( ~n9846 & n10119 ) ;
  assign n10122 = n10121 ^ n10120 ^ n7060 ;
  assign n10123 = ( ~n688 & n10118 ) | ( ~n688 & n10122 ) | ( n10118 & n10122 ) ;
  assign n10130 = n3910 ^ n2049 ^ n162 ;
  assign n10126 = n3471 ^ n2448 ^ n160 ;
  assign n10127 = ( ~n2872 & n4048 ) | ( ~n2872 & n10126 ) | ( n4048 & n10126 ) ;
  assign n10128 = ( n9119 & n9755 ) | ( n9119 & n10127 ) | ( n9755 & n10127 ) ;
  assign n10129 = ( n191 & ~n1075 ) | ( n191 & n10128 ) | ( ~n1075 & n10128 ) ;
  assign n10124 = n6252 ^ n1063 ^ n950 ;
  assign n10125 = ( n3445 & ~n6422 ) | ( n3445 & n10124 ) | ( ~n6422 & n10124 ) ;
  assign n10131 = n10130 ^ n10129 ^ n10125 ;
  assign n10132 = ( n442 & n8412 ) | ( n442 & ~n10131 ) | ( n8412 & ~n10131 ) ;
  assign n10133 = ( n7454 & n9882 ) | ( n7454 & ~n10132 ) | ( n9882 & ~n10132 ) ;
  assign n10138 = ( n1014 & n2055 ) | ( n1014 & ~n7841 ) | ( n2055 & ~n7841 ) ;
  assign n10139 = n10138 ^ n9437 ^ n4725 ;
  assign n10134 = n7055 ^ n3409 ^ n342 ;
  assign n10135 = n5609 ^ n1956 ^ n542 ;
  assign n10136 = ( n6057 & n10134 ) | ( n6057 & ~n10135 ) | ( n10134 & ~n10135 ) ;
  assign n10137 = n10136 ^ n8508 ^ n3702 ;
  assign n10140 = n10139 ^ n10137 ^ n5617 ;
  assign n10141 = ( ~n420 & n2771 ) | ( ~n420 & n7760 ) | ( n2771 & n7760 ) ;
  assign n10142 = ( n4998 & n9559 ) | ( n4998 & n10141 ) | ( n9559 & n10141 ) ;
  assign n10143 = ( ~n10133 & n10140 ) | ( ~n10133 & n10142 ) | ( n10140 & n10142 ) ;
  assign n10146 = n10048 ^ n3249 ^ n2874 ;
  assign n10144 = ( n214 & ~n2123 ) | ( n214 & n3686 ) | ( ~n2123 & n3686 ) ;
  assign n10145 = n10144 ^ n2121 ^ n1472 ;
  assign n10147 = n10146 ^ n10145 ^ n847 ;
  assign n10148 = ( n1876 & n2585 ) | ( n1876 & ~n2793 ) | ( n2585 & ~n2793 ) ;
  assign n10149 = n10148 ^ n5405 ^ n131 ;
  assign n10150 = ( n4983 & ~n5612 ) | ( n4983 & n10149 ) | ( ~n5612 & n10149 ) ;
  assign n10151 = n8936 ^ n6577 ^ n4325 ;
  assign n10152 = ( ~n4065 & n4242 ) | ( ~n4065 & n7548 ) | ( n4242 & n7548 ) ;
  assign n10153 = n10152 ^ n2904 ^ n2438 ;
  assign n10154 = n10153 ^ n7730 ^ n6960 ;
  assign n10155 = ( n7877 & n10151 ) | ( n7877 & n10154 ) | ( n10151 & n10154 ) ;
  assign n10156 = ( n1083 & ~n8010 ) | ( n1083 & n8551 ) | ( ~n8010 & n8551 ) ;
  assign n10157 = n3292 ^ n859 ^ n573 ;
  assign n10158 = ( n4864 & n5555 ) | ( n4864 & ~n10157 ) | ( n5555 & ~n10157 ) ;
  assign n10160 = n5682 ^ n4348 ^ n4345 ;
  assign n10159 = n9790 ^ n5371 ^ n4594 ;
  assign n10161 = n10160 ^ n10159 ^ n5142 ;
  assign n10162 = ( n7083 & n9430 ) | ( n7083 & n10161 ) | ( n9430 & n10161 ) ;
  assign n10163 = ( n1164 & n2804 ) | ( n1164 & ~n4670 ) | ( n2804 & ~n4670 ) ;
  assign n10178 = ( n3562 & ~n4500 ) | ( n3562 & n5339 ) | ( ~n4500 & n5339 ) ;
  assign n10175 = n2919 ^ n2485 ^ n2386 ;
  assign n10174 = n5331 ^ n2868 ^ x98 ;
  assign n10176 = n10175 ^ n10174 ^ x62 ;
  assign n10167 = ( ~n2053 & n2852 ) | ( ~n2053 & n8249 ) | ( n2852 & n8249 ) ;
  assign n10168 = n10167 ^ n3807 ^ n1836 ;
  assign n10169 = ( n3594 & n7890 ) | ( n3594 & ~n10168 ) | ( n7890 & ~n10168 ) ;
  assign n10166 = ( n3115 & n5559 ) | ( n3115 & n8896 ) | ( n5559 & n8896 ) ;
  assign n10170 = n10169 ^ n10166 ^ n3637 ;
  assign n10171 = n3729 ^ n2183 ^ n720 ;
  assign n10172 = ( n4503 & n8817 ) | ( n4503 & ~n10171 ) | ( n8817 & ~n10171 ) ;
  assign n10173 = ( n8175 & ~n10170 ) | ( n8175 & n10172 ) | ( ~n10170 & n10172 ) ;
  assign n10177 = n10176 ^ n10173 ^ n9687 ;
  assign n10164 = ( n4061 & n4789 ) | ( n4061 & n8486 ) | ( n4789 & n8486 ) ;
  assign n10165 = n10164 ^ n7126 ^ n6701 ;
  assign n10179 = n10178 ^ n10177 ^ n10165 ;
  assign n10180 = n8895 ^ n7086 ^ n2886 ;
  assign n10181 = n8341 ^ n3973 ^ n2059 ;
  assign n10182 = ( n5710 & n10180 ) | ( n5710 & n10181 ) | ( n10180 & n10181 ) ;
  assign n10183 = n10182 ^ n5175 ^ n4953 ;
  assign n10184 = n10183 ^ n9787 ^ n3440 ;
  assign n10185 = ( x24 & n1277 ) | ( x24 & ~n3629 ) | ( n1277 & ~n3629 ) ;
  assign n10186 = n10185 ^ n3190 ^ n1503 ;
  assign n10187 = n10186 ^ n3122 ^ n1812 ;
  assign n10191 = n8766 ^ n7085 ^ n4336 ;
  assign n10189 = ( ~n181 & n1388 ) | ( ~n181 & n4052 ) | ( n1388 & n4052 ) ;
  assign n10190 = ( ~x57 & n1484 ) | ( ~x57 & n10189 ) | ( n1484 & n10189 ) ;
  assign n10188 = ( ~n3929 & n6877 ) | ( ~n3929 & n9428 ) | ( n6877 & n9428 ) ;
  assign n10192 = n10191 ^ n10190 ^ n10188 ;
  assign n10193 = n9076 ^ n8963 ^ n7583 ;
  assign n10194 = ( ~n2663 & n6106 ) | ( ~n2663 & n10193 ) | ( n6106 & n10193 ) ;
  assign n10195 = ( n6220 & n8755 ) | ( n6220 & ~n10194 ) | ( n8755 & ~n10194 ) ;
  assign n10196 = n9025 ^ n2728 ^ n2154 ;
  assign n10197 = n10196 ^ n6867 ^ n5846 ;
  assign n10199 = ( n1364 & n3711 ) | ( n1364 & n8754 ) | ( n3711 & n8754 ) ;
  assign n10200 = ( ~n6546 & n8630 ) | ( ~n6546 & n10199 ) | ( n8630 & n10199 ) ;
  assign n10201 = n10200 ^ n9558 ^ n4674 ;
  assign n10198 = n3192 ^ n369 ^ n333 ;
  assign n10202 = n10201 ^ n10198 ^ n1566 ;
  assign n10203 = ( ~n5283 & n7807 ) | ( ~n5283 & n8326 ) | ( n7807 & n8326 ) ;
  assign n10204 = ( n1720 & n9388 ) | ( n1720 & n10203 ) | ( n9388 & n10203 ) ;
  assign n10205 = ( ~n10197 & n10202 ) | ( ~n10197 & n10204 ) | ( n10202 & n10204 ) ;
  assign n10208 = ( ~n1321 & n3414 ) | ( ~n1321 & n5689 ) | ( n3414 & n5689 ) ;
  assign n10206 = ( n1143 & n1414 ) | ( n1143 & n9508 ) | ( n1414 & n9508 ) ;
  assign n10207 = n10206 ^ n5826 ^ n2787 ;
  assign n10209 = n10208 ^ n10207 ^ n324 ;
  assign n10210 = ( n1492 & ~n9016 ) | ( n1492 & n10176 ) | ( ~n9016 & n10176 ) ;
  assign n10211 = ( n2469 & ~n3802 ) | ( n2469 & n3888 ) | ( ~n3802 & n3888 ) ;
  assign n10212 = ( ~n1170 & n5172 ) | ( ~n1170 & n10211 ) | ( n5172 & n10211 ) ;
  assign n10213 = ( x127 & n5487 ) | ( x127 & n8769 ) | ( n5487 & n8769 ) ;
  assign n10214 = ( ~n1748 & n10212 ) | ( ~n1748 & n10213 ) | ( n10212 & n10213 ) ;
  assign n10219 = n2374 ^ n915 ^ n466 ;
  assign n10220 = ( n658 & ~n4659 ) | ( n658 & n10219 ) | ( ~n4659 & n10219 ) ;
  assign n10215 = n5890 ^ n1829 ^ n1254 ;
  assign n10216 = ( n501 & ~n5111 ) | ( n501 & n10215 ) | ( ~n5111 & n10215 ) ;
  assign n10217 = n10216 ^ n1591 ^ x60 ;
  assign n10218 = ( ~n1053 & n3481 ) | ( ~n1053 & n10217 ) | ( n3481 & n10217 ) ;
  assign n10221 = n10220 ^ n10218 ^ n1361 ;
  assign n10222 = ( n2554 & n5983 ) | ( n2554 & ~n10221 ) | ( n5983 & ~n10221 ) ;
  assign n10223 = ( n828 & n5260 ) | ( n828 & n6148 ) | ( n5260 & n6148 ) ;
  assign n10224 = n10223 ^ n9698 ^ n3290 ;
  assign n10225 = ( n1190 & n10222 ) | ( n1190 & n10224 ) | ( n10222 & n10224 ) ;
  assign n10226 = n9109 ^ n8022 ^ n4989 ;
  assign n10227 = ( n5321 & n7947 ) | ( n5321 & ~n10226 ) | ( n7947 & ~n10226 ) ;
  assign n10228 = n8269 ^ n6229 ^ n5851 ;
  assign n10229 = n10228 ^ n4731 ^ n1879 ;
  assign n10233 = n8018 ^ n1523 ^ x88 ;
  assign n10232 = ( n3667 & n5640 ) | ( n3667 & n7845 ) | ( n5640 & n7845 ) ;
  assign n10230 = n4192 ^ n4087 ^ n3111 ;
  assign n10231 = ( n2344 & ~n3446 ) | ( n2344 & n10230 ) | ( ~n3446 & n10230 ) ;
  assign n10234 = n10233 ^ n10232 ^ n10231 ;
  assign n10235 = ( ~n1669 & n1919 ) | ( ~n1669 & n7323 ) | ( n1919 & n7323 ) ;
  assign n10243 = ( n2733 & n3737 ) | ( n2733 & ~n6896 ) | ( n3737 & ~n6896 ) ;
  assign n10241 = n8334 ^ n2124 ^ n1230 ;
  assign n10242 = ( ~n733 & n6831 ) | ( ~n733 & n10241 ) | ( n6831 & n10241 ) ;
  assign n10244 = n10243 ^ n10242 ^ n1889 ;
  assign n10245 = ( n1371 & n2401 ) | ( n1371 & ~n10244 ) | ( n2401 & ~n10244 ) ;
  assign n10237 = n3658 ^ n3117 ^ n2873 ;
  assign n10238 = n8252 ^ n4768 ^ n758 ;
  assign n10239 = n10238 ^ n9039 ^ n6605 ;
  assign n10240 = ( n1449 & n10237 ) | ( n1449 & n10239 ) | ( n10237 & n10239 ) ;
  assign n10236 = ( ~n1115 & n3275 ) | ( ~n1115 & n3318 ) | ( n3275 & n3318 ) ;
  assign n10246 = n10245 ^ n10240 ^ n10236 ;
  assign n10247 = n3383 ^ n2315 ^ n1392 ;
  assign n10248 = ( n1670 & n6591 ) | ( n1670 & ~n6817 ) | ( n6591 & ~n6817 ) ;
  assign n10249 = ( n5503 & n10247 ) | ( n5503 & ~n10248 ) | ( n10247 & ~n10248 ) ;
  assign n10250 = ( n1769 & n1943 ) | ( n1769 & ~n10249 ) | ( n1943 & ~n10249 ) ;
  assign n10258 = n2173 ^ n350 ^ n281 ;
  assign n10259 = n10258 ^ n5202 ^ n3768 ;
  assign n10260 = ( n1245 & n2468 ) | ( n1245 & n10259 ) | ( n2468 & n10259 ) ;
  assign n10261 = n10260 ^ n10026 ^ n3792 ;
  assign n10257 = ( n7463 & ~n7589 ) | ( n7463 & n10135 ) | ( ~n7589 & n10135 ) ;
  assign n10251 = n4385 ^ n4228 ^ n4014 ;
  assign n10252 = ( n1021 & ~n6224 ) | ( n1021 & n10251 ) | ( ~n6224 & n10251 ) ;
  assign n10253 = ( n1013 & ~n7144 ) | ( n1013 & n9826 ) | ( ~n7144 & n9826 ) ;
  assign n10254 = ( n7344 & ~n10252 ) | ( n7344 & n10253 ) | ( ~n10252 & n10253 ) ;
  assign n10255 = ( n1488 & n6506 ) | ( n1488 & n10254 ) | ( n6506 & n10254 ) ;
  assign n10256 = ( n3281 & ~n8412 ) | ( n3281 & n10255 ) | ( ~n8412 & n10255 ) ;
  assign n10262 = n10261 ^ n10257 ^ n10256 ;
  assign n10263 = ( n4069 & n10250 ) | ( n4069 & n10262 ) | ( n10250 & n10262 ) ;
  assign n10268 = n2385 ^ n1579 ^ n1213 ;
  assign n10269 = ( n4721 & ~n7352 ) | ( n4721 & n10268 ) | ( ~n7352 & n10268 ) ;
  assign n10265 = n1566 ^ n903 ^ n753 ;
  assign n10266 = n10265 ^ n3535 ^ n3262 ;
  assign n10264 = ( n6324 & ~n7425 ) | ( n6324 & n8352 ) | ( ~n7425 & n8352 ) ;
  assign n10267 = n10266 ^ n10264 ^ n1922 ;
  assign n10270 = n10269 ^ n10267 ^ n9070 ;
  assign n10271 = ( n2020 & ~n7808 ) | ( n2020 & n9790 ) | ( ~n7808 & n9790 ) ;
  assign n10272 = n10271 ^ n3825 ^ n1712 ;
  assign n10273 = n6570 ^ n4625 ^ n2232 ;
  assign n10274 = n4047 ^ n2246 ^ n1737 ;
  assign n10275 = ( ~n2789 & n4115 ) | ( ~n2789 & n5457 ) | ( n4115 & n5457 ) ;
  assign n10276 = ( n3387 & ~n10274 ) | ( n3387 & n10275 ) | ( ~n10274 & n10275 ) ;
  assign n10277 = n10276 ^ n8771 ^ n901 ;
  assign n10278 = n8843 ^ n8804 ^ n4275 ;
  assign n10279 = n10278 ^ n6767 ^ n770 ;
  assign n10282 = n4328 ^ n3935 ^ n916 ;
  assign n10283 = n10282 ^ n3475 ^ n1517 ;
  assign n10280 = n3636 ^ n1051 ^ n799 ;
  assign n10281 = n10280 ^ n6491 ^ n1736 ;
  assign n10284 = n10283 ^ n10281 ^ n4244 ;
  assign n10285 = ( n2636 & ~n9043 ) | ( n2636 & n9383 ) | ( ~n9043 & n9383 ) ;
  assign n10291 = ( n585 & ~n1595 ) | ( n585 & n5078 ) | ( ~n1595 & n5078 ) ;
  assign n10286 = n4725 ^ n2060 ^ n733 ;
  assign n10287 = n10286 ^ n8797 ^ n3671 ;
  assign n10288 = n7531 ^ n6671 ^ n967 ;
  assign n10289 = ( n1772 & n9545 ) | ( n1772 & ~n10288 ) | ( n9545 & ~n10288 ) ;
  assign n10290 = ( n2354 & n10287 ) | ( n2354 & n10289 ) | ( n10287 & n10289 ) ;
  assign n10292 = n10291 ^ n10290 ^ n8904 ;
  assign n10293 = ( n1973 & ~n3545 ) | ( n1973 & n5321 ) | ( ~n3545 & n5321 ) ;
  assign n10294 = n10293 ^ n8600 ^ n3831 ;
  assign n10295 = n10294 ^ n8827 ^ n685 ;
  assign n10296 = ( n1557 & n3792 ) | ( n1557 & ~n6943 ) | ( n3792 & ~n6943 ) ;
  assign n10297 = ( n2575 & n3047 ) | ( n2575 & n5049 ) | ( n3047 & n5049 ) ;
  assign n10298 = ( ~n4369 & n8322 ) | ( ~n4369 & n10297 ) | ( n8322 & n10297 ) ;
  assign n10299 = ( ~n3974 & n5047 ) | ( ~n3974 & n10298 ) | ( n5047 & n10298 ) ;
  assign n10300 = ( ~n388 & n6023 ) | ( ~n388 & n6959 ) | ( n6023 & n6959 ) ;
  assign n10301 = ( n3508 & ~n9135 ) | ( n3508 & n10300 ) | ( ~n9135 & n10300 ) ;
  assign n10302 = n10301 ^ n6820 ^ n1892 ;
  assign n10303 = n10302 ^ n8577 ^ n2883 ;
  assign n10315 = ( n2246 & n4731 ) | ( n2246 & ~n9418 ) | ( n4731 & ~n9418 ) ;
  assign n10312 = n4211 ^ n3618 ^ n261 ;
  assign n10304 = ( ~n1609 & n2091 ) | ( ~n1609 & n2281 ) | ( n2091 & n2281 ) ;
  assign n10305 = ( n1935 & n9185 ) | ( n1935 & n10304 ) | ( n9185 & n10304 ) ;
  assign n10308 = ( n1199 & n3401 ) | ( n1199 & n5381 ) | ( n3401 & n5381 ) ;
  assign n10307 = n9965 ^ n9160 ^ n758 ;
  assign n10306 = ( ~n3609 & n5363 ) | ( ~n3609 & n6360 ) | ( n5363 & n6360 ) ;
  assign n10309 = n10308 ^ n10307 ^ n10306 ;
  assign n10310 = n10309 ^ n5298 ^ n2541 ;
  assign n10311 = ( x12 & ~n10305 ) | ( x12 & n10310 ) | ( ~n10305 & n10310 ) ;
  assign n10313 = n10312 ^ n10311 ^ n2744 ;
  assign n10314 = ( ~n244 & n8463 ) | ( ~n244 & n10313 ) | ( n8463 & n10313 ) ;
  assign n10316 = n10315 ^ n10314 ^ n7646 ;
  assign n10317 = ( n5352 & n8634 ) | ( n5352 & n10316 ) | ( n8634 & n10316 ) ;
  assign n10318 = n3592 ^ n2871 ^ n1103 ;
  assign n10319 = n10318 ^ n8597 ^ n4890 ;
  assign n10320 = ( ~n2636 & n4322 ) | ( ~n2636 & n5451 ) | ( n4322 & n5451 ) ;
  assign n10321 = ( n6882 & n10319 ) | ( n6882 & ~n10320 ) | ( n10319 & ~n10320 ) ;
  assign n10322 = ( n3030 & n9787 ) | ( n3030 & ~n10321 ) | ( n9787 & ~n10321 ) ;
  assign n10323 = n7294 ^ n3763 ^ n3487 ;
  assign n10324 = n3231 ^ n2373 ^ n541 ;
  assign n10325 = ( n4778 & n8127 ) | ( n4778 & ~n10324 ) | ( n8127 & ~n10324 ) ;
  assign n10332 = n7928 ^ n3798 ^ n3597 ;
  assign n10331 = n6081 ^ n5005 ^ n1739 ;
  assign n10326 = ( ~n3702 & n4045 ) | ( ~n3702 & n5763 ) | ( n4045 & n5763 ) ;
  assign n10327 = ( n5253 & n7065 ) | ( n5253 & n10326 ) | ( n7065 & n10326 ) ;
  assign n10328 = ( ~n5690 & n9218 ) | ( ~n5690 & n10327 ) | ( n9218 & n10327 ) ;
  assign n10329 = ( n2694 & n7905 ) | ( n2694 & n10328 ) | ( n7905 & n10328 ) ;
  assign n10330 = ( n2620 & n3894 ) | ( n2620 & ~n10329 ) | ( n3894 & ~n10329 ) ;
  assign n10333 = n10332 ^ n10331 ^ n10330 ;
  assign n10334 = ( n329 & ~n2434 ) | ( n329 & n4622 ) | ( ~n2434 & n4622 ) ;
  assign n10335 = ( n2844 & n9876 ) | ( n2844 & ~n10334 ) | ( n9876 & ~n10334 ) ;
  assign n10336 = ( n1760 & ~n2228 ) | ( n1760 & n4740 ) | ( ~n2228 & n4740 ) ;
  assign n10337 = ( n716 & n2845 ) | ( n716 & n10336 ) | ( n2845 & n10336 ) ;
  assign n10338 = ( n3588 & n3903 ) | ( n3588 & n8476 ) | ( n3903 & n8476 ) ;
  assign n10339 = n1946 ^ n1760 ^ n272 ;
  assign n10340 = n3332 ^ n2317 ^ n260 ;
  assign n10341 = n10340 ^ n4633 ^ n2486 ;
  assign n10342 = ( n3426 & n10339 ) | ( n3426 & ~n10341 ) | ( n10339 & ~n10341 ) ;
  assign n10343 = ( n10337 & n10338 ) | ( n10337 & ~n10342 ) | ( n10338 & ~n10342 ) ;
  assign n10344 = n9579 ^ n8136 ^ n2574 ;
  assign n10345 = n4862 ^ n2595 ^ n2088 ;
  assign n10346 = n7600 ^ n4588 ^ n2477 ;
  assign n10347 = ( n1733 & ~n2340 ) | ( n1733 & n10346 ) | ( ~n2340 & n10346 ) ;
  assign n10348 = n6874 ^ n1175 ^ n869 ;
  assign n10349 = ( n10345 & n10347 ) | ( n10345 & n10348 ) | ( n10347 & n10348 ) ;
  assign n10351 = n550 ^ n430 ^ n359 ;
  assign n10352 = n10351 ^ n1556 ^ n304 ;
  assign n10350 = ( ~n138 & n373 ) | ( ~n138 & n6770 ) | ( n373 & n6770 ) ;
  assign n10353 = n10352 ^ n10350 ^ n6688 ;
  assign n10354 = ( n5089 & n5452 ) | ( n5089 & ~n6557 ) | ( n5452 & ~n6557 ) ;
  assign n10355 = ( n8058 & n10353 ) | ( n8058 & ~n10354 ) | ( n10353 & ~n10354 ) ;
  assign n10356 = ( n9754 & ~n10349 ) | ( n9754 & n10355 ) | ( ~n10349 & n10355 ) ;
  assign n10357 = n9386 ^ n8422 ^ n2454 ;
  assign n10359 = n6643 ^ n2358 ^ n301 ;
  assign n10360 = ( n5727 & n8954 ) | ( n5727 & n10359 ) | ( n8954 & n10359 ) ;
  assign n10358 = ( n2954 & ~n4357 ) | ( n2954 & n8185 ) | ( ~n4357 & n8185 ) ;
  assign n10361 = n10360 ^ n10358 ^ n9496 ;
  assign n10362 = ( x116 & n3088 ) | ( x116 & ~n6728 ) | ( n3088 & ~n6728 ) ;
  assign n10363 = n10362 ^ n9242 ^ n3181 ;
  assign n10364 = ( n748 & ~n2248 ) | ( n748 & n10363 ) | ( ~n2248 & n10363 ) ;
  assign n10365 = ( n561 & n8233 ) | ( n561 & ~n10006 ) | ( n8233 & ~n10006 ) ;
  assign n10366 = n10365 ^ n8842 ^ n5058 ;
  assign n10367 = n9208 ^ n4611 ^ n4592 ;
  assign n10368 = ( ~n765 & n2943 ) | ( ~n765 & n10367 ) | ( n2943 & n10367 ) ;
  assign n10369 = ( n2816 & n8155 ) | ( n2816 & n8664 ) | ( n8155 & n8664 ) ;
  assign n10370 = n10369 ^ n8863 ^ n7334 ;
  assign n10371 = ( ~n4041 & n4843 ) | ( ~n4041 & n10370 ) | ( n4843 & n10370 ) ;
  assign n10372 = ( ~n10366 & n10368 ) | ( ~n10366 & n10371 ) | ( n10368 & n10371 ) ;
  assign n10373 = ( ~n3747 & n4481 ) | ( ~n3747 & n5723 ) | ( n4481 & n5723 ) ;
  assign n10374 = n7264 ^ n5461 ^ n3357 ;
  assign n10375 = ( ~x86 & n5377 ) | ( ~x86 & n10374 ) | ( n5377 & n10374 ) ;
  assign n10376 = n10375 ^ n6570 ^ n471 ;
  assign n10377 = n10376 ^ n8692 ^ n7633 ;
  assign n10378 = ( n449 & n10373 ) | ( n449 & ~n10377 ) | ( n10373 & ~n10377 ) ;
  assign n10379 = n5682 ^ n5053 ^ n4083 ;
  assign n10380 = n7457 ^ n4050 ^ n479 ;
  assign n10381 = n10380 ^ n5743 ^ n2792 ;
  assign n10382 = n8571 ^ n6808 ^ n5722 ;
  assign n10383 = n5520 ^ n2295 ^ n2220 ;
  assign n10384 = n7990 ^ n6515 ^ n6269 ;
  assign n10385 = ( n7933 & n10383 ) | ( n7933 & n10384 ) | ( n10383 & n10384 ) ;
  assign n10386 = ( n274 & ~n1860 ) | ( n274 & n3320 ) | ( ~n1860 & n3320 ) ;
  assign n10393 = n9717 ^ n8253 ^ n423 ;
  assign n10391 = n9545 ^ n4003 ^ n2012 ;
  assign n10387 = ( ~x29 & n701 ) | ( ~x29 & n1231 ) | ( n701 & n1231 ) ;
  assign n10388 = n10387 ^ n3042 ^ n1418 ;
  assign n10389 = n10388 ^ n9967 ^ n1446 ;
  assign n10390 = ( n2195 & n3720 ) | ( n2195 & ~n10389 ) | ( n3720 & ~n10389 ) ;
  assign n10392 = n10391 ^ n10390 ^ n4432 ;
  assign n10394 = n10393 ^ n10392 ^ n4492 ;
  assign n10395 = n3606 ^ n2982 ^ n1491 ;
  assign n10396 = ( n502 & ~n1916 ) | ( n502 & n6391 ) | ( ~n1916 & n6391 ) ;
  assign n10397 = ( n3620 & n4376 ) | ( n3620 & n8131 ) | ( n4376 & n8131 ) ;
  assign n10398 = ( n10395 & n10396 ) | ( n10395 & n10397 ) | ( n10396 & n10397 ) ;
  assign n10399 = ( n2977 & ~n4952 ) | ( n2977 & n10398 ) | ( ~n4952 & n10398 ) ;
  assign n10400 = n9115 ^ n8649 ^ n4348 ;
  assign n10401 = ( n302 & n520 ) | ( n302 & ~n1283 ) | ( n520 & ~n1283 ) ;
  assign n10402 = ( n4206 & ~n8756 ) | ( n4206 & n10401 ) | ( ~n8756 & n10401 ) ;
  assign n10403 = ( n2793 & ~n3094 ) | ( n2793 & n4409 ) | ( ~n3094 & n4409 ) ;
  assign n10404 = ( n1199 & n2214 ) | ( n1199 & ~n10403 ) | ( n2214 & ~n10403 ) ;
  assign n10405 = ( n4795 & ~n10219 ) | ( n4795 & n10404 ) | ( ~n10219 & n10404 ) ;
  assign n10406 = n10405 ^ n7711 ^ n4916 ;
  assign n10407 = ( ~n1605 & n2795 ) | ( ~n1605 & n10406 ) | ( n2795 & n10406 ) ;
  assign n10408 = ( ~n2064 & n4352 ) | ( ~n2064 & n5758 ) | ( n4352 & n5758 ) ;
  assign n10409 = ( ~n4303 & n6777 ) | ( ~n4303 & n10408 ) | ( n6777 & n10408 ) ;
  assign n10410 = n10073 ^ n9315 ^ n544 ;
  assign n10411 = ( n6760 & ~n10409 ) | ( n6760 & n10410 ) | ( ~n10409 & n10410 ) ;
  assign n10412 = ( n7116 & ~n10312 ) | ( n7116 & n10411 ) | ( ~n10312 & n10411 ) ;
  assign n10413 = n10412 ^ n4398 ^ n3683 ;
  assign n10414 = n5005 ^ n4977 ^ n3414 ;
  assign n10415 = ( ~n1359 & n2327 ) | ( ~n1359 & n3740 ) | ( n2327 & n3740 ) ;
  assign n10416 = n5067 ^ n3151 ^ n206 ;
  assign n10417 = ( ~n5659 & n10415 ) | ( ~n5659 & n10416 ) | ( n10415 & n10416 ) ;
  assign n10418 = ( n1782 & n7436 ) | ( n1782 & n10417 ) | ( n7436 & n10417 ) ;
  assign n10419 = n10374 ^ n5689 ^ n2017 ;
  assign n10420 = ( n2617 & n10418 ) | ( n2617 & n10419 ) | ( n10418 & n10419 ) ;
  assign n10422 = n7557 ^ n5732 ^ n791 ;
  assign n10423 = ( n163 & n265 ) | ( n163 & n8282 ) | ( n265 & n8282 ) ;
  assign n10424 = n7541 ^ n3543 ^ n1349 ;
  assign n10425 = n10424 ^ n7712 ^ n7018 ;
  assign n10426 = ( n2843 & ~n5129 ) | ( n2843 & n10425 ) | ( ~n5129 & n10425 ) ;
  assign n10427 = ( n10422 & ~n10423 ) | ( n10422 & n10426 ) | ( ~n10423 & n10426 ) ;
  assign n10421 = n9915 ^ n7253 ^ n2231 ;
  assign n10428 = n10427 ^ n10421 ^ n10240 ;
  assign n10429 = n2594 ^ n1311 ^ n449 ;
  assign n10430 = n8209 ^ n5263 ^ n3882 ;
  assign n10431 = ( n1425 & ~n10429 ) | ( n1425 & n10430 ) | ( ~n10429 & n10430 ) ;
  assign n10432 = ( n4740 & n7904 ) | ( n4740 & ~n8745 ) | ( n7904 & ~n8745 ) ;
  assign n10433 = ( n9401 & n10431 ) | ( n9401 & n10432 ) | ( n10431 & n10432 ) ;
  assign n10434 = ( n1681 & n3345 ) | ( n1681 & n6595 ) | ( n3345 & n6595 ) ;
  assign n10435 = n1199 ^ n953 ^ x61 ;
  assign n10436 = ( ~n10433 & n10434 ) | ( ~n10433 & n10435 ) | ( n10434 & n10435 ) ;
  assign n10437 = n10436 ^ n5492 ^ n2763 ;
  assign n10441 = ( ~n2460 & n5867 ) | ( ~n2460 & n9654 ) | ( n5867 & n9654 ) ;
  assign n10442 = n10441 ^ n9548 ^ n1341 ;
  assign n10438 = ( ~x64 & n3338 ) | ( ~x64 & n4247 ) | ( n3338 & n4247 ) ;
  assign n10439 = n10438 ^ n7663 ^ n697 ;
  assign n10440 = ( n3904 & n8697 ) | ( n3904 & ~n10439 ) | ( n8697 & ~n10439 ) ;
  assign n10443 = n10442 ^ n10440 ^ n7086 ;
  assign n10446 = n4225 ^ n3797 ^ n2529 ;
  assign n10447 = n10446 ^ n3649 ^ n3609 ;
  assign n10445 = ( n803 & n2916 ) | ( n803 & n7024 ) | ( n2916 & n7024 ) ;
  assign n10444 = ( n2961 & ~n3518 ) | ( n2961 & n8397 ) | ( ~n3518 & n8397 ) ;
  assign n10448 = n10447 ^ n10445 ^ n10444 ;
  assign n10449 = ( n276 & n1993 ) | ( n276 & n7846 ) | ( n1993 & n7846 ) ;
  assign n10450 = ( n1927 & ~n3164 ) | ( n1927 & n9496 ) | ( ~n3164 & n9496 ) ;
  assign n10451 = ( n2935 & ~n7250 ) | ( n2935 & n10450 ) | ( ~n7250 & n10450 ) ;
  assign n10452 = n10451 ^ n9141 ^ n928 ;
  assign n10453 = n10452 ^ n6224 ^ n781 ;
  assign n10454 = ( n1596 & n10449 ) | ( n1596 & ~n10453 ) | ( n10449 & ~n10453 ) ;
  assign n10455 = n8786 ^ n7339 ^ n206 ;
  assign n10456 = ( ~n2234 & n10454 ) | ( ~n2234 & n10455 ) | ( n10454 & n10455 ) ;
  assign n10457 = ( n454 & n1185 ) | ( n454 & ~n7299 ) | ( n1185 & ~n7299 ) ;
  assign n10458 = n10457 ^ n3810 ^ n1753 ;
  assign n10459 = n5590 ^ n1577 ^ n631 ;
  assign n10460 = ( n6237 & n10458 ) | ( n6237 & n10459 ) | ( n10458 & n10459 ) ;
  assign n10461 = n7352 ^ n3795 ^ n963 ;
  assign n10462 = ( n2669 & n5426 ) | ( n2669 & ~n10461 ) | ( n5426 & ~n10461 ) ;
  assign n10478 = n5830 ^ n2532 ^ n1848 ;
  assign n10479 = ( n1354 & n5958 ) | ( n1354 & ~n10478 ) | ( n5958 & ~n10478 ) ;
  assign n10464 = ( ~n897 & n5097 ) | ( ~n897 & n10268 ) | ( n5097 & n10268 ) ;
  assign n10463 = ( n511 & ~n3724 ) | ( n511 & n7229 ) | ( ~n3724 & n7229 ) ;
  assign n10465 = n10464 ^ n10463 ^ n8216 ;
  assign n10466 = n10465 ^ n4944 ^ n1809 ;
  assign n10467 = ( ~n4717 & n7723 ) | ( ~n4717 & n10466 ) | ( n7723 & n10466 ) ;
  assign n10474 = n1761 ^ n1620 ^ n418 ;
  assign n10475 = n10474 ^ n9299 ^ n1608 ;
  assign n10472 = n2519 ^ n2327 ^ n1468 ;
  assign n10470 = ( n1426 & n2975 ) | ( n1426 & n3845 ) | ( n2975 & n3845 ) ;
  assign n10471 = ( ~n482 & n1301 ) | ( ~n482 & n10470 ) | ( n1301 & n10470 ) ;
  assign n10468 = ( n4871 & n8680 ) | ( n4871 & ~n9674 ) | ( n8680 & ~n9674 ) ;
  assign n10469 = n10468 ^ n10373 ^ n5004 ;
  assign n10473 = n10472 ^ n10471 ^ n10469 ;
  assign n10476 = n10475 ^ n10473 ^ n7411 ;
  assign n10477 = ( n2960 & n10467 ) | ( n2960 & ~n10476 ) | ( n10467 & ~n10476 ) ;
  assign n10480 = n10479 ^ n10477 ^ n9928 ;
  assign n10481 = ( n6115 & n10462 ) | ( n6115 & ~n10480 ) | ( n10462 & ~n10480 ) ;
  assign n10486 = ( n353 & n3108 ) | ( n353 & ~n3800 ) | ( n3108 & ~n3800 ) ;
  assign n10484 = ( n1653 & n2409 ) | ( n1653 & ~n4297 ) | ( n2409 & ~n4297 ) ;
  assign n10482 = ( n938 & n1386 ) | ( n938 & ~n2688 ) | ( n1386 & ~n2688 ) ;
  assign n10483 = ( n2555 & n4071 ) | ( n2555 & n10482 ) | ( n4071 & n10482 ) ;
  assign n10485 = n10484 ^ n10483 ^ n3729 ;
  assign n10487 = n10486 ^ n10485 ^ n2028 ;
  assign n10489 = ( n1581 & ~n1951 ) | ( n1581 & n3126 ) | ( ~n1951 & n3126 ) ;
  assign n10488 = ( ~x35 & n2106 ) | ( ~x35 & n10114 ) | ( n2106 & n10114 ) ;
  assign n10490 = n10489 ^ n10488 ^ n9506 ;
  assign n10491 = ( ~n1289 & n3294 ) | ( ~n1289 & n5913 ) | ( n3294 & n5913 ) ;
  assign n10492 = n10491 ^ n3054 ^ n2466 ;
  assign n10493 = n10492 ^ n3434 ^ n1732 ;
  assign n10494 = n6659 ^ n4186 ^ n3555 ;
  assign n10497 = ( n1593 & n6555 ) | ( n1593 & ~n10130 ) | ( n6555 & ~n10130 ) ;
  assign n10495 = ( n2410 & ~n3714 ) | ( n2410 & n8402 ) | ( ~n3714 & n8402 ) ;
  assign n10496 = ( n463 & n662 ) | ( n463 & n10495 ) | ( n662 & n10495 ) ;
  assign n10498 = n10497 ^ n10496 ^ n883 ;
  assign n10499 = n9773 ^ n9707 ^ n6305 ;
  assign n10501 = n9093 ^ n9005 ^ n4224 ;
  assign n10500 = ( n3942 & n8080 ) | ( n3942 & n9679 ) | ( n8080 & n9679 ) ;
  assign n10502 = n10501 ^ n10500 ^ n4070 ;
  assign n10503 = ( n10498 & ~n10499 ) | ( n10498 & n10502 ) | ( ~n10499 & n10502 ) ;
  assign n10508 = n6291 ^ n5943 ^ n3421 ;
  assign n10504 = ( n154 & ~n5023 ) | ( n154 & n5132 ) | ( ~n5023 & n5132 ) ;
  assign n10505 = ( ~n398 & n1214 ) | ( ~n398 & n3924 ) | ( n1214 & n3924 ) ;
  assign n10506 = ( n4499 & n10504 ) | ( n4499 & ~n10505 ) | ( n10504 & ~n10505 ) ;
  assign n10507 = n10506 ^ n3229 ^ n2202 ;
  assign n10509 = n10508 ^ n10507 ^ n10398 ;
  assign n10510 = ( x67 & n4513 ) | ( x67 & n4635 ) | ( n4513 & n4635 ) ;
  assign n10513 = n6453 ^ n4789 ^ n4217 ;
  assign n10511 = n8638 ^ n8088 ^ n7908 ;
  assign n10512 = ( ~n408 & n6092 ) | ( ~n408 & n10511 ) | ( n6092 & n10511 ) ;
  assign n10514 = n10513 ^ n10512 ^ n5895 ;
  assign n10515 = ( n221 & n3466 ) | ( n221 & n4085 ) | ( n3466 & n4085 ) ;
  assign n10516 = ( n5116 & ~n6488 ) | ( n5116 & n9764 ) | ( ~n6488 & n9764 ) ;
  assign n10517 = n10516 ^ n10383 ^ n4950 ;
  assign n10518 = n10517 ^ n4591 ^ n3100 ;
  assign n10519 = ( n4690 & n10515 ) | ( n4690 & ~n10518 ) | ( n10515 & ~n10518 ) ;
  assign n10520 = n10519 ^ n9332 ^ n1525 ;
  assign n10521 = n5399 ^ n3511 ^ n144 ;
  assign n10522 = n3711 ^ n2499 ^ n322 ;
  assign n10523 = n10522 ^ n8001 ^ n6363 ;
  assign n10524 = ( n9688 & ~n10521 ) | ( n9688 & n10523 ) | ( ~n10521 & n10523 ) ;
  assign n10525 = n1690 ^ n1459 ^ n1150 ;
  assign n10526 = ( n922 & n3602 ) | ( n922 & n10525 ) | ( n3602 & n10525 ) ;
  assign n10527 = ( n5100 & n5668 ) | ( n5100 & ~n10526 ) | ( n5668 & ~n10526 ) ;
  assign n10528 = ( n869 & n1302 ) | ( n869 & n1374 ) | ( n1302 & n1374 ) ;
  assign n10529 = n9932 ^ n7588 ^ n863 ;
  assign n10530 = ( n1366 & n10528 ) | ( n1366 & n10529 ) | ( n10528 & n10529 ) ;
  assign n10531 = n8115 ^ n5404 ^ n2705 ;
  assign n10532 = ( n3408 & ~n5263 ) | ( n3408 & n10531 ) | ( ~n5263 & n10531 ) ;
  assign n10533 = ( n1442 & n3651 ) | ( n1442 & n8042 ) | ( n3651 & n8042 ) ;
  assign n10534 = ( x116 & n10532 ) | ( x116 & ~n10533 ) | ( n10532 & ~n10533 ) ;
  assign n10535 = n10534 ^ n9771 ^ n6269 ;
  assign n10536 = n9078 ^ n8460 ^ n7688 ;
  assign n10537 = ( ~n1971 & n2703 ) | ( ~n1971 & n2954 ) | ( n2703 & n2954 ) ;
  assign n10538 = ( ~n7891 & n8582 ) | ( ~n7891 & n10537 ) | ( n8582 & n10537 ) ;
  assign n10539 = ( ~n2663 & n3042 ) | ( ~n2663 & n3621 ) | ( n3042 & n3621 ) ;
  assign n10540 = n10539 ^ n8561 ^ n4669 ;
  assign n10541 = ( n3185 & ~n6850 ) | ( n3185 & n7436 ) | ( ~n6850 & n7436 ) ;
  assign n10542 = ( n5274 & n6275 ) | ( n5274 & ~n10541 ) | ( n6275 & ~n10541 ) ;
  assign n10543 = ( n1620 & n5273 ) | ( n1620 & ~n8955 ) | ( n5273 & ~n8955 ) ;
  assign n10544 = n10543 ^ n3941 ^ n2262 ;
  assign n10545 = n7671 ^ n3184 ^ n515 ;
  assign n10547 = n8225 ^ n2924 ^ n2797 ;
  assign n10548 = n10547 ^ n4551 ^ n2333 ;
  assign n10546 = ( n584 & n3678 ) | ( n584 & n5974 ) | ( n3678 & n5974 ) ;
  assign n10549 = n10548 ^ n10546 ^ n1491 ;
  assign n10561 = n6600 ^ n2216 ^ n2206 ;
  assign n10562 = ( n2647 & ~n4450 ) | ( n2647 & n10561 ) | ( ~n4450 & n10561 ) ;
  assign n10559 = n4604 ^ n827 ^ n214 ;
  assign n10558 = ( n327 & ~n6953 ) | ( n327 & n7276 ) | ( ~n6953 & n7276 ) ;
  assign n10556 = ( n1892 & n5319 ) | ( n1892 & n6163 ) | ( n5319 & n6163 ) ;
  assign n10554 = n8953 ^ n3209 ^ n1513 ;
  assign n10551 = ( ~n698 & n738 ) | ( ~n698 & n1402 ) | ( n738 & n1402 ) ;
  assign n10552 = ( n573 & ~n6534 ) | ( n573 & n10551 ) | ( ~n6534 & n10551 ) ;
  assign n10550 = n4679 ^ n4043 ^ n2691 ;
  assign n10553 = n10552 ^ n10550 ^ n160 ;
  assign n10555 = n10554 ^ n10553 ^ n7475 ;
  assign n10557 = n10556 ^ n10555 ^ n3138 ;
  assign n10560 = n10559 ^ n10558 ^ n10557 ;
  assign n10563 = n10562 ^ n10560 ^ n1931 ;
  assign n10564 = ( n10545 & ~n10549 ) | ( n10545 & n10563 ) | ( ~n10549 & n10563 ) ;
  assign n10565 = ( n2137 & n2917 ) | ( n2137 & n6961 ) | ( n2917 & n6961 ) ;
  assign n10566 = n7897 ^ n3732 ^ n3586 ;
  assign n10567 = n10566 ^ n7692 ^ n5691 ;
  assign n10568 = ( n1443 & n2540 ) | ( n1443 & n10567 ) | ( n2540 & n10567 ) ;
  assign n10569 = ( ~n3297 & n4407 ) | ( ~n3297 & n6676 ) | ( n4407 & n6676 ) ;
  assign n10574 = ( n4585 & ~n5844 ) | ( n4585 & n6224 ) | ( ~n5844 & n6224 ) ;
  assign n10570 = n4858 ^ n4615 ^ n2345 ;
  assign n10571 = ( n1291 & ~n1441 ) | ( n1291 & n4517 ) | ( ~n1441 & n4517 ) ;
  assign n10572 = n10571 ^ n4260 ^ n1226 ;
  assign n10573 = ( n470 & ~n10570 ) | ( n470 & n10572 ) | ( ~n10570 & n10572 ) ;
  assign n10575 = n10574 ^ n10573 ^ n3643 ;
  assign n10576 = ( n6941 & n10569 ) | ( n6941 & ~n10575 ) | ( n10569 & ~n10575 ) ;
  assign n10577 = n10550 ^ n9461 ^ n416 ;
  assign n10583 = n8636 ^ n7264 ^ n2218 ;
  assign n10584 = n10583 ^ n7846 ^ n2050 ;
  assign n10581 = n6360 ^ n5086 ^ n3112 ;
  assign n10579 = ( x14 & n3196 ) | ( x14 & ~n5347 ) | ( n3196 & ~n5347 ) ;
  assign n10578 = n8926 ^ n5136 ^ n1413 ;
  assign n10580 = n10579 ^ n10578 ^ n661 ;
  assign n10582 = n10581 ^ n10580 ^ n5482 ;
  assign n10585 = n10584 ^ n10582 ^ n1604 ;
  assign n10591 = ( ~n4369 & n4672 ) | ( ~n4369 & n8560 ) | ( n4672 & n8560 ) ;
  assign n10588 = n3767 ^ n358 ^ n307 ;
  assign n10589 = ( ~n287 & n1982 ) | ( ~n287 & n10588 ) | ( n1982 & n10588 ) ;
  assign n10587 = n8402 ^ n8154 ^ n561 ;
  assign n10590 = n10589 ^ n10587 ^ n2437 ;
  assign n10586 = ( n6502 & ~n7648 ) | ( n6502 & n7727 ) | ( ~n7648 & n7727 ) ;
  assign n10592 = n10591 ^ n10590 ^ n10586 ;
  assign n10593 = n7414 ^ n4932 ^ n2344 ;
  assign n10594 = n1359 ^ n1353 ^ n1310 ;
  assign n10595 = ( n2047 & ~n7282 ) | ( n2047 & n10594 ) | ( ~n7282 & n10594 ) ;
  assign n10596 = n4517 ^ n4500 ^ n2898 ;
  assign n10597 = n10424 ^ n5708 ^ n3354 ;
  assign n10598 = ( ~n4729 & n10596 ) | ( ~n4729 & n10597 ) | ( n10596 & n10597 ) ;
  assign n10599 = ( n3039 & n6944 ) | ( n3039 & ~n10598 ) | ( n6944 & ~n10598 ) ;
  assign n10600 = ( n8868 & n10222 ) | ( n8868 & n10599 ) | ( n10222 & n10599 ) ;
  assign n10602 = n5409 ^ n3694 ^ n1536 ;
  assign n10603 = n10602 ^ n7904 ^ n284 ;
  assign n10601 = n8370 ^ n2069 ^ n1740 ;
  assign n10604 = n10603 ^ n10601 ^ n3451 ;
  assign n10605 = ( ~n284 & n2157 ) | ( ~n284 & n2300 ) | ( n2157 & n2300 ) ;
  assign n10607 = n8310 ^ n4816 ^ n3014 ;
  assign n10606 = ( ~n1915 & n4294 ) | ( ~n1915 & n10332 ) | ( n4294 & n10332 ) ;
  assign n10608 = n10607 ^ n10606 ^ n5753 ;
  assign n10609 = n10608 ^ n4749 ^ n3973 ;
  assign n10610 = ( ~n9958 & n10605 ) | ( ~n9958 & n10609 ) | ( n10605 & n10609 ) ;
  assign n10611 = n7982 ^ n5808 ^ n4699 ;
  assign n10612 = n10611 ^ n7608 ^ n1100 ;
  assign n10615 = ( n209 & n2883 ) | ( n209 & ~n3794 ) | ( n2883 & ~n3794 ) ;
  assign n10613 = n6743 ^ n3728 ^ n3276 ;
  assign n10614 = ( n3417 & n6618 ) | ( n3417 & n10613 ) | ( n6618 & n10613 ) ;
  assign n10616 = n10615 ^ n10614 ^ n3341 ;
  assign n10617 = n9163 ^ n4908 ^ n537 ;
  assign n10620 = ( n887 & ~n1758 ) | ( n887 & n10201 ) | ( ~n1758 & n10201 ) ;
  assign n10621 = n10620 ^ n3812 ^ n318 ;
  assign n10618 = n3344 ^ n2513 ^ n1975 ;
  assign n10619 = n10618 ^ n1143 ^ n749 ;
  assign n10622 = n10621 ^ n10619 ^ n10134 ;
  assign n10623 = n10622 ^ n7736 ^ n1831 ;
  assign n10624 = n10623 ^ n10397 ^ n5855 ;
  assign n10625 = ( n2256 & n10617 ) | ( n2256 & ~n10624 ) | ( n10617 & ~n10624 ) ;
  assign n10635 = n6164 ^ n4563 ^ n3524 ;
  assign n10636 = n10635 ^ n7687 ^ n5378 ;
  assign n10626 = n4249 ^ n3283 ^ n2221 ;
  assign n10627 = ( n1644 & ~n2081 ) | ( n1644 & n10626 ) | ( ~n2081 & n10626 ) ;
  assign n10628 = ( n6238 & n8745 ) | ( n6238 & ~n10627 ) | ( n8745 & ~n10627 ) ;
  assign n10629 = n10628 ^ n5737 ^ n2767 ;
  assign n10632 = n8226 ^ n5293 ^ n953 ;
  assign n10630 = ( n2582 & n2583 ) | ( n2582 & ~n5927 ) | ( n2583 & ~n5927 ) ;
  assign n10631 = ( n599 & n4752 ) | ( n599 & n10630 ) | ( n4752 & n10630 ) ;
  assign n10633 = n10632 ^ n10631 ^ n8545 ;
  assign n10634 = ( n6117 & n10629 ) | ( n6117 & ~n10633 ) | ( n10629 & ~n10633 ) ;
  assign n10637 = n10636 ^ n10634 ^ n7809 ;
  assign n10640 = n6513 ^ n4537 ^ n1245 ;
  assign n10641 = ( n2604 & n9833 ) | ( n2604 & ~n10640 ) | ( n9833 & ~n10640 ) ;
  assign n10638 = n8453 ^ n4764 ^ n1193 ;
  assign n10639 = ( ~n2232 & n2322 ) | ( ~n2232 & n10638 ) | ( n2322 & n10638 ) ;
  assign n10642 = n10641 ^ n10639 ^ n1380 ;
  assign n10643 = ( ~n4590 & n5119 ) | ( ~n4590 & n8517 ) | ( n5119 & n8517 ) ;
  assign n10644 = ( n2311 & n2750 ) | ( n2311 & n10643 ) | ( n2750 & n10643 ) ;
  assign n10645 = ( n4831 & ~n8747 ) | ( n4831 & n10644 ) | ( ~n8747 & n10644 ) ;
  assign n10646 = ( n1284 & ~n2681 ) | ( n1284 & n10645 ) | ( ~n2681 & n10645 ) ;
  assign n10647 = n6848 ^ n3925 ^ n1254 ;
  assign n10648 = ( n1566 & n5803 ) | ( n1566 & n6168 ) | ( n5803 & n6168 ) ;
  assign n10649 = ( n4909 & ~n6833 ) | ( n4909 & n10648 ) | ( ~n6833 & n10648 ) ;
  assign n10650 = ( n1820 & ~n4858 ) | ( n1820 & n5260 ) | ( ~n4858 & n5260 ) ;
  assign n10651 = n10650 ^ n8330 ^ n1031 ;
  assign n10652 = ( n3973 & n5222 ) | ( n3973 & n10651 ) | ( n5222 & n10651 ) ;
  assign n10653 = n10652 ^ n9910 ^ n3378 ;
  assign n10654 = ( n10647 & n10649 ) | ( n10647 & n10653 ) | ( n10649 & n10653 ) ;
  assign n10655 = n10654 ^ n10360 ^ n7990 ;
  assign n10656 = n10655 ^ n6636 ^ n4910 ;
  assign n10657 = ( n5390 & ~n5515 ) | ( n5390 & n6752 ) | ( ~n5515 & n6752 ) ;
  assign n10658 = ( n3515 & n6463 ) | ( n3515 & n6617 ) | ( n6463 & n6617 ) ;
  assign n10660 = n5440 ^ n1966 ^ n1537 ;
  assign n10659 = ( n832 & ~n1481 ) | ( n832 & n3264 ) | ( ~n1481 & n3264 ) ;
  assign n10661 = n10660 ^ n10659 ^ n2964 ;
  assign n10662 = ( ~x107 & n1350 ) | ( ~x107 & n6069 ) | ( n1350 & n6069 ) ;
  assign n10663 = ( n405 & n2067 ) | ( n405 & n10662 ) | ( n2067 & n10662 ) ;
  assign n10664 = ( n9986 & n10661 ) | ( n9986 & n10663 ) | ( n10661 & n10663 ) ;
  assign n10665 = ( ~x112 & n5719 ) | ( ~x112 & n10664 ) | ( n5719 & n10664 ) ;
  assign n10666 = n10665 ^ n8502 ^ n5570 ;
  assign n10667 = ( n3876 & ~n10658 ) | ( n3876 & n10666 ) | ( ~n10658 & n10666 ) ;
  assign n10670 = ( n371 & n2571 ) | ( n371 & ~n3775 ) | ( n2571 & ~n3775 ) ;
  assign n10668 = n8807 ^ n8257 ^ n6218 ;
  assign n10669 = ( n6276 & n7297 ) | ( n6276 & n10668 ) | ( n7297 & n10668 ) ;
  assign n10671 = n10670 ^ n10669 ^ n10134 ;
  assign n10672 = ( n10657 & n10667 ) | ( n10657 & n10671 ) | ( n10667 & n10671 ) ;
  assign n10673 = ( ~n1060 & n2141 ) | ( ~n1060 & n2765 ) | ( n2141 & n2765 ) ;
  assign n10674 = n10673 ^ n4831 ^ n3819 ;
  assign n10675 = n10674 ^ n9638 ^ n281 ;
  assign n10679 = n2867 ^ n501 ^ n171 ;
  assign n10680 = ( ~n6445 & n10406 ) | ( ~n6445 & n10679 ) | ( n10406 & n10679 ) ;
  assign n10676 = ( n1533 & ~n1924 ) | ( n1533 & n2913 ) | ( ~n1924 & n2913 ) ;
  assign n10677 = n10676 ^ n1612 ^ n1024 ;
  assign n10678 = n10677 ^ n975 ^ n440 ;
  assign n10681 = n10680 ^ n10678 ^ n4440 ;
  assign n10685 = ( n632 & n1279 ) | ( n632 & n2075 ) | ( n1279 & n2075 ) ;
  assign n10684 = n4510 ^ n2638 ^ n438 ;
  assign n10682 = n3856 ^ n3648 ^ n663 ;
  assign n10683 = ( n1841 & n5041 ) | ( n1841 & ~n10682 ) | ( n5041 & ~n10682 ) ;
  assign n10686 = n10685 ^ n10684 ^ n10683 ;
  assign n10687 = ( n3435 & n4856 ) | ( n3435 & n5129 ) | ( n4856 & n5129 ) ;
  assign n10688 = ( ~n2718 & n4284 ) | ( ~n2718 & n10687 ) | ( n4284 & n10687 ) ;
  assign n10689 = ( n4804 & n8105 ) | ( n4804 & n10688 ) | ( n8105 & n10688 ) ;
  assign n10693 = n7358 ^ n5690 ^ n1592 ;
  assign n10694 = n10693 ^ n9637 ^ n1380 ;
  assign n10695 = n10694 ^ n3963 ^ n234 ;
  assign n10691 = n5246 ^ n628 ^ n367 ;
  assign n10690 = n5608 ^ n1017 ^ n980 ;
  assign n10692 = n10691 ^ n10690 ^ n7146 ;
  assign n10696 = n10695 ^ n10692 ^ n4410 ;
  assign n10697 = ( ~n1844 & n4724 ) | ( ~n1844 & n4773 ) | ( n4724 & n4773 ) ;
  assign n10698 = n5049 ^ n4103 ^ n1960 ;
  assign n10699 = ( n990 & n10697 ) | ( n990 & ~n10698 ) | ( n10697 & ~n10698 ) ;
  assign n10700 = n9315 ^ n1205 ^ n1044 ;
  assign n10701 = ( n6428 & n10699 ) | ( n6428 & ~n10700 ) | ( n10699 & ~n10700 ) ;
  assign n10702 = ( n5603 & n10696 ) | ( n5603 & ~n10701 ) | ( n10696 & ~n10701 ) ;
  assign n10703 = ( n5859 & ~n7253 ) | ( n5859 & n8622 ) | ( ~n7253 & n8622 ) ;
  assign n10704 = ( n3101 & n3520 ) | ( n3101 & ~n3626 ) | ( n3520 & ~n3626 ) ;
  assign n10705 = n10704 ^ n960 ^ n321 ;
  assign n10710 = ( n1795 & ~n2622 ) | ( n1795 & n10014 ) | ( ~n2622 & n10014 ) ;
  assign n10707 = ( ~n809 & n1299 ) | ( ~n809 & n2480 ) | ( n1299 & n2480 ) ;
  assign n10706 = ( n377 & ~n9029 ) | ( n377 & n10151 ) | ( ~n9029 & n10151 ) ;
  assign n10708 = n10707 ^ n10706 ^ n375 ;
  assign n10709 = ( n1214 & n9315 ) | ( n1214 & ~n10708 ) | ( n9315 & ~n10708 ) ;
  assign n10711 = n10710 ^ n10709 ^ n1909 ;
  assign n10716 = n8038 ^ n6758 ^ n579 ;
  assign n10712 = n1136 ^ n988 ^ n891 ;
  assign n10713 = ( n8586 & n8922 ) | ( n8586 & ~n10712 ) | ( n8922 & ~n10712 ) ;
  assign n10714 = n10713 ^ n10106 ^ n7683 ;
  assign n10715 = ( x58 & ~n2831 ) | ( x58 & n10714 ) | ( ~n2831 & n10714 ) ;
  assign n10717 = n10716 ^ n10715 ^ n4464 ;
  assign n10718 = n10717 ^ n6098 ^ n2588 ;
  assign n10720 = ( ~n1911 & n2437 ) | ( ~n1911 & n5864 ) | ( n2437 & n5864 ) ;
  assign n10719 = n4874 ^ n4236 ^ n1070 ;
  assign n10721 = n10720 ^ n10719 ^ n5415 ;
  assign n10722 = n10721 ^ n10358 ^ n3380 ;
  assign n10727 = ( n2458 & ~n4699 ) | ( n2458 & n6648 ) | ( ~n4699 & n6648 ) ;
  assign n10728 = n10727 ^ n10504 ^ n5788 ;
  assign n10723 = n5462 ^ n1266 ^ x21 ;
  assign n10724 = n6743 ^ n2432 ^ n948 ;
  assign n10725 = n10724 ^ n10628 ^ n3897 ;
  assign n10726 = ( n6450 & ~n10723 ) | ( n6450 & n10725 ) | ( ~n10723 & n10725 ) ;
  assign n10729 = n10728 ^ n10726 ^ n3742 ;
  assign n10730 = ( n4424 & ~n5223 ) | ( n4424 & n6111 ) | ( ~n5223 & n6111 ) ;
  assign n10731 = n4024 ^ n2748 ^ n1644 ;
  assign n10732 = n10731 ^ n8354 ^ n6238 ;
  assign n10733 = ( ~x36 & n2645 ) | ( ~x36 & n10732 ) | ( n2645 & n10732 ) ;
  assign n10744 = ( ~n4555 & n5712 ) | ( ~n4555 & n8290 ) | ( n5712 & n8290 ) ;
  assign n10742 = n7076 ^ n3537 ^ n3442 ;
  assign n10743 = n10742 ^ n7188 ^ n5280 ;
  assign n10745 = n10744 ^ n10743 ^ n4562 ;
  assign n10739 = ( n2642 & ~n5708 ) | ( n2642 & n9733 ) | ( ~n5708 & n9733 ) ;
  assign n10740 = ( n862 & ~n3071 ) | ( n862 & n10739 ) | ( ~n3071 & n10739 ) ;
  assign n10734 = ( n1831 & ~n3126 ) | ( n1831 & n9621 ) | ( ~n3126 & n9621 ) ;
  assign n10735 = ( n4010 & n6924 ) | ( n4010 & ~n6928 ) | ( n6924 & ~n6928 ) ;
  assign n10736 = ( n9325 & n10734 ) | ( n9325 & ~n10735 ) | ( n10734 & ~n10735 ) ;
  assign n10737 = ( ~n4629 & n7808 ) | ( ~n4629 & n10736 ) | ( n7808 & n10736 ) ;
  assign n10738 = ( n9660 & ~n9704 ) | ( n9660 & n10737 ) | ( ~n9704 & n10737 ) ;
  assign n10741 = n10740 ^ n10738 ^ n7118 ;
  assign n10746 = n10745 ^ n10741 ^ n740 ;
  assign n10747 = ( n2701 & n2912 ) | ( n2701 & ~n4295 ) | ( n2912 & ~n4295 ) ;
  assign n10748 = ( n1835 & n2042 ) | ( n1835 & ~n10747 ) | ( n2042 & ~n10747 ) ;
  assign n10749 = n8643 ^ n3591 ^ n3217 ;
  assign n10750 = n10749 ^ n6753 ^ n723 ;
  assign n10751 = n10750 ^ n5747 ^ n2614 ;
  assign n10752 = n10618 ^ n3050 ^ n677 ;
  assign n10756 = ( ~n3679 & n3879 ) | ( ~n3679 & n6865 ) | ( n3879 & n6865 ) ;
  assign n10754 = ( ~n1383 & n1805 ) | ( ~n1383 & n2835 ) | ( n1805 & n2835 ) ;
  assign n10755 = n10754 ^ n6994 ^ n3113 ;
  assign n10753 = n2330 ^ n898 ^ n187 ;
  assign n10757 = n10756 ^ n10755 ^ n10753 ;
  assign n10759 = n6114 ^ n2828 ^ n1442 ;
  assign n10760 = ( n4379 & n5078 ) | ( n4379 & n10759 ) | ( n5078 & n10759 ) ;
  assign n10758 = n5220 ^ n4086 ^ n2651 ;
  assign n10761 = n10760 ^ n10758 ^ n6160 ;
  assign n10765 = n10266 ^ n3029 ^ n1265 ;
  assign n10762 = n5160 ^ n4000 ^ n2111 ;
  assign n10763 = ( n845 & n2889 ) | ( n845 & ~n10762 ) | ( n2889 & ~n10762 ) ;
  assign n10764 = n10763 ^ n10025 ^ n1641 ;
  assign n10766 = n10765 ^ n10764 ^ n6543 ;
  assign n10767 = ( n984 & n6245 ) | ( n984 & ~n9955 ) | ( n6245 & ~n9955 ) ;
  assign n10769 = ( n162 & n2879 ) | ( n162 & ~n9220 ) | ( n2879 & ~n9220 ) ;
  assign n10768 = n8981 ^ n7955 ^ n402 ;
  assign n10770 = n10769 ^ n10768 ^ n7790 ;
  assign n10773 = ( n6685 & n8320 ) | ( n6685 & n8821 ) | ( n8320 & n8821 ) ;
  assign n10774 = ( ~n6200 & n8537 ) | ( ~n6200 & n10773 ) | ( n8537 & n10773 ) ;
  assign n10775 = ( n3450 & n7615 ) | ( n3450 & n10774 ) | ( n7615 & n10774 ) ;
  assign n10771 = n8734 ^ n1329 ^ n184 ;
  assign n10772 = ( ~n8461 & n10111 ) | ( ~n8461 & n10771 ) | ( n10111 & n10771 ) ;
  assign n10776 = n10775 ^ n10772 ^ n4269 ;
  assign n10781 = n4778 ^ n4432 ^ n3198 ;
  assign n10782 = n10781 ^ n1779 ^ n514 ;
  assign n10783 = n10782 ^ n10212 ^ n3264 ;
  assign n10778 = ( n571 & ~n653 ) | ( n571 & n1698 ) | ( ~n653 & n1698 ) ;
  assign n10779 = ( ~n3385 & n3723 ) | ( ~n3385 & n10778 ) | ( n3723 & n10778 ) ;
  assign n10780 = n10779 ^ n7967 ^ n7275 ;
  assign n10777 = n7060 ^ n6753 ^ n4383 ;
  assign n10784 = n10783 ^ n10780 ^ n10777 ;
  assign n10785 = n6177 ^ n2020 ^ n1552 ;
  assign n10787 = ( n4043 & n4279 ) | ( n4043 & n8060 ) | ( n4279 & n8060 ) ;
  assign n10786 = ( n4300 & n5027 ) | ( n4300 & ~n6819 ) | ( n5027 & ~n6819 ) ;
  assign n10788 = n10787 ^ n10786 ^ n7376 ;
  assign n10789 = ( n692 & n3737 ) | ( n692 & n6892 ) | ( n3737 & n6892 ) ;
  assign n10790 = ( n4367 & ~n8735 ) | ( n4367 & n10789 ) | ( ~n8735 & n10789 ) ;
  assign n10791 = n10790 ^ n4095 ^ n3262 ;
  assign n10792 = n10791 ^ n6592 ^ n3284 ;
  assign n10793 = n8139 ^ n6016 ^ n2017 ;
  assign n10794 = n10793 ^ n8010 ^ n1180 ;
  assign n10795 = n10794 ^ n10040 ^ n2651 ;
  assign n10796 = n10795 ^ n6185 ^ n2597 ;
  assign n10797 = ( ~n3687 & n7065 ) | ( ~n3687 & n10796 ) | ( n7065 & n10796 ) ;
  assign n10798 = ( ~n10788 & n10792 ) | ( ~n10788 & n10797 ) | ( n10792 & n10797 ) ;
  assign n10799 = ( ~n1264 & n2615 ) | ( ~n1264 & n10103 ) | ( n2615 & n10103 ) ;
  assign n10804 = n7370 ^ n6656 ^ n4461 ;
  assign n10802 = n9509 ^ n8928 ^ n3377 ;
  assign n10800 = ( n4779 & n6287 ) | ( n4779 & ~n7371 ) | ( n6287 & ~n7371 ) ;
  assign n10801 = ( n4450 & n8318 ) | ( n4450 & n10800 ) | ( n8318 & n10800 ) ;
  assign n10803 = n10802 ^ n10801 ^ n3285 ;
  assign n10805 = n10804 ^ n10803 ^ n10238 ;
  assign n10809 = ( n2067 & ~n3924 ) | ( n2067 & n5254 ) | ( ~n3924 & n5254 ) ;
  assign n10810 = ( n5873 & n6652 ) | ( n5873 & ~n10809 ) | ( n6652 & ~n10809 ) ;
  assign n10811 = n10810 ^ n6994 ^ n665 ;
  assign n10806 = ( ~n2668 & n2967 ) | ( ~n2668 & n8072 ) | ( n2967 & n8072 ) ;
  assign n10807 = n10806 ^ n8383 ^ n2024 ;
  assign n10808 = n10807 ^ n8745 ^ n6810 ;
  assign n10812 = n10811 ^ n10808 ^ n3084 ;
  assign n10813 = ( n2698 & n8896 ) | ( n2698 & ~n9011 ) | ( n8896 & ~n9011 ) ;
  assign n10814 = ( ~n3524 & n4477 ) | ( ~n3524 & n7386 ) | ( n4477 & n7386 ) ;
  assign n10815 = ( n2859 & n10813 ) | ( n2859 & ~n10814 ) | ( n10813 & ~n10814 ) ;
  assign n10816 = n7929 ^ n6700 ^ n3187 ;
  assign n10817 = n10816 ^ n10534 ^ n8194 ;
  assign n10818 = ( n3086 & n5046 ) | ( n3086 & n8762 ) | ( n5046 & n8762 ) ;
  assign n10819 = n10818 ^ n2479 ^ n1624 ;
  assign n10820 = ( n1107 & n8333 ) | ( n1107 & n10819 ) | ( n8333 & n10819 ) ;
  assign n10821 = ( ~n2022 & n4750 ) | ( ~n2022 & n9622 ) | ( n4750 & n9622 ) ;
  assign n10822 = n10821 ^ n7299 ^ x23 ;
  assign n10823 = ( n2727 & n4537 ) | ( n2727 & ~n9242 ) | ( n4537 & ~n9242 ) ;
  assign n10824 = n10823 ^ n8069 ^ n7472 ;
  assign n10825 = ( n1939 & ~n5708 ) | ( n1939 & n7408 ) | ( ~n5708 & n7408 ) ;
  assign n10826 = ( n715 & n9645 ) | ( n715 & ~n10825 ) | ( n9645 & ~n10825 ) ;
  assign n10827 = n6838 ^ n5339 ^ n1815 ;
  assign n10828 = n10827 ^ n9575 ^ n1225 ;
  assign n10829 = n5696 ^ n3967 ^ n679 ;
  assign n10830 = n10829 ^ n3114 ^ n2303 ;
  assign n10831 = ( n4436 & n10828 ) | ( n4436 & ~n10830 ) | ( n10828 & ~n10830 ) ;
  assign n10832 = n10177 ^ n1735 ^ n886 ;
  assign n10833 = ( ~n4283 & n10831 ) | ( ~n4283 & n10832 ) | ( n10831 & n10832 ) ;
  assign n10834 = ( n2475 & ~n3979 ) | ( n2475 & n9888 ) | ( ~n3979 & n9888 ) ;
  assign n10835 = ( n3788 & n5102 ) | ( n3788 & n8169 ) | ( n5102 & n8169 ) ;
  assign n10836 = n6556 ^ n4635 ^ n279 ;
  assign n10837 = ( n279 & ~n5173 ) | ( n279 & n8249 ) | ( ~n5173 & n8249 ) ;
  assign n10838 = n10837 ^ n8240 ^ n2219 ;
  assign n10839 = n10838 ^ n9053 ^ n8370 ;
  assign n10850 = ( n1753 & n6271 ) | ( n1753 & ~n6294 ) | ( n6271 & ~n6294 ) ;
  assign n10851 = ( n1961 & ~n6444 ) | ( n1961 & n8648 ) | ( ~n6444 & n8648 ) ;
  assign n10852 = ( n10501 & ~n10850 ) | ( n10501 & n10851 ) | ( ~n10850 & n10851 ) ;
  assign n10848 = n1721 ^ n594 ^ n462 ;
  assign n10849 = n10848 ^ n8218 ^ n1284 ;
  assign n10844 = n8063 ^ n4202 ^ n1671 ;
  assign n10845 = ( n1322 & ~n3856 ) | ( n1322 & n10844 ) | ( ~n3856 & n10844 ) ;
  assign n10842 = n4233 ^ n2918 ^ n2853 ;
  assign n10843 = ( n1420 & n6623 ) | ( n1420 & ~n10842 ) | ( n6623 & ~n10842 ) ;
  assign n10846 = n10845 ^ n10843 ^ n1521 ;
  assign n10840 = n3413 ^ n3113 ^ n2368 ;
  assign n10841 = n10840 ^ n8228 ^ n6136 ;
  assign n10847 = n10846 ^ n10841 ^ n756 ;
  assign n10853 = n10852 ^ n10849 ^ n10847 ;
  assign n10854 = ( n10836 & n10839 ) | ( n10836 & n10853 ) | ( n10839 & n10853 ) ;
  assign n10859 = ( n320 & ~n4952 ) | ( n320 & n7229 ) | ( ~n4952 & n7229 ) ;
  assign n10856 = ( ~n4952 & n5815 ) | ( ~n4952 & n7358 ) | ( n5815 & n7358 ) ;
  assign n10855 = ( ~x68 & n9139 ) | ( ~x68 & n9270 ) | ( n9139 & n9270 ) ;
  assign n10857 = n10856 ^ n10855 ^ n8652 ;
  assign n10858 = ( n3019 & n8588 ) | ( n3019 & n10857 ) | ( n8588 & n10857 ) ;
  assign n10860 = n10859 ^ n10858 ^ n2379 ;
  assign n10864 = ( n1275 & ~n3591 ) | ( n1275 & n3904 ) | ( ~n3591 & n3904 ) ;
  assign n10861 = n4315 ^ n3842 ^ n3779 ;
  assign n10862 = n10861 ^ n8099 ^ n4789 ;
  assign n10863 = ( n2054 & ~n2967 ) | ( n2054 & n10862 ) | ( ~n2967 & n10862 ) ;
  assign n10865 = n10864 ^ n10863 ^ n925 ;
  assign n10866 = ( ~n177 & n787 ) | ( ~n177 & n6641 ) | ( n787 & n6641 ) ;
  assign n10867 = ( n2937 & n3163 ) | ( n2937 & n3174 ) | ( n3163 & n3174 ) ;
  assign n10868 = n10867 ^ n9141 ^ n7482 ;
  assign n10869 = ( n4584 & ~n10866 ) | ( n4584 & n10868 ) | ( ~n10866 & n10868 ) ;
  assign n10870 = ( n6987 & n7434 ) | ( n6987 & n10869 ) | ( n7434 & n10869 ) ;
  assign n10871 = n10870 ^ n5503 ^ n1701 ;
  assign n10872 = n2747 ^ n2317 ^ x35 ;
  assign n10873 = ( ~n8129 & n10726 ) | ( ~n8129 & n10872 ) | ( n10726 & n10872 ) ;
  assign n10882 = n5541 ^ n1986 ^ n1529 ;
  assign n10880 = n1773 ^ n1653 ^ n517 ;
  assign n10878 = n9412 ^ n5272 ^ n5167 ;
  assign n10877 = n8931 ^ n5958 ^ n3989 ;
  assign n10879 = n10878 ^ n10877 ^ n8013 ;
  assign n10881 = n10880 ^ n10879 ^ x28 ;
  assign n10874 = n4031 ^ n2232 ^ n1778 ;
  assign n10875 = ( n974 & ~n1136 ) | ( n974 & n2079 ) | ( ~n1136 & n2079 ) ;
  assign n10876 = ( ~n4866 & n10874 ) | ( ~n4866 & n10875 ) | ( n10874 & n10875 ) ;
  assign n10883 = n10882 ^ n10881 ^ n10876 ;
  assign n10884 = n5805 ^ n3912 ^ n727 ;
  assign n10885 = ( n1286 & n4046 ) | ( n1286 & n4167 ) | ( n4046 & n4167 ) ;
  assign n10886 = ( ~n4894 & n10884 ) | ( ~n4894 & n10885 ) | ( n10884 & n10885 ) ;
  assign n10887 = n10886 ^ n9096 ^ n4078 ;
  assign n10888 = ( ~n10222 & n10324 ) | ( ~n10222 & n10887 ) | ( n10324 & n10887 ) ;
  assign n10889 = ( n974 & n1761 ) | ( n974 & ~n2304 ) | ( n1761 & ~n2304 ) ;
  assign n10890 = n10889 ^ n7452 ^ n2735 ;
  assign n10891 = n7711 ^ n5744 ^ n1777 ;
  assign n10892 = ( n2261 & n6399 ) | ( n2261 & n10891 ) | ( n6399 & n10891 ) ;
  assign n10893 = n10892 ^ n4045 ^ n1268 ;
  assign n10894 = ( n5002 & ~n10890 ) | ( n5002 & n10893 ) | ( ~n10890 & n10893 ) ;
  assign n10895 = n4067 ^ n1897 ^ n1094 ;
  assign n10896 = n10895 ^ n8913 ^ n3163 ;
  assign n10897 = n7590 ^ n3353 ^ n3036 ;
  assign n10898 = ( n854 & n6133 ) | ( n854 & n10897 ) | ( n6133 & n10897 ) ;
  assign n10899 = ( n3475 & n3667 ) | ( n3475 & ~n4790 ) | ( n3667 & ~n4790 ) ;
  assign n10905 = ( n571 & n6210 ) | ( n571 & n7498 ) | ( n6210 & n7498 ) ;
  assign n10906 = n10905 ^ n9498 ^ n1648 ;
  assign n10903 = ( n2987 & ~n3035 ) | ( n2987 & n3620 ) | ( ~n3035 & n3620 ) ;
  assign n10902 = n6678 ^ n5556 ^ n872 ;
  assign n10904 = n10903 ^ n10902 ^ n6791 ;
  assign n10900 = ( x45 & n2889 ) | ( x45 & n3969 ) | ( n2889 & n3969 ) ;
  assign n10901 = ( n5058 & n7782 ) | ( n5058 & n10900 ) | ( n7782 & n10900 ) ;
  assign n10907 = n10906 ^ n10904 ^ n10901 ;
  assign n10908 = ( ~n743 & n1183 ) | ( ~n743 & n5232 ) | ( n1183 & n5232 ) ;
  assign n10909 = n10908 ^ n7168 ^ n5646 ;
  assign n10910 = ( n528 & n7819 ) | ( n528 & ~n10909 ) | ( n7819 & ~n10909 ) ;
  assign n10911 = ( n554 & ~n1024 ) | ( n554 & n3167 ) | ( ~n1024 & n3167 ) ;
  assign n10912 = ( n681 & n1669 ) | ( n681 & n5230 ) | ( n1669 & n5230 ) ;
  assign n10913 = n10912 ^ n8017 ^ n3318 ;
  assign n10914 = n6529 ^ n4858 ^ n1500 ;
  assign n10915 = n10914 ^ n7346 ^ n4751 ;
  assign n10916 = ( x75 & ~n10768 ) | ( x75 & n10915 ) | ( ~n10768 & n10915 ) ;
  assign n10917 = ( ~n10911 & n10913 ) | ( ~n10911 & n10916 ) | ( n10913 & n10916 ) ;
  assign n10918 = ( ~n8570 & n10910 ) | ( ~n8570 & n10917 ) | ( n10910 & n10917 ) ;
  assign n10919 = n8792 ^ n6689 ^ n2567 ;
  assign n10920 = n5580 ^ n4638 ^ n711 ;
  assign n10921 = n10920 ^ n3923 ^ n2731 ;
  assign n10923 = n7316 ^ n5350 ^ n4645 ;
  assign n10922 = ( n1048 & n2356 ) | ( n1048 & ~n3569 ) | ( n2356 & ~n3569 ) ;
  assign n10924 = n10923 ^ n10922 ^ n9008 ;
  assign n10926 = n3373 ^ n1372 ^ n484 ;
  assign n10927 = n10926 ^ n5010 ^ n4204 ;
  assign n10925 = ( n1106 & n1749 ) | ( n1106 & ~n3080 ) | ( n1749 & ~n3080 ) ;
  assign n10928 = n10927 ^ n10925 ^ n4861 ;
  assign n10929 = ( ~n1164 & n3545 ) | ( ~n1164 & n8240 ) | ( n3545 & n8240 ) ;
  assign n10930 = ( n1455 & n2748 ) | ( n1455 & ~n2760 ) | ( n2748 & ~n2760 ) ;
  assign n10931 = ( n2757 & n5340 ) | ( n2757 & n6150 ) | ( n5340 & n6150 ) ;
  assign n10932 = n10931 ^ n5113 ^ n252 ;
  assign n10933 = n8511 ^ n2750 ^ n1979 ;
  assign n10934 = ( n675 & ~n6119 ) | ( n675 & n10933 ) | ( ~n6119 & n10933 ) ;
  assign n10935 = ( n984 & n1794 ) | ( n984 & n10934 ) | ( n1794 & n10934 ) ;
  assign n10936 = ( n2241 & n4266 ) | ( n2241 & ~n6999 ) | ( n4266 & ~n6999 ) ;
  assign n10937 = ( n6554 & n6580 ) | ( n6554 & n10936 ) | ( n6580 & n10936 ) ;
  assign n10938 = ( n7957 & n10099 ) | ( n7957 & n10937 ) | ( n10099 & n10937 ) ;
  assign n10939 = n10938 ^ n8648 ^ n7869 ;
  assign n10940 = n4098 ^ n3420 ^ n301 ;
  assign n10941 = n10940 ^ n4860 ^ n2565 ;
  assign n10942 = ( n5048 & n8004 ) | ( n5048 & ~n10941 ) | ( n8004 & ~n10941 ) ;
  assign n10946 = ( n2273 & ~n4731 ) | ( n2273 & n5867 ) | ( ~n4731 & n5867 ) ;
  assign n10944 = ( ~n2308 & n9121 ) | ( ~n2308 & n10085 ) | ( n9121 & n10085 ) ;
  assign n10943 = n8941 ^ n3940 ^ n1804 ;
  assign n10945 = n10944 ^ n10943 ^ n4215 ;
  assign n10947 = n10946 ^ n10945 ^ n1309 ;
  assign n10949 = ( x87 & n829 ) | ( x87 & n1354 ) | ( n829 & n1354 ) ;
  assign n10950 = ( n1249 & ~n5409 ) | ( n1249 & n10949 ) | ( ~n5409 & n10949 ) ;
  assign n10948 = n9803 ^ n4595 ^ n1138 ;
  assign n10951 = n10950 ^ n10948 ^ n10396 ;
  assign n10952 = ( n962 & ~n3276 ) | ( n962 & n9871 ) | ( ~n3276 & n9871 ) ;
  assign n10953 = ( ~n6972 & n9354 ) | ( ~n6972 & n10952 ) | ( n9354 & n10952 ) ;
  assign n10954 = ( ~n141 & n5559 ) | ( ~n141 & n6496 ) | ( n5559 & n6496 ) ;
  assign n10955 = n10954 ^ n4904 ^ n3130 ;
  assign n10964 = ( n629 & ~n3536 ) | ( n629 & n5402 ) | ( ~n3536 & n5402 ) ;
  assign n10965 = ( n651 & n788 ) | ( n651 & n10964 ) | ( n788 & n10964 ) ;
  assign n10961 = ( ~n1242 & n7473 ) | ( ~n1242 & n8027 ) | ( n7473 & n8027 ) ;
  assign n10962 = n10961 ^ n4949 ^ n1410 ;
  assign n10960 = n7953 ^ n4936 ^ n1637 ;
  assign n10963 = n10962 ^ n10960 ^ n1305 ;
  assign n10966 = n10965 ^ n10963 ^ n6971 ;
  assign n10956 = n5172 ^ n3839 ^ n2228 ;
  assign n10957 = n8355 ^ n7809 ^ n3857 ;
  assign n10958 = ( n1274 & n5630 ) | ( n1274 & n6505 ) | ( n5630 & n6505 ) ;
  assign n10959 = ( n10956 & n10957 ) | ( n10956 & ~n10958 ) | ( n10957 & ~n10958 ) ;
  assign n10967 = n10966 ^ n10959 ^ n10621 ;
  assign n10968 = n10967 ^ n8061 ^ n5645 ;
  assign n10969 = ( ~x78 & n209 ) | ( ~x78 & n429 ) | ( n209 & n429 ) ;
  assign n10970 = ( ~x24 & n2029 ) | ( ~x24 & n2726 ) | ( n2029 & n2726 ) ;
  assign n10971 = ( n2024 & n8247 ) | ( n2024 & ~n10970 ) | ( n8247 & ~n10970 ) ;
  assign n10972 = ( n7129 & n10969 ) | ( n7129 & n10971 ) | ( n10969 & n10971 ) ;
  assign n10973 = n10472 ^ n3654 ^ n3189 ;
  assign n10974 = ( n515 & ~n4080 ) | ( n515 & n10973 ) | ( ~n4080 & n10973 ) ;
  assign n10975 = ( n9617 & ~n10972 ) | ( n9617 & n10974 ) | ( ~n10972 & n10974 ) ;
  assign n10979 = ( x22 & n1784 ) | ( x22 & n8717 ) | ( n1784 & n8717 ) ;
  assign n10976 = n6162 ^ n3574 ^ n1790 ;
  assign n10977 = ( n2713 & n5390 ) | ( n2713 & ~n10976 ) | ( n5390 & ~n10976 ) ;
  assign n10978 = n10977 ^ n6018 ^ n4922 ;
  assign n10980 = n10979 ^ n10978 ^ n1323 ;
  assign n10981 = n10980 ^ n10484 ^ n3667 ;
  assign n10982 = ( n7886 & n9212 ) | ( n7886 & n10913 ) | ( n9212 & n10913 ) ;
  assign n10986 = ( n2066 & n7154 ) | ( n2066 & ~n9011 ) | ( n7154 & ~n9011 ) ;
  assign n10983 = n6685 ^ n5830 ^ n5472 ;
  assign n10984 = ( n4432 & n4522 ) | ( n4432 & ~n10983 ) | ( n4522 & ~n10983 ) ;
  assign n10985 = ( n2757 & n3213 ) | ( n2757 & n10984 ) | ( n3213 & n10984 ) ;
  assign n10987 = n10986 ^ n10985 ^ n1230 ;
  assign n10988 = n10196 ^ n6245 ^ n1977 ;
  assign n10989 = ( n1493 & ~n1612 ) | ( n1493 & n10988 ) | ( ~n1612 & n10988 ) ;
  assign n10990 = n10989 ^ n7010 ^ n5931 ;
  assign n10992 = n9666 ^ n4576 ^ n290 ;
  assign n10991 = n8899 ^ n5259 ^ n2398 ;
  assign n10993 = n10992 ^ n10991 ^ n7287 ;
  assign n11000 = ( ~n828 & n1189 ) | ( ~n828 & n1276 ) | ( n1189 & n1276 ) ;
  assign n11001 = ( n1714 & ~n3464 ) | ( n1714 & n3581 ) | ( ~n3464 & n3581 ) ;
  assign n11002 = ( n1389 & ~n11000 ) | ( n1389 & n11001 ) | ( ~n11000 & n11001 ) ;
  assign n11003 = n11002 ^ n4101 ^ n1167 ;
  assign n10997 = n9666 ^ n7711 ^ x84 ;
  assign n10998 = n10997 ^ n9698 ^ n279 ;
  assign n10999 = ( n4823 & ~n9491 ) | ( n4823 & n10998 ) | ( ~n9491 & n10998 ) ;
  assign n11004 = n11003 ^ n10999 ^ n3233 ;
  assign n11005 = n7907 ^ n5350 ^ n4157 ;
  assign n11006 = n11005 ^ n4146 ^ n3641 ;
  assign n11007 = ( ~n638 & n11004 ) | ( ~n638 & n11006 ) | ( n11004 & n11006 ) ;
  assign n10994 = ( n4731 & n8163 ) | ( n4731 & ~n10464 ) | ( n8163 & ~n10464 ) ;
  assign n10995 = n8796 ^ n4459 ^ n2278 ;
  assign n10996 = ( n6509 & ~n10994 ) | ( n6509 & n10995 ) | ( ~n10994 & n10995 ) ;
  assign n11008 = n11007 ^ n10996 ^ n4715 ;
  assign n11009 = ( n9591 & n10993 ) | ( n9591 & ~n11008 ) | ( n10993 & ~n11008 ) ;
  assign n11012 = ( ~n1096 & n6235 ) | ( ~n1096 & n7544 ) | ( n6235 & n7544 ) ;
  assign n11013 = ( n1437 & n4110 ) | ( n1437 & n11012 ) | ( n4110 & n11012 ) ;
  assign n11011 = ( n3036 & ~n7823 ) | ( n3036 & n9520 ) | ( ~n7823 & n9520 ) ;
  assign n11010 = ( n1769 & n5428 ) | ( n1769 & ~n5980 ) | ( n5428 & ~n5980 ) ;
  assign n11014 = n11013 ^ n11011 ^ n11010 ;
  assign n11015 = n9077 ^ n4052 ^ n1075 ;
  assign n11016 = n10940 ^ n10336 ^ n8220 ;
  assign n11017 = ( n1363 & n3519 ) | ( n1363 & ~n11016 ) | ( n3519 & ~n11016 ) ;
  assign n11018 = ( ~n2765 & n11015 ) | ( ~n2765 & n11017 ) | ( n11015 & n11017 ) ;
  assign n11022 = ( n641 & ~n2304 ) | ( n641 & n5638 ) | ( ~n2304 & n5638 ) ;
  assign n11023 = ( x73 & n2459 ) | ( x73 & ~n11022 ) | ( n2459 & ~n11022 ) ;
  assign n11019 = n4096 ^ n3174 ^ n1653 ;
  assign n11020 = n11019 ^ n8161 ^ n1448 ;
  assign n11021 = ( n4183 & ~n5652 ) | ( n4183 & n11020 ) | ( ~n5652 & n11020 ) ;
  assign n11024 = n11023 ^ n11021 ^ n3108 ;
  assign n11027 = n8331 ^ n5810 ^ n5601 ;
  assign n11025 = n6230 ^ n3926 ^ n2693 ;
  assign n11026 = ( ~n4824 & n9269 ) | ( ~n4824 & n11025 ) | ( n9269 & n11025 ) ;
  assign n11028 = n11027 ^ n11026 ^ n2092 ;
  assign n11029 = ( n1319 & ~n6411 ) | ( n1319 & n9659 ) | ( ~n6411 & n9659 ) ;
  assign n11030 = n11029 ^ n7561 ^ n3036 ;
  assign n11038 = ( n882 & ~n2037 ) | ( n882 & n5052 ) | ( ~n2037 & n5052 ) ;
  assign n11036 = n8292 ^ n4770 ^ n1665 ;
  assign n11033 = ( n1181 & n1513 ) | ( n1181 & ~n2768 ) | ( n1513 & ~n2768 ) ;
  assign n11034 = n11033 ^ n9430 ^ n2220 ;
  assign n11035 = ( n752 & n5883 ) | ( n752 & ~n11034 ) | ( n5883 & ~n11034 ) ;
  assign n11037 = n11036 ^ n11035 ^ n9078 ;
  assign n11031 = n9513 ^ n9475 ^ n8739 ;
  assign n11032 = n11031 ^ n10861 ^ n5583 ;
  assign n11039 = n11038 ^ n11037 ^ n11032 ;
  assign n11046 = ( n1641 & n1840 ) | ( n1641 & ~n3633 ) | ( n1840 & ~n3633 ) ;
  assign n11047 = n11046 ^ n6971 ^ n2429 ;
  assign n11040 = ( n2075 & n4169 ) | ( n2075 & n7207 ) | ( n4169 & n7207 ) ;
  assign n11041 = ( n2660 & n5783 ) | ( n2660 & n11040 ) | ( n5783 & n11040 ) ;
  assign n11042 = n7830 ^ n5869 ^ n5316 ;
  assign n11043 = ( n1799 & n2767 ) | ( n1799 & n7041 ) | ( n2767 & n7041 ) ;
  assign n11044 = ( n2070 & n11042 ) | ( n2070 & ~n11043 ) | ( n11042 & ~n11043 ) ;
  assign n11045 = ( n3513 & ~n11041 ) | ( n3513 & n11044 ) | ( ~n11041 & n11044 ) ;
  assign n11048 = n11047 ^ n11045 ^ n10375 ;
  assign n11057 = ( n176 & ~n3616 ) | ( n176 & n6825 ) | ( ~n3616 & n6825 ) ;
  assign n11050 = n6344 ^ n4131 ^ n204 ;
  assign n11049 = n8931 ^ n4981 ^ n3847 ;
  assign n11051 = n11050 ^ n11049 ^ n4383 ;
  assign n11052 = ( ~n2577 & n2972 ) | ( ~n2577 & n9222 ) | ( n2972 & n9222 ) ;
  assign n11053 = n6618 ^ n2013 ^ n1025 ;
  assign n11054 = ( ~n2134 & n9472 ) | ( ~n2134 & n11053 ) | ( n9472 & n11053 ) ;
  assign n11055 = ( n972 & n7277 ) | ( n972 & n11054 ) | ( n7277 & n11054 ) ;
  assign n11056 = ( ~n11051 & n11052 ) | ( ~n11051 & n11055 ) | ( n11052 & n11055 ) ;
  assign n11058 = n11057 ^ n11056 ^ n3645 ;
  assign n11062 = n7004 ^ n3023 ^ x52 ;
  assign n11060 = ( n834 & n1067 ) | ( n834 & n1635 ) | ( n1067 & n1635 ) ;
  assign n11059 = n6209 ^ n3420 ^ n1581 ;
  assign n11061 = n11060 ^ n11059 ^ n535 ;
  assign n11063 = n11062 ^ n11061 ^ n9054 ;
  assign n11064 = ( n6520 & ~n7628 ) | ( n6520 & n8881 ) | ( ~n7628 & n8881 ) ;
  assign n11065 = ( n3811 & ~n5418 ) | ( n3811 & n11064 ) | ( ~n5418 & n11064 ) ;
  assign n11074 = n5993 ^ n1628 ^ n1596 ;
  assign n11073 = ( ~n187 & n1666 ) | ( ~n187 & n4683 ) | ( n1666 & n4683 ) ;
  assign n11066 = n4239 ^ n3913 ^ n2206 ;
  assign n11069 = n4325 ^ n3033 ^ n3024 ;
  assign n11067 = n5229 ^ n2327 ^ n554 ;
  assign n11068 = n11067 ^ n2932 ^ n2177 ;
  assign n11070 = n11069 ^ n11068 ^ n259 ;
  assign n11071 = ( ~n8595 & n11066 ) | ( ~n8595 & n11070 ) | ( n11066 & n11070 ) ;
  assign n11072 = ( n1081 & ~n5716 ) | ( n1081 & n11071 ) | ( ~n5716 & n11071 ) ;
  assign n11075 = n11074 ^ n11073 ^ n11072 ;
  assign n11076 = ( n2299 & n5160 ) | ( n2299 & n11075 ) | ( n5160 & n11075 ) ;
  assign n11082 = n8115 ^ n3639 ^ n741 ;
  assign n11081 = ( n5157 & ~n6741 ) | ( n5157 & n10152 ) | ( ~n6741 & n10152 ) ;
  assign n11079 = ( n5112 & n6631 ) | ( n5112 & ~n10107 ) | ( n6631 & ~n10107 ) ;
  assign n11077 = n5732 ^ n4111 ^ n2815 ;
  assign n11078 = ( n5311 & n7832 ) | ( n5311 & n11077 ) | ( n7832 & n11077 ) ;
  assign n11080 = n11079 ^ n11078 ^ n7692 ;
  assign n11083 = n11082 ^ n11081 ^ n11080 ;
  assign n11084 = n2374 ^ n1136 ^ n189 ;
  assign n11085 = n3129 ^ n1423 ^ n1153 ;
  assign n11086 = ( ~n3489 & n11084 ) | ( ~n3489 & n11085 ) | ( n11084 & n11085 ) ;
  assign n11087 = n1111 ^ n153 ^ x126 ;
  assign n11088 = ( n3971 & ~n4651 ) | ( n3971 & n11087 ) | ( ~n4651 & n11087 ) ;
  assign n11089 = n11088 ^ n9574 ^ n3613 ;
  assign n11090 = n11089 ^ n7752 ^ n4859 ;
  assign n11093 = ( n2685 & ~n4440 ) | ( n2685 & n5271 ) | ( ~n4440 & n5271 ) ;
  assign n11092 = n6866 ^ n5459 ^ n1165 ;
  assign n11094 = n11093 ^ n11092 ^ n8298 ;
  assign n11091 = ( n1650 & ~n5334 ) | ( n1650 & n5665 ) | ( ~n5334 & n5665 ) ;
  assign n11095 = n11094 ^ n11091 ^ n1863 ;
  assign n11098 = n6301 ^ n2874 ^ n2561 ;
  assign n11099 = n11098 ^ n6565 ^ n1572 ;
  assign n11096 = n3122 ^ n2335 ^ n470 ;
  assign n11097 = ( n3534 & ~n9903 ) | ( n3534 & n11096 ) | ( ~n9903 & n11096 ) ;
  assign n11100 = n11099 ^ n11097 ^ n7358 ;
  assign n11101 = ( x25 & n4314 ) | ( x25 & n5429 ) | ( n4314 & n5429 ) ;
  assign n11102 = n11101 ^ n10236 ^ n2334 ;
  assign n11103 = n5747 ^ n3446 ^ n1259 ;
  assign n11104 = n11103 ^ n6359 ^ n3072 ;
  assign n11105 = ( n10658 & ~n11040 ) | ( n10658 & n11104 ) | ( ~n11040 & n11104 ) ;
  assign n11106 = ( ~n4311 & n7694 ) | ( ~n4311 & n9724 ) | ( n7694 & n9724 ) ;
  assign n11107 = n11106 ^ n6350 ^ n4219 ;
  assign n11108 = n11107 ^ n10937 ^ n205 ;
  assign n11109 = ( ~n5013 & n5497 ) | ( ~n5013 & n7495 ) | ( n5497 & n7495 ) ;
  assign n11110 = ( ~n1248 & n2349 ) | ( ~n1248 & n4770 ) | ( n2349 & n4770 ) ;
  assign n11111 = n11110 ^ n4587 ^ n1449 ;
  assign n11112 = n11111 ^ n6991 ^ n2935 ;
  assign n11113 = ( n2228 & ~n11109 ) | ( n2228 & n11112 ) | ( ~n11109 & n11112 ) ;
  assign n11114 = n10035 ^ n9712 ^ n6208 ;
  assign n11115 = n11114 ^ n6737 ^ n6660 ;
  assign n11116 = ( n8565 & ~n11113 ) | ( n8565 & n11115 ) | ( ~n11113 & n11115 ) ;
  assign n11117 = ( n608 & n1514 ) | ( n608 & ~n9229 ) | ( n1514 & ~n9229 ) ;
  assign n11118 = n11117 ^ n8238 ^ n7484 ;
  assign n11119 = n9479 ^ n1498 ^ n211 ;
  assign n11120 = n10193 ^ n8175 ^ n1230 ;
  assign n11121 = ( n11118 & n11119 ) | ( n11118 & n11120 ) | ( n11119 & n11120 ) ;
  assign n11122 = n6972 ^ n5823 ^ n3367 ;
  assign n11123 = ( ~n1080 & n3372 ) | ( ~n1080 & n8768 ) | ( n3372 & n8768 ) ;
  assign n11124 = n11123 ^ n8133 ^ n3974 ;
  assign n11125 = ( n1505 & n3728 ) | ( n1505 & n8008 ) | ( n3728 & n8008 ) ;
  assign n11126 = ( n2232 & ~n5463 ) | ( n2232 & n11125 ) | ( ~n5463 & n11125 ) ;
  assign n11127 = ( ~n1983 & n7772 ) | ( ~n1983 & n11126 ) | ( n7772 & n11126 ) ;
  assign n11128 = ( n11122 & n11124 ) | ( n11122 & n11127 ) | ( n11124 & n11127 ) ;
  assign n11129 = n9937 ^ n6428 ^ n2919 ;
  assign n11130 = n11129 ^ n5078 ^ n2608 ;
  assign n11131 = ( x31 & n731 ) | ( x31 & ~n9810 ) | ( n731 & ~n9810 ) ;
  assign n11132 = ( n3714 & n11130 ) | ( n3714 & n11131 ) | ( n11130 & n11131 ) ;
  assign n11133 = ( n714 & ~n2687 ) | ( n714 & n3379 ) | ( ~n2687 & n3379 ) ;
  assign n11134 = ( n681 & n3091 ) | ( n681 & ~n4215 ) | ( n3091 & ~n4215 ) ;
  assign n11135 = ( n8041 & n9867 ) | ( n8041 & n11134 ) | ( n9867 & n11134 ) ;
  assign n11136 = ( n608 & n7214 ) | ( n608 & n11135 ) | ( n7214 & n11135 ) ;
  assign n11137 = ( n2853 & ~n9404 ) | ( n2853 & n9587 ) | ( ~n9404 & n9587 ) ;
  assign n11138 = ( n9818 & ~n11136 ) | ( n9818 & n11137 ) | ( ~n11136 & n11137 ) ;
  assign n11139 = ( n1218 & ~n4729 ) | ( n1218 & n5859 ) | ( ~n4729 & n5859 ) ;
  assign n11140 = n11139 ^ n10410 ^ n6794 ;
  assign n11141 = ( ~n2428 & n4933 ) | ( ~n2428 & n7074 ) | ( n4933 & n7074 ) ;
  assign n11142 = n11141 ^ n5293 ^ n4795 ;
  assign n11143 = ( n4961 & n8058 ) | ( n4961 & ~n11142 ) | ( n8058 & ~n11142 ) ;
  assign n11144 = ( ~n382 & n9522 ) | ( ~n382 & n11143 ) | ( n9522 & n11143 ) ;
  assign n11145 = ( ~n4512 & n6344 ) | ( ~n4512 & n9423 ) | ( n6344 & n9423 ) ;
  assign n11146 = n11145 ^ n3889 ^ n383 ;
  assign n11147 = n11146 ^ n9188 ^ n3056 ;
  assign n11148 = n4813 ^ n4398 ^ n3786 ;
  assign n11149 = n11148 ^ n6008 ^ n5862 ;
  assign n11156 = n5538 ^ n3922 ^ n1584 ;
  assign n11157 = ( n2046 & ~n5357 ) | ( n2046 & n9265 ) | ( ~n5357 & n9265 ) ;
  assign n11158 = ( n3373 & n8186 ) | ( n3373 & ~n11157 ) | ( n8186 & ~n11157 ) ;
  assign n11159 = ( n4041 & ~n11156 ) | ( n4041 & n11158 ) | ( ~n11156 & n11158 ) ;
  assign n11150 = ( n2010 & n2530 ) | ( n2010 & n5118 ) | ( n2530 & n5118 ) ;
  assign n11151 = n11150 ^ n3245 ^ n920 ;
  assign n11152 = n5572 ^ n903 ^ n599 ;
  assign n11153 = n11152 ^ n5139 ^ n186 ;
  assign n11154 = n11153 ^ n10339 ^ n2898 ;
  assign n11155 = ( n8127 & ~n11151 ) | ( n8127 & n11154 ) | ( ~n11151 & n11154 ) ;
  assign n11160 = n11159 ^ n11155 ^ n5772 ;
  assign n11162 = ( n2760 & n4329 ) | ( n2760 & n6414 ) | ( n4329 & n6414 ) ;
  assign n11161 = ( n287 & n1084 ) | ( n287 & ~n6317 ) | ( n1084 & ~n6317 ) ;
  assign n11163 = n11162 ^ n11161 ^ n10369 ;
  assign n11164 = ( n5492 & ~n6589 ) | ( n5492 & n7371 ) | ( ~n6589 & n7371 ) ;
  assign n11165 = n11164 ^ n11145 ^ n5721 ;
  assign n11177 = n4822 ^ n1806 ^ n169 ;
  assign n11178 = n11177 ^ n5972 ^ n1535 ;
  assign n11179 = n11178 ^ n6443 ^ n3747 ;
  assign n11171 = n7031 ^ n5035 ^ n959 ;
  assign n11172 = n11171 ^ n8761 ^ n2670 ;
  assign n11173 = ( n368 & n2364 ) | ( n368 & n3284 ) | ( n2364 & n3284 ) ;
  assign n11174 = n9334 ^ n4172 ^ n1561 ;
  assign n11175 = ( n1786 & n11173 ) | ( n1786 & ~n11174 ) | ( n11173 & ~n11174 ) ;
  assign n11176 = ( n254 & n11172 ) | ( n254 & ~n11175 ) | ( n11172 & ~n11175 ) ;
  assign n11168 = ( n1680 & n6149 ) | ( n1680 & ~n9836 ) | ( n6149 & ~n9836 ) ;
  assign n11169 = n11168 ^ n9854 ^ n5857 ;
  assign n11166 = n4069 ^ n2396 ^ n2019 ;
  assign n11167 = ( n4663 & n10288 ) | ( n4663 & n11166 ) | ( n10288 & n11166 ) ;
  assign n11170 = n11169 ^ n11167 ^ n5968 ;
  assign n11180 = n11179 ^ n11176 ^ n11170 ;
  assign n11181 = ( n1983 & ~n3353 ) | ( n1983 & n5212 ) | ( ~n3353 & n5212 ) ;
  assign n11182 = ( n1564 & ~n2838 ) | ( n1564 & n9728 ) | ( ~n2838 & n9728 ) ;
  assign n11183 = ( n5184 & n11181 ) | ( n5184 & ~n11182 ) | ( n11181 & ~n11182 ) ;
  assign n11184 = ( n2661 & n7314 ) | ( n2661 & n11183 ) | ( n7314 & n11183 ) ;
  assign n11187 = n5956 ^ n3584 ^ n2375 ;
  assign n11188 = ( n412 & n7701 ) | ( n412 & n11187 ) | ( n7701 & n11187 ) ;
  assign n11185 = n2983 ^ n2290 ^ n1717 ;
  assign n11186 = ( ~n6643 & n9658 ) | ( ~n6643 & n11185 ) | ( n9658 & n11185 ) ;
  assign n11189 = n11188 ^ n11186 ^ n3605 ;
  assign n11190 = ( ~n2959 & n4335 ) | ( ~n2959 & n11189 ) | ( n4335 & n11189 ) ;
  assign n11193 = n10258 ^ n7498 ^ n6727 ;
  assign n11191 = ( n1596 & ~n2553 ) | ( n1596 & n7472 ) | ( ~n2553 & n7472 ) ;
  assign n11192 = ( n1777 & ~n2305 ) | ( n1777 & n11191 ) | ( ~n2305 & n11191 ) ;
  assign n11194 = n11193 ^ n11192 ^ n6001 ;
  assign n11195 = ( ~n1673 & n2341 ) | ( ~n1673 & n2904 ) | ( n2341 & n2904 ) ;
  assign n11196 = ( ~n4524 & n5903 ) | ( ~n4524 & n6708 ) | ( n5903 & n6708 ) ;
  assign n11197 = ( ~n3848 & n11195 ) | ( ~n3848 & n11196 ) | ( n11195 & n11196 ) ;
  assign n11198 = ( n5419 & ~n10434 ) | ( n5419 & n11197 ) | ( ~n10434 & n11197 ) ;
  assign n11199 = ( n7912 & n8489 ) | ( n7912 & ~n10245 ) | ( n8489 & ~n10245 ) ;
  assign n11200 = ( n3129 & ~n5918 ) | ( n3129 & n6308 ) | ( ~n5918 & n6308 ) ;
  assign n11201 = ( n5895 & ~n8661 ) | ( n5895 & n11200 ) | ( ~n8661 & n11200 ) ;
  assign n11202 = n11201 ^ n8844 ^ n3701 ;
  assign n11203 = ( n2286 & ~n10908 ) | ( n2286 & n11202 ) | ( ~n10908 & n11202 ) ;
  assign n11204 = ( n990 & n1934 ) | ( n990 & n7432 ) | ( n1934 & n7432 ) ;
  assign n11205 = n11204 ^ n9024 ^ n3799 ;
  assign n11206 = n11205 ^ n9434 ^ n3202 ;
  assign n11207 = ( n617 & ~n2656 ) | ( n617 & n8378 ) | ( ~n2656 & n8378 ) ;
  assign n11208 = ( n2802 & n3042 ) | ( n2802 & ~n8040 ) | ( n3042 & ~n8040 ) ;
  assign n11209 = n11208 ^ n5555 ^ n5478 ;
  assign n11210 = ( ~n3868 & n9413 ) | ( ~n3868 & n11209 ) | ( n9413 & n11209 ) ;
  assign n11216 = ( n189 & n4198 ) | ( n189 & ~n6329 ) | ( n4198 & ~n6329 ) ;
  assign n11211 = ( n685 & n6077 ) | ( n685 & ~n10501 ) | ( n6077 & ~n10501 ) ;
  assign n11212 = n11211 ^ n2042 ^ n1671 ;
  assign n11213 = ( ~n2537 & n7410 ) | ( ~n2537 & n11212 ) | ( n7410 & n11212 ) ;
  assign n11214 = n11213 ^ n9573 ^ n4207 ;
  assign n11215 = n11214 ^ n10712 ^ n4030 ;
  assign n11217 = n11216 ^ n11215 ^ n790 ;
  assign n11218 = ( n1291 & n4512 ) | ( n1291 & ~n11217 ) | ( n4512 & ~n11217 ) ;
  assign n11219 = ( ~n11207 & n11210 ) | ( ~n11207 & n11218 ) | ( n11210 & n11218 ) ;
  assign n11220 = ( n3803 & n7638 ) | ( n3803 & n9347 ) | ( n7638 & n9347 ) ;
  assign n11221 = n11220 ^ n8828 ^ n3671 ;
  assign n11222 = n2914 ^ n913 ^ n446 ;
  assign n11223 = ( n2067 & n4365 ) | ( n2067 & n4500 ) | ( n4365 & n4500 ) ;
  assign n11224 = n5904 ^ n4142 ^ n3207 ;
  assign n11225 = ( ~n2657 & n11223 ) | ( ~n2657 & n11224 ) | ( n11223 & n11224 ) ;
  assign n11226 = ( n2619 & n11222 ) | ( n2619 & ~n11225 ) | ( n11222 & ~n11225 ) ;
  assign n11227 = ( n1449 & n4772 ) | ( n1449 & ~n9226 ) | ( n4772 & ~n9226 ) ;
  assign n11228 = n8192 ^ n4381 ^ n3154 ;
  assign n11229 = ( n3991 & n10370 ) | ( n3991 & ~n11228 ) | ( n10370 & ~n11228 ) ;
  assign n11231 = ( ~n704 & n6457 ) | ( ~n704 & n7997 ) | ( n6457 & n7997 ) ;
  assign n11230 = n10427 ^ n9652 ^ n4861 ;
  assign n11232 = n11231 ^ n11230 ^ n10512 ;
  assign n11233 = ( ~n979 & n10176 ) | ( ~n979 & n11232 ) | ( n10176 & n11232 ) ;
  assign n11234 = n10403 ^ n9683 ^ n3647 ;
  assign n11235 = ( x24 & n2309 ) | ( x24 & n11234 ) | ( n2309 & n11234 ) ;
  assign n11236 = n11235 ^ n10676 ^ n1421 ;
  assign n11237 = n4515 ^ n3106 ^ x40 ;
  assign n11239 = n9687 ^ n6080 ^ n2654 ;
  assign n11238 = n6776 ^ n3204 ^ n244 ;
  assign n11240 = n11239 ^ n11238 ^ n9116 ;
  assign n11241 = ( n3248 & n4392 ) | ( n3248 & n4674 ) | ( n4392 & n4674 ) ;
  assign n11243 = n9366 ^ n9006 ^ n3490 ;
  assign n11242 = ( n6315 & ~n6724 ) | ( n6315 & n10693 ) | ( ~n6724 & n10693 ) ;
  assign n11244 = n11243 ^ n11242 ^ n6952 ;
  assign n11245 = ( n8211 & ~n11241 ) | ( n8211 & n11244 ) | ( ~n11241 & n11244 ) ;
  assign n11246 = ( n11237 & n11240 ) | ( n11237 & ~n11245 ) | ( n11240 & ~n11245 ) ;
  assign n11247 = n3272 ^ n2914 ^ n963 ;
  assign n11248 = ( n4273 & n5297 ) | ( n4273 & n11247 ) | ( n5297 & n11247 ) ;
  assign n11249 = ( n8183 & n11246 ) | ( n8183 & ~n11248 ) | ( n11246 & ~n11248 ) ;
  assign n11250 = n3765 ^ n1528 ^ n463 ;
  assign n11251 = ( ~n6620 & n7997 ) | ( ~n6620 & n11250 ) | ( n7997 & n11250 ) ;
  assign n11252 = n8551 ^ n7113 ^ n1430 ;
  assign n11253 = ( n3120 & n8395 ) | ( n3120 & n11252 ) | ( n8395 & n11252 ) ;
  assign n11254 = ( ~n9782 & n11251 ) | ( ~n9782 & n11253 ) | ( n11251 & n11253 ) ;
  assign n11260 = n5028 ^ n4511 ^ n906 ;
  assign n11258 = ( n730 & n1175 ) | ( n730 & n2171 ) | ( n1175 & n2171 ) ;
  assign n11255 = ( n576 & n4796 ) | ( n576 & ~n6539 ) | ( n4796 & ~n6539 ) ;
  assign n11256 = n9031 ^ n4420 ^ n1627 ;
  assign n11257 = ( n4095 & ~n11255 ) | ( n4095 & n11256 ) | ( ~n11255 & n11256 ) ;
  assign n11259 = n11258 ^ n11257 ^ n4546 ;
  assign n11261 = n11260 ^ n11259 ^ n7728 ;
  assign n11262 = n9091 ^ n4407 ^ n2415 ;
  assign n11263 = n8411 ^ n5356 ^ n3939 ;
  assign n11264 = ( n4393 & n11262 ) | ( n4393 & n11263 ) | ( n11262 & n11263 ) ;
  assign n11265 = ( n238 & n10723 ) | ( n238 & ~n11264 ) | ( n10723 & ~n11264 ) ;
  assign n11266 = ( n666 & n1637 ) | ( n666 & n1769 ) | ( n1637 & n1769 ) ;
  assign n11267 = ( ~n2124 & n5605 ) | ( ~n2124 & n7897 ) | ( n5605 & n7897 ) ;
  assign n11268 = ( ~n2176 & n5545 ) | ( ~n2176 & n11267 ) | ( n5545 & n11267 ) ;
  assign n11269 = ( ~n5968 & n11266 ) | ( ~n5968 & n11268 ) | ( n11266 & n11268 ) ;
  assign n11270 = n6425 ^ n5029 ^ n4351 ;
  assign n11271 = n11270 ^ n1837 ^ n956 ;
  assign n11272 = ( ~n5360 & n7347 ) | ( ~n5360 & n11271 ) | ( n7347 & n11271 ) ;
  assign n11273 = n5963 ^ n3067 ^ n149 ;
  assign n11274 = ( n6891 & ~n11272 ) | ( n6891 & n11273 ) | ( ~n11272 & n11273 ) ;
  assign n11275 = n11023 ^ n10851 ^ n4110 ;
  assign n11276 = n9595 ^ n5359 ^ n5142 ;
  assign n11277 = ( ~n10477 & n11275 ) | ( ~n10477 & n11276 ) | ( n11275 & n11276 ) ;
  assign n11284 = ( x88 & n6100 ) | ( x88 & n10515 ) | ( n6100 & n10515 ) ;
  assign n11283 = n8658 ^ n3301 ^ n1228 ;
  assign n11279 = n9725 ^ n2513 ^ n581 ;
  assign n11278 = ( ~n5356 & n6298 ) | ( ~n5356 & n7071 ) | ( n6298 & n7071 ) ;
  assign n11280 = n11279 ^ n11278 ^ n755 ;
  assign n11281 = n11280 ^ n10109 ^ n9388 ;
  assign n11282 = n11281 ^ n9872 ^ n3290 ;
  assign n11285 = n11284 ^ n11283 ^ n11282 ;
  assign n11286 = n7988 ^ n6440 ^ n963 ;
  assign n11287 = n11286 ^ n3734 ^ n3416 ;
  assign n11288 = ( n4859 & ~n5780 ) | ( n4859 & n11287 ) | ( ~n5780 & n11287 ) ;
  assign n11289 = ( ~n5584 & n11285 ) | ( ~n5584 & n11288 ) | ( n11285 & n11288 ) ;
  assign n11292 = ( n4653 & n4818 ) | ( n4653 & ~n7264 ) | ( n4818 & ~n7264 ) ;
  assign n11293 = n11292 ^ n4109 ^ n3800 ;
  assign n11291 = n4434 ^ n2878 ^ n709 ;
  assign n11294 = n11293 ^ n11291 ^ n4481 ;
  assign n11290 = n4707 ^ n2194 ^ n1577 ;
  assign n11295 = n11294 ^ n11290 ^ n5807 ;
  assign n11296 = n10949 ^ n7471 ^ n5388 ;
  assign n11297 = n8963 ^ n5281 ^ n2082 ;
  assign n11298 = n11297 ^ n1207 ^ n872 ;
  assign n11303 = n9269 ^ n4522 ^ n1771 ;
  assign n11299 = n7060 ^ n7023 ^ n1641 ;
  assign n11300 = n11299 ^ n9380 ^ n7426 ;
  assign n11301 = n11300 ^ n4678 ^ n3719 ;
  assign n11302 = ( n4309 & n7123 ) | ( n4309 & ~n11301 ) | ( n7123 & ~n11301 ) ;
  assign n11304 = n11303 ^ n11302 ^ n9489 ;
  assign n11305 = ( n602 & ~n11298 ) | ( n602 & n11304 ) | ( ~n11298 & n11304 ) ;
  assign n11306 = ( n2964 & ~n4146 ) | ( n2964 & n6298 ) | ( ~n4146 & n6298 ) ;
  assign n11307 = n3248 ^ n1732 ^ n800 ;
  assign n11308 = ( n1069 & n3134 ) | ( n1069 & n3652 ) | ( n3134 & n3652 ) ;
  assign n11309 = ( n8650 & n11307 ) | ( n8650 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11310 = ( n3397 & n11306 ) | ( n3397 & n11309 ) | ( n11306 & n11309 ) ;
  assign n11311 = ( ~n443 & n6738 ) | ( ~n443 & n7005 ) | ( n6738 & n7005 ) ;
  assign n11312 = ( n1026 & n11310 ) | ( n1026 & ~n11311 ) | ( n11310 & ~n11311 ) ;
  assign n11313 = ( n1429 & n5418 ) | ( n1429 & ~n8348 ) | ( n5418 & ~n8348 ) ;
  assign n11314 = n11313 ^ n7620 ^ n3502 ;
  assign n11315 = ( n3288 & n10573 ) | ( n3288 & n11314 ) | ( n10573 & n11314 ) ;
  assign n11316 = n11315 ^ n10922 ^ n5124 ;
  assign n11317 = n9078 ^ n6434 ^ n5403 ;
  assign n11318 = ( n451 & n831 ) | ( n451 & n6322 ) | ( n831 & n6322 ) ;
  assign n11319 = ( ~n463 & n3901 ) | ( ~n463 & n3981 ) | ( n3901 & n3981 ) ;
  assign n11320 = n11319 ^ n2421 ^ n1829 ;
  assign n11321 = ( n9301 & n11318 ) | ( n9301 & n11320 ) | ( n11318 & n11320 ) ;
  assign n11322 = ( n2458 & ~n11317 ) | ( n2458 & n11321 ) | ( ~n11317 & n11321 ) ;
  assign n11323 = n10665 ^ n4023 ^ n1013 ;
  assign n11324 = ( ~n4036 & n5710 ) | ( ~n4036 & n11323 ) | ( n5710 & n11323 ) ;
  assign n11325 = ( x76 & ~n1376 ) | ( x76 & n2504 ) | ( ~n1376 & n2504 ) ;
  assign n11329 = ( ~n2484 & n3995 ) | ( ~n2484 & n5151 ) | ( n3995 & n5151 ) ;
  assign n11330 = ( n1952 & ~n4386 ) | ( n1952 & n11329 ) | ( ~n4386 & n11329 ) ;
  assign n11331 = n11330 ^ n5447 ^ n1076 ;
  assign n11326 = n5150 ^ n2274 ^ x26 ;
  assign n11327 = n8562 ^ n3501 ^ n1411 ;
  assign n11328 = ( n7816 & n11326 ) | ( n7816 & ~n11327 ) | ( n11326 & ~n11327 ) ;
  assign n11332 = n11331 ^ n11328 ^ n11047 ;
  assign n11333 = n10087 ^ n3490 ^ n3223 ;
  assign n11336 = ( ~n413 & n2597 ) | ( ~n413 & n4846 ) | ( n2597 & n4846 ) ;
  assign n11334 = ( n3379 & ~n5297 ) | ( n3379 & n10473 ) | ( ~n5297 & n10473 ) ;
  assign n11335 = n11334 ^ n4298 ^ n262 ;
  assign n11337 = n11336 ^ n11335 ^ n9314 ;
  assign n11338 = ( x91 & ~n4342 ) | ( x91 & n5483 ) | ( ~n4342 & n5483 ) ;
  assign n11339 = ( n1701 & n10168 ) | ( n1701 & n11338 ) | ( n10168 & n11338 ) ;
  assign n11340 = ( n2600 & ~n9085 ) | ( n2600 & n11339 ) | ( ~n9085 & n11339 ) ;
  assign n11341 = n11340 ^ n4374 ^ n196 ;
  assign n11342 = ( n536 & ~n715 ) | ( n536 & n1629 ) | ( ~n715 & n1629 ) ;
  assign n11343 = n11342 ^ n1636 ^ n690 ;
  assign n11344 = ( n3493 & n6691 ) | ( n3493 & ~n11343 ) | ( n6691 & ~n11343 ) ;
  assign n11345 = n11344 ^ n6543 ^ n597 ;
  assign n11346 = n10336 ^ n5770 ^ n1173 ;
  assign n11347 = ( n6123 & ~n7834 ) | ( n6123 & n9396 ) | ( ~n7834 & n9396 ) ;
  assign n11348 = ( n4570 & ~n8653 ) | ( n4570 & n11347 ) | ( ~n8653 & n11347 ) ;
  assign n11349 = ( n5829 & n11346 ) | ( n5829 & n11348 ) | ( n11346 & n11348 ) ;
  assign n11350 = n10241 ^ n2745 ^ n1902 ;
  assign n11351 = n11350 ^ n5932 ^ n1025 ;
  assign n11352 = ( ~n429 & n1776 ) | ( ~n429 & n8919 ) | ( n1776 & n8919 ) ;
  assign n11353 = ( n4831 & n11351 ) | ( n4831 & n11352 ) | ( n11351 & n11352 ) ;
  assign n11354 = ( n956 & n4711 ) | ( n956 & ~n5266 ) | ( n4711 & ~n5266 ) ;
  assign n11355 = ( n528 & n10419 ) | ( n528 & ~n11354 ) | ( n10419 & ~n11354 ) ;
  assign n11356 = ( n3783 & ~n11353 ) | ( n3783 & n11355 ) | ( ~n11353 & n11355 ) ;
  assign n11357 = n9575 ^ n8431 ^ n4621 ;
  assign n11358 = ( n2141 & n5887 ) | ( n2141 & ~n11357 ) | ( n5887 & ~n11357 ) ;
  assign n11359 = ( ~n1692 & n2136 ) | ( ~n1692 & n11358 ) | ( n2136 & n11358 ) ;
  assign n11360 = ( n3112 & n11356 ) | ( n3112 & ~n11359 ) | ( n11356 & ~n11359 ) ;
  assign n11361 = ( n5189 & n7887 ) | ( n5189 & ~n9643 ) | ( n7887 & ~n9643 ) ;
  assign n11367 = n8782 ^ n2261 ^ n1083 ;
  assign n11364 = ( n628 & ~n2150 ) | ( n628 & n5592 ) | ( ~n2150 & n5592 ) ;
  assign n11365 = n11364 ^ n6870 ^ n2783 ;
  assign n11362 = ( ~x13 & n1298 ) | ( ~x13 & n9434 ) | ( n1298 & n9434 ) ;
  assign n11363 = ( ~n7189 & n7469 ) | ( ~n7189 & n11362 ) | ( n7469 & n11362 ) ;
  assign n11366 = n11365 ^ n11363 ^ n6074 ;
  assign n11368 = n11367 ^ n11366 ^ n3780 ;
  assign n11369 = ( n696 & n992 ) | ( n696 & n6017 ) | ( n992 & n6017 ) ;
  assign n11370 = ( n620 & n2943 ) | ( n620 & ~n6045 ) | ( n2943 & ~n6045 ) ;
  assign n11371 = n2018 ^ n1157 ^ n238 ;
  assign n11372 = n11371 ^ n8040 ^ n7294 ;
  assign n11373 = n11372 ^ n2137 ^ n363 ;
  assign n11374 = ( n11369 & n11370 ) | ( n11369 & ~n11373 ) | ( n11370 & ~n11373 ) ;
  assign n11375 = n11374 ^ n5886 ^ n4353 ;
  assign n11376 = n9872 ^ n1907 ^ n1068 ;
  assign n11377 = n4762 ^ n2342 ^ n743 ;
  assign n11378 = ( ~n5796 & n11376 ) | ( ~n5796 & n11377 ) | ( n11376 & n11377 ) ;
  assign n11379 = n11378 ^ n6373 ^ n5610 ;
  assign n11382 = n3457 ^ n707 ^ n474 ;
  assign n11383 = n8953 ^ n4654 ^ n1661 ;
  assign n11384 = ( ~n3441 & n11382 ) | ( ~n3441 & n11383 ) | ( n11382 & n11383 ) ;
  assign n11380 = ( n5386 & ~n9340 ) | ( n5386 & n10537 ) | ( ~n9340 & n10537 ) ;
  assign n11381 = n11380 ^ n7022 ^ n5566 ;
  assign n11385 = n11384 ^ n11381 ^ n3887 ;
  assign n11386 = ( n5131 & n9631 ) | ( n5131 & n9728 ) | ( n9631 & n9728 ) ;
  assign n11387 = ( n5528 & ~n7265 ) | ( n5528 & n8597 ) | ( ~n7265 & n8597 ) ;
  assign n11388 = ( n5643 & ~n9650 ) | ( n5643 & n11387 ) | ( ~n9650 & n11387 ) ;
  assign n11389 = n10965 ^ n9145 ^ n5301 ;
  assign n11390 = ( n1339 & n8844 ) | ( n1339 & n11389 ) | ( n8844 & n11389 ) ;
  assign n11391 = n9059 ^ n5849 ^ n2942 ;
  assign n11392 = ( n844 & ~n3163 ) | ( n844 & n3368 ) | ( ~n3163 & n3368 ) ;
  assign n11393 = ( n1739 & n9525 ) | ( n1739 & n10124 ) | ( n9525 & n10124 ) ;
  assign n11394 = ( ~n6771 & n11392 ) | ( ~n6771 & n11393 ) | ( n11392 & n11393 ) ;
  assign n11395 = ( n2723 & n11391 ) | ( n2723 & n11394 ) | ( n11391 & n11394 ) ;
  assign n11396 = ( ~n554 & n1449 ) | ( ~n554 & n11395 ) | ( n1449 & n11395 ) ;
  assign n11397 = ( n10698 & n11390 ) | ( n10698 & ~n11396 ) | ( n11390 & ~n11396 ) ;
  assign n11398 = ( n297 & n940 ) | ( n297 & n2488 ) | ( n940 & n2488 ) ;
  assign n11399 = ( n8328 & ~n8544 ) | ( n8328 & n11398 ) | ( ~n8544 & n11398 ) ;
  assign n11400 = ( n3112 & ~n7458 ) | ( n3112 & n10110 ) | ( ~n7458 & n10110 ) ;
  assign n11401 = ( n3333 & n3849 ) | ( n3333 & ~n11400 ) | ( n3849 & ~n11400 ) ;
  assign n11402 = ( n8558 & n10264 ) | ( n8558 & n11401 ) | ( n10264 & n11401 ) ;
  assign n11403 = n11402 ^ n3292 ^ n2903 ;
  assign n11404 = ( n2042 & ~n4364 ) | ( n2042 & n4757 ) | ( ~n4364 & n4757 ) ;
  assign n11405 = n11404 ^ n7333 ^ n2877 ;
  assign n11406 = n8064 ^ n2661 ^ n1485 ;
  assign n11415 = n4015 ^ n3453 ^ n426 ;
  assign n11411 = ( ~n637 & n3391 ) | ( ~n637 & n5449 ) | ( n3391 & n5449 ) ;
  assign n11412 = ( n2354 & ~n5769 ) | ( n2354 & n11411 ) | ( ~n5769 & n11411 ) ;
  assign n11413 = n11412 ^ n7781 ^ n2478 ;
  assign n11410 = n8934 ^ n7022 ^ n3679 ;
  assign n11407 = ( n2076 & ~n3784 ) | ( n2076 & n10594 ) | ( ~n3784 & n10594 ) ;
  assign n11408 = n11407 ^ n6256 ^ x104 ;
  assign n11409 = ( n5800 & ~n7087 ) | ( n5800 & n11408 ) | ( ~n7087 & n11408 ) ;
  assign n11414 = n11413 ^ n11410 ^ n11409 ;
  assign n11416 = n11415 ^ n11414 ^ n6425 ;
  assign n11417 = ( n1601 & n11406 ) | ( n1601 & ~n11416 ) | ( n11406 & ~n11416 ) ;
  assign n11419 = n4325 ^ n2217 ^ n1854 ;
  assign n11418 = n8873 ^ n6709 ^ n1894 ;
  assign n11420 = n11419 ^ n11418 ^ n2580 ;
  assign n11421 = ( n6849 & n7414 ) | ( n6849 & n11420 ) | ( n7414 & n11420 ) ;
  assign n11426 = n6222 ^ n4165 ^ n201 ;
  assign n11427 = ( n1402 & ~n3376 ) | ( n1402 & n5889 ) | ( ~n3376 & n5889 ) ;
  assign n11428 = n9103 ^ n2418 ^ n1744 ;
  assign n11429 = ( ~n1601 & n6866 ) | ( ~n1601 & n9908 ) | ( n6866 & n9908 ) ;
  assign n11430 = n4124 ^ n1427 ^ x4 ;
  assign n11431 = ( n11428 & n11429 ) | ( n11428 & ~n11430 ) | ( n11429 & ~n11430 ) ;
  assign n11432 = ( n589 & n11427 ) | ( n589 & n11431 ) | ( n11427 & n11431 ) ;
  assign n11433 = ( ~n523 & n3524 ) | ( ~n523 & n11432 ) | ( n3524 & n11432 ) ;
  assign n11434 = ( n1082 & ~n11426 ) | ( n1082 & n11433 ) | ( ~n11426 & n11433 ) ;
  assign n11422 = ( ~n1587 & n3829 ) | ( ~n1587 & n6765 ) | ( n3829 & n6765 ) ;
  assign n11423 = n11422 ^ n2398 ^ n1358 ;
  assign n11424 = n11423 ^ n6305 ^ n1011 ;
  assign n11425 = n11424 ^ n11287 ^ n10072 ;
  assign n11435 = n11434 ^ n11425 ^ n1373 ;
  assign n11436 = ( n1022 & n2221 ) | ( n1022 & ~n3740 ) | ( n2221 & ~n3740 ) ;
  assign n11437 = ( n1679 & n6187 ) | ( n1679 & ~n10809 ) | ( n6187 & ~n10809 ) ;
  assign n11438 = n11437 ^ n970 ^ n712 ;
  assign n11439 = n3357 ^ n2607 ^ n1336 ;
  assign n11440 = ( n2814 & ~n11438 ) | ( n2814 & n11439 ) | ( ~n11438 & n11439 ) ;
  assign n11442 = n6697 ^ n2376 ^ n793 ;
  assign n11441 = ( ~n2776 & n3061 ) | ( ~n2776 & n3107 ) | ( n3061 & n3107 ) ;
  assign n11443 = n11442 ^ n11441 ^ n5801 ;
  assign n11444 = n11443 ^ n6588 ^ n4954 ;
  assign n11445 = n11444 ^ n10419 ^ n4592 ;
  assign n11446 = n11445 ^ n9502 ^ n6894 ;
  assign n11452 = n2476 ^ n1902 ^ n925 ;
  assign n11449 = n4608 ^ n4064 ^ n2022 ;
  assign n11450 = n11449 ^ n9115 ^ n8079 ;
  assign n11451 = ( ~n4002 & n5743 ) | ( ~n4002 & n11450 ) | ( n5743 & n11450 ) ;
  assign n11447 = n8130 ^ n4105 ^ n217 ;
  assign n11448 = n11447 ^ n4674 ^ n2545 ;
  assign n11453 = n11452 ^ n11451 ^ n11448 ;
  assign n11457 = ( ~n6118 & n6776 ) | ( ~n6118 & n9506 ) | ( n6776 & n9506 ) ;
  assign n11455 = n4704 ^ n4070 ^ n1937 ;
  assign n11454 = ( n3644 & ~n5521 ) | ( n3644 & n10242 ) | ( ~n5521 & n10242 ) ;
  assign n11456 = n11455 ^ n11454 ^ n10003 ;
  assign n11458 = n11457 ^ n11456 ^ n4633 ;
  assign n11459 = n7754 ^ n5593 ^ n5529 ;
  assign n11460 = n11459 ^ n9066 ^ n1704 ;
  assign n11461 = ( n626 & n640 ) | ( n626 & ~n1927 ) | ( n640 & ~n1927 ) ;
  assign n11462 = ( n205 & ~n8735 ) | ( n205 & n11461 ) | ( ~n8735 & n11461 ) ;
  assign n11463 = ( n4124 & n11362 ) | ( n4124 & n11462 ) | ( n11362 & n11462 ) ;
  assign n11468 = ( n302 & n642 ) | ( n302 & n1111 ) | ( n642 & n1111 ) ;
  assign n11467 = n5035 ^ n3130 ^ x50 ;
  assign n11469 = n11468 ^ n11467 ^ n4048 ;
  assign n11470 = ( ~n547 & n5980 ) | ( ~n547 & n11469 ) | ( n5980 & n11469 ) ;
  assign n11464 = n7099 ^ n4157 ^ n3470 ;
  assign n11465 = ( ~n847 & n7510 ) | ( ~n847 & n8250 ) | ( n7510 & n8250 ) ;
  assign n11466 = ( n1642 & ~n11464 ) | ( n1642 & n11465 ) | ( ~n11464 & n11465 ) ;
  assign n11471 = n11470 ^ n11466 ^ n5044 ;
  assign n11473 = n5589 ^ n5023 ^ n200 ;
  assign n11472 = n8829 ^ n8827 ^ n1783 ;
  assign n11474 = n11473 ^ n11472 ^ n2887 ;
  assign n11479 = ( ~n1808 & n3393 ) | ( ~n1808 & n4254 ) | ( n3393 & n4254 ) ;
  assign n11480 = n11479 ^ n4556 ^ n528 ;
  assign n11481 = n11480 ^ n7022 ^ n1798 ;
  assign n11477 = n3017 ^ n2795 ^ n1584 ;
  assign n11478 = ( n1063 & n1346 ) | ( n1063 & n11477 ) | ( n1346 & n11477 ) ;
  assign n11482 = n11481 ^ n11478 ^ n4555 ;
  assign n11475 = ( n141 & ~n1309 ) | ( n141 & n3440 ) | ( ~n1309 & n3440 ) ;
  assign n11476 = ( n3712 & ~n7425 ) | ( n3712 & n11475 ) | ( ~n7425 & n11475 ) ;
  assign n11483 = n11482 ^ n11476 ^ n3944 ;
  assign n11491 = ( n1042 & ~n4878 ) | ( n1042 & n9163 ) | ( ~n4878 & n9163 ) ;
  assign n11489 = ( n3293 & n4080 ) | ( n3293 & n5617 ) | ( n4080 & n5617 ) ;
  assign n11490 = ( ~n1390 & n3563 ) | ( ~n1390 & n11489 ) | ( n3563 & n11489 ) ;
  assign n11484 = ( ~n651 & n3333 ) | ( ~n651 & n7190 ) | ( n3333 & n7190 ) ;
  assign n11485 = ( n3568 & n3574 ) | ( n3568 & n11484 ) | ( n3574 & n11484 ) ;
  assign n11486 = ( ~n3707 & n6769 ) | ( ~n3707 & n8688 ) | ( n6769 & n8688 ) ;
  assign n11487 = n11486 ^ n3821 ^ n2307 ;
  assign n11488 = ( n5743 & n11485 ) | ( n5743 & ~n11487 ) | ( n11485 & ~n11487 ) ;
  assign n11492 = n11491 ^ n11490 ^ n11488 ;
  assign n11493 = ( n240 & n2038 ) | ( n240 & ~n2586 ) | ( n2038 & ~n2586 ) ;
  assign n11494 = ( n6786 & ~n10626 ) | ( n6786 & n11493 ) | ( ~n10626 & n11493 ) ;
  assign n11495 = ( n1264 & n1845 ) | ( n1264 & n4382 ) | ( n1845 & n4382 ) ;
  assign n11496 = n11495 ^ n9563 ^ n4030 ;
  assign n11497 = ( ~n3924 & n11494 ) | ( ~n3924 & n11496 ) | ( n11494 & n11496 ) ;
  assign n11498 = ( n3001 & n7375 ) | ( n3001 & n8283 ) | ( n7375 & n8283 ) ;
  assign n11499 = ( n2687 & n10891 ) | ( n2687 & n11498 ) | ( n10891 & n11498 ) ;
  assign n11500 = n11499 ^ n5969 ^ n2835 ;
  assign n11501 = ( n2598 & n2692 ) | ( n2598 & ~n8918 ) | ( n2692 & ~n8918 ) ;
  assign n11502 = ( n4149 & ~n9389 ) | ( n4149 & n11501 ) | ( ~n9389 & n11501 ) ;
  assign n11507 = n7986 ^ n4114 ^ n1772 ;
  assign n11504 = n1700 ^ n1578 ^ n1480 ;
  assign n11505 = ( ~n229 & n4907 ) | ( ~n229 & n11504 ) | ( n4907 & n11504 ) ;
  assign n11503 = ( n1276 & n6899 ) | ( n1276 & ~n8627 ) | ( n6899 & ~n8627 ) ;
  assign n11506 = n11505 ^ n11503 ^ n5704 ;
  assign n11508 = n11507 ^ n11506 ^ n2797 ;
  assign n11509 = n4863 ^ n3196 ^ n2288 ;
  assign n11510 = ( n4159 & n4752 ) | ( n4159 & ~n11509 ) | ( n4752 & ~n11509 ) ;
  assign n11511 = ( n6157 & n6237 ) | ( n6157 & n11510 ) | ( n6237 & n11510 ) ;
  assign n11512 = n11511 ^ n10819 ^ n10571 ;
  assign n11513 = ( n3165 & ~n5210 ) | ( n3165 & n5763 ) | ( ~n5210 & n5763 ) ;
  assign n11514 = n11513 ^ n6752 ^ n4414 ;
  assign n11515 = n10603 ^ n7005 ^ n2158 ;
  assign n11516 = n10814 ^ n8457 ^ n6084 ;
  assign n11517 = ( n11514 & n11515 ) | ( n11514 & ~n11516 ) | ( n11515 & ~n11516 ) ;
  assign n11518 = n7298 ^ n2889 ^ n1668 ;
  assign n11519 = ( n1052 & ~n2245 ) | ( n1052 & n5987 ) | ( ~n2245 & n5987 ) ;
  assign n11520 = n11519 ^ n9126 ^ n6501 ;
  assign n11521 = n11520 ^ n9315 ^ n2665 ;
  assign n11522 = ( n816 & ~n1983 ) | ( n816 & n9658 ) | ( ~n1983 & n9658 ) ;
  assign n11523 = n6640 ^ n1101 ^ n523 ;
  assign n11524 = ( n3963 & n11522 ) | ( n3963 & n11523 ) | ( n11522 & n11523 ) ;
  assign n11525 = n1322 ^ n892 ^ n749 ;
  assign n11526 = ( ~n9060 & n11524 ) | ( ~n9060 & n11525 ) | ( n11524 & n11525 ) ;
  assign n11527 = ( ~n261 & n8161 ) | ( ~n261 & n10265 ) | ( n8161 & n10265 ) ;
  assign n11528 = n11527 ^ n11159 ^ x12 ;
  assign n11529 = ( ~n159 & n2401 ) | ( ~n159 & n7854 ) | ( n2401 & n7854 ) ;
  assign n11530 = n11529 ^ n8252 ^ n1237 ;
  assign n11531 = n11530 ^ n11514 ^ n1079 ;
  assign n11532 = ( ~n9440 & n11528 ) | ( ~n9440 & n11531 ) | ( n11528 & n11531 ) ;
  assign n11533 = ( n902 & ~n1257 ) | ( n902 & n6825 ) | ( ~n1257 & n6825 ) ;
  assign n11534 = n6129 ^ n6051 ^ n2010 ;
  assign n11535 = ( ~n1707 & n2375 ) | ( ~n1707 & n11534 ) | ( n2375 & n11534 ) ;
  assign n11536 = ( n653 & n1013 ) | ( n653 & ~n6018 ) | ( n1013 & ~n6018 ) ;
  assign n11537 = ( n11533 & ~n11535 ) | ( n11533 & n11536 ) | ( ~n11535 & n11536 ) ;
  assign n11538 = n10635 ^ n5477 ^ n3338 ;
  assign n11539 = ( ~n3647 & n11462 ) | ( ~n3647 & n11538 ) | ( n11462 & n11538 ) ;
  assign n11540 = n11259 ^ n3866 ^ n1313 ;
  assign n11541 = n9498 ^ n7889 ^ n3550 ;
  assign n11542 = n11541 ^ n9186 ^ n2962 ;
  assign n11543 = n11542 ^ n8632 ^ n5394 ;
  assign n11544 = n11035 ^ n5368 ^ n3184 ;
  assign n11545 = n9145 ^ n5953 ^ n4194 ;
  assign n11546 = n4772 ^ n4334 ^ n1512 ;
  assign n11547 = ( n921 & n6734 ) | ( n921 & ~n11546 ) | ( n6734 & ~n11546 ) ;
  assign n11548 = n11005 ^ n4280 ^ n430 ;
  assign n11549 = ( n11545 & ~n11547 ) | ( n11545 & n11548 ) | ( ~n11547 & n11548 ) ;
  assign n11550 = ( n7543 & ~n11544 ) | ( n7543 & n11549 ) | ( ~n11544 & n11549 ) ;
  assign n11551 = ( n2309 & n4116 ) | ( n2309 & n5421 ) | ( n4116 & n5421 ) ;
  assign n11552 = n11551 ^ n10253 ^ n3067 ;
  assign n11553 = n11552 ^ n7407 ^ n6277 ;
  assign n11554 = ( n2081 & n5390 ) | ( n2081 & ~n5418 ) | ( n5390 & ~n5418 ) ;
  assign n11555 = n11554 ^ n2974 ^ n1739 ;
  assign n11556 = ( n1667 & ~n2111 ) | ( n1667 & n7614 ) | ( ~n2111 & n7614 ) ;
  assign n11557 = ( n5153 & n6573 ) | ( n5153 & n11556 ) | ( n6573 & n11556 ) ;
  assign n11558 = n11557 ^ n11441 ^ n337 ;
  assign n11559 = ( n2718 & n2826 ) | ( n2718 & n7146 ) | ( n2826 & n7146 ) ;
  assign n11560 = ( n706 & n900 ) | ( n706 & ~n1714 ) | ( n900 & ~n1714 ) ;
  assign n11561 = n11560 ^ n7048 ^ n1350 ;
  assign n11563 = ( ~n2857 & n8117 ) | ( ~n2857 & n9051 ) | ( n8117 & n9051 ) ;
  assign n11564 = n11563 ^ n9887 ^ n1493 ;
  assign n11565 = n11564 ^ n3533 ^ n2885 ;
  assign n11562 = n10080 ^ n5740 ^ n1917 ;
  assign n11566 = n11565 ^ n11562 ^ n8827 ;
  assign n11567 = ( ~n2945 & n5131 ) | ( ~n2945 & n6487 ) | ( n5131 & n6487 ) ;
  assign n11568 = n4088 ^ n2229 ^ n1871 ;
  assign n11569 = n11568 ^ n10383 ^ n2810 ;
  assign n11570 = n4141 ^ n2712 ^ n444 ;
  assign n11571 = ( n11567 & n11569 ) | ( n11567 & ~n11570 ) | ( n11569 & ~n11570 ) ;
  assign n11572 = ( n3869 & ~n6042 ) | ( n3869 & n7369 ) | ( ~n6042 & n7369 ) ;
  assign n11573 = ( n7231 & n11571 ) | ( n7231 & n11572 ) | ( n11571 & n11572 ) ;
  assign n11574 = n7336 ^ n4244 ^ n3939 ;
  assign n11575 = n11574 ^ n4593 ^ n2799 ;
  assign n11576 = n11575 ^ n3358 ^ n3041 ;
  assign n11577 = ( n1207 & n1927 ) | ( n1207 & ~n4661 ) | ( n1927 & ~n4661 ) ;
  assign n11578 = n11577 ^ n3696 ^ n275 ;
  assign n11579 = ( n482 & n6733 ) | ( n482 & n11578 ) | ( n6733 & n11578 ) ;
  assign n11580 = n10984 ^ n6561 ^ n5045 ;
  assign n11581 = n9882 ^ n4636 ^ n3019 ;
  assign n11582 = ( n1678 & n3347 ) | ( n1678 & ~n11581 ) | ( n3347 & ~n11581 ) ;
  assign n11583 = ( n1204 & ~n7516 ) | ( n1204 & n11582 ) | ( ~n7516 & n11582 ) ;
  assign n11584 = n11583 ^ n6835 ^ n4660 ;
  assign n11585 = ( ~n1759 & n11580 ) | ( ~n1759 & n11584 ) | ( n11580 & n11584 ) ;
  assign n11586 = ( n2222 & n4858 ) | ( n2222 & n5541 ) | ( n4858 & n5541 ) ;
  assign n11587 = ( n5578 & n6302 ) | ( n5578 & n11586 ) | ( n6302 & n11586 ) ;
  assign n11588 = n7776 ^ n6469 ^ n163 ;
  assign n11589 = n11588 ^ n9389 ^ n2859 ;
  assign n11590 = ( n1654 & ~n11587 ) | ( n1654 & n11589 ) | ( ~n11587 & n11589 ) ;
  assign n11591 = ( n4607 & n5976 ) | ( n4607 & n5979 ) | ( n5976 & n5979 ) ;
  assign n11592 = ( n5073 & ~n7008 ) | ( n5073 & n11591 ) | ( ~n7008 & n11591 ) ;
  assign n11593 = ( n835 & n4518 ) | ( n835 & n8029 ) | ( n4518 & n8029 ) ;
  assign n11594 = n6828 ^ n990 ^ n591 ;
  assign n11595 = ( n3202 & n3794 ) | ( n3202 & ~n11594 ) | ( n3794 & ~n11594 ) ;
  assign n11596 = ( ~n2832 & n6155 ) | ( ~n2832 & n11207 ) | ( n6155 & n11207 ) ;
  assign n11597 = n3315 ^ n408 ^ n342 ;
  assign n11598 = n11597 ^ n10020 ^ n1808 ;
  assign n11599 = ( x47 & n427 ) | ( x47 & ~n11598 ) | ( n427 & ~n11598 ) ;
  assign n11600 = ( x19 & n6948 ) | ( x19 & ~n11599 ) | ( n6948 & ~n11599 ) ;
  assign n11601 = ( n713 & ~n11596 ) | ( n713 & n11600 ) | ( ~n11596 & n11600 ) ;
  assign n11605 = n9321 ^ n2970 ^ x90 ;
  assign n11602 = ( x32 & n3414 ) | ( x32 & n10884 ) | ( n3414 & n10884 ) ;
  assign n11603 = ( ~n2383 & n3541 ) | ( ~n2383 & n4605 ) | ( n3541 & n4605 ) ;
  assign n11604 = ( n2253 & n11602 ) | ( n2253 & n11603 ) | ( n11602 & n11603 ) ;
  assign n11606 = n11605 ^ n11604 ^ n9857 ;
  assign n11607 = ( n882 & n5412 ) | ( n882 & n6831 ) | ( n5412 & n6831 ) ;
  assign n11608 = ( n4150 & n8222 ) | ( n4150 & n11607 ) | ( n8222 & n11607 ) ;
  assign n11609 = n11608 ^ n9805 ^ n302 ;
  assign n11610 = ( n721 & n3969 ) | ( n721 & ~n4915 ) | ( n3969 & ~n4915 ) ;
  assign n11611 = n11610 ^ n5417 ^ n3349 ;
  assign n11612 = ( n3960 & n4254 ) | ( n3960 & ~n6890 ) | ( n4254 & ~n6890 ) ;
  assign n11613 = n11612 ^ n5706 ^ n1775 ;
  assign n11614 = ( n8538 & ~n10083 ) | ( n8538 & n11613 ) | ( ~n10083 & n11613 ) ;
  assign n11615 = n6317 ^ n3407 ^ n3003 ;
  assign n11616 = ( n1334 & n10416 ) | ( n1334 & n11615 ) | ( n10416 & n11615 ) ;
  assign n11617 = n11616 ^ n9544 ^ n2092 ;
  assign n11618 = n7538 ^ n5565 ^ n3788 ;
  assign n11619 = ( n1325 & ~n7938 ) | ( n1325 & n11618 ) | ( ~n7938 & n11618 ) ;
  assign n11620 = ( n913 & n3160 ) | ( n913 & n11619 ) | ( n3160 & n11619 ) ;
  assign n11621 = ( ~n1199 & n3690 ) | ( ~n1199 & n6990 ) | ( n3690 & n6990 ) ;
  assign n11622 = n11621 ^ n6910 ^ n1902 ;
  assign n11623 = ( n1293 & n3723 ) | ( n1293 & ~n9548 ) | ( n3723 & ~n9548 ) ;
  assign n11624 = ( n6184 & ~n11622 ) | ( n6184 & n11623 ) | ( ~n11622 & n11623 ) ;
  assign n11625 = ( ~n7424 & n7461 ) | ( ~n7424 & n11624 ) | ( n7461 & n11624 ) ;
  assign n11626 = n9391 ^ n8932 ^ n6777 ;
  assign n11627 = ( n769 & n2844 ) | ( n769 & ~n11626 ) | ( n2844 & ~n11626 ) ;
  assign n11628 = n11472 ^ n8145 ^ n4961 ;
  assign n11629 = ( n889 & ~n1866 ) | ( n889 & n7470 ) | ( ~n1866 & n7470 ) ;
  assign n11630 = n11340 ^ n7363 ^ n1261 ;
  assign n11631 = ( n11118 & n11629 ) | ( n11118 & n11630 ) | ( n11629 & n11630 ) ;
  assign n11632 = ( n2529 & n2995 ) | ( n2529 & n3850 ) | ( n2995 & n3850 ) ;
  assign n11633 = n11632 ^ n8783 ^ n7572 ;
  assign n11640 = ( n3956 & ~n5133 ) | ( n3956 & n8758 ) | ( ~n5133 & n8758 ) ;
  assign n11641 = n11640 ^ n10216 ^ n9487 ;
  assign n11638 = n4910 ^ n4037 ^ n1917 ;
  assign n11637 = n10264 ^ n10059 ^ n3060 ;
  assign n11634 = ( n2223 & n7560 ) | ( n2223 & ~n8145 ) | ( n7560 & ~n8145 ) ;
  assign n11635 = ( ~n819 & n7951 ) | ( ~n819 & n11634 ) | ( n7951 & n11634 ) ;
  assign n11636 = n11635 ^ n10889 ^ n372 ;
  assign n11639 = n11638 ^ n11637 ^ n11636 ;
  assign n11642 = n11641 ^ n11639 ^ n5635 ;
  assign n11643 = n11642 ^ n8885 ^ n421 ;
  assign n11645 = n10109 ^ n8981 ^ n6927 ;
  assign n11644 = ( n4275 & n7187 ) | ( n4275 & n10964 ) | ( n7187 & n10964 ) ;
  assign n11646 = n11645 ^ n11644 ^ n2809 ;
  assign n11647 = n11646 ^ n7566 ^ n2735 ;
  assign n11650 = n4736 ^ n3408 ^ n2136 ;
  assign n11648 = n8866 ^ n5404 ^ x42 ;
  assign n11649 = n11648 ^ n5981 ^ n4108 ;
  assign n11651 = n11650 ^ n11649 ^ n10727 ;
  assign n11652 = n6910 ^ n2528 ^ n235 ;
  assign n11653 = n11652 ^ n5690 ^ n1934 ;
  assign n11654 = ( n5022 & ~n8129 ) | ( n5022 & n11653 ) | ( ~n8129 & n11653 ) ;
  assign n11655 = ( n283 & n5646 ) | ( n283 & ~n11654 ) | ( n5646 & ~n11654 ) ;
  assign n11656 = ( n2991 & n3689 ) | ( n2991 & ~n11655 ) | ( n3689 & ~n11655 ) ;
  assign n11657 = ( ~n7099 & n7405 ) | ( ~n7099 & n10152 ) | ( n7405 & n10152 ) ;
  assign n11658 = ( n3439 & ~n9001 ) | ( n3439 & n11657 ) | ( ~n9001 & n11657 ) ;
  assign n11659 = n11658 ^ n8856 ^ n1894 ;
  assign n11660 = n9483 ^ n7632 ^ n387 ;
  assign n11661 = n11660 ^ n4711 ^ n573 ;
  assign n11662 = n11088 ^ n2791 ^ n1735 ;
  assign n11663 = n11662 ^ n3728 ^ n2772 ;
  assign n11664 = ( ~n2528 & n6653 ) | ( ~n2528 & n7113 ) | ( n6653 & n7113 ) ;
  assign n11665 = n8253 ^ n4269 ^ n1081 ;
  assign n11666 = ( n2990 & n9640 ) | ( n2990 & ~n11665 ) | ( n9640 & ~n11665 ) ;
  assign n11667 = ( n676 & n11664 ) | ( n676 & n11666 ) | ( n11664 & n11666 ) ;
  assign n11668 = n11667 ^ n1434 ^ n997 ;
  assign n11669 = n11668 ^ n4687 ^ n2014 ;
  assign n11670 = ( n8575 & n11663 ) | ( n8575 & ~n11669 ) | ( n11663 & ~n11669 ) ;
  assign n11671 = ( ~n6104 & n11661 ) | ( ~n6104 & n11670 ) | ( n11661 & n11670 ) ;
  assign n11673 = n9728 ^ n7703 ^ n1662 ;
  assign n11672 = ( n1536 & ~n5826 ) | ( n1536 & n8417 ) | ( ~n5826 & n8417 ) ;
  assign n11674 = n11673 ^ n11672 ^ n9176 ;
  assign n11676 = ( n1833 & n3313 ) | ( n1833 & n11266 ) | ( n3313 & n11266 ) ;
  assign n11677 = n2393 ^ n2162 ^ n1568 ;
  assign n11678 = n3743 ^ n1923 ^ n1893 ;
  assign n11679 = ( ~n3407 & n11677 ) | ( ~n3407 & n11678 ) | ( n11677 & n11678 ) ;
  assign n11680 = ( n10425 & n11676 ) | ( n10425 & ~n11679 ) | ( n11676 & ~n11679 ) ;
  assign n11681 = ( n375 & ~n5797 ) | ( n375 & n11680 ) | ( ~n5797 & n11680 ) ;
  assign n11675 = ( n3752 & n5061 ) | ( n3752 & n10348 ) | ( n5061 & n10348 ) ;
  assign n11682 = n11681 ^ n11675 ^ n5794 ;
  assign n11683 = ( ~n3228 & n7260 ) | ( ~n3228 & n9894 ) | ( n7260 & n9894 ) ;
  assign n11684 = ( n1120 & ~n7565 ) | ( n1120 & n10882 ) | ( ~n7565 & n10882 ) ;
  assign n11685 = ( n936 & n8851 ) | ( n936 & ~n11684 ) | ( n8851 & ~n11684 ) ;
  assign n11686 = n6887 ^ n6475 ^ n5891 ;
  assign n11687 = ( ~n4171 & n7821 ) | ( ~n4171 & n11686 ) | ( n7821 & n11686 ) ;
  assign n11688 = n11657 ^ n4293 ^ n2511 ;
  assign n11689 = n9643 ^ n2366 ^ n778 ;
  assign n11690 = ( n8250 & n8795 ) | ( n8250 & ~n11689 ) | ( n8795 & ~n11689 ) ;
  assign n11696 = ( n2788 & ~n3803 ) | ( n2788 & n8069 ) | ( ~n3803 & n8069 ) ;
  assign n11697 = ( n3343 & n5090 ) | ( n3343 & ~n11696 ) | ( n5090 & ~n11696 ) ;
  assign n11698 = n11697 ^ n9877 ^ n879 ;
  assign n11699 = n11698 ^ n11174 ^ n1708 ;
  assign n11700 = ( ~n479 & n3200 ) | ( ~n479 & n4403 ) | ( n3200 & n4403 ) ;
  assign n11701 = ( n1261 & n6175 ) | ( n1261 & n11700 ) | ( n6175 & n11700 ) ;
  assign n11702 = ( n1811 & n3450 ) | ( n1811 & n11701 ) | ( n3450 & n11701 ) ;
  assign n11703 = n11702 ^ n9974 ^ n4497 ;
  assign n11704 = n3935 ^ n3879 ^ n2806 ;
  assign n11705 = n11704 ^ n6162 ^ n5793 ;
  assign n11706 = n11705 ^ n3233 ^ n804 ;
  assign n11707 = n11706 ^ n4241 ^ x62 ;
  assign n11708 = ( n11699 & n11703 ) | ( n11699 & n11707 ) | ( n11703 & n11707 ) ;
  assign n11691 = n4691 ^ n972 ^ n273 ;
  assign n11692 = n11691 ^ n593 ^ n573 ;
  assign n11693 = ( n1096 & n4464 ) | ( n1096 & n11306 ) | ( n4464 & n11306 ) ;
  assign n11694 = ( n1070 & ~n5972 ) | ( n1070 & n7829 ) | ( ~n5972 & n7829 ) ;
  assign n11695 = ( ~n11692 & n11693 ) | ( ~n11692 & n11694 ) | ( n11693 & n11694 ) ;
  assign n11709 = n11708 ^ n11695 ^ n5653 ;
  assign n11711 = n10914 ^ n5181 ^ n3103 ;
  assign n11710 = ( n3606 & ~n5783 ) | ( n3606 & n10587 ) | ( ~n5783 & n10587 ) ;
  assign n11712 = n11711 ^ n11710 ^ n11376 ;
  assign n11713 = ( n2728 & ~n4141 ) | ( n2728 & n11712 ) | ( ~n4141 & n11712 ) ;
  assign n11714 = ( n556 & n4621 ) | ( n556 & n9347 ) | ( n4621 & n9347 ) ;
  assign n11715 = n11714 ^ n3080 ^ n2083 ;
  assign n11718 = n7853 ^ n7635 ^ n3240 ;
  assign n11719 = ( n3324 & n11013 ) | ( n3324 & ~n11718 ) | ( n11013 & ~n11718 ) ;
  assign n11716 = ( n3056 & ~n4220 ) | ( n3056 & n10665 ) | ( ~n4220 & n10665 ) ;
  assign n11717 = ( n4561 & ~n11068 ) | ( n4561 & n11716 ) | ( ~n11068 & n11716 ) ;
  assign n11720 = n11719 ^ n11717 ^ n7274 ;
  assign n11721 = ( ~n4773 & n10119 ) | ( ~n4773 & n11720 ) | ( n10119 & n11720 ) ;
  assign n11722 = ( n2411 & n8267 ) | ( n2411 & n11721 ) | ( n8267 & n11721 ) ;
  assign n11723 = ( ~n1712 & n11715 ) | ( ~n1712 & n11722 ) | ( n11715 & n11722 ) ;
  assign n11724 = ( n449 & n2761 ) | ( n449 & ~n11723 ) | ( n2761 & ~n11723 ) ;
  assign n11729 = n7547 ^ n3272 ^ n586 ;
  assign n11725 = ( n1156 & ~n4578 ) | ( n1156 & n8568 ) | ( ~n4578 & n8568 ) ;
  assign n11726 = ( n1281 & n8233 ) | ( n1281 & ~n11725 ) | ( n8233 & ~n11725 ) ;
  assign n11727 = n11726 ^ n2641 ^ n244 ;
  assign n11728 = ( n4945 & n7370 ) | ( n4945 & n11727 ) | ( n7370 & n11727 ) ;
  assign n11730 = n11729 ^ n11728 ^ n4869 ;
  assign n11731 = n6660 ^ n3748 ^ n653 ;
  assign n11732 = ( n1558 & ~n9889 ) | ( n1558 & n11731 ) | ( ~n9889 & n11731 ) ;
  assign n11733 = ( n3697 & ~n7003 ) | ( n3697 & n11732 ) | ( ~n7003 & n11732 ) ;
  assign n11734 = n11733 ^ n6442 ^ n1158 ;
  assign n11737 = n10936 ^ n7452 ^ n6070 ;
  assign n11735 = n4939 ^ n306 ^ n303 ;
  assign n11736 = ( ~n1021 & n3524 ) | ( ~n1021 & n11735 ) | ( n3524 & n11735 ) ;
  assign n11738 = n11737 ^ n11736 ^ n8356 ;
  assign n11739 = n11738 ^ n11383 ^ n2281 ;
  assign n11740 = n6940 ^ n2603 ^ n2138 ;
  assign n11741 = ( n1491 & n5668 ) | ( n1491 & n5726 ) | ( n5668 & n5726 ) ;
  assign n11742 = ( n3326 & n4101 ) | ( n3326 & ~n5639 ) | ( n4101 & ~n5639 ) ;
  assign n11743 = n6366 ^ n5236 ^ n2517 ;
  assign n11744 = ( ~n1400 & n11742 ) | ( ~n1400 & n11743 ) | ( n11742 & n11743 ) ;
  assign n11745 = ( n9046 & n11741 ) | ( n9046 & n11744 ) | ( n11741 & n11744 ) ;
  assign n11746 = ( ~n3120 & n5013 ) | ( ~n3120 & n9942 ) | ( n5013 & n9942 ) ;
  assign n11747 = ( n11740 & ~n11745 ) | ( n11740 & n11746 ) | ( ~n11745 & n11746 ) ;
  assign n11748 = ( n1980 & n4386 ) | ( n1980 & n11747 ) | ( n4386 & n11747 ) ;
  assign n11749 = ( n457 & ~n3045 ) | ( n457 & n3785 ) | ( ~n3045 & n3785 ) ;
  assign n11750 = ( n1985 & n3077 ) | ( n1985 & ~n5522 ) | ( n3077 & ~n5522 ) ;
  assign n11751 = ( ~n409 & n11749 ) | ( ~n409 & n11750 ) | ( n11749 & n11750 ) ;
  assign n11752 = n10467 ^ n8077 ^ n1950 ;
  assign n11754 = n9438 ^ n7419 ^ n4597 ;
  assign n11753 = ( ~n4967 & n7033 ) | ( ~n4967 & n7687 ) | ( n7033 & n7687 ) ;
  assign n11755 = n11754 ^ n11753 ^ n10841 ;
  assign n11756 = ( n1773 & n6905 ) | ( n1773 & ~n10644 ) | ( n6905 & ~n10644 ) ;
  assign n11757 = ( n898 & n2206 ) | ( n898 & n10094 ) | ( n2206 & n10094 ) ;
  assign n11758 = ( x125 & ~n1078 ) | ( x125 & n2891 ) | ( ~n1078 & n2891 ) ;
  assign n11759 = ( n2264 & ~n4599 ) | ( n2264 & n11758 ) | ( ~n4599 & n11758 ) ;
  assign n11763 = n2808 ^ n2199 ^ n1381 ;
  assign n11764 = ( n2301 & n3539 ) | ( n2301 & ~n11763 ) | ( n3539 & ~n11763 ) ;
  assign n11765 = ( n1125 & ~n2698 ) | ( n1125 & n11764 ) | ( ~n2698 & n11764 ) ;
  assign n11760 = ( n1056 & n8137 ) | ( n1056 & n9351 ) | ( n8137 & n9351 ) ;
  assign n11761 = n11760 ^ n9612 ^ n2116 ;
  assign n11762 = ( n1982 & n6898 ) | ( n1982 & n11761 ) | ( n6898 & n11761 ) ;
  assign n11766 = n11765 ^ n11762 ^ n5547 ;
  assign n11767 = ( ~n5190 & n8066 ) | ( ~n5190 & n8677 ) | ( n8066 & n8677 ) ;
  assign n11768 = ( ~n769 & n2672 ) | ( ~n769 & n4447 ) | ( n2672 & n4447 ) ;
  assign n11769 = ( n2258 & n2617 ) | ( n2258 & ~n3557 ) | ( n2617 & ~n3557 ) ;
  assign n11770 = n11769 ^ n7455 ^ n479 ;
  assign n11771 = ( ~n148 & n2505 ) | ( ~n148 & n8007 ) | ( n2505 & n8007 ) ;
  assign n11772 = n11771 ^ n1680 ^ n858 ;
  assign n11773 = ( n4653 & ~n8652 ) | ( n4653 & n11772 ) | ( ~n8652 & n11772 ) ;
  assign n11774 = ( n10651 & n11770 ) | ( n10651 & n11773 ) | ( n11770 & n11773 ) ;
  assign n11775 = ( n11767 & n11768 ) | ( n11767 & ~n11774 ) | ( n11768 & ~n11774 ) ;
  assign n11780 = n8625 ^ n2629 ^ n131 ;
  assign n11778 = ( n2704 & n4265 ) | ( n2704 & ~n4578 ) | ( n4265 & ~n4578 ) ;
  assign n11779 = ( n9646 & n11017 ) | ( n9646 & n11778 ) | ( n11017 & n11778 ) ;
  assign n11776 = ( ~n4860 & n4862 ) | ( ~n4860 & n11714 ) | ( n4862 & n11714 ) ;
  assign n11777 = ( ~n4514 & n9972 ) | ( ~n4514 & n11776 ) | ( n9972 & n11776 ) ;
  assign n11781 = n11780 ^ n11779 ^ n11777 ;
  assign n11786 = ( n699 & ~n7774 ) | ( n699 & n9683 ) | ( ~n7774 & n9683 ) ;
  assign n11784 = ( x16 & n1261 ) | ( x16 & n4210 ) | ( n1261 & n4210 ) ;
  assign n11782 = n7693 ^ n6956 ^ n6760 ;
  assign n11783 = n11782 ^ n6301 ^ n1381 ;
  assign n11785 = n11784 ^ n11783 ^ n6775 ;
  assign n11787 = n11786 ^ n11785 ^ n1355 ;
  assign n11788 = ( n3271 & ~n4184 ) | ( n3271 & n11787 ) | ( ~n4184 & n11787 ) ;
  assign n11791 = n9187 ^ n8171 ^ n3289 ;
  assign n11789 = n10927 ^ n3811 ^ n1474 ;
  assign n11790 = ( ~n1460 & n10790 ) | ( ~n1460 & n11789 ) | ( n10790 & n11789 ) ;
  assign n11792 = n11791 ^ n11790 ^ n8645 ;
  assign n11793 = ( n321 & n4193 ) | ( n321 & ~n7428 ) | ( n4193 & ~n7428 ) ;
  assign n11794 = ( n2585 & n6972 ) | ( n2585 & ~n11793 ) | ( n6972 & ~n11793 ) ;
  assign n11795 = ( n1930 & n8597 ) | ( n1930 & n10513 ) | ( n8597 & n10513 ) ;
  assign n11797 = n9391 ^ n6573 ^ n1010 ;
  assign n11796 = n8702 ^ n8407 ^ n1043 ;
  assign n11798 = n11797 ^ n11796 ^ n11096 ;
  assign n11799 = ( n11794 & n11795 ) | ( n11794 & n11798 ) | ( n11795 & n11798 ) ;
  assign n11800 = n11799 ^ n3587 ^ n2802 ;
  assign n11801 = n11800 ^ n11189 ^ n640 ;
  assign n11802 = ( n1040 & ~n3243 ) | ( n1040 & n4965 ) | ( ~n3243 & n4965 ) ;
  assign n11803 = n11802 ^ n4526 ^ n507 ;
  assign n11804 = n8102 ^ n4973 ^ n4085 ;
  assign n11805 = n11059 ^ n1847 ^ n1187 ;
  assign n11806 = ( n562 & ~n4701 ) | ( n562 & n11805 ) | ( ~n4701 & n11805 ) ;
  assign n11807 = ( n4766 & ~n6954 ) | ( n4766 & n11806 ) | ( ~n6954 & n11806 ) ;
  assign n11809 = ( n802 & ~n7633 ) | ( n802 & n10442 ) | ( ~n7633 & n10442 ) ;
  assign n11808 = ( n733 & ~n7821 ) | ( n733 & n9863 ) | ( ~n7821 & n9863 ) ;
  assign n11810 = n11809 ^ n11808 ^ n6514 ;
  assign n11811 = n9130 ^ n2283 ^ n1842 ;
  assign n11812 = n11811 ^ n5815 ^ n5252 ;
  assign n11813 = ( ~n952 & n1143 ) | ( ~n952 & n11377 ) | ( n1143 & n11377 ) ;
  assign n11814 = ( n1012 & n7036 ) | ( n1012 & ~n11813 ) | ( n7036 & ~n11813 ) ;
  assign n11815 = ( ~n804 & n3854 ) | ( ~n804 & n4843 ) | ( n3854 & n4843 ) ;
  assign n11816 = ( n1583 & n4299 ) | ( n1583 & n11815 ) | ( n4299 & n11815 ) ;
  assign n11817 = ( ~x1 & n392 ) | ( ~x1 & n9884 ) | ( n392 & n9884 ) ;
  assign n11818 = ( n3392 & ~n6392 ) | ( n3392 & n11817 ) | ( ~n6392 & n11817 ) ;
  assign n11826 = ( ~x18 & n152 ) | ( ~x18 & n2641 ) | ( n152 & n2641 ) ;
  assign n11823 = ( n2061 & n6554 ) | ( n2061 & ~n8112 ) | ( n6554 & ~n8112 ) ;
  assign n11824 = ( n2962 & ~n5090 ) | ( n2962 & n11823 ) | ( ~n5090 & n11823 ) ;
  assign n11825 = n11824 ^ n7408 ^ n3109 ;
  assign n11819 = ( n257 & n2606 ) | ( n257 & ~n3540 ) | ( n2606 & ~n3540 ) ;
  assign n11820 = n11819 ^ n2705 ^ n513 ;
  assign n11821 = ( n900 & ~n4102 ) | ( n900 & n11820 ) | ( ~n4102 & n11820 ) ;
  assign n11822 = ( n6806 & ~n9415 ) | ( n6806 & n11821 ) | ( ~n9415 & n11821 ) ;
  assign n11827 = n11826 ^ n11825 ^ n11822 ;
  assign n11829 = ( n699 & n1450 ) | ( n699 & n3047 ) | ( n1450 & n3047 ) ;
  assign n11830 = ( n1252 & ~n9891 ) | ( n1252 & n11829 ) | ( ~n9891 & n11829 ) ;
  assign n11831 = ( n5635 & n7222 ) | ( n5635 & n11830 ) | ( n7222 & n11830 ) ;
  assign n11828 = ( n3702 & ~n5198 ) | ( n3702 & n6162 ) | ( ~n5198 & n6162 ) ;
  assign n11832 = n11831 ^ n11828 ^ n4002 ;
  assign n11833 = ( n781 & ~n5329 ) | ( n781 & n11704 ) | ( ~n5329 & n11704 ) ;
  assign n11838 = ( n535 & ~n5209 ) | ( n535 & n8340 ) | ( ~n5209 & n8340 ) ;
  assign n11834 = ( ~n307 & n2181 ) | ( ~n307 & n3081 ) | ( n2181 & n3081 ) ;
  assign n11835 = ( n3614 & n3634 ) | ( n3614 & n11834 ) | ( n3634 & n11834 ) ;
  assign n11836 = ( ~n3301 & n5810 ) | ( ~n3301 & n7833 ) | ( n5810 & n7833 ) ;
  assign n11837 = ( n6486 & n11835 ) | ( n6486 & n11836 ) | ( n11835 & n11836 ) ;
  assign n11839 = n11838 ^ n11837 ^ n3466 ;
  assign n11840 = n9050 ^ n6986 ^ n2101 ;
  assign n11841 = ( n946 & n9551 ) | ( n946 & ~n11840 ) | ( n9551 & ~n11840 ) ;
  assign n11849 = n3241 ^ n3204 ^ n2386 ;
  assign n11847 = ( n777 & n2116 ) | ( n777 & n4673 ) | ( n2116 & n4673 ) ;
  assign n11848 = n11847 ^ n10771 ^ n9469 ;
  assign n11842 = ( n4636 & n5284 ) | ( n4636 & ~n9008 ) | ( n5284 & ~n9008 ) ;
  assign n11843 = n11842 ^ n11749 ^ n2829 ;
  assign n11844 = ( ~n2877 & n3714 ) | ( ~n2877 & n11843 ) | ( n3714 & n11843 ) ;
  assign n11845 = ( ~n2465 & n6796 ) | ( ~n2465 & n11844 ) | ( n6796 & n11844 ) ;
  assign n11846 = n11845 ^ n3549 ^ n2927 ;
  assign n11850 = n11849 ^ n11848 ^ n11846 ;
  assign n11856 = n3584 ^ n2636 ^ n137 ;
  assign n11852 = ( n933 & n4189 ) | ( n933 & ~n11238 ) | ( n4189 & ~n11238 ) ;
  assign n11853 = ( n10468 & n10789 ) | ( n10468 & n11852 ) | ( n10789 & n11852 ) ;
  assign n11851 = ( ~n1879 & n3060 ) | ( ~n1879 & n8782 ) | ( n3060 & n8782 ) ;
  assign n11854 = n11853 ^ n11851 ^ n2441 ;
  assign n11855 = n11854 ^ n10392 ^ n5255 ;
  assign n11857 = n11856 ^ n11855 ^ n7585 ;
  assign n11860 = ( ~n1504 & n2021 ) | ( ~n1504 & n3648 ) | ( n2021 & n3648 ) ;
  assign n11858 = ( n3388 & n7970 ) | ( n3388 & ~n9469 ) | ( n7970 & ~n9469 ) ;
  assign n11859 = ( n372 & n8641 ) | ( n372 & n11858 ) | ( n8641 & n11858 ) ;
  assign n11861 = n11860 ^ n11859 ^ n4014 ;
  assign n11862 = ( ~x39 & n2725 ) | ( ~x39 & n3373 ) | ( n2725 & n3373 ) ;
  assign n11863 = ( n8392 & n9946 ) | ( n8392 & ~n11862 ) | ( n9946 & ~n11862 ) ;
  assign n11864 = ( n3770 & n6059 ) | ( n3770 & n6726 ) | ( n6059 & n6726 ) ;
  assign n11865 = ( n2749 & n5348 ) | ( n2749 & n11864 ) | ( n5348 & n11864 ) ;
  assign n11867 = ( n4348 & n5180 ) | ( n4348 & n5400 ) | ( n5180 & n5400 ) ;
  assign n11866 = n7243 ^ n3540 ^ n1088 ;
  assign n11868 = n11867 ^ n11866 ^ n1929 ;
  assign n11871 = n10690 ^ n8782 ^ n4701 ;
  assign n11872 = ( x42 & ~n5233 ) | ( x42 & n11871 ) | ( ~n5233 & n11871 ) ;
  assign n11873 = n11872 ^ n2495 ^ n318 ;
  assign n11869 = n5994 ^ n2972 ^ n2182 ;
  assign n11870 = n11869 ^ n6460 ^ n3742 ;
  assign n11874 = n11873 ^ n11870 ^ n2266 ;
  assign n11876 = ( n727 & n5732 ) | ( n727 & n8821 ) | ( n5732 & n8821 ) ;
  assign n11875 = n10827 ^ n8525 ^ n5255 ;
  assign n11877 = n11876 ^ n11875 ^ n11366 ;
  assign n11879 = ( n7267 & n9200 ) | ( n7267 & ~n9707 ) | ( n9200 & ~n9707 ) ;
  assign n11878 = n6075 ^ n5505 ^ n1770 ;
  assign n11880 = n11879 ^ n11878 ^ x121 ;
  assign n11882 = ( n1085 & ~n2089 ) | ( n1085 & n2144 ) | ( ~n2089 & n2144 ) ;
  assign n11883 = n11882 ^ n6135 ^ n818 ;
  assign n11889 = ( n3959 & n4625 ) | ( n3959 & ~n10444 ) | ( n4625 & ~n10444 ) ;
  assign n11884 = n7714 ^ n6325 ^ n3363 ;
  assign n11885 = n11884 ^ n3934 ^ n2572 ;
  assign n11886 = ( ~n746 & n2452 ) | ( ~n746 & n11885 ) | ( n2452 & n11885 ) ;
  assign n11887 = ( n7093 & ~n11245 ) | ( n7093 & n11886 ) | ( ~n11245 & n11886 ) ;
  assign n11888 = n11887 ^ n10120 ^ n8450 ;
  assign n11890 = n11889 ^ n11888 ^ n3904 ;
  assign n11891 = ( ~n8315 & n11883 ) | ( ~n8315 & n11890 ) | ( n11883 & n11890 ) ;
  assign n11881 = ( n626 & n1050 ) | ( n626 & n6949 ) | ( n1050 & n6949 ) ;
  assign n11892 = n11891 ^ n11881 ^ n9956 ;
  assign n11899 = ( ~n8058 & n11371 ) | ( ~n8058 & n11516 ) | ( n11371 & n11516 ) ;
  assign n11895 = n11560 ^ n7831 ^ n2589 ;
  assign n11893 = n2068 ^ n1781 ^ n565 ;
  assign n11894 = n11893 ^ n9858 ^ n1602 ;
  assign n11896 = n11895 ^ n11894 ^ n9441 ;
  assign n11897 = n11896 ^ n10390 ^ n10224 ;
  assign n11898 = ( n6769 & n11849 ) | ( n6769 & ~n11897 ) | ( n11849 & ~n11897 ) ;
  assign n11900 = n11899 ^ n11898 ^ n959 ;
  assign n11901 = n7743 ^ n7317 ^ n6475 ;
  assign n11902 = ( n8253 & ~n10431 ) | ( n8253 & n11901 ) | ( ~n10431 & n11901 ) ;
  assign n11903 = ( ~n1169 & n1712 ) | ( ~n1169 & n6321 ) | ( n1712 & n6321 ) ;
  assign n11904 = ( ~n6520 & n10874 ) | ( ~n6520 & n11903 ) | ( n10874 & n11903 ) ;
  assign n11905 = ( n838 & n3588 ) | ( n838 & n11904 ) | ( n3588 & n11904 ) ;
  assign n11906 = n9229 ^ n2502 ^ n1270 ;
  assign n11907 = n11906 ^ n3194 ^ n1764 ;
  assign n11910 = n5783 ^ n3531 ^ n3387 ;
  assign n11908 = n11765 ^ n4516 ^ n3829 ;
  assign n11909 = n11908 ^ n9068 ^ n3788 ;
  assign n11911 = n11910 ^ n11909 ^ n1047 ;
  assign n11912 = ( n10714 & n11907 ) | ( n10714 & n11911 ) | ( n11907 & n11911 ) ;
  assign n11913 = ( n1727 & n6404 ) | ( n1727 & n6913 ) | ( n6404 & n6913 ) ;
  assign n11914 = ( n8479 & ~n8686 ) | ( n8479 & n11913 ) | ( ~n8686 & n11913 ) ;
  assign n11916 = n5742 ^ n5696 ^ n3170 ;
  assign n11915 = ( ~n3752 & n4952 ) | ( ~n3752 & n8200 ) | ( n4952 & n8200 ) ;
  assign n11917 = n11916 ^ n11915 ^ n1670 ;
  assign n11918 = ( n7344 & n11914 ) | ( n7344 & ~n11917 ) | ( n11914 & ~n11917 ) ;
  assign n11928 = ( n3432 & n7008 ) | ( n3432 & n10353 ) | ( n7008 & n10353 ) ;
  assign n11926 = ( n3801 & ~n4248 ) | ( n3801 & n4627 ) | ( ~n4248 & n4627 ) ;
  assign n11925 = n10438 ^ n2861 ^ n915 ;
  assign n11927 = n11926 ^ n11925 ^ n5692 ;
  assign n11919 = ( n1805 & n3691 ) | ( n1805 & ~n10167 ) | ( n3691 & ~n10167 ) ;
  assign n11920 = ( ~n5713 & n6869 ) | ( ~n5713 & n7654 ) | ( n6869 & n7654 ) ;
  assign n11921 = ( ~n9226 & n11919 ) | ( ~n9226 & n11920 ) | ( n11919 & n11920 ) ;
  assign n11922 = n3586 ^ n1638 ^ n525 ;
  assign n11923 = ( n10713 & ~n11040 ) | ( n10713 & n11922 ) | ( ~n11040 & n11922 ) ;
  assign n11924 = ( ~n9098 & n11921 ) | ( ~n9098 & n11923 ) | ( n11921 & n11923 ) ;
  assign n11929 = n11928 ^ n11927 ^ n11924 ;
  assign n11930 = ( x67 & n3624 ) | ( x67 & n4750 ) | ( n3624 & n4750 ) ;
  assign n11937 = ( n5862 & n5980 ) | ( n5862 & ~n7132 ) | ( n5980 & ~n7132 ) ;
  assign n11934 = n5728 ^ n4729 ^ n4433 ;
  assign n11932 = n4483 ^ n318 ^ n254 ;
  assign n11933 = n11932 ^ n8696 ^ n1450 ;
  assign n11935 = n11934 ^ n11933 ^ n5753 ;
  assign n11931 = ( n1470 & n4410 ) | ( n1470 & n5463 ) | ( n4410 & n5463 ) ;
  assign n11936 = n11935 ^ n11933 ^ n11931 ;
  assign n11938 = n11937 ^ n11936 ^ n5514 ;
  assign n11941 = n7912 ^ n1039 ^ n184 ;
  assign n11942 = n11941 ^ n7966 ^ n6079 ;
  assign n11939 = ( n1173 & n4572 ) | ( n1173 & ~n9806 ) | ( n4572 & ~n9806 ) ;
  assign n11940 = ( n2325 & ~n4558 ) | ( n2325 & n11939 ) | ( ~n4558 & n11939 ) ;
  assign n11943 = n11942 ^ n11940 ^ n9868 ;
  assign n11947 = ( n4827 & n7585 ) | ( n4827 & ~n11932 ) | ( n7585 & ~n11932 ) ;
  assign n11948 = ( n452 & ~n2540 ) | ( n452 & n8099 ) | ( ~n2540 & n8099 ) ;
  assign n11949 = ( ~n7678 & n11947 ) | ( ~n7678 & n11948 ) | ( n11947 & n11948 ) ;
  assign n11945 = n7024 ^ n2875 ^ n1365 ;
  assign n11944 = ( n6761 & n9222 ) | ( n6761 & ~n9917 ) | ( n9222 & ~n9917 ) ;
  assign n11946 = n11945 ^ n11944 ^ n992 ;
  assign n11950 = n11949 ^ n11946 ^ n3049 ;
  assign n11951 = n11950 ^ n7547 ^ n857 ;
  assign n11952 = n11092 ^ n5968 ^ n1905 ;
  assign n11953 = n11952 ^ n8756 ^ n7795 ;
  assign n11954 = ( n1931 & n3328 ) | ( n1931 & n11953 ) | ( n3328 & n11953 ) ;
  assign n11955 = n9089 ^ n6556 ^ n3666 ;
  assign n11956 = ( n5787 & n9414 ) | ( n5787 & ~n9924 ) | ( n9414 & ~n9924 ) ;
  assign n11957 = ( n11658 & ~n11955 ) | ( n11658 & n11956 ) | ( ~n11955 & n11956 ) ;
  assign n11958 = ( ~n212 & n10963 ) | ( ~n212 & n11957 ) | ( n10963 & n11957 ) ;
  assign n11959 = n11958 ^ n7922 ^ n146 ;
  assign n11960 = n4628 ^ n4249 ^ n2872 ;
  assign n11961 = ( n3332 & ~n11418 ) | ( n3332 & n11960 ) | ( ~n11418 & n11960 ) ;
  assign n11962 = n11961 ^ n8775 ^ n5161 ;
  assign n11964 = n6114 ^ n3865 ^ n3728 ;
  assign n11963 = ( ~n736 & n4357 ) | ( ~n736 & n5566 ) | ( n4357 & n5566 ) ;
  assign n11965 = n11964 ^ n11963 ^ n161 ;
  assign n11966 = ( ~n4541 & n8854 ) | ( ~n4541 & n11965 ) | ( n8854 & n11965 ) ;
  assign n11967 = ( x110 & ~n2052 ) | ( x110 & n9587 ) | ( ~n2052 & n9587 ) ;
  assign n11968 = ( ~n2606 & n5858 ) | ( ~n2606 & n11967 ) | ( n5858 & n11967 ) ;
  assign n11969 = ( n2660 & ~n5350 ) | ( n2660 & n5522 ) | ( ~n5350 & n5522 ) ;
  assign n11970 = ( ~n2666 & n4324 ) | ( ~n2666 & n4811 ) | ( n4324 & n4811 ) ;
  assign n11971 = ( n6928 & n11969 ) | ( n6928 & ~n11970 ) | ( n11969 & ~n11970 ) ;
  assign n11975 = n7447 ^ n4339 ^ n252 ;
  assign n11976 = ( n2341 & ~n10763 ) | ( n2341 & n11975 ) | ( ~n10763 & n11975 ) ;
  assign n11973 = ( n4927 & n6237 ) | ( n4927 & ~n8561 ) | ( n6237 & ~n8561 ) ;
  assign n11972 = ( ~n2337 & n3848 ) | ( ~n2337 & n11363 ) | ( n3848 & n11363 ) ;
  assign n11974 = n11973 ^ n11972 ^ n5123 ;
  assign n11977 = n11976 ^ n11974 ^ n9001 ;
  assign n11978 = n4011 ^ n2631 ^ n2476 ;
  assign n11979 = ( n1037 & n11428 ) | ( n1037 & ~n11978 ) | ( n11428 & ~n11978 ) ;
  assign n11987 = ( n6876 & ~n7832 ) | ( n6876 & n8396 ) | ( ~n7832 & n8396 ) ;
  assign n11988 = ( n814 & n10142 ) | ( n814 & n11987 ) | ( n10142 & n11987 ) ;
  assign n11985 = n1679 ^ n855 ^ n624 ;
  assign n11982 = n3978 ^ n2704 ^ n798 ;
  assign n11981 = ( ~n772 & n1400 ) | ( ~n772 & n3275 ) | ( n1400 & n3275 ) ;
  assign n11980 = n6292 ^ n304 ^ n177 ;
  assign n11983 = n11982 ^ n11981 ^ n11980 ;
  assign n11984 = n11983 ^ n10649 ^ n2576 ;
  assign n11986 = n11985 ^ n11984 ^ n3053 ;
  assign n11989 = n11988 ^ n11986 ^ n1097 ;
  assign n11990 = n3022 ^ n1142 ^ n209 ;
  assign n11991 = n11990 ^ n7646 ^ x84 ;
  assign n11992 = ( ~n1936 & n6107 ) | ( ~n1936 & n9224 ) | ( n6107 & n9224 ) ;
  assign n11993 = n10697 ^ n4950 ^ n290 ;
  assign n11994 = n11278 ^ n10880 ^ n804 ;
  assign n11995 = ( n2091 & n2896 ) | ( n2091 & n3349 ) | ( n2896 & n3349 ) ;
  assign n11996 = ( ~n5678 & n11994 ) | ( ~n5678 & n11995 ) | ( n11994 & n11995 ) ;
  assign n11997 = ( ~n559 & n11993 ) | ( ~n559 & n11996 ) | ( n11993 & n11996 ) ;
  assign n11998 = ( n831 & n2829 ) | ( n831 & ~n10275 ) | ( n2829 & ~n10275 ) ;
  assign n11999 = ( n1547 & ~n4449 ) | ( n1547 & n9711 ) | ( ~n4449 & n9711 ) ;
  assign n12000 = n11999 ^ n8306 ^ n2885 ;
  assign n12001 = ( ~n1489 & n11998 ) | ( ~n1489 & n12000 ) | ( n11998 & n12000 ) ;
  assign n12002 = ( n2928 & ~n11997 ) | ( n2928 & n12001 ) | ( ~n11997 & n12001 ) ;
  assign n12003 = ( n3589 & n5436 ) | ( n3589 & n12002 ) | ( n5436 & n12002 ) ;
  assign n12004 = n4352 ^ n1234 ^ n181 ;
  assign n12005 = ( ~x22 & n8064 ) | ( ~x22 & n12004 ) | ( n8064 & n12004 ) ;
  assign n12006 = ( n7683 & ~n10100 ) | ( n7683 & n12005 ) | ( ~n10100 & n12005 ) ;
  assign n12007 = ( n3806 & n7041 ) | ( n3806 & n8095 ) | ( n7041 & n8095 ) ;
  assign n12008 = n9145 ^ n3239 ^ n1821 ;
  assign n12009 = ( ~n1144 & n11982 ) | ( ~n1144 & n12008 ) | ( n11982 & n12008 ) ;
  assign n12010 = ( n430 & n5228 ) | ( n430 & n7945 ) | ( n5228 & n7945 ) ;
  assign n12011 = n2142 ^ n2099 ^ n1553 ;
  assign n12012 = ( n5492 & n9003 ) | ( n5492 & n12011 ) | ( n9003 & n12011 ) ;
  assign n12013 = ( n1956 & n4542 ) | ( n1956 & n12012 ) | ( n4542 & n12012 ) ;
  assign n12014 = ( ~n11130 & n12010 ) | ( ~n11130 & n12013 ) | ( n12010 & n12013 ) ;
  assign n12015 = n6064 ^ n5279 ^ n3793 ;
  assign n12016 = ( n829 & ~n7747 ) | ( n829 & n12015 ) | ( ~n7747 & n12015 ) ;
  assign n12017 = n2998 ^ n1645 ^ n1547 ;
  assign n12018 = n6617 ^ n4818 ^ n4662 ;
  assign n12019 = ( ~n1272 & n9500 ) | ( ~n1272 & n12018 ) | ( n9500 & n12018 ) ;
  assign n12020 = ( n5526 & n12017 ) | ( n5526 & n12019 ) | ( n12017 & n12019 ) ;
  assign n12021 = ( ~n1782 & n12016 ) | ( ~n1782 & n12020 ) | ( n12016 & n12020 ) ;
  assign n12022 = ( n4481 & n6752 ) | ( n4481 & n6941 ) | ( n6752 & n6941 ) ;
  assign n12023 = n12022 ^ n10969 ^ n8818 ;
  assign n12026 = ( ~n905 & n8058 ) | ( ~n905 & n9278 ) | ( n8058 & n9278 ) ;
  assign n12024 = n11426 ^ n10466 ^ n2562 ;
  assign n12025 = n12024 ^ n10910 ^ n6447 ;
  assign n12027 = n12026 ^ n12025 ^ n1887 ;
  assign n12028 = ( n1877 & n6655 ) | ( n1877 & n7671 ) | ( n6655 & n7671 ) ;
  assign n12029 = ( ~n995 & n3361 ) | ( ~n995 & n12028 ) | ( n3361 & n12028 ) ;
  assign n12030 = n10191 ^ n4376 ^ n4275 ;
  assign n12031 = ( ~n612 & n12029 ) | ( ~n612 & n12030 ) | ( n12029 & n12030 ) ;
  assign n12032 = ( ~n5999 & n6012 ) | ( ~n5999 & n10938 ) | ( n6012 & n10938 ) ;
  assign n12034 = n7099 ^ n6822 ^ n4052 ;
  assign n12033 = n10878 ^ n9401 ^ n5263 ;
  assign n12035 = n12034 ^ n12033 ^ n10855 ;
  assign n12036 = n9629 ^ n6262 ^ n2128 ;
  assign n12037 = n12036 ^ n10266 ^ n273 ;
  assign n12038 = n6830 ^ n4153 ^ n2303 ;
  assign n12039 = n12038 ^ n10193 ^ n8695 ;
  assign n12040 = ( n2466 & n6248 ) | ( n2466 & ~n12039 ) | ( n6248 & ~n12039 ) ;
  assign n12041 = ( n6047 & n12037 ) | ( n6047 & ~n12040 ) | ( n12037 & ~n12040 ) ;
  assign n12042 = n7598 ^ n2642 ^ n1908 ;
  assign n12043 = ( ~n5854 & n8754 ) | ( ~n5854 & n12042 ) | ( n8754 & n12042 ) ;
  assign n12044 = n4584 ^ n1653 ^ n1612 ;
  assign n12045 = n12044 ^ n3155 ^ n903 ;
  assign n12046 = n9264 ^ n6773 ^ n3617 ;
  assign n12047 = ( n7597 & ~n12045 ) | ( n7597 & n12046 ) | ( ~n12045 & n12046 ) ;
  assign n12048 = n12047 ^ n9053 ^ n8332 ;
  assign n12049 = n11556 ^ n7522 ^ n3357 ;
  assign n12055 = n10340 ^ n7114 ^ n1600 ;
  assign n12051 = ( n137 & n894 ) | ( n137 & ~n4932 ) | ( n894 & ~n4932 ) ;
  assign n12052 = ( n464 & ~n7494 ) | ( n464 & n12051 ) | ( ~n7494 & n12051 ) ;
  assign n12053 = n12052 ^ n5922 ^ x89 ;
  assign n12054 = n12053 ^ n6320 ^ n1787 ;
  assign n12050 = n9065 ^ n7098 ^ n6397 ;
  assign n12056 = n12055 ^ n12054 ^ n12050 ;
  assign n12057 = ( n417 & n7158 ) | ( n417 & ~n12056 ) | ( n7158 & ~n12056 ) ;
  assign n12058 = ( n409 & n503 ) | ( n409 & n2161 ) | ( n503 & n2161 ) ;
  assign n12059 = ( n4604 & ~n7251 ) | ( n4604 & n12058 ) | ( ~n7251 & n12058 ) ;
  assign n12060 = ( n8160 & n11245 ) | ( n8160 & n12059 ) | ( n11245 & n12059 ) ;
  assign n12061 = ( n2859 & ~n3668 ) | ( n2859 & n4775 ) | ( ~n3668 & n4775 ) ;
  assign n12066 = n9658 ^ n5256 ^ n1156 ;
  assign n12067 = ( ~n890 & n1008 ) | ( ~n890 & n12066 ) | ( n1008 & n12066 ) ;
  assign n12065 = n8283 ^ n5727 ^ n2834 ;
  assign n12063 = ( ~n3353 & n5476 ) | ( ~n3353 & n7939 ) | ( n5476 & n7939 ) ;
  assign n12062 = ( n2826 & n5601 ) | ( n2826 & n6869 ) | ( n5601 & n6869 ) ;
  assign n12064 = n12063 ^ n12062 ^ n10754 ;
  assign n12068 = n12067 ^ n12065 ^ n12064 ;
  assign n12069 = ( n8670 & ~n12061 ) | ( n8670 & n12068 ) | ( ~n12061 & n12068 ) ;
  assign n12070 = n8245 ^ n8060 ^ n6217 ;
  assign n12071 = ( ~n1380 & n1922 ) | ( ~n1380 & n12070 ) | ( n1922 & n12070 ) ;
  assign n12072 = ( n5058 & ~n6894 ) | ( n5058 & n12071 ) | ( ~n6894 & n12071 ) ;
  assign n12073 = ( n1649 & ~n3425 ) | ( n1649 & n12072 ) | ( ~n3425 & n12072 ) ;
  assign n12074 = n6003 ^ n2737 ^ n2431 ;
  assign n12075 = n12074 ^ n4976 ^ n1767 ;
  assign n12078 = ( n971 & ~n5345 ) | ( n971 & n6439 ) | ( ~n5345 & n6439 ) ;
  assign n12076 = ( n1954 & n7651 ) | ( n1954 & ~n10264 ) | ( n7651 & ~n10264 ) ;
  assign n12077 = ( n998 & ~n10353 ) | ( n998 & n12076 ) | ( ~n10353 & n12076 ) ;
  assign n12079 = n12078 ^ n12077 ^ n10189 ;
  assign n12080 = ( n5233 & n9283 ) | ( n5233 & ~n12079 ) | ( n9283 & ~n12079 ) ;
  assign n12081 = n11557 ^ n2351 ^ n729 ;
  assign n12082 = ( n1011 & ~n1510 ) | ( n1011 & n4026 ) | ( ~n1510 & n4026 ) ;
  assign n12083 = n11715 ^ n8396 ^ n2387 ;
  assign n12084 = ( n7818 & n12082 ) | ( n7818 & ~n12083 ) | ( n12082 & ~n12083 ) ;
  assign n12085 = ( n4527 & n7202 ) | ( n4527 & ~n12084 ) | ( n7202 & ~n12084 ) ;
  assign n12086 = ( ~n833 & n3761 ) | ( ~n833 & n7262 ) | ( n3761 & n7262 ) ;
  assign n12089 = ( x30 & n1794 ) | ( x30 & n3316 ) | ( n1794 & n3316 ) ;
  assign n12090 = n12089 ^ n6314 ^ n1643 ;
  assign n12091 = n12090 ^ n11123 ^ n4019 ;
  assign n12087 = n7780 ^ n2654 ^ n2568 ;
  assign n12088 = ( ~n931 & n8730 ) | ( ~n931 & n12087 ) | ( n8730 & n12087 ) ;
  assign n12092 = n12091 ^ n12088 ^ n706 ;
  assign n12093 = ( n5706 & n6359 ) | ( n5706 & n10844 ) | ( n6359 & n10844 ) ;
  assign n12107 = ( ~n137 & n614 ) | ( ~n137 & n4953 ) | ( n614 & n4953 ) ;
  assign n12108 = ( ~n3989 & n5624 ) | ( ~n3989 & n6660 ) | ( n5624 & n6660 ) ;
  assign n12109 = ( n2914 & ~n12107 ) | ( n2914 & n12108 ) | ( ~n12107 & n12108 ) ;
  assign n12110 = n12109 ^ n9689 ^ n921 ;
  assign n12094 = ( n2629 & n8633 ) | ( n2629 & n10690 ) | ( n8633 & n10690 ) ;
  assign n12095 = ( ~n4207 & n5174 ) | ( ~n4207 & n12094 ) | ( n5174 & n12094 ) ;
  assign n12096 = n12095 ^ n4303 ^ n3385 ;
  assign n12100 = ( x98 & ~n1610 ) | ( x98 & n1835 ) | ( ~n1610 & n1835 ) ;
  assign n12101 = ( ~n947 & n2766 ) | ( ~n947 & n12100 ) | ( n2766 & n12100 ) ;
  assign n12102 = ( n7186 & n8456 ) | ( n7186 & ~n12101 ) | ( n8456 & ~n12101 ) ;
  assign n12103 = n12102 ^ n10071 ^ n8295 ;
  assign n12104 = ( n350 & n6410 ) | ( n350 & ~n12103 ) | ( n6410 & ~n12103 ) ;
  assign n12097 = n3936 ^ n1396 ^ n767 ;
  assign n12098 = n12097 ^ n10913 ^ n3950 ;
  assign n12099 = ( ~n3908 & n11870 ) | ( ~n3908 & n12098 ) | ( n11870 & n12098 ) ;
  assign n12105 = n12104 ^ n12099 ^ n4364 ;
  assign n12106 = ( n5554 & n12096 ) | ( n5554 & ~n12105 ) | ( n12096 & ~n12105 ) ;
  assign n12111 = n12110 ^ n12106 ^ n875 ;
  assign n12112 = n6227 ^ n5144 ^ n1620 ;
  assign n12113 = n12112 ^ n10724 ^ n4313 ;
  assign n12114 = ( n182 & n4777 ) | ( n182 & ~n8358 ) | ( n4777 & ~n8358 ) ;
  assign n12115 = ( ~n191 & n2388 ) | ( ~n191 & n2771 ) | ( n2388 & n2771 ) ;
  assign n12116 = n12115 ^ n10282 ^ n2129 ;
  assign n12117 = ( n10658 & n12114 ) | ( n10658 & ~n12116 ) | ( n12114 & ~n12116 ) ;
  assign n12118 = n11666 ^ n6019 ^ n5967 ;
  assign n12119 = n12118 ^ n10877 ^ n1952 ;
  assign n12120 = ( ~n2498 & n6558 ) | ( ~n2498 & n12119 ) | ( n6558 & n12119 ) ;
  assign n12121 = n3667 ^ n2901 ^ n1636 ;
  assign n12122 = ( n989 & n4488 ) | ( n989 & ~n5025 ) | ( n4488 & ~n5025 ) ;
  assign n12123 = ( n8863 & ~n12121 ) | ( n8863 & n12122 ) | ( ~n12121 & n12122 ) ;
  assign n12124 = ( n4041 & n6356 ) | ( n4041 & n12123 ) | ( n6356 & n12123 ) ;
  assign n12126 = n3936 ^ n2404 ^ n201 ;
  assign n12125 = n9774 ^ n5067 ^ n3849 ;
  assign n12127 = n12126 ^ n12125 ^ n5239 ;
  assign n12128 = ( n3889 & ~n7755 ) | ( n3889 & n10945 ) | ( ~n7755 & n10945 ) ;
  assign n12129 = n6189 ^ n2907 ^ n470 ;
  assign n12130 = ( n1871 & n10199 ) | ( n1871 & n11618 ) | ( n10199 & n11618 ) ;
  assign n12131 = n11680 ^ n3523 ^ n2511 ;
  assign n12133 = n5138 ^ n1888 ^ n540 ;
  assign n12132 = n2945 ^ n435 ^ n207 ;
  assign n12134 = n12133 ^ n12132 ^ n2012 ;
  assign n12135 = n3112 ^ n1910 ^ n638 ;
  assign n12136 = n12135 ^ n2492 ^ n487 ;
  assign n12137 = n12136 ^ n4104 ^ n2365 ;
  assign n12138 = ( n1343 & n3909 ) | ( n1343 & ~n11407 ) | ( n3909 & ~n11407 ) ;
  assign n12139 = ( n10137 & n12137 ) | ( n10137 & ~n12138 ) | ( n12137 & ~n12138 ) ;
  assign n12140 = ( n3925 & n12134 ) | ( n3925 & n12139 ) | ( n12134 & n12139 ) ;
  assign n12141 = ( n12130 & n12131 ) | ( n12130 & n12140 ) | ( n12131 & n12140 ) ;
  assign n12142 = n8688 ^ n4003 ^ n741 ;
  assign n12143 = ( n859 & n7715 ) | ( n859 & ~n12142 ) | ( n7715 & ~n12142 ) ;
  assign n12144 = ( n8900 & n10175 ) | ( n8900 & n12143 ) | ( n10175 & n12143 ) ;
  assign n12150 = ( n1547 & n4344 ) | ( n1547 & n5378 ) | ( n4344 & n5378 ) ;
  assign n12151 = ( n1791 & ~n5337 ) | ( n1791 & n12150 ) | ( ~n5337 & n12150 ) ;
  assign n12145 = ( ~n2673 & n3756 ) | ( ~n2673 & n11019 ) | ( n3756 & n11019 ) ;
  assign n12146 = n12145 ^ n11166 ^ n1796 ;
  assign n12147 = ( n577 & n1213 ) | ( n577 & n3882 ) | ( n1213 & n3882 ) ;
  assign n12148 = ( n4580 & ~n8690 ) | ( n4580 & n12147 ) | ( ~n8690 & n12147 ) ;
  assign n12149 = ( n4527 & n12146 ) | ( n4527 & ~n12148 ) | ( n12146 & ~n12148 ) ;
  assign n12152 = n12151 ^ n12149 ^ n8998 ;
  assign n12156 = ( n2081 & n2444 ) | ( n2081 & n7374 ) | ( n2444 & n7374 ) ;
  assign n12153 = n10035 ^ n3129 ^ n768 ;
  assign n12154 = n12153 ^ n8061 ^ n1156 ;
  assign n12155 = ( n4104 & n4145 ) | ( n4104 & n12154 ) | ( n4145 & n12154 ) ;
  assign n12157 = n12156 ^ n12155 ^ n10403 ;
  assign n12160 = n4354 ^ n4021 ^ n677 ;
  assign n12158 = ( x110 & n534 ) | ( x110 & n4176 ) | ( n534 & n4176 ) ;
  assign n12159 = ( n664 & n5058 ) | ( n664 & ~n12158 ) | ( n5058 & ~n12158 ) ;
  assign n12161 = n12160 ^ n12159 ^ n3227 ;
  assign n12165 = n5039 ^ n4618 ^ n2111 ;
  assign n12163 = ( n4597 & n5826 ) | ( n4597 & n9574 ) | ( n5826 & n9574 ) ;
  assign n12162 = n9268 ^ n3517 ^ n2403 ;
  assign n12164 = n12163 ^ n12162 ^ n8506 ;
  assign n12166 = n12165 ^ n12164 ^ n9017 ;
  assign n12167 = n10521 ^ n8257 ^ n411 ;
  assign n12168 = n12167 ^ n9289 ^ n8576 ;
  assign n12169 = ( n4160 & ~n9181 ) | ( n4160 & n12168 ) | ( ~n9181 & n12168 ) ;
  assign n12170 = n3477 ^ n1360 ^ n238 ;
  assign n12171 = ( n3268 & n6110 ) | ( n3268 & n12170 ) | ( n6110 & n12170 ) ;
  assign n12172 = ( n1412 & n1789 ) | ( n1412 & ~n6803 ) | ( n1789 & ~n6803 ) ;
  assign n12173 = n12172 ^ n9358 ^ n7388 ;
  assign n12174 = n12173 ^ n1490 ^ n1437 ;
  assign n12175 = ( n11017 & ~n12171 ) | ( n11017 & n12174 ) | ( ~n12171 & n12174 ) ;
  assign n12176 = n6044 ^ n4608 ^ n161 ;
  assign n12178 = n7996 ^ n4424 ^ n1278 ;
  assign n12177 = n10241 ^ n7297 ^ n1438 ;
  assign n12179 = n12178 ^ n12177 ^ n10026 ;
  assign n12180 = ( n6047 & n9891 ) | ( n6047 & n12179 ) | ( n9891 & n12179 ) ;
  assign n12184 = n3808 ^ n2787 ^ n2481 ;
  assign n12181 = ( n5317 & ~n6148 ) | ( n5317 & n10844 ) | ( ~n6148 & n10844 ) ;
  assign n12182 = n12181 ^ n4744 ^ n3107 ;
  assign n12183 = n12182 ^ n10589 ^ n6082 ;
  assign n12185 = n12184 ^ n12183 ^ n2949 ;
  assign n12186 = ( ~n3439 & n3824 ) | ( ~n3439 & n12185 ) | ( n3824 & n12185 ) ;
  assign n12187 = n12186 ^ n7206 ^ n3285 ;
  assign n12188 = ( n11686 & ~n12180 ) | ( n11686 & n12187 ) | ( ~n12180 & n12187 ) ;
  assign n12189 = n11718 ^ n7841 ^ n4669 ;
  assign n12190 = ( n1358 & n2039 ) | ( n1358 & ~n4891 ) | ( n2039 & ~n4891 ) ;
  assign n12191 = n12190 ^ n11677 ^ n1556 ;
  assign n12192 = ( n1062 & ~n3007 ) | ( n1062 & n6170 ) | ( ~n3007 & n6170 ) ;
  assign n12193 = ( n6341 & ~n11237 ) | ( n6341 & n12192 ) | ( ~n11237 & n12192 ) ;
  assign n12194 = ( n1301 & n2658 ) | ( n1301 & n3501 ) | ( n2658 & n3501 ) ;
  assign n12195 = n12194 ^ n5903 ^ n2666 ;
  assign n12196 = ( n9761 & ~n12193 ) | ( n9761 & n12195 ) | ( ~n12193 & n12195 ) ;
  assign n12197 = ( n627 & n9623 ) | ( n627 & ~n12196 ) | ( n9623 & ~n12196 ) ;
  assign n12198 = n12197 ^ n12148 ^ n3773 ;
  assign n12199 = n9696 ^ n5965 ^ n2092 ;
  assign n12200 = n11348 ^ n4484 ^ n2861 ;
  assign n12201 = ( n7389 & ~n8617 ) | ( n7389 & n8749 ) | ( ~n8617 & n8749 ) ;
  assign n12202 = n9225 ^ n1812 ^ n1062 ;
  assign n12205 = n11168 ^ n6023 ^ n1650 ;
  assign n12203 = n10867 ^ n8005 ^ n6982 ;
  assign n12204 = n12203 ^ n2408 ^ n974 ;
  assign n12206 = n12205 ^ n12204 ^ n1214 ;
  assign n12207 = n12206 ^ n7355 ^ n6381 ;
  assign n12208 = ( n5303 & n7134 ) | ( n5303 & n9772 ) | ( n7134 & n9772 ) ;
  assign n12209 = ( n175 & n3004 ) | ( n175 & n6788 ) | ( n3004 & n6788 ) ;
  assign n12211 = n6880 ^ n5734 ^ n1132 ;
  assign n12210 = ( n4407 & n6759 ) | ( n4407 & ~n9928 ) | ( n6759 & ~n9928 ) ;
  assign n12212 = n12211 ^ n12210 ^ n218 ;
  assign n12213 = n9573 ^ n3949 ^ n2183 ;
  assign n12214 = ( ~n1301 & n3811 ) | ( ~n1301 & n9256 ) | ( n3811 & n9256 ) ;
  assign n12215 = n12214 ^ n5171 ^ n600 ;
  assign n12216 = ( ~n1684 & n8009 ) | ( ~n1684 & n9775 ) | ( n8009 & n9775 ) ;
  assign n12217 = n12216 ^ n3676 ^ n394 ;
  assign n12218 = n12217 ^ n4084 ^ n1528 ;
  assign n12219 = n12218 ^ n3182 ^ n1163 ;
  assign n12220 = ( n12213 & n12215 ) | ( n12213 & n12219 ) | ( n12215 & n12219 ) ;
  assign n12221 = n4393 ^ n2458 ^ n1427 ;
  assign n12222 = ( x69 & ~n2308 ) | ( x69 & n12221 ) | ( ~n2308 & n12221 ) ;
  assign n12223 = ( n2990 & n11485 ) | ( n2990 & n12222 ) | ( n11485 & n12222 ) ;
  assign n12224 = ( ~n3705 & n5974 ) | ( ~n3705 & n9053 ) | ( n5974 & n9053 ) ;
  assign n12225 = ( n684 & n8996 ) | ( n684 & ~n12224 ) | ( n8996 & ~n12224 ) ;
  assign n12226 = n12225 ^ n10641 ^ n3953 ;
  assign n12227 = ( n5770 & n7839 ) | ( n5770 & ~n12226 ) | ( n7839 & ~n12226 ) ;
  assign n12228 = ( ~n1938 & n5504 ) | ( ~n1938 & n6366 ) | ( n5504 & n6366 ) ;
  assign n12229 = ( n2620 & n4469 ) | ( n2620 & n12228 ) | ( n4469 & n12228 ) ;
  assign n12230 = n12229 ^ n8783 ^ n8562 ;
  assign n12231 = n6054 ^ n3290 ^ n326 ;
  assign n12233 = n8073 ^ n6786 ^ n6039 ;
  assign n12232 = n11972 ^ n11002 ^ n3989 ;
  assign n12234 = n12233 ^ n12232 ^ n7382 ;
  assign n12235 = ( n948 & n6585 ) | ( n948 & ~n12012 ) | ( n6585 & ~n12012 ) ;
  assign n12236 = ( n1206 & n1224 ) | ( n1206 & ~n12235 ) | ( n1224 & ~n12235 ) ;
  assign n12237 = ( n12231 & ~n12234 ) | ( n12231 & n12236 ) | ( ~n12234 & n12236 ) ;
  assign n12245 = ( n1754 & n4659 ) | ( n1754 & ~n5199 ) | ( n4659 & ~n5199 ) ;
  assign n12241 = ( ~n1738 & n6495 ) | ( ~n1738 & n7420 ) | ( n6495 & n7420 ) ;
  assign n12240 = ( n5589 & n5754 ) | ( n5589 & ~n6366 ) | ( n5754 & ~n6366 ) ;
  assign n12242 = n12241 ^ n12240 ^ n4455 ;
  assign n12243 = ( x48 & ~n7097 ) | ( x48 & n12242 ) | ( ~n7097 & n12242 ) ;
  assign n12238 = n8474 ^ n5428 ^ n3592 ;
  assign n12239 = ( n8569 & n10704 ) | ( n8569 & ~n12238 ) | ( n10704 & ~n12238 ) ;
  assign n12244 = n12243 ^ n12239 ^ n6327 ;
  assign n12246 = n12245 ^ n12244 ^ n9451 ;
  assign n12247 = n2779 ^ n2130 ^ n1859 ;
  assign n12248 = n12247 ^ n2810 ^ n685 ;
  assign n12249 = n12248 ^ n9093 ^ n1967 ;
  assign n12250 = n12249 ^ n9451 ^ n3982 ;
  assign n12251 = n12250 ^ n10786 ^ n7674 ;
  assign n12252 = ( n609 & n2393 ) | ( n609 & n12251 ) | ( n2393 & n12251 ) ;
  assign n12253 = n5107 ^ n4207 ^ n148 ;
  assign n12254 = n9455 ^ n5219 ^ n1056 ;
  assign n12255 = ( ~n2051 & n12253 ) | ( ~n2051 & n12254 ) | ( n12253 & n12254 ) ;
  assign n12257 = n6882 ^ n2091 ^ n1271 ;
  assign n12256 = n7544 ^ n3425 ^ n2450 ;
  assign n12258 = n12257 ^ n12256 ^ n7681 ;
  assign n12259 = ( n5520 & n11741 ) | ( n5520 & ~n12258 ) | ( n11741 & ~n12258 ) ;
  assign n12261 = ( n3654 & n4977 ) | ( n3654 & ~n6200 ) | ( n4977 & ~n6200 ) ;
  assign n12260 = n8575 ^ n8176 ^ n4794 ;
  assign n12262 = n12261 ^ n12260 ^ n9189 ;
  assign n12265 = ( ~n2262 & n3873 ) | ( ~n2262 & n4458 ) | ( n3873 & n4458 ) ;
  assign n12263 = n3949 ^ n1234 ^ n295 ;
  assign n12264 = ( n5228 & ~n6579 ) | ( n5228 & n12263 ) | ( ~n6579 & n12263 ) ;
  assign n12266 = n12265 ^ n12264 ^ n9892 ;
  assign n12267 = ( n5978 & ~n8891 ) | ( n5978 & n10867 ) | ( ~n8891 & n10867 ) ;
  assign n12268 = ( n9425 & n9861 ) | ( n9425 & ~n12267 ) | ( n9861 & ~n12267 ) ;
  assign n12269 = ( n2357 & n2522 ) | ( n2357 & n7996 ) | ( n2522 & n7996 ) ;
  assign n12270 = ( n4288 & n7482 ) | ( n4288 & n12269 ) | ( n7482 & n12269 ) ;
  assign n12271 = ( n4568 & n7764 ) | ( n4568 & n12270 ) | ( n7764 & n12270 ) ;
  assign n12272 = ( ~n4133 & n8040 ) | ( ~n4133 & n12271 ) | ( n8040 & n12271 ) ;
  assign n12273 = n8175 ^ n2273 ^ n1636 ;
  assign n12274 = n8984 ^ n2343 ^ n1660 ;
  assign n12275 = ( n2242 & n8496 ) | ( n2242 & ~n11352 ) | ( n8496 & ~n11352 ) ;
  assign n12276 = ( ~n4055 & n8099 ) | ( ~n4055 & n12275 ) | ( n8099 & n12275 ) ;
  assign n12277 = ( ~x38 & x76 ) | ( ~x38 & n12276 ) | ( x76 & n12276 ) ;
  assign n12278 = n3088 ^ n2911 ^ n1452 ;
  assign n12279 = n12278 ^ n10508 ^ n1555 ;
  assign n12280 = ( ~n12274 & n12277 ) | ( ~n12274 & n12279 ) | ( n12277 & n12279 ) ;
  assign n12281 = n6020 ^ n3340 ^ n1882 ;
  assign n12282 = n11153 ^ n4321 ^ n1427 ;
  assign n12283 = ( n7048 & n12281 ) | ( n7048 & n12282 ) | ( n12281 & n12282 ) ;
  assign n12284 = ( n2009 & ~n3491 ) | ( n2009 & n3581 ) | ( ~n3491 & n3581 ) ;
  assign n12285 = ( n187 & n2893 ) | ( n187 & n12284 ) | ( n2893 & n12284 ) ;
  assign n12286 = n12285 ^ n11387 ^ n4187 ;
  assign n12287 = n7638 ^ n2189 ^ n2005 ;
  assign n12288 = n3718 ^ n3309 ^ n1345 ;
  assign n12289 = ( ~n459 & n12287 ) | ( ~n459 & n12288 ) | ( n12287 & n12288 ) ;
  assign n12290 = ( n4218 & n12286 ) | ( n4218 & n12289 ) | ( n12286 & n12289 ) ;
  assign n12297 = ( n2883 & ~n5813 ) | ( n2883 & n9831 ) | ( ~n5813 & n9831 ) ;
  assign n12293 = n7759 ^ n3543 ^ n424 ;
  assign n12294 = n12293 ^ n5674 ^ n4513 ;
  assign n12295 = n12294 ^ n9204 ^ n9068 ;
  assign n12291 = ( n4701 & n6142 ) | ( n4701 & n7454 ) | ( n6142 & n7454 ) ;
  assign n12292 = ( ~n549 & n11557 ) | ( ~n549 & n12291 ) | ( n11557 & n12291 ) ;
  assign n12296 = n12295 ^ n12292 ^ n3037 ;
  assign n12298 = n12297 ^ n12296 ^ n6458 ;
  assign n12299 = ( n6308 & n8738 ) | ( n6308 & n9024 ) | ( n8738 & n9024 ) ;
  assign n12300 = n11567 ^ n4238 ^ n399 ;
  assign n12301 = ( n4289 & n4346 ) | ( n4289 & ~n12300 ) | ( n4346 & ~n12300 ) ;
  assign n12302 = n12301 ^ n9392 ^ n9117 ;
  assign n12303 = n12302 ^ n4520 ^ n2540 ;
  assign n12304 = n12303 ^ n11035 ^ n4284 ;
  assign n12312 = n11779 ^ n8452 ^ n5736 ;
  assign n12305 = ( n3227 & ~n4796 ) | ( n3227 & n10387 ) | ( ~n4796 & n10387 ) ;
  assign n12306 = ( ~n1195 & n7852 ) | ( ~n1195 & n12305 ) | ( n7852 & n12305 ) ;
  assign n12307 = n12306 ^ n4482 ^ n751 ;
  assign n12308 = ( n2191 & n5079 ) | ( n2191 & n6734 ) | ( n5079 & n6734 ) ;
  assign n12309 = n4504 ^ n4083 ^ n3639 ;
  assign n12310 = ( n1157 & ~n12308 ) | ( n1157 & n12309 ) | ( ~n12308 & n12309 ) ;
  assign n12311 = ( n5938 & n12307 ) | ( n5938 & n12310 ) | ( n12307 & n12310 ) ;
  assign n12313 = n12312 ^ n12311 ^ n1673 ;
  assign n12314 = n7953 ^ n2099 ^ n479 ;
  assign n12315 = ( ~n9579 & n10819 ) | ( ~n9579 & n12314 ) | ( n10819 & n12314 ) ;
  assign n12318 = n5303 ^ n3473 ^ n1146 ;
  assign n12317 = n10431 ^ n7754 ^ n4790 ;
  assign n12316 = n5692 ^ n3700 ^ n878 ;
  assign n12319 = n12318 ^ n12317 ^ n12316 ;
  assign n12320 = n10017 ^ n5163 ^ n3749 ;
  assign n12321 = ( ~n1804 & n5255 ) | ( ~n1804 & n12320 ) | ( n5255 & n12320 ) ;
  assign n12322 = ( n5609 & n10090 ) | ( n5609 & n12321 ) | ( n10090 & n12321 ) ;
  assign n12324 = ( n3830 & n6252 ) | ( n3830 & ~n6552 ) | ( n6252 & ~n6552 ) ;
  assign n12325 = n7006 ^ n5777 ^ n5470 ;
  assign n12326 = ( ~n5475 & n12324 ) | ( ~n5475 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12323 = n6748 ^ n5686 ^ n1809 ;
  assign n12327 = n12326 ^ n12323 ^ n1001 ;
  assign n12328 = n11621 ^ n6199 ^ n5194 ;
  assign n12335 = ( n3701 & n4565 ) | ( n3701 & n8647 ) | ( n4565 & n8647 ) ;
  assign n12334 = ( ~n1555 & n4024 ) | ( ~n1555 & n9796 ) | ( n4024 & n9796 ) ;
  assign n12332 = ( n2524 & n5213 ) | ( n2524 & ~n11186 ) | ( n5213 & ~n11186 ) ;
  assign n12329 = n9794 ^ n8375 ^ n4070 ;
  assign n12330 = n8938 ^ n8912 ^ n7925 ;
  assign n12331 = ( n2526 & ~n12329 ) | ( n2526 & n12330 ) | ( ~n12329 & n12330 ) ;
  assign n12333 = n12332 ^ n12331 ^ n7620 ;
  assign n12336 = n12335 ^ n12334 ^ n12333 ;
  assign n12357 = n11811 ^ n8849 ^ n8238 ;
  assign n12353 = n5295 ^ n3943 ^ n3932 ;
  assign n12352 = ( ~x80 & n1776 ) | ( ~x80 & n3463 ) | ( n1776 & n3463 ) ;
  assign n12354 = n12353 ^ n12352 ^ n1858 ;
  assign n12355 = n10878 ^ n7753 ^ n1593 ;
  assign n12356 = ( n3226 & n12354 ) | ( n3226 & n12355 ) | ( n12354 & n12355 ) ;
  assign n12349 = n2407 ^ n433 ^ n359 ;
  assign n12350 = ( n2748 & n7725 ) | ( n2748 & ~n8565 ) | ( n7725 & ~n8565 ) ;
  assign n12351 = ( n3363 & ~n12349 ) | ( n3363 & n12350 ) | ( ~n12349 & n12350 ) ;
  assign n12358 = n12357 ^ n12356 ^ n12351 ;
  assign n12337 = ( n2012 & ~n5304 ) | ( n2012 & n8569 ) | ( ~n5304 & n8569 ) ;
  assign n12338 = n5518 ^ n5209 ^ n3997 ;
  assign n12339 = ( n1056 & n2105 ) | ( n1056 & ~n7908 ) | ( n2105 & ~n7908 ) ;
  assign n12340 = n12339 ^ n4529 ^ n519 ;
  assign n12341 = ( n6100 & n12338 ) | ( n6100 & ~n12340 ) | ( n12338 & ~n12340 ) ;
  assign n12344 = n6146 ^ n5140 ^ n803 ;
  assign n12343 = n8717 ^ n6974 ^ n6340 ;
  assign n12345 = n12344 ^ n12343 ^ n12260 ;
  assign n12342 = n5281 ^ n2872 ^ n2474 ;
  assign n12346 = n12345 ^ n12342 ^ n10012 ;
  assign n12347 = n12346 ^ n11767 ^ n5527 ;
  assign n12348 = ( n12337 & ~n12341 ) | ( n12337 & n12347 ) | ( ~n12341 & n12347 ) ;
  assign n12359 = n12358 ^ n12348 ^ n7666 ;
  assign n12360 = ( n368 & ~n396 ) | ( n368 & n5761 ) | ( ~n396 & n5761 ) ;
  assign n12361 = ( n5428 & n8512 ) | ( n5428 & n12360 ) | ( n8512 & n12360 ) ;
  assign n12362 = n10241 ^ n8556 ^ n7779 ;
  assign n12363 = ( n4037 & ~n7037 ) | ( n4037 & n11001 ) | ( ~n7037 & n11001 ) ;
  assign n12367 = ( n1298 & n2511 ) | ( n1298 & n7811 ) | ( n2511 & n7811 ) ;
  assign n12364 = n4158 ^ n2080 ^ n243 ;
  assign n12365 = ( n6865 & n9673 ) | ( n6865 & ~n10223 ) | ( n9673 & ~n10223 ) ;
  assign n12366 = ( n5320 & ~n12364 ) | ( n5320 & n12365 ) | ( ~n12364 & n12365 ) ;
  assign n12368 = n12367 ^ n12366 ^ n599 ;
  assign n12369 = ( n5620 & ~n8039 ) | ( n5620 & n12368 ) | ( ~n8039 & n12368 ) ;
  assign n12370 = n7090 ^ n6878 ^ n2585 ;
  assign n12373 = ( n707 & n1708 ) | ( n707 & n12247 ) | ( n1708 & n12247 ) ;
  assign n12371 = n8077 ^ n2664 ^ n490 ;
  assign n12372 = n12371 ^ n6622 ^ n691 ;
  assign n12374 = n12373 ^ n12372 ^ n592 ;
  assign n12375 = ( ~n7340 & n12370 ) | ( ~n7340 & n12374 ) | ( n12370 & n12374 ) ;
  assign n12376 = ( n5946 & ~n10489 ) | ( n5946 & n11393 ) | ( ~n10489 & n11393 ) ;
  assign n12377 = n12376 ^ n7274 ^ n6069 ;
  assign n12378 = ( n2605 & ~n11055 ) | ( n2605 & n12377 ) | ( ~n11055 & n12377 ) ;
  assign n12379 = ( ~n5486 & n9093 ) | ( ~n5486 & n9291 ) | ( n9093 & n9291 ) ;
  assign n12380 = ( n6965 & n10021 ) | ( n6965 & n12379 ) | ( n10021 & n12379 ) ;
  assign n12381 = n10249 ^ n10043 ^ n5211 ;
  assign n12382 = n10768 ^ n5194 ^ n3241 ;
  assign n12386 = n6574 ^ n1562 ^ n1111 ;
  assign n12384 = n2302 ^ x76 ^ x46 ;
  assign n12385 = ( n6609 & n9011 ) | ( n6609 & n12384 ) | ( n9011 & n12384 ) ;
  assign n12383 = n11621 ^ n5074 ^ n4770 ;
  assign n12387 = n12386 ^ n12385 ^ n12383 ;
  assign n12388 = n12387 ^ n9884 ^ n4821 ;
  assign n12389 = n12388 ^ n9747 ^ n4983 ;
  assign n12390 = n11449 ^ n6358 ^ n4170 ;
  assign n12391 = ( ~n2813 & n12074 ) | ( ~n2813 & n12390 ) | ( n12074 & n12390 ) ;
  assign n12392 = ( n160 & n3938 ) | ( n160 & ~n12391 ) | ( n3938 & ~n12391 ) ;
  assign n12393 = ( n6657 & n10502 ) | ( n6657 & n12392 ) | ( n10502 & n12392 ) ;
  assign n12394 = n5387 ^ n4469 ^ n2626 ;
  assign n12395 = ( n6649 & ~n10829 ) | ( n6649 & n12394 ) | ( ~n10829 & n12394 ) ;
  assign n12396 = ( n569 & n2462 ) | ( n569 & ~n11173 ) | ( n2462 & ~n11173 ) ;
  assign n12397 = ( n3144 & n4994 ) | ( n3144 & ~n12396 ) | ( n4994 & ~n12396 ) ;
  assign n12398 = ( ~n8523 & n12309 ) | ( ~n8523 & n12397 ) | ( n12309 & n12397 ) ;
  assign n12402 = n10940 ^ n10345 ^ n7325 ;
  assign n12399 = ( n1500 & n2408 ) | ( n1500 & n3071 ) | ( n2408 & n3071 ) ;
  assign n12400 = ( n1473 & n11372 ) | ( n1473 & ~n12399 ) | ( n11372 & ~n12399 ) ;
  assign n12401 = n12400 ^ n10198 ^ n6009 ;
  assign n12403 = n12402 ^ n12401 ^ n10522 ;
  assign n12404 = ( ~n6296 & n6513 ) | ( ~n6296 & n7474 ) | ( n6513 & n7474 ) ;
  assign n12405 = ( n3242 & n7352 ) | ( n3242 & ~n12404 ) | ( n7352 & ~n12404 ) ;
  assign n12406 = n10489 ^ n6856 ^ n558 ;
  assign n12407 = n12406 ^ n5997 ^ n3718 ;
  assign n12408 = ( n7958 & n12405 ) | ( n7958 & n12407 ) | ( n12405 & n12407 ) ;
  assign n12409 = n12408 ^ n12143 ^ n11175 ;
  assign n12410 = ( n3217 & n9389 ) | ( n3217 & ~n11223 ) | ( n9389 & ~n11223 ) ;
  assign n12411 = n12410 ^ n7647 ^ n3139 ;
  assign n12412 = n8902 ^ n5848 ^ n3631 ;
  assign n12413 = ( n3258 & ~n8250 ) | ( n3258 & n11582 ) | ( ~n8250 & n11582 ) ;
  assign n12414 = n7134 ^ n971 ^ n163 ;
  assign n12415 = ( n1603 & ~n2376 ) | ( n1603 & n12414 ) | ( ~n2376 & n12414 ) ;
  assign n12416 = n12285 ^ n5208 ^ n4556 ;
  assign n12417 = ( ~n11569 & n12415 ) | ( ~n11569 & n12416 ) | ( n12415 & n12416 ) ;
  assign n12418 = ( n2995 & n4821 ) | ( n2995 & n9093 ) | ( n4821 & n9093 ) ;
  assign n12419 = ( n6372 & n7727 ) | ( n6372 & ~n11538 ) | ( n7727 & ~n11538 ) ;
  assign n12420 = n4717 ^ n1079 ^ n397 ;
  assign n12421 = n12420 ^ n10077 ^ n402 ;
  assign n12422 = ( ~n1945 & n12419 ) | ( ~n1945 & n12421 ) | ( n12419 & n12421 ) ;
  assign n12423 = n12422 ^ n8148 ^ n7531 ;
  assign n12424 = n12017 ^ n11794 ^ n10193 ;
  assign n12425 = n12424 ^ n10961 ^ n3239 ;
  assign n12433 = ( ~n673 & n1201 ) | ( ~n673 & n5915 ) | ( n1201 & n5915 ) ;
  assign n12429 = n7548 ^ n5216 ^ n151 ;
  assign n12430 = n3620 ^ n1715 ^ n232 ;
  assign n12431 = ( ~n3843 & n12429 ) | ( ~n3843 & n12430 ) | ( n12429 & n12430 ) ;
  assign n12426 = ( n199 & n935 ) | ( n199 & n6933 ) | ( n935 & n6933 ) ;
  assign n12427 = ( n666 & n9228 ) | ( n666 & ~n12426 ) | ( n9228 & ~n12426 ) ;
  assign n12428 = ( n1542 & ~n12351 ) | ( n1542 & n12427 ) | ( ~n12351 & n12427 ) ;
  assign n12432 = n12431 ^ n12428 ^ n4214 ;
  assign n12434 = n12433 ^ n12432 ^ n2632 ;
  assign n12435 = ( ~n8760 & n8792 ) | ( ~n8760 & n10107 ) | ( n8792 & n10107 ) ;
  assign n12436 = ( x11 & n2588 ) | ( x11 & ~n12435 ) | ( n2588 & ~n12435 ) ;
  assign n12437 = ( ~n7312 & n9733 ) | ( ~n7312 & n12436 ) | ( n9733 & n12436 ) ;
  assign n12444 = n4158 ^ n2644 ^ n1369 ;
  assign n12442 = n10321 ^ n6898 ^ n4577 ;
  assign n12443 = ( n2957 & ~n7577 ) | ( n2957 & n12442 ) | ( ~n7577 & n12442 ) ;
  assign n12440 = n2212 ^ n2030 ^ x98 ;
  assign n12438 = n9124 ^ n2757 ^ n745 ;
  assign n12439 = n12438 ^ n7168 ^ n4235 ;
  assign n12441 = n12440 ^ n12439 ^ n9591 ;
  assign n12445 = n12444 ^ n12443 ^ n12441 ;
  assign n12450 = n6505 ^ n4435 ^ n130 ;
  assign n12446 = ( n666 & n4818 ) | ( n666 & n7403 ) | ( n4818 & n7403 ) ;
  assign n12447 = n5911 ^ n3240 ^ n2758 ;
  assign n12448 = ( n1124 & n3005 ) | ( n1124 & n12447 ) | ( n3005 & n12447 ) ;
  assign n12449 = ( n5225 & n12446 ) | ( n5225 & n12448 ) | ( n12446 & n12448 ) ;
  assign n12451 = n12450 ^ n12449 ^ n12407 ;
  assign n12452 = n11822 ^ n9319 ^ n1156 ;
  assign n12454 = ( ~n4774 & n7105 ) | ( ~n4774 & n7589 ) | ( n7105 & n7589 ) ;
  assign n12453 = n5842 ^ n3365 ^ n2235 ;
  assign n12455 = n12454 ^ n12453 ^ n8115 ;
  assign n12456 = ( n2050 & n10121 ) | ( n2050 & ~n10450 ) | ( n10121 & ~n10450 ) ;
  assign n12457 = ( ~n969 & n4313 ) | ( ~n969 & n12456 ) | ( n4313 & n12456 ) ;
  assign n12458 = n10396 ^ n9775 ^ n7296 ;
  assign n12459 = ( n11410 & n12457 ) | ( n11410 & ~n12458 ) | ( n12457 & ~n12458 ) ;
  assign n12460 = ( n6002 & n7884 ) | ( n6002 & ~n9877 ) | ( n7884 & ~n9877 ) ;
  assign n12461 = n9166 ^ n6319 ^ n3456 ;
  assign n12462 = ( n3297 & n10127 ) | ( n3297 & ~n12461 ) | ( n10127 & ~n12461 ) ;
  assign n12466 = ( ~n3198 & n5349 ) | ( ~n3198 & n5689 ) | ( n5349 & n5689 ) ;
  assign n12463 = n6119 ^ n3095 ^ n1352 ;
  assign n12464 = n12463 ^ n10561 ^ n1975 ;
  assign n12465 = ( ~n2802 & n4561 ) | ( ~n2802 & n12464 ) | ( n4561 & n12464 ) ;
  assign n12467 = n12466 ^ n12465 ^ n5742 ;
  assign n12471 = n10515 ^ n8905 ^ n1814 ;
  assign n12468 = ( n974 & n1673 ) | ( n974 & ~n7885 ) | ( n1673 & ~n7885 ) ;
  assign n12469 = ( ~n1295 & n3779 ) | ( ~n1295 & n12468 ) | ( n3779 & n12468 ) ;
  assign n12470 = ( ~n4307 & n10505 ) | ( ~n4307 & n12469 ) | ( n10505 & n12469 ) ;
  assign n12472 = n12471 ^ n12470 ^ n1988 ;
  assign n12473 = n4340 ^ n2666 ^ x111 ;
  assign n12474 = ( n3598 & ~n4283 ) | ( n3598 & n5612 ) | ( ~n4283 & n5612 ) ;
  assign n12475 = ( ~n7754 & n12473 ) | ( ~n7754 & n12474 ) | ( n12473 & n12474 ) ;
  assign n12476 = n10348 ^ n9800 ^ n766 ;
  assign n12478 = n6127 ^ n5695 ^ n4779 ;
  assign n12479 = n5314 ^ n4576 ^ n301 ;
  assign n12480 = ( n415 & n12478 ) | ( n415 & ~n12479 ) | ( n12478 & ~n12479 ) ;
  assign n12481 = ( ~n5164 & n5394 ) | ( ~n5164 & n12480 ) | ( n5394 & n12480 ) ;
  assign n12482 = n12481 ^ n5130 ^ n1894 ;
  assign n12477 = n4756 ^ n2925 ^ n2586 ;
  assign n12483 = n12482 ^ n12477 ^ n3359 ;
  assign n12484 = ( n12475 & n12476 ) | ( n12475 & n12483 ) | ( n12476 & n12483 ) ;
  assign n12485 = n10297 ^ n3154 ^ n326 ;
  assign n12486 = n12485 ^ n12341 ^ n8481 ;
  assign n12487 = ( n1676 & n1761 ) | ( n1676 & ~n3363 ) | ( n1761 & ~n3363 ) ;
  assign n12488 = ( n423 & n4648 ) | ( n423 & ~n12487 ) | ( n4648 & ~n12487 ) ;
  assign n12489 = ( n1463 & n10483 ) | ( n1463 & n12488 ) | ( n10483 & n12488 ) ;
  assign n12492 = ( n174 & ~n1840 ) | ( n174 & n4675 ) | ( ~n1840 & n4675 ) ;
  assign n12490 = ( n941 & ~n3502 ) | ( n941 & n7621 ) | ( ~n3502 & n7621 ) ;
  assign n12491 = ( n1896 & n5386 ) | ( n1896 & n12490 ) | ( n5386 & n12490 ) ;
  assign n12493 = n12492 ^ n12491 ^ n2147 ;
  assign n12494 = ( n4902 & ~n12384 ) | ( n4902 & n12493 ) | ( ~n12384 & n12493 ) ;
  assign n12495 = n4640 ^ n1798 ^ n1540 ;
  assign n12496 = ( n937 & ~n5823 ) | ( n937 & n12495 ) | ( ~n5823 & n12495 ) ;
  assign n12497 = ( n1529 & ~n4216 ) | ( n1529 & n12496 ) | ( ~n4216 & n12496 ) ;
  assign n12498 = ( n411 & ~n9530 ) | ( n411 & n11340 ) | ( ~n9530 & n11340 ) ;
  assign n12499 = ( n4037 & n5037 ) | ( n4037 & ~n12498 ) | ( n5037 & ~n12498 ) ;
  assign n12500 = ( ~n12494 & n12497 ) | ( ~n12494 & n12499 ) | ( n12497 & n12499 ) ;
  assign n12501 = ( n5279 & ~n6819 ) | ( n5279 & n9555 ) | ( ~n6819 & n9555 ) ;
  assign n12502 = ( ~n1600 & n5491 ) | ( ~n1600 & n7783 ) | ( n5491 & n7783 ) ;
  assign n12503 = ( n1694 & n6301 ) | ( n1694 & n9791 ) | ( n6301 & n9791 ) ;
  assign n12504 = n12503 ^ n6436 ^ n1660 ;
  assign n12505 = ( n2390 & ~n11650 ) | ( n2390 & n12504 ) | ( ~n11650 & n12504 ) ;
  assign n12509 = ( n3126 & n3221 ) | ( n3126 & ~n3619 ) | ( n3221 & ~n3619 ) ;
  assign n12508 = n8593 ^ n7123 ^ n4148 ;
  assign n12506 = ( n1853 & n2765 ) | ( n1853 & ~n10219 ) | ( n2765 & ~n10219 ) ;
  assign n12507 = n12506 ^ n2824 ^ n2092 ;
  assign n12510 = n12509 ^ n12508 ^ n12507 ;
  assign n12511 = ( n1449 & ~n5266 ) | ( n1449 & n7759 ) | ( ~n5266 & n7759 ) ;
  assign n12512 = ( n1162 & n10936 ) | ( n1162 & n12511 ) | ( n10936 & n12511 ) ;
  assign n12514 = n6109 ^ n2864 ^ n1108 ;
  assign n12513 = ( ~n2848 & n5425 ) | ( ~n2848 & n8329 ) | ( n5425 & n8329 ) ;
  assign n12515 = n12514 ^ n12513 ^ n270 ;
  assign n12518 = ( n974 & n6462 ) | ( n974 & n8207 ) | ( n6462 & n8207 ) ;
  assign n12516 = n6545 ^ n4181 ^ n1333 ;
  assign n12517 = n12516 ^ n5957 ^ n4412 ;
  assign n12519 = n12518 ^ n12517 ^ n5862 ;
  assign n12520 = ( ~n6258 & n7423 ) | ( ~n6258 & n8199 ) | ( n7423 & n8199 ) ;
  assign n12521 = ( ~n6064 & n7339 ) | ( ~n6064 & n7378 ) | ( n7339 & n7378 ) ;
  assign n12522 = ( n3353 & ~n6063 ) | ( n3353 & n8716 ) | ( ~n6063 & n8716 ) ;
  assign n12523 = ( n7569 & n11040 ) | ( n7569 & ~n12522 ) | ( n11040 & ~n12522 ) ;
  assign n12524 = n12523 ^ n8780 ^ n7199 ;
  assign n12525 = n12524 ^ n8382 ^ n3436 ;
  assign n12535 = n4919 ^ n2743 ^ n2724 ;
  assign n12536 = n5001 ^ n4461 ^ n4140 ;
  assign n12537 = ( n7776 & n12535 ) | ( n7776 & ~n12536 ) | ( n12535 & ~n12536 ) ;
  assign n12538 = ( n916 & n5151 ) | ( n916 & ~n12537 ) | ( n5151 & ~n12537 ) ;
  assign n12532 = ( n1343 & ~n5068 ) | ( n1343 & n5665 ) | ( ~n5068 & n5665 ) ;
  assign n12533 = n12532 ^ n4050 ^ n3113 ;
  assign n12526 = n3525 ^ n2633 ^ n2387 ;
  assign n12527 = ( n6120 & n12353 ) | ( n6120 & n12526 ) | ( n12353 & n12526 ) ;
  assign n12528 = ( n6074 & n6532 ) | ( n6074 & n12527 ) | ( n6532 & n12527 ) ;
  assign n12529 = n9954 ^ n9193 ^ n6690 ;
  assign n12530 = n12529 ^ n7572 ^ n4572 ;
  assign n12531 = ( ~n5266 & n12528 ) | ( ~n5266 & n12530 ) | ( n12528 & n12530 ) ;
  assign n12534 = n12533 ^ n12531 ^ n1421 ;
  assign n12539 = n12538 ^ n12534 ^ n3301 ;
  assign n12540 = n4865 ^ n3779 ^ n1450 ;
  assign n12541 = n11475 ^ n2772 ^ n2355 ;
  assign n12542 = n12541 ^ n12012 ^ n4331 ;
  assign n12543 = ( n8254 & ~n12540 ) | ( n8254 & n12542 ) | ( ~n12540 & n12542 ) ;
  assign n12549 = ( n780 & ~n827 ) | ( n780 & n8905 ) | ( ~n827 & n8905 ) ;
  assign n12547 = n8167 ^ n4599 ^ x28 ;
  assign n12548 = n12547 ^ n2435 ^ n165 ;
  assign n12545 = ( n856 & n2499 ) | ( n856 & ~n2780 ) | ( n2499 & ~n2780 ) ;
  assign n12544 = n3647 ^ n2856 ^ n1275 ;
  assign n12546 = n12545 ^ n12544 ^ n9068 ;
  assign n12550 = n12549 ^ n12548 ^ n12546 ;
  assign n12551 = n12096 ^ n6430 ^ n4699 ;
  assign n12553 = ( n4115 & ~n5482 ) | ( n4115 & n6581 ) | ( ~n5482 & n6581 ) ;
  assign n12552 = ( ~n1691 & n4313 ) | ( ~n1691 & n10365 ) | ( n4313 & n10365 ) ;
  assign n12554 = n12553 ^ n12552 ^ n6218 ;
  assign n12560 = n8105 ^ n5506 ^ n5013 ;
  assign n12555 = ( n4090 & ~n4093 ) | ( n4090 & n7010 ) | ( ~n4093 & n7010 ) ;
  assign n12556 = ( ~n5329 & n7886 ) | ( ~n5329 & n12555 ) | ( n7886 & n12555 ) ;
  assign n12557 = ( n4365 & n7502 ) | ( n4365 & n12556 ) | ( n7502 & n12556 ) ;
  assign n12558 = ( n1546 & n8634 ) | ( n1546 & ~n9702 ) | ( n8634 & ~n9702 ) ;
  assign n12559 = ( n1034 & ~n12557 ) | ( n1034 & n12558 ) | ( ~n12557 & n12558 ) ;
  assign n12561 = n12560 ^ n12559 ^ n3002 ;
  assign n12562 = n4172 ^ n2058 ^ n1035 ;
  assign n12563 = n5385 ^ n3507 ^ n957 ;
  assign n12564 = n12563 ^ n4157 ^ n1145 ;
  assign n12565 = ( n1407 & n8008 ) | ( n1407 & ~n12564 ) | ( n8008 & ~n12564 ) ;
  assign n12566 = n12565 ^ n2623 ^ n1242 ;
  assign n12567 = ( n10543 & ~n12562 ) | ( n10543 & n12566 ) | ( ~n12562 & n12566 ) ;
  assign n12574 = ( n906 & n5684 ) | ( n906 & ~n7780 ) | ( n5684 & ~n7780 ) ;
  assign n12575 = ( n2766 & ~n3067 ) | ( n2766 & n12182 ) | ( ~n3067 & n12182 ) ;
  assign n12576 = ( x45 & n2241 ) | ( x45 & ~n5483 ) | ( n2241 & ~n5483 ) ;
  assign n12577 = n12576 ^ n7108 ^ n4610 ;
  assign n12578 = ( n12574 & ~n12575 ) | ( n12574 & n12577 ) | ( ~n12575 & n12577 ) ;
  assign n12573 = n6333 ^ n1246 ^ n532 ;
  assign n12568 = n11769 ^ n6832 ^ n5991 ;
  assign n12569 = ( n454 & n1597 ) | ( n454 & ~n5896 ) | ( n1597 & ~n5896 ) ;
  assign n12570 = n12569 ^ n5973 ^ n1732 ;
  assign n12571 = ( n3551 & n12568 ) | ( n3551 & n12570 ) | ( n12568 & n12570 ) ;
  assign n12572 = n12571 ^ n3647 ^ n2889 ;
  assign n12579 = n12578 ^ n12573 ^ n12572 ;
  assign n12580 = n11640 ^ n6799 ^ n2649 ;
  assign n12581 = n4759 ^ n2010 ^ n982 ;
  assign n12582 = ( n2318 & n3387 ) | ( n2318 & ~n10391 ) | ( n3387 & ~n10391 ) ;
  assign n12583 = ( n1956 & n12581 ) | ( n1956 & n12582 ) | ( n12581 & n12582 ) ;
  assign n12584 = ( n4027 & n12580 ) | ( n4027 & ~n12583 ) | ( n12580 & ~n12583 ) ;
  assign n12591 = ( n5050 & n9287 ) | ( n5050 & n12042 ) | ( n9287 & n12042 ) ;
  assign n12590 = ( n3136 & n5187 ) | ( n3136 & n8580 ) | ( n5187 & n8580 ) ;
  assign n12585 = ( n4462 & ~n8007 ) | ( n4462 & n12193 ) | ( ~n8007 & n12193 ) ;
  assign n12586 = n6819 ^ n3879 ^ n1949 ;
  assign n12587 = ( ~n5864 & n12585 ) | ( ~n5864 & n12586 ) | ( n12585 & n12586 ) ;
  assign n12588 = ( ~n1719 & n10754 ) | ( ~n1719 & n12587 ) | ( n10754 & n12587 ) ;
  assign n12589 = n12588 ^ n10781 ^ n4789 ;
  assign n12592 = n12591 ^ n12590 ^ n12589 ;
  assign n12593 = ( n5117 & n9356 ) | ( n5117 & n11799 ) | ( n9356 & n11799 ) ;
  assign n12594 = n9630 ^ n5970 ^ n5538 ;
  assign n12595 = n4873 ^ n1103 ^ n574 ;
  assign n12596 = n12595 ^ n9173 ^ n3728 ;
  assign n12597 = n12596 ^ n7700 ^ n1265 ;
  assign n12598 = n12597 ^ n5281 ^ n237 ;
  assign n12599 = n7445 ^ n5934 ^ n2493 ;
  assign n12600 = ( n494 & n2487 ) | ( n494 & ~n4237 ) | ( n2487 & ~n4237 ) ;
  assign n12601 = ( n1107 & n4858 ) | ( n1107 & ~n12600 ) | ( n4858 & ~n12600 ) ;
  assign n12602 = ( n4468 & n7195 ) | ( n4468 & ~n12601 ) | ( n7195 & ~n12601 ) ;
  assign n12603 = ( ~n926 & n1995 ) | ( ~n926 & n2449 ) | ( n1995 & n2449 ) ;
  assign n12604 = n9711 ^ n6705 ^ n4630 ;
  assign n12605 = n12604 ^ n10291 ^ n6434 ;
  assign n12606 = ( n9213 & n12603 ) | ( n9213 & n12605 ) | ( n12603 & n12605 ) ;
  assign n12607 = ( n11931 & n12602 ) | ( n11931 & n12606 ) | ( n12602 & n12606 ) ;
  assign n12609 = ( ~n417 & n1670 ) | ( ~n417 & n3442 ) | ( n1670 & n3442 ) ;
  assign n12608 = n9777 ^ n7355 ^ n2850 ;
  assign n12610 = n12609 ^ n12608 ^ n9100 ;
  assign n12611 = n12610 ^ n7457 ^ n2439 ;
  assign n12613 = ( n1330 & ~n3904 ) | ( n1330 & n6425 ) | ( ~n3904 & n6425 ) ;
  assign n12612 = ( n5340 & n9218 ) | ( n5340 & ~n11288 ) | ( n9218 & ~n11288 ) ;
  assign n12614 = n12613 ^ n12612 ^ n1801 ;
  assign n12616 = n7673 ^ n5042 ^ n4388 ;
  assign n12615 = ( n3070 & n5439 ) | ( n3070 & n9496 ) | ( n5439 & n9496 ) ;
  assign n12617 = n12616 ^ n12615 ^ n1612 ;
  assign n12618 = ( n3653 & n6463 ) | ( n3653 & ~n12617 ) | ( n6463 & ~n12617 ) ;
  assign n12619 = ( n3939 & n7814 ) | ( n3939 & n8333 ) | ( n7814 & n8333 ) ;
  assign n12621 = n7457 ^ n5213 ^ n1268 ;
  assign n12620 = n12108 ^ n9498 ^ n5162 ;
  assign n12622 = n12621 ^ n12620 ^ n986 ;
  assign n12632 = n10607 ^ n6276 ^ n3663 ;
  assign n12631 = n4104 ^ n1987 ^ n1333 ;
  assign n12627 = ( ~n282 & n4467 ) | ( ~n282 & n11860 ) | ( n4467 & n11860 ) ;
  assign n12624 = n9081 ^ n8282 ^ n5909 ;
  assign n12623 = n9803 ^ n7240 ^ n5366 ;
  assign n12625 = n12624 ^ n12623 ^ n3125 ;
  assign n12626 = n12625 ^ n7370 ^ n2057 ;
  assign n12628 = n12627 ^ n12626 ^ n1355 ;
  assign n12629 = ( ~n4624 & n9425 ) | ( ~n4624 & n12628 ) | ( n9425 & n12628 ) ;
  assign n12630 = ( n3006 & n4432 ) | ( n3006 & ~n12629 ) | ( n4432 & ~n12629 ) ;
  assign n12633 = n12632 ^ n12631 ^ n12630 ;
  assign n12634 = n5971 ^ n4621 ^ n1135 ;
  assign n12635 = n9985 ^ n7036 ^ n2487 ;
  assign n12636 = ( n8419 & n8563 ) | ( n8419 & n12635 ) | ( n8563 & n12635 ) ;
  assign n12637 = n11156 ^ n5251 ^ n355 ;
  assign n12638 = ( n6705 & ~n8877 ) | ( n6705 & n12637 ) | ( ~n8877 & n12637 ) ;
  assign n12639 = ( n3627 & n12636 ) | ( n3627 & n12638 ) | ( n12636 & n12638 ) ;
  assign n12640 = ( ~n6816 & n10126 ) | ( ~n6816 & n12639 ) | ( n10126 & n12639 ) ;
  assign n12641 = ( ~n3353 & n12634 ) | ( ~n3353 & n12640 ) | ( n12634 & n12640 ) ;
  assign n12642 = ( ~n2663 & n2681 ) | ( ~n2663 & n8825 ) | ( n2681 & n8825 ) ;
  assign n12643 = n12642 ^ n5180 ^ n3062 ;
  assign n12644 = ( ~n968 & n1692 ) | ( ~n968 & n12643 ) | ( n1692 & n12643 ) ;
  assign n12645 = ( ~n2603 & n4325 ) | ( ~n2603 & n12644 ) | ( n4325 & n12644 ) ;
  assign n12646 = ( n8648 & n10036 ) | ( n8648 & n12645 ) | ( n10036 & n12645 ) ;
  assign n12647 = n8837 ^ n4822 ^ n2572 ;
  assign n12648 = n6633 ^ n4759 ^ n862 ;
  assign n12649 = ( n1934 & ~n6754 ) | ( n1934 & n12648 ) | ( ~n6754 & n12648 ) ;
  assign n12650 = ( n3234 & ~n12647 ) | ( n3234 & n12649 ) | ( ~n12647 & n12649 ) ;
  assign n12651 = ( n1900 & ~n2174 ) | ( n1900 & n6161 ) | ( ~n2174 & n6161 ) ;
  assign n12652 = n12651 ^ n12371 ^ n8750 ;
  assign n12653 = n12652 ^ n10083 ^ n2037 ;
  assign n12654 = ( n447 & ~n4205 ) | ( n447 & n4496 ) | ( ~n4205 & n4496 ) ;
  assign n12655 = ( n5921 & ~n9003 ) | ( n5921 & n12654 ) | ( ~n9003 & n12654 ) ;
  assign n12656 = ( n241 & n5975 ) | ( n241 & n8732 ) | ( n5975 & n8732 ) ;
  assign n12657 = ( n9527 & n10083 ) | ( n9527 & ~n12656 ) | ( n10083 & ~n12656 ) ;
  assign n12658 = ( n5237 & n8008 ) | ( n5237 & n12278 ) | ( n8008 & n12278 ) ;
  assign n12663 = ( n2009 & ~n2722 ) | ( n2009 & n5840 ) | ( ~n2722 & n5840 ) ;
  assign n12664 = ( n1142 & ~n2831 ) | ( n1142 & n3733 ) | ( ~n2831 & n3733 ) ;
  assign n12665 = n12664 ^ n6295 ^ n5317 ;
  assign n12666 = ( n3404 & n7424 ) | ( n3404 & ~n12665 ) | ( n7424 & ~n12665 ) ;
  assign n12667 = ( n10848 & n12663 ) | ( n10848 & ~n12666 ) | ( n12663 & ~n12666 ) ;
  assign n12661 = n7808 ^ n4093 ^ n1543 ;
  assign n12660 = n7928 ^ n4193 ^ n3351 ;
  assign n12659 = ( ~n645 & n3242 ) | ( ~n645 & n11811 ) | ( n3242 & n11811 ) ;
  assign n12662 = n12661 ^ n12660 ^ n12659 ;
  assign n12668 = n12667 ^ n12662 ^ n10151 ;
  assign n12669 = ( n12657 & ~n12658 ) | ( n12657 & n12668 ) | ( ~n12658 & n12668 ) ;
  assign n12670 = ( n2962 & n8660 ) | ( n2962 & ~n12052 ) | ( n8660 & ~n12052 ) ;
  assign n12671 = n12670 ^ n4122 ^ n1872 ;
  assign n12672 = ( ~n7102 & n7870 ) | ( ~n7102 & n12671 ) | ( n7870 & n12671 ) ;
  assign n12673 = ( ~n6403 & n11217 ) | ( ~n6403 & n12672 ) | ( n11217 & n12672 ) ;
  assign n12674 = ( n10484 & n10845 ) | ( n10484 & ~n11164 ) | ( n10845 & ~n11164 ) ;
  assign n12675 = ( n968 & ~n2904 ) | ( n968 & n7581 ) | ( ~n2904 & n7581 ) ;
  assign n12676 = ( n290 & n562 ) | ( n290 & n2628 ) | ( n562 & n2628 ) ;
  assign n12677 = n12676 ^ n9673 ^ n7576 ;
  assign n12678 = ( n10215 & n11346 ) | ( n10215 & ~n12677 ) | ( n11346 & ~n12677 ) ;
  assign n12679 = ( n12609 & n12675 ) | ( n12609 & n12678 ) | ( n12675 & n12678 ) ;
  assign n12680 = n11745 ^ n9520 ^ n518 ;
  assign n12681 = n12680 ^ n11441 ^ n5696 ;
  assign n12682 = ( n1285 & ~n2993 ) | ( n1285 & n3786 ) | ( ~n2993 & n3786 ) ;
  assign n12683 = ( n374 & n11575 ) | ( n374 & ~n12682 ) | ( n11575 & ~n12682 ) ;
  assign n12684 = n12683 ^ n4053 ^ n2694 ;
  assign n12685 = ( n7260 & n8393 ) | ( n7260 & n12684 ) | ( n8393 & n12684 ) ;
  assign n12686 = n7011 ^ n3652 ^ n1171 ;
  assign n12687 = ( n4637 & ~n8263 ) | ( n4637 & n12686 ) | ( ~n8263 & n12686 ) ;
  assign n12688 = ( n4722 & n4886 ) | ( n4722 & ~n5042 ) | ( n4886 & ~n5042 ) ;
  assign n12689 = ( n3755 & n6899 ) | ( n3755 & ~n12688 ) | ( n6899 & ~n12688 ) ;
  assign n12690 = ( n255 & n1543 ) | ( n255 & n4314 ) | ( n1543 & n4314 ) ;
  assign n12691 = n11001 ^ n2692 ^ n1639 ;
  assign n12692 = n10572 ^ n4093 ^ n3034 ;
  assign n12693 = n12692 ^ n10146 ^ n1455 ;
  assign n12694 = ( n3149 & n6014 ) | ( n3149 & n12693 ) | ( n6014 & n12693 ) ;
  assign n12695 = ( ~n12690 & n12691 ) | ( ~n12690 & n12694 ) | ( n12691 & n12694 ) ;
  assign n12696 = n6207 ^ n2347 ^ n637 ;
  assign n12697 = n12253 ^ n10090 ^ n3827 ;
  assign n12699 = n6234 ^ n5924 ^ n2384 ;
  assign n12698 = n7887 ^ n1488 ^ n1430 ;
  assign n12700 = n12699 ^ n12698 ^ n987 ;
  assign n12701 = ( n718 & n1295 ) | ( n718 & ~n1594 ) | ( n1295 & ~n1594 ) ;
  assign n12702 = ( n2571 & ~n9713 ) | ( n2571 & n12701 ) | ( ~n9713 & n12701 ) ;
  assign n12703 = n12601 ^ n8662 ^ n1001 ;
  assign n12705 = ( n1199 & n2394 ) | ( n1199 & ~n4561 ) | ( n2394 & ~n4561 ) ;
  assign n12704 = n6960 ^ n5027 ^ n1743 ;
  assign n12706 = n12705 ^ n12704 ^ n7260 ;
  assign n12707 = n10699 ^ n5853 ^ n1279 ;
  assign n12708 = ( n319 & ~n343 ) | ( n319 & n1101 ) | ( ~n343 & n1101 ) ;
  assign n12709 = ( n956 & n8922 ) | ( n956 & n12708 ) | ( n8922 & n12708 ) ;
  assign n12710 = n12709 ^ n12170 ^ n10106 ;
  assign n12711 = n12710 ^ n12125 ^ n9791 ;
  assign n12712 = n4627 ^ n3671 ^ n3334 ;
  assign n12713 = ( x102 & ~n2491 ) | ( x102 & n5326 ) | ( ~n2491 & n5326 ) ;
  assign n12714 = ( n2309 & n3699 ) | ( n2309 & ~n12713 ) | ( n3699 & ~n12713 ) ;
  assign n12715 = n12714 ^ n7180 ^ n2801 ;
  assign n12716 = ( n6453 & n10676 ) | ( n6453 & n12715 ) | ( n10676 & n12715 ) ;
  assign n12717 = n12716 ^ n5939 ^ n2111 ;
  assign n12718 = ( n5436 & ~n11638 ) | ( n5436 & n12717 ) | ( ~n11638 & n12717 ) ;
  assign n12719 = n4150 ^ n887 ^ n621 ;
  assign n12720 = n12719 ^ n5522 ^ n4047 ;
  assign n12721 = ( ~n9516 & n12718 ) | ( ~n9516 & n12720 ) | ( n12718 & n12720 ) ;
  assign n12722 = ( ~n917 & n12712 ) | ( ~n917 & n12721 ) | ( n12712 & n12721 ) ;
  assign n12723 = ( n938 & n5538 ) | ( n938 & n8260 ) | ( n5538 & n8260 ) ;
  assign n12724 = n12723 ^ n8740 ^ n513 ;
  assign n12725 = ( n3879 & ~n5712 ) | ( n3879 & n5759 ) | ( ~n5712 & n5759 ) ;
  assign n12726 = n12725 ^ n6516 ^ n2560 ;
  assign n12727 = n12726 ^ n5479 ^ n2507 ;
  assign n12728 = n9007 ^ n5709 ^ n3392 ;
  assign n12729 = n12728 ^ n10238 ^ n9068 ;
  assign n12730 = ( n2139 & n2824 ) | ( n2139 & ~n5580 ) | ( n2824 & ~n5580 ) ;
  assign n12731 = ( n1892 & ~n5095 ) | ( n1892 & n12730 ) | ( ~n5095 & n12730 ) ;
  assign n12732 = n10208 ^ n7908 ^ n1799 ;
  assign n12733 = ( n2020 & n3393 ) | ( n2020 & n7187 ) | ( n3393 & n7187 ) ;
  assign n12734 = ( ~n641 & n2275 ) | ( ~n641 & n12733 ) | ( n2275 & n12733 ) ;
  assign n12735 = ( ~n3475 & n12732 ) | ( ~n3475 & n12734 ) | ( n12732 & n12734 ) ;
  assign n12736 = ( n1478 & n2359 ) | ( n1478 & ~n5455 ) | ( n2359 & ~n5455 ) ;
  assign n12737 = n12736 ^ n10112 ^ n8055 ;
  assign n12738 = ( n3985 & n5409 ) | ( n3985 & n8769 ) | ( n5409 & n8769 ) ;
  assign n12739 = n12738 ^ n4659 ^ n2366 ;
  assign n12740 = n12739 ^ n8331 ^ n5173 ;
  assign n12741 = ( ~n2763 & n11536 ) | ( ~n2763 & n12740 ) | ( n11536 & n12740 ) ;
  assign n12744 = n7897 ^ n3210 ^ n532 ;
  assign n12745 = n12744 ^ n6068 ^ n1693 ;
  assign n12746 = ( n4871 & n8919 ) | ( n4871 & ~n12745 ) | ( n8919 & ~n12745 ) ;
  assign n12742 = ( n633 & ~n2319 ) | ( n633 & n6531 ) | ( ~n2319 & n6531 ) ;
  assign n12743 = n12742 ^ n11692 ^ n960 ;
  assign n12747 = n12746 ^ n12743 ^ n12158 ;
  assign n12752 = ( n4438 & ~n7300 ) | ( n4438 & n12394 ) | ( ~n7300 & n12394 ) ;
  assign n12748 = n12575 ^ n8072 ^ n793 ;
  assign n12749 = ( n1962 & n10172 ) | ( n1962 & n12748 ) | ( n10172 & n12748 ) ;
  assign n12750 = n10844 ^ n7015 ^ n2685 ;
  assign n12751 = ( n6893 & ~n12749 ) | ( n6893 & n12750 ) | ( ~n12749 & n12750 ) ;
  assign n12753 = n12752 ^ n12751 ^ n8427 ;
  assign n12755 = ( n2060 & n2513 ) | ( n2060 & ~n5219 ) | ( n2513 & ~n5219 ) ;
  assign n12756 = n12755 ^ n5266 ^ n2268 ;
  assign n12754 = n4444 ^ n2559 ^ n2377 ;
  assign n12757 = n12756 ^ n12754 ^ n3058 ;
  assign n12758 = n11503 ^ n8853 ^ n3552 ;
  assign n12759 = n10416 ^ n9525 ^ n3655 ;
  assign n12760 = ( n7760 & n10583 ) | ( n7760 & n12759 ) | ( n10583 & n12759 ) ;
  assign n12761 = n12760 ^ n11693 ^ n1929 ;
  assign n12762 = n9150 ^ n5102 ^ n1076 ;
  assign n12763 = ( n1196 & n1290 ) | ( n1196 & n3101 ) | ( n1290 & n3101 ) ;
  assign n12764 = n12763 ^ n3782 ^ n2883 ;
  assign n12765 = n9739 ^ n7163 ^ n3148 ;
  assign n12766 = ( n190 & n1004 ) | ( n190 & ~n1105 ) | ( n1004 & ~n1105 ) ;
  assign n12767 = ( ~n417 & n4422 ) | ( ~n417 & n7347 ) | ( n4422 & n7347 ) ;
  assign n12768 = n12767 ^ n7481 ^ n569 ;
  assign n12769 = ( n4419 & n12766 ) | ( n4419 & ~n12768 ) | ( n12766 & ~n12768 ) ;
  assign n12770 = ( n12764 & ~n12765 ) | ( n12764 & n12769 ) | ( ~n12765 & n12769 ) ;
  assign n12771 = ( n1460 & n2427 ) | ( n1460 & n4667 ) | ( n2427 & n4667 ) ;
  assign n12772 = ( n4265 & n9476 ) | ( n4265 & ~n12771 ) | ( n9476 & ~n12771 ) ;
  assign n12774 = n4892 ^ n2891 ^ n1798 ;
  assign n12773 = ( n1874 & n4549 ) | ( n1874 & ~n9882 ) | ( n4549 & ~n9882 ) ;
  assign n12775 = n12774 ^ n12773 ^ n10863 ;
  assign n12776 = ( n8994 & n10320 ) | ( n8994 & ~n10475 ) | ( n10320 & ~n10475 ) ;
  assign n12777 = n8475 ^ n3123 ^ n2689 ;
  assign n12778 = ( ~n5654 & n7476 ) | ( ~n5654 & n12777 ) | ( n7476 & n12777 ) ;
  assign n12780 = n3738 ^ n1946 ^ n1286 ;
  assign n12781 = n12780 ^ n4243 ^ n3496 ;
  assign n12779 = ( n2522 & n2529 ) | ( n2522 & n7092 ) | ( n2529 & n7092 ) ;
  assign n12782 = n12781 ^ n12779 ^ n7096 ;
  assign n12784 = n4353 ^ n1788 ^ n1000 ;
  assign n12785 = ( n593 & n1927 ) | ( n593 & n12784 ) | ( n1927 & n12784 ) ;
  assign n12783 = ( n1070 & ~n1611 ) | ( n1070 & n9967 ) | ( ~n1611 & n9967 ) ;
  assign n12786 = n12785 ^ n12783 ^ n2596 ;
  assign n12790 = n11240 ^ n6537 ^ n3400 ;
  assign n12788 = ( n5103 & ~n6134 ) | ( n5103 & n8347 ) | ( ~n6134 & n8347 ) ;
  assign n12787 = ( n9889 & ~n10274 ) | ( n9889 & n12055 ) | ( ~n10274 & n12055 ) ;
  assign n12789 = n12788 ^ n12787 ^ n6105 ;
  assign n12791 = n12790 ^ n12789 ^ n12710 ;
  assign n12792 = ( ~n1886 & n3443 ) | ( ~n1886 & n4805 ) | ( n3443 & n4805 ) ;
  assign n12793 = ( ~n708 & n12632 ) | ( ~n708 & n12792 ) | ( n12632 & n12792 ) ;
  assign n12794 = n11696 ^ n11082 ^ x59 ;
  assign n12795 = n3144 ^ n3043 ^ n146 ;
  assign n12796 = ( n5234 & n10255 ) | ( n5234 & ~n12795 ) | ( n10255 & ~n12795 ) ;
  assign n12800 = n2111 ^ n1851 ^ n1699 ;
  assign n12799 = ( n6741 & ~n8450 ) | ( n6741 & n12275 ) | ( ~n8450 & n12275 ) ;
  assign n12797 = ( n129 & n7251 ) | ( n129 & ~n10470 ) | ( n7251 & ~n10470 ) ;
  assign n12798 = n12797 ^ n7009 ^ n3626 ;
  assign n12801 = n12800 ^ n12799 ^ n12798 ;
  assign n12802 = ( n3855 & n12796 ) | ( n3855 & ~n12801 ) | ( n12796 & ~n12801 ) ;
  assign n12803 = ( n136 & n12794 ) | ( n136 & ~n12802 ) | ( n12794 & ~n12802 ) ;
  assign n12804 = n3715 ^ n1220 ^ n576 ;
  assign n12805 = ( n4020 & n6836 ) | ( n4020 & ~n12804 ) | ( n6836 & ~n12804 ) ;
  assign n12806 = n12805 ^ n4768 ^ n1244 ;
  assign n12807 = n12806 ^ n9092 ^ n4999 ;
  assign n12808 = n12807 ^ n11926 ^ n388 ;
  assign n12809 = ( n1199 & n4865 ) | ( n1199 & n12808 ) | ( n4865 & n12808 ) ;
  assign n12811 = ( n246 & ~n1686 ) | ( n246 & n8238 ) | ( ~n1686 & n8238 ) ;
  assign n12810 = n7230 ^ n5161 ^ n990 ;
  assign n12812 = n12811 ^ n12810 ^ n7618 ;
  assign n12819 = ( n647 & n3792 ) | ( n647 & ~n5229 ) | ( n3792 & ~n5229 ) ;
  assign n12820 = ( n2178 & ~n2445 ) | ( n2178 & n12819 ) | ( ~n2445 & n12819 ) ;
  assign n12821 = n12820 ^ n11382 ^ n5190 ;
  assign n12814 = n6134 ^ n3334 ^ n309 ;
  assign n12815 = ( n3846 & n3884 ) | ( n3846 & ~n5176 ) | ( n3884 & ~n5176 ) ;
  assign n12816 = n12815 ^ n12017 ^ n10555 ;
  assign n12817 = n12816 ^ n2080 ^ n532 ;
  assign n12818 = ( ~n10638 & n12814 ) | ( ~n10638 & n12817 ) | ( n12814 & n12817 ) ;
  assign n12813 = ( n5086 & n8950 ) | ( n5086 & n12544 ) | ( n8950 & n12544 ) ;
  assign n12822 = n12821 ^ n12818 ^ n12813 ;
  assign n12826 = n4973 ^ n4344 ^ n2190 ;
  assign n12823 = n5418 ^ n2781 ^ n300 ;
  assign n12824 = n12823 ^ n10387 ^ n9567 ;
  assign n12825 = ( n829 & n3657 ) | ( n829 & ~n12824 ) | ( n3657 & ~n12824 ) ;
  assign n12827 = n12826 ^ n12825 ^ n8906 ;
  assign n12828 = n5101 ^ n3995 ^ n1539 ;
  assign n12829 = ( n248 & n3636 ) | ( n248 & ~n12828 ) | ( n3636 & ~n12828 ) ;
  assign n12830 = ( n1039 & ~n2400 ) | ( n1039 & n5034 ) | ( ~n2400 & n5034 ) ;
  assign n12831 = ( n11941 & n12829 ) | ( n11941 & ~n12830 ) | ( n12829 & ~n12830 ) ;
  assign n12832 = n12831 ^ n12302 ^ n1969 ;
  assign n12833 = ( x35 & n905 ) | ( x35 & n6952 ) | ( n905 & n6952 ) ;
  assign n12838 = n11062 ^ n2185 ^ n1142 ;
  assign n12834 = ( ~n166 & n1606 ) | ( ~n166 & n12642 ) | ( n1606 & n12642 ) ;
  assign n12835 = ( n3223 & n3845 ) | ( n3223 & ~n6057 ) | ( n3845 & ~n6057 ) ;
  assign n12836 = n8109 ^ n1848 ^ n202 ;
  assign n12837 = ( n12834 & ~n12835 ) | ( n12834 & n12836 ) | ( ~n12835 & n12836 ) ;
  assign n12839 = n12838 ^ n12837 ^ n12777 ;
  assign n12840 = ( n7252 & n12456 ) | ( n7252 & n12839 ) | ( n12456 & n12839 ) ;
  assign n12841 = ( n9818 & ~n12833 ) | ( n9818 & n12840 ) | ( ~n12833 & n12840 ) ;
  assign n12842 = ( n3562 & n12832 ) | ( n3562 & ~n12841 ) | ( n12832 & ~n12841 ) ;
  assign n12843 = n6526 ^ n1573 ^ x62 ;
  assign n12844 = n12843 ^ n7154 ^ n3717 ;
  assign n12845 = n12844 ^ n1817 ^ n1018 ;
  assign n12846 = n5774 ^ n3634 ^ n2532 ;
  assign n12847 = ( n289 & n9407 ) | ( n289 & ~n10056 ) | ( n9407 & ~n10056 ) ;
  assign n12848 = ( n1240 & ~n12846 ) | ( n1240 & n12847 ) | ( ~n12846 & n12847 ) ;
  assign n12849 = n7839 ^ n6049 ^ n2804 ;
  assign n12850 = ( n12350 & n12848 ) | ( n12350 & n12849 ) | ( n12848 & n12849 ) ;
  assign n12851 = ( ~n11722 & n12845 ) | ( ~n11722 & n12850 ) | ( n12845 & n12850 ) ;
  assign n12852 = ( n223 & ~n531 ) | ( n223 & n10885 ) | ( ~n531 & n10885 ) ;
  assign n12853 = n12852 ^ n7292 ^ n1339 ;
  assign n12854 = ( n1218 & ~n12514 ) | ( n1218 & n12853 ) | ( ~n12514 & n12853 ) ;
  assign n12855 = ( n8125 & n8654 ) | ( n8125 & n12854 ) | ( n8654 & n12854 ) ;
  assign n12856 = n3714 ^ n1636 ^ n1395 ;
  assign n12857 = n12856 ^ n7303 ^ n4417 ;
  assign n12858 = ( ~n2620 & n3887 ) | ( ~n2620 & n7758 ) | ( n3887 & n7758 ) ;
  assign n12860 = ( n726 & n1590 ) | ( n726 & ~n9558 ) | ( n1590 & ~n9558 ) ;
  assign n12859 = n7933 ^ n3730 ^ n553 ;
  assign n12861 = n12860 ^ n12859 ^ n10525 ;
  assign n12864 = n5259 ^ n4863 ^ n1360 ;
  assign n12862 = ( n3650 & n9232 ) | ( n3650 & n12364 ) | ( n9232 & n12364 ) ;
  assign n12863 = ( n4044 & ~n11136 ) | ( n4044 & n12862 ) | ( ~n11136 & n12862 ) ;
  assign n12865 = n12864 ^ n12863 ^ n11594 ;
  assign n12866 = n5060 ^ n3768 ^ n1290 ;
  assign n12868 = n6487 ^ n3858 ^ n302 ;
  assign n12869 = ( n2437 & n11125 ) | ( n2437 & ~n12868 ) | ( n11125 & ~n12868 ) ;
  assign n12867 = n9238 ^ n5314 ^ n4658 ;
  assign n12870 = n12869 ^ n12867 ^ n5374 ;
  assign n12871 = ( n7816 & n12866 ) | ( n7816 & ~n12870 ) | ( n12866 & ~n12870 ) ;
  assign n12872 = n11571 ^ n9929 ^ x66 ;
  assign n12882 = ( n584 & n2733 ) | ( n584 & n4273 ) | ( n2733 & n4273 ) ;
  assign n12881 = ( n1227 & n2269 ) | ( n1227 & ~n9471 ) | ( n2269 & ~n9471 ) ;
  assign n12879 = ( ~n1639 & n4622 ) | ( ~n1639 & n9253 ) | ( n4622 & n9253 ) ;
  assign n12880 = ( ~n9329 & n10643 ) | ( ~n9329 & n12879 ) | ( n10643 & n12879 ) ;
  assign n12883 = n12882 ^ n12881 ^ n12880 ;
  assign n12876 = ( n581 & n924 ) | ( n581 & ~n3934 ) | ( n924 & ~n3934 ) ;
  assign n12875 = ( n2409 & n6422 ) | ( n2409 & n7143 ) | ( n6422 & n7143 ) ;
  assign n12877 = n12876 ^ n12875 ^ n1979 ;
  assign n12873 = n12569 ^ n6895 ^ n5736 ;
  assign n12874 = n12873 ^ n1573 ^ n1041 ;
  assign n12878 = n12877 ^ n12874 ^ n581 ;
  assign n12884 = n12883 ^ n12878 ^ n8645 ;
  assign n12885 = ( ~n2304 & n4514 ) | ( ~n2304 & n7246 ) | ( n4514 & n7246 ) ;
  assign n12886 = n12885 ^ n11567 ^ n2080 ;
  assign n12887 = ( n3058 & n4410 ) | ( n3058 & n6106 ) | ( n4410 & n6106 ) ;
  assign n12888 = n12887 ^ n5621 ^ n4245 ;
  assign n12889 = n4562 ^ n2943 ^ n2105 ;
  assign n12890 = ( n4459 & n7672 ) | ( n4459 & n12889 ) | ( n7672 & n12889 ) ;
  assign n12891 = ( n277 & n12888 ) | ( n277 & n12890 ) | ( n12888 & n12890 ) ;
  assign n12892 = n11797 ^ n9541 ^ n5728 ;
  assign n12893 = ( n1298 & n8904 ) | ( n1298 & ~n12892 ) | ( n8904 & ~n12892 ) ;
  assign n12895 = ( n2841 & n3870 ) | ( n2841 & ~n5385 ) | ( n3870 & ~n5385 ) ;
  assign n12894 = n11297 ^ n3937 ^ n2348 ;
  assign n12896 = n12895 ^ n12894 ^ n530 ;
  assign n12897 = ( n4515 & n10241 ) | ( n4515 & n11266 ) | ( n10241 & n11266 ) ;
  assign n12898 = ( n4635 & ~n12896 ) | ( n4635 & n12897 ) | ( ~n12896 & n12897 ) ;
  assign n12899 = ( n3350 & n3384 ) | ( n3350 & n7034 ) | ( n3384 & n7034 ) ;
  assign n12900 = n12899 ^ n3205 ^ n1394 ;
  assign n12906 = ( n3024 & ~n3239 ) | ( n3024 & n6218 ) | ( ~n3239 & n6218 ) ;
  assign n12904 = ( ~n1542 & n3560 ) | ( ~n1542 & n10211 ) | ( n3560 & n10211 ) ;
  assign n12905 = n12904 ^ n6595 ^ n3194 ;
  assign n12901 = n5913 ^ n3449 ^ n1438 ;
  assign n12902 = n12901 ^ n5650 ^ n2507 ;
  assign n12903 = n12902 ^ n6741 ^ n2113 ;
  assign n12907 = n12906 ^ n12905 ^ n12903 ;
  assign n12910 = n12214 ^ n11789 ^ n405 ;
  assign n12908 = ( n2485 & n3130 ) | ( n2485 & ~n6311 ) | ( n3130 & ~n6311 ) ;
  assign n12909 = n12908 ^ n5564 ^ n4782 ;
  assign n12911 = n12910 ^ n12909 ^ n8444 ;
  assign n12912 = ( ~n12900 & n12907 ) | ( ~n12900 & n12911 ) | ( n12907 & n12911 ) ;
  assign n12913 = ( n961 & n3185 ) | ( n961 & n5892 ) | ( n3185 & n5892 ) ;
  assign n12914 = ( n9524 & n10914 ) | ( n9524 & n12913 ) | ( n10914 & n12913 ) ;
  assign n12915 = n9678 ^ n2592 ^ n1050 ;
  assign n12916 = ( n1161 & n1733 ) | ( n1161 & ~n12915 ) | ( n1733 & ~n12915 ) ;
  assign n12917 = n12916 ^ n12483 ^ n11760 ;
  assign n12920 = n12856 ^ n2827 ^ n663 ;
  assign n12921 = n12920 ^ n12087 ^ n3788 ;
  assign n12918 = ( n638 & n1834 ) | ( n638 & n3855 ) | ( n1834 & n3855 ) ;
  assign n12919 = n12918 ^ n7172 ^ n4392 ;
  assign n12922 = n12921 ^ n12919 ^ n4284 ;
  assign n12923 = ( n260 & n5864 ) | ( n260 & ~n12922 ) | ( n5864 & ~n12922 ) ;
  assign n12924 = ( ~n2842 & n2889 ) | ( ~n2842 & n6958 ) | ( n2889 & n6958 ) ;
  assign n12925 = ( n5963 & n6500 ) | ( n5963 & n8299 ) | ( n6500 & n8299 ) ;
  assign n12926 = ( ~n1716 & n12924 ) | ( ~n1716 & n12925 ) | ( n12924 & n12925 ) ;
  assign n12927 = n12926 ^ n11470 ^ x77 ;
  assign n12928 = ( n4546 & ~n8293 ) | ( n4546 & n12927 ) | ( ~n8293 & n12927 ) ;
  assign n12929 = n3878 ^ n2759 ^ n1059 ;
  assign n12930 = ( n1563 & n8503 ) | ( n1563 & ~n12929 ) | ( n8503 & ~n12929 ) ;
  assign n12931 = ( ~n947 & n6325 ) | ( ~n947 & n12930 ) | ( n6325 & n12930 ) ;
  assign n12934 = ( n5802 & n6337 ) | ( n5802 & ~n9041 ) | ( n6337 & ~n9041 ) ;
  assign n12935 = n12934 ^ n12391 ^ n8524 ;
  assign n12936 = n8576 ^ n8564 ^ n298 ;
  assign n12937 = ( n4059 & n12935 ) | ( n4059 & ~n12936 ) | ( n12935 & ~n12936 ) ;
  assign n12932 = ( n1505 & n2477 ) | ( n1505 & ~n7142 ) | ( n2477 & ~n7142 ) ;
  assign n12933 = ( n5616 & n11634 ) | ( n5616 & n12932 ) | ( n11634 & n12932 ) ;
  assign n12938 = n12937 ^ n12933 ^ n7460 ;
  assign n12939 = ( x98 & n5418 ) | ( x98 & ~n10423 ) | ( n5418 & ~n10423 ) ;
  assign n12940 = ( n6119 & ~n12588 ) | ( n6119 & n12939 ) | ( ~n12588 & n12939 ) ;
  assign n12941 = n7558 ^ n2514 ^ n433 ;
  assign n12942 = n12941 ^ n5153 ^ n4971 ;
  assign n12943 = ( n252 & n7699 ) | ( n252 & ~n12942 ) | ( n7699 & ~n12942 ) ;
  assign n12944 = n12943 ^ n5647 ^ n3976 ;
  assign n12945 = n12944 ^ n4238 ^ n1708 ;
  assign n12946 = n12945 ^ n10291 ^ n1828 ;
  assign n12947 = ( x24 & n1033 ) | ( x24 & n12895 ) | ( n1033 & n12895 ) ;
  assign n12948 = n12947 ^ n7539 ^ n4429 ;
  assign n12949 = ( n1661 & n1767 ) | ( n1661 & n4738 ) | ( n1767 & n4738 ) ;
  assign n12950 = n4762 ^ n4517 ^ n1017 ;
  assign n12951 = ( n11538 & n12949 ) | ( n11538 & ~n12950 ) | ( n12949 & ~n12950 ) ;
  assign n12952 = ( n1562 & n7002 ) | ( n1562 & ~n12951 ) | ( n7002 & ~n12951 ) ;
  assign n12953 = ( n1606 & ~n3506 ) | ( n1606 & n4976 ) | ( ~n3506 & n4976 ) ;
  assign n12954 = n12953 ^ n1893 ^ n1852 ;
  assign n12955 = n11214 ^ n1133 ^ n998 ;
  assign n12956 = ( n7034 & ~n12954 ) | ( n7034 & n12955 ) | ( ~n12954 & n12955 ) ;
  assign n12957 = ( n1269 & n6081 ) | ( n1269 & n8217 ) | ( n6081 & n8217 ) ;
  assign n12958 = n1693 ^ n1375 ^ n822 ;
  assign n12959 = n12958 ^ n7459 ^ n3572 ;
  assign n12960 = n12959 ^ n4044 ^ n3324 ;
  assign n12961 = ( n5066 & ~n5926 ) | ( n5066 & n8100 ) | ( ~n5926 & n8100 ) ;
  assign n12965 = ( n2617 & n9099 ) | ( n2617 & ~n11068 ) | ( n9099 & ~n11068 ) ;
  assign n12962 = ( n675 & ~n2903 ) | ( n675 & n8963 ) | ( ~n2903 & n8963 ) ;
  assign n12963 = n12962 ^ n8480 ^ n1083 ;
  assign n12964 = ( ~n5415 & n8988 ) | ( ~n5415 & n12963 ) | ( n8988 & n12963 ) ;
  assign n12966 = n12965 ^ n12964 ^ n3156 ;
  assign n12967 = ( ~n1341 & n1863 ) | ( ~n1341 & n12966 ) | ( n1863 & n12966 ) ;
  assign n12968 = ( n680 & n12961 ) | ( n680 & n12967 ) | ( n12961 & n12967 ) ;
  assign n12969 = ( ~n1133 & n3975 ) | ( ~n1133 & n12968 ) | ( n3975 & n12968 ) ;
  assign n12979 = n6660 ^ n2170 ^ n593 ;
  assign n12974 = n4455 ^ n3552 ^ n2366 ;
  assign n12975 = n2602 ^ n1607 ^ n1299 ;
  assign n12976 = n12975 ^ n8107 ^ n4571 ;
  assign n12977 = ( n8717 & ~n12974 ) | ( n8717 & n12976 ) | ( ~n12974 & n12976 ) ;
  assign n12978 = n12977 ^ n6824 ^ n236 ;
  assign n12971 = n3451 ^ n3314 ^ n665 ;
  assign n12970 = n4339 ^ n3482 ^ n2407 ;
  assign n12972 = n12971 ^ n12970 ^ n3560 ;
  assign n12973 = n12972 ^ n9003 ^ n6838 ;
  assign n12980 = n12979 ^ n12978 ^ n12973 ;
  assign n12981 = ( n464 & n3064 ) | ( n464 & ~n10936 ) | ( n3064 & ~n10936 ) ;
  assign n12982 = n12981 ^ n8005 ^ n812 ;
  assign n12983 = n12982 ^ n11239 ^ n2812 ;
  assign n12984 = ( n1482 & n2210 ) | ( n1482 & ~n4398 ) | ( n2210 & ~n4398 ) ;
  assign n12985 = n12984 ^ n6966 ^ n6744 ;
  assign n12989 = ( n2178 & ~n4586 ) | ( n2178 & n7146 ) | ( ~n4586 & n7146 ) ;
  assign n12986 = ( n5333 & n7171 ) | ( n5333 & ~n7763 ) | ( n7171 & ~n7763 ) ;
  assign n12987 = ( n447 & n3670 ) | ( n447 & n7176 ) | ( n3670 & n7176 ) ;
  assign n12988 = ( n1141 & ~n12986 ) | ( n1141 & n12987 ) | ( ~n12986 & n12987 ) ;
  assign n12990 = n12989 ^ n12988 ^ n8020 ;
  assign n12991 = ( n336 & ~n5283 ) | ( n336 & n10365 ) | ( ~n5283 & n10365 ) ;
  assign n12992 = n7583 ^ n5213 ^ n2845 ;
  assign n12993 = ( ~n2283 & n7567 ) | ( ~n2283 & n12992 ) | ( n7567 & n12992 ) ;
  assign n12994 = n4936 ^ n3506 ^ n2376 ;
  assign n12995 = ( n2635 & ~n7895 ) | ( n2635 & n12994 ) | ( ~n7895 & n12994 ) ;
  assign n12996 = n12995 ^ n2068 ^ n596 ;
  assign n12997 = ( ~n808 & n7057 ) | ( ~n808 & n8771 ) | ( n7057 & n8771 ) ;
  assign n13000 = n5394 ^ n2337 ^ n1587 ;
  assign n13001 = n13000 ^ n7377 ^ n2595 ;
  assign n12998 = n9384 ^ n3788 ^ n2376 ;
  assign n12999 = ( n3781 & ~n4127 ) | ( n3781 & n12998 ) | ( ~n4127 & n12998 ) ;
  assign n13002 = n13001 ^ n12999 ^ n3384 ;
  assign n13003 = ( n5601 & n7311 ) | ( n5601 & n10743 ) | ( n7311 & n10743 ) ;
  assign n13006 = ( n4438 & ~n4935 ) | ( n4438 & n5177 ) | ( ~n4935 & n5177 ) ;
  assign n13007 = ( n2523 & n3216 ) | ( n2523 & ~n8520 ) | ( n3216 & ~n8520 ) ;
  assign n13008 = ( n3423 & n13006 ) | ( n3423 & n13007 ) | ( n13006 & n13007 ) ;
  assign n13005 = ( n365 & ~n9353 ) | ( n365 & n12553 ) | ( ~n9353 & n12553 ) ;
  assign n13009 = n13008 ^ n13005 ^ n9512 ;
  assign n13010 = n13009 ^ n7323 ^ n370 ;
  assign n13004 = ( n2276 & ~n11038 ) | ( n2276 & n12788 ) | ( ~n11038 & n12788 ) ;
  assign n13011 = n13010 ^ n13004 ^ n6369 ;
  assign n13012 = n11835 ^ n3561 ^ x4 ;
  assign n13013 = ( n1265 & ~n3668 ) | ( n1265 & n6142 ) | ( ~n3668 & n6142 ) ;
  assign n13014 = ( n7251 & n13012 ) | ( n7251 & ~n13013 ) | ( n13012 & ~n13013 ) ;
  assign n13027 = n10318 ^ n7557 ^ n1457 ;
  assign n13021 = n12663 ^ n4878 ^ n804 ;
  assign n13022 = n10096 ^ n3013 ^ n475 ;
  assign n13023 = n13022 ^ n6582 ^ n3489 ;
  assign n13024 = ( n5114 & ~n13021 ) | ( n5114 & n13023 ) | ( ~n13021 & n13023 ) ;
  assign n13025 = n13024 ^ n9959 ^ n9955 ;
  assign n13020 = ( n3444 & n6552 ) | ( n3444 & n6686 ) | ( n6552 & n6686 ) ;
  assign n13026 = n13025 ^ n13020 ^ n4843 ;
  assign n13015 = ( n777 & ~n3862 ) | ( n777 & n11292 ) | ( ~n3862 & n11292 ) ;
  assign n13016 = ( ~n2314 & n7495 ) | ( ~n2314 & n13015 ) | ( n7495 & n13015 ) ;
  assign n13017 = n8447 ^ n3141 ^ n1566 ;
  assign n13018 = ( ~n1334 & n6967 ) | ( ~n1334 & n13017 ) | ( n6967 & n13017 ) ;
  assign n13019 = ( n7386 & n13016 ) | ( n7386 & ~n13018 ) | ( n13016 & ~n13018 ) ;
  assign n13028 = n13027 ^ n13026 ^ n13019 ;
  assign n13032 = ( n4023 & n4567 ) | ( n4023 & n4805 ) | ( n4567 & n4805 ) ;
  assign n13033 = ( n10499 & ~n11662 ) | ( n10499 & n13032 ) | ( ~n11662 & n13032 ) ;
  assign n13029 = n9024 ^ n5274 ^ n3568 ;
  assign n13030 = n13029 ^ n9014 ^ n3120 ;
  assign n13031 = ( n1156 & n5041 ) | ( n1156 & n13030 ) | ( n5041 & n13030 ) ;
  assign n13034 = n13033 ^ n13031 ^ n11088 ;
  assign n13035 = ( ~n7263 & n9776 ) | ( ~n7263 & n12999 ) | ( n9776 & n12999 ) ;
  assign n13036 = n9201 ^ n7585 ^ n1923 ;
  assign n13037 = n13036 ^ n3098 ^ x35 ;
  assign n13038 = ( ~n12238 & n13035 ) | ( ~n12238 & n13037 ) | ( n13035 & n13037 ) ;
  assign n13039 = ( n771 & n2925 ) | ( n771 & ~n5064 ) | ( n2925 & ~n5064 ) ;
  assign n13040 = ( n1678 & n3530 ) | ( n1678 & n13039 ) | ( n3530 & n13039 ) ;
  assign n13045 = n2900 ^ n797 ^ n643 ;
  assign n13041 = ( n838 & ~n2263 ) | ( n838 & n3882 ) | ( ~n2263 & n3882 ) ;
  assign n13042 = n11449 ^ n4973 ^ n4228 ;
  assign n13043 = ( ~n6432 & n13041 ) | ( ~n6432 & n13042 ) | ( n13041 & n13042 ) ;
  assign n13044 = n13043 ^ n8064 ^ n2117 ;
  assign n13046 = n13045 ^ n13044 ^ n9776 ;
  assign n13047 = n13046 ^ n12347 ^ n4822 ;
  assign n13048 = ( ~n890 & n3314 ) | ( ~n890 & n9985 ) | ( n3314 & n9985 ) ;
  assign n13049 = ( ~n3642 & n3964 ) | ( ~n3642 & n13048 ) | ( n3964 & n13048 ) ;
  assign n13050 = ( n3271 & n5883 ) | ( n3271 & ~n13049 ) | ( n5883 & ~n13049 ) ;
  assign n13051 = ( n938 & ~n9119 ) | ( n938 & n9255 ) | ( ~n9119 & n9255 ) ;
  assign n13052 = n13051 ^ n2529 ^ n1783 ;
  assign n13053 = ( n1824 & ~n1932 ) | ( n1824 & n6825 ) | ( ~n1932 & n6825 ) ;
  assign n13054 = n13053 ^ n5295 ^ n2386 ;
  assign n13055 = ( n4573 & ~n6076 ) | ( n4573 & n7673 ) | ( ~n6076 & n7673 ) ;
  assign n13056 = ( n2959 & ~n13054 ) | ( n2959 & n13055 ) | ( ~n13054 & n13055 ) ;
  assign n13059 = n8340 ^ n6064 ^ n3235 ;
  assign n13057 = ( n11418 & n11515 ) | ( n11418 & n12190 ) | ( n11515 & n12190 ) ;
  assign n13058 = ( ~n3205 & n4160 ) | ( ~n3205 & n13057 ) | ( n4160 & n13057 ) ;
  assign n13060 = n13059 ^ n13058 ^ n2006 ;
  assign n13070 = ( ~n3699 & n8191 ) | ( ~n3699 & n12705 ) | ( n8191 & n12705 ) ;
  assign n13066 = n10365 ^ n1012 ^ n413 ;
  assign n13067 = n13066 ^ n10409 ^ n3728 ;
  assign n13068 = n13067 ^ n9032 ^ n4023 ;
  assign n13069 = ( n3329 & n8651 ) | ( n3329 & ~n13068 ) | ( n8651 & ~n13068 ) ;
  assign n13062 = ( n1299 & n2821 ) | ( n1299 & n5391 ) | ( n2821 & n5391 ) ;
  assign n13063 = n13062 ^ n11575 ^ n11562 ;
  assign n13061 = n11736 ^ n7695 ^ n4010 ;
  assign n13064 = n13063 ^ n13061 ^ n720 ;
  assign n13065 = ( n2694 & n10696 ) | ( n2694 & ~n13064 ) | ( n10696 & ~n13064 ) ;
  assign n13071 = n13070 ^ n13069 ^ n13065 ;
  assign n13072 = n3995 ^ n2207 ^ n812 ;
  assign n13073 = ( n899 & n2657 ) | ( n899 & n11475 ) | ( n2657 & n11475 ) ;
  assign n13074 = ( n147 & ~n13072 ) | ( n147 & n13073 ) | ( ~n13072 & n13073 ) ;
  assign n13075 = n13074 ^ n10011 ^ n5387 ;
  assign n13076 = ( n9128 & n12847 ) | ( n9128 & n13075 ) | ( n12847 & n13075 ) ;
  assign n13077 = ( n2502 & n7436 ) | ( n2502 & ~n10444 ) | ( n7436 & ~n10444 ) ;
  assign n13078 = n13077 ^ n8876 ^ n4122 ;
  assign n13079 = ( ~n1899 & n7149 ) | ( ~n1899 & n13078 ) | ( n7149 & n13078 ) ;
  assign n13082 = n8694 ^ n7667 ^ n5287 ;
  assign n13080 = ( n4352 & n4720 ) | ( n4352 & ~n5155 ) | ( n4720 & ~n5155 ) ;
  assign n13081 = ( ~n2007 & n6572 ) | ( ~n2007 & n13080 ) | ( n6572 & n13080 ) ;
  assign n13083 = n13082 ^ n13081 ^ n12773 ;
  assign n13084 = ( ~n2149 & n8967 ) | ( ~n2149 & n13083 ) | ( n8967 & n13083 ) ;
  assign n13085 = n10683 ^ n8880 ^ n7779 ;
  assign n13086 = ( n9782 & n12849 ) | ( n9782 & ~n13085 ) | ( n12849 & ~n13085 ) ;
  assign n13089 = ( x96 & ~n3852 ) | ( x96 & n6163 ) | ( ~n3852 & n6163 ) ;
  assign n13087 = n10739 ^ n7251 ^ n209 ;
  assign n13088 = ( n6014 & ~n10111 ) | ( n6014 & n13087 ) | ( ~n10111 & n13087 ) ;
  assign n13090 = n13089 ^ n13088 ^ n5612 ;
  assign n13093 = n12586 ^ n10243 ^ n6451 ;
  assign n13094 = n13093 ^ n4052 ^ n1534 ;
  assign n13091 = n3597 ^ n2425 ^ n2231 ;
  assign n13092 = n13091 ^ n12182 ^ n1034 ;
  assign n13095 = n13094 ^ n13092 ^ n1054 ;
  assign n13096 = n13095 ^ n5671 ^ n5135 ;
  assign n13097 = n13096 ^ n11952 ^ n11228 ;
  assign n13107 = ( n302 & ~n4821 ) | ( n302 & n12342 ) | ( ~n4821 & n12342 ) ;
  assign n13098 = ( n4134 & ~n8412 ) | ( n4134 & n11967 ) | ( ~n8412 & n11967 ) ;
  assign n13099 = n13098 ^ n8668 ^ n1932 ;
  assign n13100 = n13099 ^ n11362 ^ n11067 ;
  assign n13101 = n5948 ^ n5123 ^ n3767 ;
  assign n13102 = n13101 ^ n8569 ^ n4714 ;
  assign n13103 = n13102 ^ n5586 ^ n4510 ;
  assign n13104 = ( ~n9727 & n11947 ) | ( ~n9727 & n13103 ) | ( n11947 & n13103 ) ;
  assign n13105 = ( n3291 & n13100 ) | ( n3291 & ~n13104 ) | ( n13100 & ~n13104 ) ;
  assign n13106 = ( n5831 & n13006 ) | ( n5831 & ~n13105 ) | ( n13006 & ~n13105 ) ;
  assign n13108 = n13107 ^ n13106 ^ n10137 ;
  assign n13109 = n6282 ^ n5393 ^ n2349 ;
  assign n13110 = n13109 ^ n7418 ^ n5838 ;
  assign n13111 = n12155 ^ n11503 ^ n6344 ;
  assign n13112 = ( n1885 & n7026 ) | ( n1885 & ~n13111 ) | ( n7026 & ~n13111 ) ;
  assign n13114 = ( ~n997 & n1066 ) | ( ~n997 & n2097 ) | ( n1066 & n2097 ) ;
  assign n13115 = ( n3169 & n5051 ) | ( n3169 & ~n13114 ) | ( n5051 & ~n13114 ) ;
  assign n13113 = n12755 ^ n6571 ^ x1 ;
  assign n13116 = n13115 ^ n13113 ^ n11308 ;
  assign n13117 = ( n3295 & n9963 ) | ( n3295 & n13116 ) | ( n9963 & n13116 ) ;
  assign n13120 = ( n7112 & n8349 ) | ( n7112 & n8807 ) | ( n8349 & n8807 ) ;
  assign n13118 = n5900 ^ n5393 ^ n2817 ;
  assign n13119 = n13118 ^ n3219 ^ n946 ;
  assign n13121 = n13120 ^ n13119 ^ n8244 ;
  assign n13122 = n11037 ^ n4849 ^ n4040 ;
  assign n13123 = ( n5372 & n7493 ) | ( n5372 & n9816 ) | ( n7493 & n9816 ) ;
  assign n13124 = n13123 ^ n8763 ^ n7592 ;
  assign n13125 = ( n1604 & n6341 ) | ( n1604 & n13124 ) | ( n6341 & n13124 ) ;
  assign n13126 = ( ~n1666 & n5479 ) | ( ~n1666 & n13125 ) | ( n5479 & n13125 ) ;
  assign n13127 = ( n3304 & ~n8810 ) | ( n3304 & n12823 ) | ( ~n8810 & n12823 ) ;
  assign n13128 = n13127 ^ n9634 ^ n3464 ;
  assign n13130 = ( ~n775 & n4209 ) | ( ~n775 & n5549 ) | ( n4209 & n5549 ) ;
  assign n13129 = ( n1560 & n5879 ) | ( n1560 & ~n6288 ) | ( n5879 & ~n6288 ) ;
  assign n13131 = n13130 ^ n13129 ^ n11602 ;
  assign n13141 = ( ~n2467 & n5067 ) | ( ~n2467 & n8729 ) | ( n5067 & n8729 ) ;
  assign n13142 = ( n4715 & n4757 ) | ( n4715 & n13141 ) | ( n4757 & n13141 ) ;
  assign n13138 = n6838 ^ n4812 ^ n2712 ;
  assign n13139 = ( n6896 & n8393 ) | ( n6896 & n10965 ) | ( n8393 & n10965 ) ;
  assign n13140 = ( n1906 & ~n13138 ) | ( n1906 & n13139 ) | ( ~n13138 & n13139 ) ;
  assign n13143 = n13142 ^ n13140 ^ x47 ;
  assign n13137 = n12335 ^ n9959 ^ n2353 ;
  assign n13132 = ( n3965 & n7489 ) | ( n3965 & n10152 ) | ( n7489 & n10152 ) ;
  assign n13133 = n13132 ^ n11477 ^ n2279 ;
  assign n13134 = n13133 ^ n3582 ^ n3338 ;
  assign n13135 = n13134 ^ n6341 ^ n1274 ;
  assign n13136 = ( ~n4536 & n9656 ) | ( ~n4536 & n13135 ) | ( n9656 & n13135 ) ;
  assign n13144 = n13143 ^ n13137 ^ n13136 ;
  assign n13145 = ( n947 & n6917 ) | ( n947 & ~n9678 ) | ( n6917 & ~n9678 ) ;
  assign n13146 = ( n1406 & ~n7109 ) | ( n1406 & n13145 ) | ( ~n7109 & n13145 ) ;
  assign n13147 = ( n4734 & ~n7070 ) | ( n4734 & n13146 ) | ( ~n7070 & n13146 ) ;
  assign n13148 = n9589 ^ n3134 ^ n1517 ;
  assign n13155 = ( ~n882 & n10707 ) | ( ~n882 & n11903 ) | ( n10707 & n11903 ) ;
  assign n13151 = n2133 ^ n1421 ^ n993 ;
  assign n13152 = ( n4411 & n8449 ) | ( n4411 & ~n13151 ) | ( n8449 & ~n13151 ) ;
  assign n13153 = n13152 ^ n5726 ^ n3444 ;
  assign n13150 = n8136 ^ n5822 ^ n4093 ;
  assign n13154 = n13153 ^ n13150 ^ n6293 ;
  assign n13156 = n13155 ^ n13154 ^ n586 ;
  assign n13149 = ( n6360 & n6595 ) | ( n6360 & n7823 ) | ( n6595 & n7823 ) ;
  assign n13157 = n13156 ^ n13149 ^ n3270 ;
  assign n13158 = n6359 ^ n5265 ^ n1198 ;
  assign n13160 = n10588 ^ n3976 ^ n1081 ;
  assign n13161 = ( n1588 & n6500 ) | ( n1588 & ~n13160 ) | ( n6500 & ~n13160 ) ;
  assign n13159 = ( n3456 & ~n4736 ) | ( n3456 & n5958 ) | ( ~n4736 & n5958 ) ;
  assign n13162 = n13161 ^ n13159 ^ n6276 ;
  assign n13163 = ( n3508 & n4516 ) | ( n3508 & n10710 ) | ( n4516 & n10710 ) ;
  assign n13164 = n13163 ^ n11313 ^ n6050 ;
  assign n13165 = ( x11 & n1739 ) | ( x11 & n2469 ) | ( n1739 & n2469 ) ;
  assign n13166 = ( n679 & n2523 ) | ( n679 & n13165 ) | ( n2523 & n13165 ) ;
  assign n13167 = ( ~n2712 & n4651 ) | ( ~n2712 & n12719 ) | ( n4651 & n12719 ) ;
  assign n13175 = n9530 ^ n3433 ^ n2632 ;
  assign n13168 = ( ~n3773 & n8778 ) | ( ~n3773 & n9741 ) | ( n8778 & n9741 ) ;
  assign n13169 = n13168 ^ n2097 ^ n1017 ;
  assign n13170 = n10756 ^ n6429 ^ n3084 ;
  assign n13171 = ( ~n309 & n462 ) | ( ~n309 & n12962 ) | ( n462 & n12962 ) ;
  assign n13172 = ( n1855 & n3060 ) | ( n1855 & n13171 ) | ( n3060 & n13171 ) ;
  assign n13173 = ( n13169 & n13170 ) | ( n13169 & n13172 ) | ( n13170 & n13172 ) ;
  assign n13174 = ( ~n2203 & n7795 ) | ( ~n2203 & n13173 ) | ( n7795 & n13173 ) ;
  assign n13176 = n13175 ^ n13174 ^ n1700 ;
  assign n13177 = ( n3229 & n5191 ) | ( n3229 & ~n7688 ) | ( n5191 & ~n7688 ) ;
  assign n13178 = n13177 ^ n11854 ^ n247 ;
  assign n13179 = n13178 ^ n10501 ^ n1690 ;
  assign n13180 = ( n4742 & ~n8031 ) | ( n4742 & n12671 ) | ( ~n8031 & n12671 ) ;
  assign n13181 = n13180 ^ n10843 ^ n6717 ;
  assign n13182 = ( ~n2348 & n2843 ) | ( ~n2348 & n7375 ) | ( n2843 & n7375 ) ;
  assign n13183 = ( n1015 & ~n2971 ) | ( n1015 & n3546 ) | ( ~n2971 & n3546 ) ;
  assign n13184 = n13183 ^ n6652 ^ n820 ;
  assign n13185 = ( n1755 & ~n5567 ) | ( n1755 & n9239 ) | ( ~n5567 & n9239 ) ;
  assign n13186 = ( ~n5884 & n13184 ) | ( ~n5884 & n13185 ) | ( n13184 & n13185 ) ;
  assign n13187 = n2971 ^ n2406 ^ n1007 ;
  assign n13190 = n3860 ^ n2794 ^ n2429 ;
  assign n13189 = n6574 ^ n5885 ^ n4482 ;
  assign n13188 = n4310 ^ n3206 ^ n615 ;
  assign n13191 = n13190 ^ n13189 ^ n13188 ;
  assign n13192 = ( n4712 & n13187 ) | ( n4712 & ~n13191 ) | ( n13187 & ~n13191 ) ;
  assign n13193 = ( n1710 & n5617 ) | ( n1710 & n11380 ) | ( n5617 & n11380 ) ;
  assign n13194 = ( n262 & ~n328 ) | ( n262 & n1864 ) | ( ~n328 & n1864 ) ;
  assign n13195 = ( ~n5229 & n8004 ) | ( ~n5229 & n9828 ) | ( n8004 & n9828 ) ;
  assign n13196 = ( n9011 & n13194 ) | ( n9011 & ~n13195 ) | ( n13194 & ~n13195 ) ;
  assign n13197 = n10716 ^ n10324 ^ n1887 ;
  assign n13198 = n13197 ^ n3329 ^ n2635 ;
  assign n13199 = ( ~n334 & n5746 ) | ( ~n334 & n13198 ) | ( n5746 & n13198 ) ;
  assign n13200 = n12927 ^ n7041 ^ n5664 ;
  assign n13201 = ( n260 & n3347 ) | ( n260 & n10107 ) | ( n3347 & n10107 ) ;
  assign n13202 = n13201 ^ n9545 ^ n3022 ;
  assign n13204 = ( n236 & ~n3276 ) | ( n236 & n9238 ) | ( ~n3276 & n9238 ) ;
  assign n13203 = n5842 ^ n5123 ^ n2711 ;
  assign n13205 = n13204 ^ n13203 ^ x4 ;
  assign n13206 = n5776 ^ n5109 ^ n3404 ;
  assign n13207 = ( n7983 & n13000 ) | ( n7983 & n13206 ) | ( n13000 & n13206 ) ;
  assign n13208 = ( n3085 & n13205 ) | ( n3085 & ~n13207 ) | ( n13205 & ~n13207 ) ;
  assign n13209 = ( n1624 & n12414 ) | ( n1624 & ~n12935 ) | ( n12414 & ~n12935 ) ;
  assign n13210 = ( n6017 & n13208 ) | ( n6017 & ~n13209 ) | ( n13208 & ~n13209 ) ;
  assign n13211 = n8487 ^ n3975 ^ n790 ;
  assign n13212 = ( n256 & n8294 ) | ( n256 & ~n13211 ) | ( n8294 & ~n13211 ) ;
  assign n13213 = ( ~n2764 & n10964 ) | ( ~n2764 & n13212 ) | ( n10964 & n13212 ) ;
  assign n13214 = ( n681 & n1709 ) | ( n681 & n5560 ) | ( n1709 & n5560 ) ;
  assign n13215 = ( n1820 & n5203 ) | ( n1820 & ~n13214 ) | ( n5203 & ~n13214 ) ;
  assign n13216 = n13215 ^ n4623 ^ n1163 ;
  assign n13217 = n13216 ^ n11669 ^ n2542 ;
  assign n13220 = n8295 ^ n6062 ^ n5400 ;
  assign n13218 = ( n454 & ~n5572 ) | ( n454 & n8088 ) | ( ~n5572 & n8088 ) ;
  assign n13219 = n13218 ^ n10429 ^ n827 ;
  assign n13221 = n13220 ^ n13219 ^ n12435 ;
  assign n13222 = n13221 ^ n3148 ^ n1930 ;
  assign n13229 = n6892 ^ n1639 ^ n547 ;
  assign n13227 = n6246 ^ n3703 ^ n3172 ;
  assign n13228 = n13227 ^ n7120 ^ n1117 ;
  assign n13223 = n8782 ^ n7902 ^ n5657 ;
  assign n13224 = n13223 ^ n7541 ^ n959 ;
  assign n13225 = n13224 ^ n8899 ^ n4292 ;
  assign n13226 = ( n1346 & ~n2025 ) | ( n1346 & n13225 ) | ( ~n2025 & n13225 ) ;
  assign n13230 = n13229 ^ n13228 ^ n13226 ;
  assign n13231 = n9345 ^ n6664 ^ n3930 ;
  assign n13232 = n8396 ^ n4177 ^ n426 ;
  assign n13233 = n7529 ^ n7230 ^ n6334 ;
  assign n13234 = ( n1402 & n13232 ) | ( n1402 & n13233 ) | ( n13232 & n13233 ) ;
  assign n13235 = n13234 ^ n6927 ^ n5341 ;
  assign n13237 = ( n1056 & n5715 ) | ( n1056 & n9143 ) | ( n5715 & n9143 ) ;
  assign n13236 = n10516 ^ n8501 ^ n6105 ;
  assign n13238 = n13237 ^ n13236 ^ n2011 ;
  assign n13239 = ( n5809 & n12206 ) | ( n5809 & n13238 ) | ( n12206 & n13238 ) ;
  assign n13240 = ( n6868 & n10466 ) | ( n6868 & n13239 ) | ( n10466 & n13239 ) ;
  assign n13241 = ( n994 & n5173 ) | ( n994 & ~n7261 ) | ( n5173 & ~n7261 ) ;
  assign n13242 = ( n2557 & n3774 ) | ( n2557 & ~n13241 ) | ( n3774 & ~n13241 ) ;
  assign n13243 = ( n2055 & n2432 ) | ( n2055 & n7829 ) | ( n2432 & n7829 ) ;
  assign n13244 = n13243 ^ n12763 ^ n8753 ;
  assign n13245 = ( n3435 & ~n6116 ) | ( n3435 & n11350 ) | ( ~n6116 & n11350 ) ;
  assign n13246 = ( ~n10882 & n13244 ) | ( ~n10882 & n13245 ) | ( n13244 & n13245 ) ;
  assign n13247 = ( n7485 & n11866 ) | ( n7485 & ~n13246 ) | ( n11866 & ~n13246 ) ;
  assign n13248 = n9205 ^ n8356 ^ n6395 ;
  assign n13251 = ( n2314 & n3697 ) | ( n2314 & n5301 ) | ( n3697 & n5301 ) ;
  assign n13249 = ( n1534 & ~n3190 ) | ( n1534 & n7670 ) | ( ~n3190 & n7670 ) ;
  assign n13250 = ( n8838 & ~n10226 ) | ( n8838 & n13249 ) | ( ~n10226 & n13249 ) ;
  assign n13252 = n13251 ^ n13250 ^ n1707 ;
  assign n13253 = n4249 ^ n791 ^ x105 ;
  assign n13254 = n13253 ^ n10256 ^ n2121 ;
  assign n13255 = n10418 ^ n6326 ^ n5556 ;
  assign n13256 = n13255 ^ n9579 ^ n6648 ;
  assign n13257 = n13256 ^ n11882 ^ n5074 ;
  assign n13258 = ( n319 & n1950 ) | ( n319 & ~n2856 ) | ( n1950 & ~n2856 ) ;
  assign n13259 = n13258 ^ n4740 ^ n4073 ;
  assign n13260 = ( n2028 & n3698 ) | ( n2028 & ~n13259 ) | ( n3698 & ~n13259 ) ;
  assign n13261 = ( n825 & n4478 ) | ( n825 & n5631 ) | ( n4478 & n5631 ) ;
  assign n13262 = ( n10937 & ~n11786 ) | ( n10937 & n13261 ) | ( ~n11786 & n13261 ) ;
  assign n13263 = ( n4979 & ~n5970 ) | ( n4979 & n13262 ) | ( ~n5970 & n13262 ) ;
  assign n13264 = ( n4659 & n6496 ) | ( n4659 & ~n12487 ) | ( n6496 & ~n12487 ) ;
  assign n13265 = ( n1563 & n1596 ) | ( n1563 & n9924 ) | ( n1596 & n9924 ) ;
  assign n13266 = ( n7017 & ~n13264 ) | ( n7017 & n13265 ) | ( ~n13264 & n13265 ) ;
  assign n13267 = n11344 ^ n4607 ^ n1488 ;
  assign n13273 = ( n1570 & n5592 ) | ( n1570 & ~n9738 ) | ( n5592 & ~n9738 ) ;
  assign n13271 = n2641 ^ n2564 ^ n1966 ;
  assign n13272 = n13271 ^ n7642 ^ n6936 ;
  assign n13274 = n13273 ^ n13272 ^ n4678 ;
  assign n13269 = n12340 ^ n10321 ^ n8242 ;
  assign n13270 = ( n7479 & n13138 ) | ( n7479 & ~n13269 ) | ( n13138 & ~n13269 ) ;
  assign n13268 = ( n2565 & n2882 ) | ( n2565 & n9168 ) | ( n2882 & n9168 ) ;
  assign n13275 = n13274 ^ n13270 ^ n13268 ;
  assign n13277 = n7270 ^ n6469 ^ n665 ;
  assign n13276 = n9256 ^ n4163 ^ n3275 ;
  assign n13278 = n13277 ^ n13276 ^ n4770 ;
  assign n13279 = ( n3941 & ~n5059 ) | ( n3941 & n6175 ) | ( ~n5059 & n6175 ) ;
  assign n13280 = n13279 ^ n2557 ^ n890 ;
  assign n13281 = n13280 ^ n3502 ^ n3189 ;
  assign n13282 = ( n813 & ~n8013 ) | ( n813 & n9243 ) | ( ~n8013 & n9243 ) ;
  assign n13287 = n4030 ^ n1773 ^ n796 ;
  assign n13283 = n7150 ^ n4878 ^ n2531 ;
  assign n13284 = ( n2449 & n5510 ) | ( n2449 & n13283 ) | ( n5510 & n13283 ) ;
  assign n13285 = ( x25 & n8866 ) | ( x25 & n13284 ) | ( n8866 & n13284 ) ;
  assign n13286 = n13285 ^ n8647 ^ n7539 ;
  assign n13288 = n13287 ^ n13286 ^ n5990 ;
  assign n13289 = ( n10161 & n13282 ) | ( n10161 & ~n13288 ) | ( n13282 & ~n13288 ) ;
  assign n13290 = n13289 ^ n8601 ^ n3748 ;
  assign n13291 = n7322 ^ n2941 ^ n2694 ;
  assign n13292 = n11660 ^ n6075 ^ n4470 ;
  assign n13293 = ( n545 & n1444 ) | ( n545 & ~n13292 ) | ( n1444 & ~n13292 ) ;
  assign n13294 = ( n3856 & n13291 ) | ( n3856 & ~n13293 ) | ( n13291 & ~n13293 ) ;
  assign n13295 = n9660 ^ n7570 ^ n7229 ;
  assign n13296 = n3454 ^ n970 ^ n837 ;
  assign n13297 = n13296 ^ n8851 ^ n1973 ;
  assign n13298 = n9151 ^ n8502 ^ n6120 ;
  assign n13299 = ( n2918 & n5860 ) | ( n2918 & n13298 ) | ( n5860 & n13298 ) ;
  assign n13300 = n9139 ^ n7891 ^ n6325 ;
  assign n13301 = ( n2113 & n5028 ) | ( n2113 & ~n7306 ) | ( n5028 & ~n7306 ) ;
  assign n13302 = ( n3729 & ~n4313 ) | ( n3729 & n9138 ) | ( ~n4313 & n9138 ) ;
  assign n13303 = ( n8250 & n13301 ) | ( n8250 & ~n13302 ) | ( n13301 & ~n13302 ) ;
  assign n13306 = ( n2399 & n2812 ) | ( n2399 & ~n6271 ) | ( n2812 & ~n6271 ) ;
  assign n13307 = n13306 ^ n5814 ^ n5773 ;
  assign n13305 = ( ~n2695 & n2961 ) | ( ~n2695 & n12137 ) | ( n2961 & n12137 ) ;
  assign n13304 = ( n5352 & n7299 ) | ( n5352 & ~n11778 ) | ( n7299 & ~n11778 ) ;
  assign n13308 = n13307 ^ n13305 ^ n13304 ;
  assign n13309 = ( n1215 & n5775 ) | ( n1215 & ~n12159 ) | ( n5775 & ~n12159 ) ;
  assign n13311 = ( n6253 & ~n8324 ) | ( n6253 & n8854 ) | ( ~n8324 & n8854 ) ;
  assign n13310 = n5450 ^ n1818 ^ n545 ;
  assign n13312 = n13311 ^ n13310 ^ n2994 ;
  assign n13313 = n13312 ^ n8063 ^ n1076 ;
  assign n13316 = n3506 ^ n3204 ^ n2315 ;
  assign n13314 = n11597 ^ n1037 ^ n507 ;
  assign n13315 = n13314 ^ n5509 ^ n4967 ;
  assign n13317 = n13316 ^ n13315 ^ n2633 ;
  assign n13318 = ( n1408 & n2489 ) | ( n1408 & ~n3253 ) | ( n2489 & ~n3253 ) ;
  assign n13319 = n13318 ^ n6885 ^ n6092 ;
  assign n13320 = ( n3282 & n3502 ) | ( n3282 & ~n9062 ) | ( n3502 & ~n9062 ) ;
  assign n13321 = n12805 ^ n7579 ^ n4856 ;
  assign n13323 = n9182 ^ n2341 ^ n1721 ;
  assign n13322 = ( n950 & n2758 ) | ( n950 & n4444 ) | ( n2758 & n4444 ) ;
  assign n13324 = n13323 ^ n13322 ^ n2316 ;
  assign n13325 = ( n1840 & n7172 ) | ( n1840 & ~n13324 ) | ( n7172 & ~n13324 ) ;
  assign n13326 = ( n799 & ~n4515 ) | ( n799 & n13325 ) | ( ~n4515 & n13325 ) ;
  assign n13329 = ( n3761 & n6676 ) | ( n3761 & ~n9665 ) | ( n6676 & ~n9665 ) ;
  assign n13327 = n3747 ^ n649 ^ x119 ;
  assign n13328 = ( ~n243 & n7503 ) | ( ~n243 & n13327 ) | ( n7503 & n13327 ) ;
  assign n13330 = n13329 ^ n13328 ^ n11852 ;
  assign n13331 = n13330 ^ n10502 ^ n4077 ;
  assign n13334 = n3982 ^ n2599 ^ n1551 ;
  assign n13332 = ( n1632 & n2215 ) | ( n1632 & n4180 ) | ( n2215 & n4180 ) ;
  assign n13333 = ( n1547 & n6313 ) | ( n1547 & n13332 ) | ( n6313 & n13332 ) ;
  assign n13335 = n13334 ^ n13333 ^ n5620 ;
  assign n13336 = n10569 ^ n7032 ^ n6792 ;
  assign n13337 = n13336 ^ n7990 ^ n2897 ;
  assign n13338 = n10786 ^ n2456 ^ n992 ;
  assign n13339 = n13338 ^ n12661 ^ n9735 ;
  assign n13340 = ( n2087 & n6632 ) | ( n2087 & n11698 ) | ( n6632 & n11698 ) ;
  assign n13341 = ( n8805 & n12773 ) | ( n8805 & ~n13340 ) | ( n12773 & ~n13340 ) ;
  assign n13342 = ( n4818 & n13339 ) | ( n4818 & n13341 ) | ( n13339 & n13341 ) ;
  assign n13343 = ( n6759 & n9193 ) | ( n6759 & ~n10615 ) | ( n9193 & ~n10615 ) ;
  assign n13344 = ( n1883 & n7024 ) | ( n1883 & n11313 ) | ( n7024 & n11313 ) ;
  assign n13345 = n13344 ^ n11664 ^ n2906 ;
  assign n13346 = n10759 ^ n4803 ^ n1162 ;
  assign n13347 = ( n2647 & ~n10492 ) | ( n2647 & n11820 ) | ( ~n10492 & n11820 ) ;
  assign n13348 = ( n3816 & ~n9494 ) | ( n3816 & n13347 ) | ( ~n9494 & n13347 ) ;
  assign n13349 = ( ~n4352 & n13346 ) | ( ~n4352 & n13348 ) | ( n13346 & n13348 ) ;
  assign n13350 = n13091 ^ n7832 ^ n1299 ;
  assign n13351 = ( n609 & n12190 ) | ( n609 & ~n13350 ) | ( n12190 & ~n13350 ) ;
  assign n13352 = n9516 ^ n6995 ^ n192 ;
  assign n13353 = n13352 ^ n11828 ^ n5493 ;
  assign n13354 = ( n1179 & ~n5211 ) | ( n1179 & n13353 ) | ( ~n5211 & n13353 ) ;
  assign n13356 = n9185 ^ n5456 ^ n410 ;
  assign n13357 = ( n1434 & ~n3903 ) | ( n1434 & n13356 ) | ( ~n3903 & n13356 ) ;
  assign n13358 = n13357 ^ n6157 ^ n1631 ;
  assign n13355 = ( n4408 & ~n9504 ) | ( n4408 & n10200 ) | ( ~n9504 & n10200 ) ;
  assign n13359 = n13358 ^ n13355 ^ n4458 ;
  assign n13360 = ( n143 & n401 ) | ( n143 & n3739 ) | ( n401 & n3739 ) ;
  assign n13361 = n10627 ^ n7191 ^ n7106 ;
  assign n13362 = ( n1484 & n13360 ) | ( n1484 & n13361 ) | ( n13360 & n13361 ) ;
  assign n13363 = n11826 ^ n4838 ^ n2291 ;
  assign n13364 = ( n5388 & n11237 ) | ( n5388 & n13363 ) | ( n11237 & n13363 ) ;
  assign n13371 = ( n452 & ~n5367 ) | ( n452 & n8634 ) | ( ~n5367 & n8634 ) ;
  assign n13372 = n6276 ^ n5954 ^ n559 ;
  assign n13373 = ( n4828 & n13371 ) | ( n4828 & ~n13372 ) | ( n13371 & ~n13372 ) ;
  assign n13368 = ( n1030 & ~n3809 ) | ( n1030 & n4093 ) | ( ~n3809 & n4093 ) ;
  assign n13369 = n13368 ^ n3925 ^ n3611 ;
  assign n13370 = ( n7588 & n10204 ) | ( n7588 & n13369 ) | ( n10204 & n13369 ) ;
  assign n13366 = ( n5269 & n10663 ) | ( n5269 & ~n12602 ) | ( n10663 & ~n12602 ) ;
  assign n13365 = n12900 ^ n1769 ^ n1145 ;
  assign n13367 = n13366 ^ n13365 ^ n11879 ;
  assign n13374 = n13373 ^ n13370 ^ n13367 ;
  assign n13375 = ( n789 & n2317 ) | ( n789 & n10051 ) | ( n2317 & n10051 ) ;
  assign n13376 = n13375 ^ n3303 ^ x89 ;
  assign n13377 = ( n1837 & n7360 ) | ( n1837 & ~n13376 ) | ( n7360 & ~n13376 ) ;
  assign n13378 = ( ~x15 & n365 ) | ( ~x15 & n4831 ) | ( n365 & n4831 ) ;
  assign n13379 = ( n1950 & n3978 ) | ( n1950 & n7808 ) | ( n3978 & n7808 ) ;
  assign n13380 = ( n2976 & n13378 ) | ( n2976 & n13379 ) | ( n13378 & n13379 ) ;
  assign n13381 = n8591 ^ n6302 ^ n948 ;
  assign n13382 = ( ~n366 & n2797 ) | ( ~n366 & n13381 ) | ( n2797 & n13381 ) ;
  assign n13383 = ( ~n3055 & n8653 ) | ( ~n3055 & n13382 ) | ( n8653 & n13382 ) ;
  assign n13384 = ( ~n5353 & n13380 ) | ( ~n5353 & n13383 ) | ( n13380 & n13383 ) ;
  assign n13385 = ( ~n6930 & n7762 ) | ( ~n6930 & n13384 ) | ( n7762 & n13384 ) ;
  assign n13386 = n13330 ^ n6125 ^ n1672 ;
  assign n13387 = ( ~n4361 & n8938 ) | ( ~n4361 & n13386 ) | ( n8938 & n13386 ) ;
  assign n13388 = n13016 ^ n7683 ^ n4819 ;
  assign n13389 = n11441 ^ n6820 ^ n1202 ;
  assign n13390 = n13389 ^ n13366 ^ n6351 ;
  assign n13391 = n8662 ^ n8401 ^ n2281 ;
  assign n13392 = ( ~n13388 & n13390 ) | ( ~n13388 & n13391 ) | ( n13390 & n13391 ) ;
  assign n13393 = ( n5505 & n13387 ) | ( n5505 & ~n13392 ) | ( n13387 & ~n13392 ) ;
  assign n13394 = n6944 ^ n1096 ^ n896 ;
  assign n13395 = n13394 ^ n11727 ^ n1629 ;
  assign n13396 = n13053 ^ n7576 ^ n2817 ;
  assign n13397 = ( ~n2803 & n12139 ) | ( ~n2803 & n13396 ) | ( n12139 & n13396 ) ;
  assign n13398 = n9248 ^ n5587 ^ n1523 ;
  assign n13399 = ( n5119 & n6598 ) | ( n5119 & ~n13398 ) | ( n6598 & ~n13398 ) ;
  assign n13400 = n9321 ^ n9078 ^ n2735 ;
  assign n13401 = n11719 ^ n2859 ^ n959 ;
  assign n13402 = ( n1021 & ~n4359 ) | ( n1021 & n13401 ) | ( ~n4359 & n13401 ) ;
  assign n13403 = ( ~n1034 & n2097 ) | ( ~n1034 & n12203 ) | ( n2097 & n12203 ) ;
  assign n13404 = ( n6417 & n9684 ) | ( n6417 & ~n12371 ) | ( n9684 & ~n12371 ) ;
  assign n13405 = ( ~n13402 & n13403 ) | ( ~n13402 & n13404 ) | ( n13403 & n13404 ) ;
  assign n13406 = n13405 ^ n4490 ^ n977 ;
  assign n13407 = ( n9922 & n13400 ) | ( n9922 & ~n13406 ) | ( n13400 & ~n13406 ) ;
  assign n13412 = n6223 ^ n5625 ^ n1190 ;
  assign n13413 = ( n6169 & ~n10531 ) | ( n6169 & n13412 ) | ( ~n10531 & n13412 ) ;
  assign n13410 = n8220 ^ n1608 ^ n228 ;
  assign n13408 = ( n842 & n1730 ) | ( n842 & ~n4079 ) | ( n1730 & ~n4079 ) ;
  assign n13409 = n13408 ^ n10484 ^ n9169 ;
  assign n13411 = n13410 ^ n13409 ^ n9299 ;
  assign n13414 = n13413 ^ n13411 ^ n8005 ;
  assign n13415 = ( n11002 & ~n11915 ) | ( n11002 & n13414 ) | ( ~n11915 & n13414 ) ;
  assign n13424 = n6159 ^ n3701 ^ n1845 ;
  assign n13425 = ( ~n1201 & n7697 ) | ( ~n1201 & n13424 ) | ( n7697 & n13424 ) ;
  assign n13426 = ( n3134 & n4897 ) | ( n3134 & n13425 ) | ( n4897 & n13425 ) ;
  assign n13417 = n3833 ^ n2844 ^ x9 ;
  assign n13416 = ( n1289 & ~n3892 ) | ( n1289 & n5020 ) | ( ~n3892 & n5020 ) ;
  assign n13418 = n13417 ^ n13416 ^ n5466 ;
  assign n13419 = ( n6565 & n9078 ) | ( n6565 & n9406 ) | ( n9078 & n9406 ) ;
  assign n13420 = ( n3671 & n5247 ) | ( n3671 & n13419 ) | ( n5247 & n13419 ) ;
  assign n13421 = ( n600 & n11050 ) | ( n600 & ~n13420 ) | ( n11050 & ~n13420 ) ;
  assign n13422 = ( n6225 & n6983 ) | ( n6225 & ~n13421 ) | ( n6983 & ~n13421 ) ;
  assign n13423 = ( n2916 & n13418 ) | ( n2916 & ~n13422 ) | ( n13418 & ~n13422 ) ;
  assign n13427 = n13426 ^ n13423 ^ n8637 ;
  assign n13428 = ( ~n4720 & n5189 ) | ( ~n4720 & n11271 ) | ( n5189 & n11271 ) ;
  assign n13429 = n8058 ^ n6023 ^ n4354 ;
  assign n13430 = ( n1341 & n4907 ) | ( n1341 & n13429 ) | ( n4907 & n13429 ) ;
  assign n13431 = n13430 ^ n6731 ^ n1028 ;
  assign n13434 = ( n706 & n3745 ) | ( n706 & n8820 ) | ( n3745 & n8820 ) ;
  assign n13432 = ( n1671 & n1692 ) | ( n1671 & ~n7668 ) | ( n1692 & ~n7668 ) ;
  assign n13433 = n13432 ^ n8760 ^ n1733 ;
  assign n13435 = n13434 ^ n13433 ^ n5390 ;
  assign n13436 = ( n2501 & ~n3594 ) | ( n2501 & n6291 ) | ( ~n3594 & n6291 ) ;
  assign n13437 = n13436 ^ n12915 ^ n11006 ;
  assign n13438 = ( n13204 & n13392 ) | ( n13204 & ~n13437 ) | ( n13392 & ~n13437 ) ;
  assign n13439 = n6454 ^ n5581 ^ n1855 ;
  assign n13440 = ( n7978 & n10863 ) | ( n7978 & n13439 ) | ( n10863 & n13439 ) ;
  assign n13441 = ( n687 & ~n3532 ) | ( n687 & n13440 ) | ( ~n3532 & n13440 ) ;
  assign n13442 = n10329 ^ n3071 ^ n2860 ;
  assign n13443 = n13054 ^ n3822 ^ n2017 ;
  assign n13451 = ( n3052 & n3232 ) | ( n3052 & ~n11050 ) | ( n3232 & ~n11050 ) ;
  assign n13450 = ( n959 & n9196 ) | ( n959 & ~n9223 ) | ( n9196 & ~n9223 ) ;
  assign n13448 = ( n931 & n2916 ) | ( n931 & ~n4652 ) | ( n2916 & ~n4652 ) ;
  assign n13445 = ( n1907 & n3788 ) | ( n1907 & ~n9592 ) | ( n3788 & ~n9592 ) ;
  assign n13446 = ( ~n7217 & n13274 ) | ( ~n7217 & n13445 ) | ( n13274 & n13445 ) ;
  assign n13447 = n13446 ^ n2796 ^ n1010 ;
  assign n13444 = n12514 ^ n12414 ^ n7412 ;
  assign n13449 = n13448 ^ n13447 ^ n13444 ;
  assign n13452 = n13451 ^ n13450 ^ n13449 ;
  assign n13453 = n11547 ^ n8626 ^ n2742 ;
  assign n13454 = n8351 ^ n1850 ^ n1490 ;
  assign n13455 = ( ~n1055 & n7113 ) | ( ~n1055 & n13454 ) | ( n7113 & n13454 ) ;
  assign n13456 = n13455 ^ n6760 ^ n2526 ;
  assign n13457 = ( ~n2283 & n3848 ) | ( ~n2283 & n8573 ) | ( n3848 & n8573 ) ;
  assign n13458 = ( ~n12848 & n13456 ) | ( ~n12848 & n13457 ) | ( n13456 & n13457 ) ;
  assign n13459 = ( x35 & n2314 ) | ( x35 & ~n13291 ) | ( n2314 & ~n13291 ) ;
  assign n13460 = ( ~n3637 & n6038 ) | ( ~n3637 & n13459 ) | ( n6038 & n13459 ) ;
  assign n13461 = ( ~n1435 & n5476 ) | ( ~n1435 & n10126 ) | ( n5476 & n10126 ) ;
  assign n13462 = n13461 ^ n9004 ^ n2017 ;
  assign n13463 = n10040 ^ n8335 ^ n3153 ;
  assign n13464 = n13463 ^ n10560 ^ n5713 ;
  assign n13469 = n9772 ^ n6635 ^ n1080 ;
  assign n13465 = n7900 ^ n5530 ^ n1500 ;
  assign n13466 = n13465 ^ n6531 ^ n4218 ;
  assign n13467 = n13466 ^ n4258 ^ n1588 ;
  assign n13468 = ( n1783 & ~n7031 ) | ( n1783 & n13467 ) | ( ~n7031 & n13467 ) ;
  assign n13470 = n13469 ^ n13468 ^ n9686 ;
  assign n13471 = ( n5870 & n9138 ) | ( n5870 & ~n13470 ) | ( n9138 & ~n13470 ) ;
  assign n13472 = ( n1006 & n5822 ) | ( n1006 & ~n6403 ) | ( n5822 & ~n6403 ) ;
  assign n13473 = ( n4660 & n6271 ) | ( n4660 & ~n13472 ) | ( n6271 & ~n13472 ) ;
  assign n13482 = n5975 ^ n5920 ^ n3734 ;
  assign n13483 = ( n830 & n2250 ) | ( n830 & n2512 ) | ( n2250 & n2512 ) ;
  assign n13484 = n13483 ^ n5690 ^ n252 ;
  assign n13485 = n13484 ^ n12616 ^ n5806 ;
  assign n13486 = ( ~n769 & n13482 ) | ( ~n769 & n13485 ) | ( n13482 & n13485 ) ;
  assign n13479 = ( n2061 & n2599 ) | ( n2061 & ~n10800 ) | ( n2599 & ~n10800 ) ;
  assign n13480 = n13479 ^ n9955 ^ n5416 ;
  assign n13478 = n9255 ^ n3291 ^ n251 ;
  assign n13481 = n13480 ^ n13478 ^ n2334 ;
  assign n13474 = n9775 ^ n1026 ^ n898 ;
  assign n13475 = n13474 ^ n8855 ^ n8703 ;
  assign n13476 = n13475 ^ n3521 ^ n1440 ;
  assign n13477 = ( n5815 & n7289 ) | ( n5815 & ~n13476 ) | ( n7289 & ~n13476 ) ;
  assign n13487 = n13486 ^ n13481 ^ n13477 ;
  assign n13488 = ( n2079 & n8695 ) | ( n2079 & n11422 ) | ( n8695 & n11422 ) ;
  assign n13489 = n13488 ^ n6403 ^ n5974 ;
  assign n13496 = n3641 ^ n2961 ^ n1889 ;
  assign n13494 = n10126 ^ n8365 ^ n5125 ;
  assign n13490 = ( n2768 & n5373 ) | ( n2768 & ~n8837 ) | ( n5373 & ~n8837 ) ;
  assign n13491 = n13490 ^ n2198 ^ n1403 ;
  assign n13492 = n13491 ^ n12780 ^ n6889 ;
  assign n13493 = ( n428 & n8362 ) | ( n428 & n13492 ) | ( n8362 & n13492 ) ;
  assign n13495 = n13494 ^ n13493 ^ n11051 ;
  assign n13497 = n13496 ^ n13495 ^ n2379 ;
  assign n13498 = ( n4384 & ~n5035 ) | ( n4384 & n11934 ) | ( ~n5035 & n11934 ) ;
  assign n13499 = ( n5284 & ~n12507 ) | ( n5284 & n13498 ) | ( ~n12507 & n13498 ) ;
  assign n13500 = n13499 ^ n4240 ^ n3162 ;
  assign n13501 = n9015 ^ n5424 ^ n4452 ;
  assign n13502 = ( n5470 & n12402 ) | ( n5470 & ~n13501 ) | ( n12402 & ~n13501 ) ;
  assign n13503 = ( n1373 & n2098 ) | ( n1373 & n2772 ) | ( n2098 & n2772 ) ;
  assign n13504 = n13503 ^ n3819 ^ n1578 ;
  assign n13505 = ( ~n4000 & n6513 ) | ( ~n4000 & n13504 ) | ( n6513 & n13504 ) ;
  assign n13506 = ( n1473 & n5357 ) | ( n1473 & n7823 ) | ( n5357 & n7823 ) ;
  assign n13507 = ( ~n7722 & n13505 ) | ( ~n7722 & n13506 ) | ( n13505 & n13506 ) ;
  assign n13508 = n13507 ^ n7343 ^ n2517 ;
  assign n13509 = ( n8801 & n11268 ) | ( n8801 & ~n13508 ) | ( n11268 & ~n13508 ) ;
  assign n13510 = ( n3951 & n7452 ) | ( n3951 & ~n11054 ) | ( n7452 & ~n11054 ) ;
  assign n13511 = ( n651 & n9460 ) | ( n651 & ~n13510 ) | ( n9460 & ~n13510 ) ;
  assign n13512 = n13511 ^ n6306 ^ n2766 ;
  assign n13513 = n13512 ^ n5495 ^ n4861 ;
  assign n13514 = ( n4773 & n4885 ) | ( n4773 & n7944 ) | ( n4885 & n7944 ) ;
  assign n13515 = n13514 ^ n4764 ^ n2380 ;
  assign n13516 = ( n575 & ~n1683 ) | ( n575 & n13515 ) | ( ~n1683 & n13515 ) ;
  assign n13517 = n13516 ^ n10909 ^ n1912 ;
  assign n13519 = ( ~n4435 & n6068 ) | ( ~n4435 & n10464 ) | ( n6068 & n10464 ) ;
  assign n13518 = n13067 ^ n10029 ^ n3581 ;
  assign n13520 = n13519 ^ n13518 ^ n3857 ;
  assign n13523 = ( n2097 & n11934 ) | ( n2097 & ~n12479 ) | ( n11934 & ~n12479 ) ;
  assign n13524 = n13523 ^ n4642 ^ n2253 ;
  assign n13525 = ( n6118 & n9067 ) | ( n6118 & n13524 ) | ( n9067 & n13524 ) ;
  assign n13521 = ( n7262 & ~n9484 ) | ( n7262 & n11012 ) | ( ~n9484 & n11012 ) ;
  assign n13522 = ( n4875 & n5746 ) | ( n4875 & n13521 ) | ( n5746 & n13521 ) ;
  assign n13526 = n13525 ^ n13522 ^ n621 ;
  assign n13527 = ( n2259 & n7609 ) | ( n2259 & ~n11197 ) | ( n7609 & ~n11197 ) ;
  assign n13528 = ( n357 & n3449 ) | ( n357 & ~n13527 ) | ( n3449 & ~n13527 ) ;
  assign n13529 = ( n955 & n5321 ) | ( n955 & ~n9492 ) | ( n5321 & ~n9492 ) ;
  assign n13530 = ( ~n6756 & n9974 ) | ( ~n6756 & n13529 ) | ( n9974 & n13529 ) ;
  assign n13531 = ( ~n1155 & n6616 ) | ( ~n1155 & n11524 ) | ( n6616 & n11524 ) ;
  assign n13532 = ( n1536 & n3234 ) | ( n1536 & n4360 ) | ( n3234 & n4360 ) ;
  assign n13533 = n13532 ^ n3097 ^ n651 ;
  assign n13534 = n13533 ^ n4409 ^ n569 ;
  assign n13535 = ( ~n13512 & n13531 ) | ( ~n13512 & n13534 ) | ( n13531 & n13534 ) ;
  assign n13536 = n2796 ^ n2542 ^ n774 ;
  assign n13537 = n13536 ^ n12890 ^ n2407 ;
  assign n13538 = ( n10173 & n11570 ) | ( n10173 & n13537 ) | ( n11570 & n13537 ) ;
  assign n13539 = ( n1448 & ~n4080 ) | ( n1448 & n13538 ) | ( ~n4080 & n13538 ) ;
  assign n13540 = ( n399 & n2260 ) | ( n399 & ~n4443 ) | ( n2260 & ~n4443 ) ;
  assign n13541 = n5563 ^ n1354 ^ n1197 ;
  assign n13542 = ( n11003 & n13540 ) | ( n11003 & ~n13541 ) | ( n13540 & ~n13541 ) ;
  assign n13543 = ( n3504 & n6994 ) | ( n3504 & n10626 ) | ( n6994 & n10626 ) ;
  assign n13544 = n13543 ^ n12000 ^ n634 ;
  assign n13545 = ( n1862 & n7729 ) | ( n1862 & n13544 ) | ( n7729 & n13544 ) ;
  assign n13546 = n10468 ^ n6023 ^ n2766 ;
  assign n13547 = ( n1373 & n3164 ) | ( n1373 & n13546 ) | ( n3164 & n13546 ) ;
  assign n13548 = ( n1036 & n4691 ) | ( n1036 & n5361 ) | ( n4691 & n5361 ) ;
  assign n13549 = n13548 ^ n7416 ^ n4910 ;
  assign n13550 = ( n1867 & n3113 ) | ( n1867 & n7809 ) | ( n3113 & n7809 ) ;
  assign n13551 = n13550 ^ n3582 ^ n2827 ;
  assign n13555 = ( n2505 & n4551 ) | ( n2505 & n13091 ) | ( n4551 & n13091 ) ;
  assign n13556 = ( n2669 & n12090 ) | ( n2669 & n13555 ) | ( n12090 & n13555 ) ;
  assign n13553 = ( n3005 & n3539 ) | ( n3005 & n3834 ) | ( n3539 & n3834 ) ;
  assign n13552 = n12661 ^ n9464 ^ n5595 ;
  assign n13554 = n13553 ^ n13552 ^ n9651 ;
  assign n13557 = n13556 ^ n13554 ^ n9924 ;
  assign n13558 = n2994 ^ n1793 ^ n404 ;
  assign n13559 = ( ~n926 & n3957 ) | ( ~n926 & n13558 ) | ( n3957 & n13558 ) ;
  assign n13560 = ( ~x34 & n8459 ) | ( ~x34 & n11840 ) | ( n8459 & n11840 ) ;
  assign n13561 = n13560 ^ n4129 ^ n390 ;
  assign n13562 = ( n2093 & n13559 ) | ( n2093 & n13561 ) | ( n13559 & n13561 ) ;
  assign n13563 = ( n6272 & n6979 ) | ( n6272 & n7405 ) | ( n6979 & n7405 ) ;
  assign n13564 = n5202 ^ n3584 ^ n1360 ;
  assign n13565 = n13564 ^ n9800 ^ n9400 ;
  assign n13568 = ( n1047 & n2328 ) | ( n1047 & n4982 ) | ( n2328 & n4982 ) ;
  assign n13566 = ( ~n1816 & n5383 ) | ( ~n1816 & n7105 ) | ( n5383 & n7105 ) ;
  assign n13567 = n13566 ^ n11630 ^ n811 ;
  assign n13569 = n13568 ^ n13567 ^ n434 ;
  assign n13570 = ( ~n13563 & n13565 ) | ( ~n13563 & n13569 ) | ( n13565 & n13569 ) ;
  assign n13571 = ( ~n5312 & n8746 ) | ( ~n5312 & n12089 ) | ( n8746 & n12089 ) ;
  assign n13572 = n7328 ^ n5843 ^ n4016 ;
  assign n13573 = ( n8325 & n13571 ) | ( n8325 & ~n13572 ) | ( n13571 & ~n13572 ) ;
  assign n13574 = n13258 ^ n12503 ^ n5204 ;
  assign n13578 = n3647 ^ n2719 ^ n1211 ;
  assign n13579 = n13578 ^ n7917 ^ n5248 ;
  assign n13580 = ( n1185 & ~n7335 ) | ( n1185 & n13579 ) | ( ~n7335 & n13579 ) ;
  assign n13576 = n8813 ^ n3561 ^ x6 ;
  assign n13577 = ( ~n7449 & n8461 ) | ( ~n7449 & n13576 ) | ( n8461 & n13576 ) ;
  assign n13575 = n10915 ^ n6722 ^ n1122 ;
  assign n13581 = n13580 ^ n13577 ^ n13575 ;
  assign n13582 = ( ~n512 & n523 ) | ( ~n512 & n8569 ) | ( n523 & n8569 ) ;
  assign n13583 = n8474 ^ n2511 ^ n2368 ;
  assign n13584 = ( n3770 & n3903 ) | ( n3770 & n13583 ) | ( n3903 & n13583 ) ;
  assign n13593 = ( x107 & n5763 ) | ( x107 & n9117 ) | ( n5763 & n9117 ) ;
  assign n13587 = ( n562 & n660 ) | ( n562 & ~n7511 ) | ( n660 & ~n7511 ) ;
  assign n13588 = n13587 ^ n8064 ^ n7577 ;
  assign n13589 = n3841 ^ n2335 ^ n1241 ;
  assign n13590 = ( n711 & n11082 ) | ( n711 & ~n13589 ) | ( n11082 & ~n13589 ) ;
  assign n13591 = ( ~n6990 & n8749 ) | ( ~n6990 & n13590 ) | ( n8749 & n13590 ) ;
  assign n13592 = ( n826 & n13588 ) | ( n826 & n13591 ) | ( n13588 & n13591 ) ;
  assign n13585 = n11640 ^ n6830 ^ n5696 ;
  assign n13586 = n13585 ^ n4691 ^ n1611 ;
  assign n13594 = n13593 ^ n13592 ^ n13586 ;
  assign n13595 = ( x36 & n2067 ) | ( x36 & ~n13310 ) | ( n2067 & ~n13310 ) ;
  assign n13596 = n12426 ^ n8803 ^ n5323 ;
  assign n13597 = ( n11449 & n13595 ) | ( n11449 & ~n13596 ) | ( n13595 & ~n13596 ) ;
  assign n13598 = ( n8079 & ~n8553 ) | ( n8079 & n12024 ) | ( ~n8553 & n12024 ) ;
  assign n13599 = ( n1577 & n6863 ) | ( n1577 & ~n13421 ) | ( n6863 & ~n13421 ) ;
  assign n13600 = ( n4475 & n13598 ) | ( n4475 & n13599 ) | ( n13598 & n13599 ) ;
  assign n13601 = n13383 ^ n11011 ^ x44 ;
  assign n13602 = ( ~n4015 & n11506 ) | ( ~n4015 & n13601 ) | ( n11506 & n13601 ) ;
  assign n13603 = ( n1736 & n2232 ) | ( n1736 & n8290 ) | ( n2232 & n8290 ) ;
  assign n13604 = ( ~n4194 & n5596 ) | ( ~n4194 & n11754 ) | ( n5596 & n11754 ) ;
  assign n13611 = n11151 ^ n7031 ^ n2302 ;
  assign n13607 = n8075 ^ n4641 ^ n4573 ;
  assign n13608 = ( ~n259 & n2409 ) | ( ~n259 & n3547 ) | ( n2409 & n3547 ) ;
  assign n13609 = ( ~n8802 & n9235 ) | ( ~n8802 & n13608 ) | ( n9235 & n13608 ) ;
  assign n13610 = ( n4661 & n13607 ) | ( n4661 & n13609 ) | ( n13607 & n13609 ) ;
  assign n13612 = n13611 ^ n13610 ^ n2563 ;
  assign n13605 = n12929 ^ n9676 ^ n7352 ;
  assign n13606 = n13605 ^ n2982 ^ n816 ;
  assign n13613 = n13612 ^ n13606 ^ n831 ;
  assign n13614 = n11152 ^ n4415 ^ n3226 ;
  assign n13615 = ( ~n912 & n2040 ) | ( ~n912 & n9091 ) | ( n2040 & n9091 ) ;
  assign n13616 = ( n1925 & ~n13614 ) | ( n1925 & n13615 ) | ( ~n13614 & n13615 ) ;
  assign n13617 = ( x119 & n722 ) | ( x119 & ~n9772 ) | ( n722 & ~n9772 ) ;
  assign n13618 = ( n2520 & ~n6140 ) | ( n2520 & n11819 ) | ( ~n6140 & n11819 ) ;
  assign n13619 = ( n1310 & n13617 ) | ( n1310 & n13618 ) | ( n13617 & n13618 ) ;
  assign n13620 = n13619 ^ n12453 ^ n8912 ;
  assign n13621 = n10128 ^ n8925 ^ n4034 ;
  assign n13622 = ( n11684 & n13620 ) | ( n11684 & ~n13621 ) | ( n13620 & ~n13621 ) ;
  assign n13623 = ( n2459 & n4767 ) | ( n2459 & n6852 ) | ( n4767 & n6852 ) ;
  assign n13624 = n11020 ^ n10308 ^ n2474 ;
  assign n13625 = n10645 ^ n9175 ^ n5555 ;
  assign n13626 = n4217 ^ n1900 ^ n775 ;
  assign n13627 = ( n1833 & n6293 ) | ( n1833 & n13626 ) | ( n6293 & n13626 ) ;
  assign n13628 = n13627 ^ n8590 ^ n6943 ;
  assign n13634 = ( ~n473 & n1252 ) | ( ~n473 & n1949 ) | ( n1252 & n1949 ) ;
  assign n13635 = n13634 ^ n10054 ^ n5316 ;
  assign n13631 = ( n170 & n8249 ) | ( n170 & n12879 ) | ( n8249 & n12879 ) ;
  assign n13632 = n13631 ^ n7339 ^ n1097 ;
  assign n13633 = ( n290 & n9192 ) | ( n290 & n13632 ) | ( n9192 & n13632 ) ;
  assign n13636 = n13635 ^ n13633 ^ n3016 ;
  assign n13629 = ( n3622 & n4101 ) | ( n3622 & ~n6830 ) | ( n4101 & ~n6830 ) ;
  assign n13630 = n13629 ^ n11567 ^ n8499 ;
  assign n13637 = n13636 ^ n13630 ^ n10346 ;
  assign n13638 = ( n2213 & n4625 ) | ( n2213 & ~n11330 ) | ( n4625 & ~n11330 ) ;
  assign n13639 = n13638 ^ n9620 ^ x17 ;
  assign n13641 = n8778 ^ n6649 ^ n5689 ;
  assign n13640 = ( n1180 & n3831 ) | ( n1180 & n8796 ) | ( n3831 & n8796 ) ;
  assign n13642 = n13641 ^ n13640 ^ n6488 ;
  assign n13643 = ( ~n10351 & n12317 ) | ( ~n10351 & n13642 ) | ( n12317 & n13642 ) ;
  assign n13644 = n11915 ^ n11263 ^ n5854 ;
  assign n13646 = n7336 ^ n6432 ^ n4624 ;
  assign n13645 = ( n433 & ~n2570 ) | ( n433 & n3770 ) | ( ~n2570 & n3770 ) ;
  assign n13647 = n13646 ^ n13645 ^ n5102 ;
  assign n13648 = ( n7641 & ~n13644 ) | ( n7641 & n13647 ) | ( ~n13644 & n13647 ) ;
  assign n13649 = ( n1325 & n4332 ) | ( n1325 & n13648 ) | ( n4332 & n13648 ) ;
  assign n13650 = ( n10048 & n10756 ) | ( n10048 & ~n13649 ) | ( n10756 & ~n13649 ) ;
  assign n13651 = ( ~n1879 & n8463 ) | ( ~n1879 & n13170 ) | ( n8463 & n13170 ) ;
  assign n13652 = ( ~n3138 & n6807 ) | ( ~n3138 & n13651 ) | ( n6807 & n13651 ) ;
  assign n13653 = n6049 ^ n4436 ^ n3917 ;
  assign n13654 = ( n280 & n4307 ) | ( n280 & ~n13653 ) | ( n4307 & ~n13653 ) ;
  assign n13655 = n8836 ^ n7918 ^ n838 ;
  assign n13656 = ( n7674 & n13654 ) | ( n7674 & n13655 ) | ( n13654 & n13655 ) ;
  assign n13657 = ( n990 & n3443 ) | ( n990 & n13656 ) | ( n3443 & n13656 ) ;
  assign n13663 = ( n1764 & ~n3076 ) | ( n1764 & n4882 ) | ( ~n3076 & n4882 ) ;
  assign n13660 = ( n6537 & n9403 ) | ( n6537 & ~n10191 ) | ( n9403 & ~n10191 ) ;
  assign n13661 = ( ~n2096 & n3140 ) | ( ~n2096 & n13660 ) | ( n3140 & n13660 ) ;
  assign n13658 = ( n2236 & ~n4165 ) | ( n2236 & n11177 ) | ( ~n4165 & n11177 ) ;
  assign n13659 = ( n11222 & n12732 ) | ( n11222 & n13658 ) | ( n12732 & n13658 ) ;
  assign n13662 = n13661 ^ n13659 ^ n9531 ;
  assign n13664 = n13663 ^ n13662 ^ n10846 ;
  assign n13665 = n10477 ^ n6443 ^ n4955 ;
  assign n13671 = n4806 ^ n4010 ^ n225 ;
  assign n13669 = n7961 ^ n6458 ^ n6383 ;
  assign n13670 = n13669 ^ n8012 ^ x115 ;
  assign n13666 = ( n4375 & n9774 ) | ( n4375 & n12133 ) | ( n9774 & n12133 ) ;
  assign n13667 = n13666 ^ n10868 ^ n5106 ;
  assign n13668 = n13667 ^ n6301 ^ n5699 ;
  assign n13672 = n13671 ^ n13670 ^ n13668 ;
  assign n13673 = ( ~n4945 & n10912 ) | ( ~n4945 & n10976 ) | ( n10912 & n10976 ) ;
  assign n13674 = ( ~n738 & n1311 ) | ( ~n738 & n6308 ) | ( n1311 & n6308 ) ;
  assign n13675 = n13674 ^ n8544 ^ n2997 ;
  assign n13676 = ( n1022 & ~n11498 ) | ( n1022 & n13675 ) | ( ~n11498 & n13675 ) ;
  assign n13677 = n9999 ^ n9200 ^ n7705 ;
  assign n13678 = n13677 ^ n9437 ^ n3366 ;
  assign n13679 = ( n352 & ~n2418 ) | ( n352 & n13678 ) | ( ~n2418 & n13678 ) ;
  assign n13686 = ( n290 & n1252 ) | ( n290 & ~n5109 ) | ( n1252 & ~n5109 ) ;
  assign n13687 = n13686 ^ n11669 ^ n229 ;
  assign n13688 = ( ~n4374 & n12704 ) | ( ~n4374 & n13687 ) | ( n12704 & n13687 ) ;
  assign n13690 = ( n2930 & ~n6460 ) | ( n2930 & n10130 ) | ( ~n6460 & n10130 ) ;
  assign n13681 = ( ~n1072 & n4170 ) | ( ~n1072 & n12320 ) | ( n4170 & n12320 ) ;
  assign n13689 = n13681 ^ n7294 ^ n1301 ;
  assign n13691 = n13690 ^ n13689 ^ n5908 ;
  assign n13692 = ( n7126 & n13688 ) | ( n7126 & n13691 ) | ( n13688 & n13691 ) ;
  assign n13680 = ( n4253 & n6963 ) | ( n4253 & ~n9761 ) | ( n6963 & ~n9761 ) ;
  assign n13682 = n13681 ^ n9019 ^ n1223 ;
  assign n13683 = ( n1424 & n13680 ) | ( n1424 & n13682 ) | ( n13680 & n13682 ) ;
  assign n13684 = n9149 ^ n5600 ^ n2026 ;
  assign n13685 = ( n8807 & ~n13683 ) | ( n8807 & n13684 ) | ( ~n13683 & n13684 ) ;
  assign n13693 = n13692 ^ n13685 ^ n6371 ;
  assign n13695 = ( n5770 & ~n10451 ) | ( n5770 & n10545 ) | ( ~n10451 & n10545 ) ;
  assign n13694 = n9316 ^ n6432 ^ n267 ;
  assign n13696 = n13695 ^ n13694 ^ n7564 ;
  assign n13697 = ( ~n3363 & n4432 ) | ( ~n3363 & n5144 ) | ( n4432 & n5144 ) ;
  assign n13698 = ( n5596 & n11575 ) | ( n5596 & ~n13697 ) | ( n11575 & ~n13697 ) ;
  assign n13699 = n13698 ^ n6807 ^ n2973 ;
  assign n13700 = ( n1007 & n3069 ) | ( n1007 & n5231 ) | ( n3069 & n5231 ) ;
  assign n13701 = ( x38 & n5399 ) | ( x38 & ~n13700 ) | ( n5399 & ~n13700 ) ;
  assign n13702 = ( n697 & ~n11855 ) | ( n697 & n13701 ) | ( ~n11855 & n13701 ) ;
  assign n13708 = ( n2604 & ~n6329 ) | ( n2604 & n9855 ) | ( ~n6329 & n9855 ) ;
  assign n13704 = ( ~n950 & n1082 ) | ( ~n950 & n2279 ) | ( n1082 & n2279 ) ;
  assign n13705 = ( n2910 & n12780 ) | ( n2910 & ~n13704 ) | ( n12780 & ~n13704 ) ;
  assign n13706 = ( n1213 & ~n2834 ) | ( n1213 & n13705 ) | ( ~n2834 & n13705 ) ;
  assign n13703 = ( n1126 & ~n4172 ) | ( n1126 & n7783 ) | ( ~n4172 & n7783 ) ;
  assign n13707 = n13706 ^ n13703 ^ n11854 ;
  assign n13709 = n13708 ^ n13707 ^ n6396 ;
  assign n13710 = n10679 ^ n3394 ^ n304 ;
  assign n13711 = n13710 ^ n5101 ^ n4862 ;
  assign n13712 = n13711 ^ n11990 ^ n6357 ;
  assign n13714 = n12719 ^ n9013 ^ n5217 ;
  assign n13715 = n13714 ^ n9683 ^ n2762 ;
  assign n13713 = n7084 ^ n6267 ^ n2378 ;
  assign n13716 = n13715 ^ n13713 ^ n3455 ;
  assign n13717 = n9931 ^ n7949 ^ n2745 ;
  assign n13718 = ( n4152 & n10098 ) | ( n4152 & n13717 ) | ( n10098 & n13717 ) ;
  assign n13720 = n9678 ^ n4104 ^ n589 ;
  assign n13719 = ( n1617 & ~n1847 ) | ( n1617 & n11580 ) | ( ~n1847 & n11580 ) ;
  assign n13721 = n13720 ^ n13719 ^ n243 ;
  assign n13722 = ( n931 & n1185 ) | ( n931 & n1280 ) | ( n1185 & n1280 ) ;
  assign n13723 = ( n644 & n11336 ) | ( n644 & n13722 ) | ( n11336 & n13722 ) ;
  assign n13724 = n13723 ^ n5982 ^ n4226 ;
  assign n13725 = n13724 ^ n7574 ^ n1563 ;
  assign n13726 = n8417 ^ n6556 ^ n6460 ;
  assign n13727 = ( n3942 & n7163 ) | ( n3942 & n13726 ) | ( n7163 & n13726 ) ;
  assign n13730 = ( n4927 & n7591 ) | ( n4927 & n7997 ) | ( n7591 & n7997 ) ;
  assign n13731 = ( n737 & ~n12044 ) | ( n737 & n13730 ) | ( ~n12044 & n13730 ) ;
  assign n13729 = ( n794 & n4823 ) | ( n794 & ~n12440 ) | ( n4823 & ~n12440 ) ;
  assign n13728 = n12145 ^ n10043 ^ n8899 ;
  assign n13732 = n13731 ^ n13729 ^ n13728 ;
  assign n13733 = ( n2864 & ~n5969 ) | ( n2864 & n13732 ) | ( ~n5969 & n13732 ) ;
  assign n13734 = ( ~n2044 & n3068 ) | ( ~n2044 & n5524 ) | ( n3068 & n5524 ) ;
  assign n13735 = ( ~n1816 & n5327 ) | ( ~n1816 & n7063 ) | ( n5327 & n7063 ) ;
  assign n13736 = ( n1403 & n13734 ) | ( n1403 & ~n13735 ) | ( n13734 & ~n13735 ) ;
  assign n13737 = ( n433 & n6313 ) | ( n433 & n10023 ) | ( n6313 & n10023 ) ;
  assign n13738 = ( ~n6748 & n9796 ) | ( ~n6748 & n13737 ) | ( n9796 & n13737 ) ;
  assign n13745 = ( ~n2912 & n7276 ) | ( ~n2912 & n12241 ) | ( n7276 & n12241 ) ;
  assign n13739 = ( n7347 & ~n8499 ) | ( n7347 & n10369 ) | ( ~n8499 & n10369 ) ;
  assign n13740 = n13739 ^ n8029 ^ n7022 ;
  assign n13741 = ( n219 & n2511 ) | ( n219 & ~n3946 ) | ( n2511 & ~n3946 ) ;
  assign n13742 = n13741 ^ n2583 ^ n252 ;
  assign n13743 = ( n9728 & n12233 ) | ( n9728 & ~n13742 ) | ( n12233 & ~n13742 ) ;
  assign n13744 = ( n8150 & ~n13740 ) | ( n8150 & n13743 ) | ( ~n13740 & n13743 ) ;
  assign n13746 = n13745 ^ n13744 ^ n484 ;
  assign n13747 = ( n729 & ~n1911 ) | ( n729 & n9898 ) | ( ~n1911 & n9898 ) ;
  assign n13748 = n10765 ^ n4783 ^ n780 ;
  assign n13749 = n13748 ^ n12337 ^ n8948 ;
  assign n13750 = ( n1486 & n8501 ) | ( n1486 & ~n12654 ) | ( n8501 & ~n12654 ) ;
  assign n13751 = n13750 ^ n10621 ^ n1305 ;
  assign n13752 = ( n3196 & n13749 ) | ( n3196 & ~n13751 ) | ( n13749 & ~n13751 ) ;
  assign n13753 = ( n2845 & n4747 ) | ( n2845 & ~n10636 ) | ( n4747 & ~n10636 ) ;
  assign n13754 = ( n579 & n9748 ) | ( n579 & n10202 ) | ( n9748 & n10202 ) ;
  assign n13755 = ( n1301 & n3069 ) | ( n1301 & ~n4831 ) | ( n3069 & ~n4831 ) ;
  assign n13756 = ( n2018 & n4925 ) | ( n2018 & n13755 ) | ( n4925 & n13755 ) ;
  assign n13757 = n6715 ^ n2327 ^ n1226 ;
  assign n13758 = ( x105 & n3136 ) | ( x105 & n13757 ) | ( n3136 & n13757 ) ;
  assign n13759 = ( n8500 & ~n13756 ) | ( n8500 & n13758 ) | ( ~n13756 & n13758 ) ;
  assign n13760 = n13759 ^ n2532 ^ n141 ;
  assign n13762 = ( ~n2020 & n5222 ) | ( ~n2020 & n10908 ) | ( n5222 & n10908 ) ;
  assign n13761 = n8066 ^ n6974 ^ x44 ;
  assign n13763 = n13762 ^ n13761 ^ n234 ;
  assign n13765 = n4995 ^ n3178 ^ n135 ;
  assign n13766 = n13765 ^ n4162 ^ n3407 ;
  assign n13764 = ( ~n2859 & n2948 ) | ( ~n2859 & n10670 ) | ( n2948 & n10670 ) ;
  assign n13767 = n13766 ^ n13764 ^ n12428 ;
  assign n13768 = ( n453 & ~n8801 ) | ( n453 & n12623 ) | ( ~n8801 & n12623 ) ;
  assign n13770 = n11769 ^ n2561 ^ n2528 ;
  assign n13769 = ( n4499 & n8487 ) | ( n4499 & n9490 ) | ( n8487 & n9490 ) ;
  assign n13771 = n13770 ^ n13769 ^ n9897 ;
  assign n13772 = n13771 ^ n13220 ^ n6915 ;
  assign n13773 = n5795 ^ n1169 ^ n499 ;
  assign n13774 = n4591 ^ n4325 ^ n961 ;
  assign n13775 = ( ~n3306 & n4734 ) | ( ~n3306 & n13774 ) | ( n4734 & n13774 ) ;
  assign n13776 = n13775 ^ n7339 ^ n5567 ;
  assign n13777 = ( n5334 & ~n10999 ) | ( n5334 & n13776 ) | ( ~n10999 & n13776 ) ;
  assign n13781 = ( n2931 & ~n3268 ) | ( n2931 & n13273 ) | ( ~n3268 & n13273 ) ;
  assign n13778 = n2831 ^ n2303 ^ n1580 ;
  assign n13779 = ( ~n5505 & n9046 ) | ( ~n5505 & n13778 ) | ( n9046 & n13778 ) ;
  assign n13780 = ( n5895 & ~n11919 ) | ( n5895 & n13779 ) | ( ~n11919 & n13779 ) ;
  assign n13782 = n13781 ^ n13780 ^ n9398 ;
  assign n13783 = ( n13773 & ~n13777 ) | ( n13773 & n13782 ) | ( ~n13777 & n13782 ) ;
  assign n13784 = ( n810 & n2870 ) | ( n810 & n4278 ) | ( n2870 & n4278 ) ;
  assign n13785 = n10106 ^ n6346 ^ n1913 ;
  assign n13786 = n13785 ^ n3515 ^ n1522 ;
  assign n13787 = n13786 ^ n13430 ^ n7675 ;
  assign n13788 = ( ~n12790 & n13784 ) | ( ~n12790 & n13787 ) | ( n13784 & n13787 ) ;
  assign n13791 = ( n2111 & n7174 ) | ( n2111 & ~n10351 ) | ( n7174 & ~n10351 ) ;
  assign n13789 = ( ~n1704 & n2159 ) | ( ~n1704 & n12581 ) | ( n2159 & n12581 ) ;
  assign n13790 = ( n5646 & ~n7017 ) | ( n5646 & n13789 ) | ( ~n7017 & n13789 ) ;
  assign n13792 = n13791 ^ n13790 ^ n3258 ;
  assign n13793 = ( n5841 & ~n8632 ) | ( n5841 & n10771 ) | ( ~n8632 & n10771 ) ;
  assign n13794 = ( n494 & n3849 ) | ( n494 & ~n13793 ) | ( n3849 & ~n13793 ) ;
  assign n13795 = n13705 ^ n8191 ^ n440 ;
  assign n13796 = ( n7345 & ~n11109 ) | ( n7345 & n13795 ) | ( ~n11109 & n13795 ) ;
  assign n13797 = n13796 ^ n7896 ^ n2013 ;
  assign n13798 = n5837 ^ n2849 ^ n646 ;
  assign n13799 = ( n3676 & ~n7964 ) | ( n3676 & n13798 ) | ( ~n7964 & n13798 ) ;
  assign n13800 = ( n1410 & ~n13797 ) | ( n1410 & n13799 ) | ( ~n13797 & n13799 ) ;
  assign n13801 = ( ~n2005 & n3159 ) | ( ~n2005 & n5528 ) | ( n3159 & n5528 ) ;
  assign n13802 = ( n3150 & n6189 ) | ( n3150 & n13801 ) | ( n6189 & n13801 ) ;
  assign n13803 = n3728 ^ n3515 ^ n1070 ;
  assign n13804 = n13803 ^ n3554 ^ x103 ;
  assign n13805 = n13804 ^ n8094 ^ n7313 ;
  assign n13806 = ( n287 & n6303 ) | ( n287 & ~n11266 ) | ( n6303 & ~n11266 ) ;
  assign n13807 = n13806 ^ n5847 ^ n4171 ;
  assign n13808 = ( n10856 & ~n12987 ) | ( n10856 & n13807 ) | ( ~n12987 & n13807 ) ;
  assign n13809 = ( n9575 & n9974 ) | ( n9575 & ~n13808 ) | ( n9974 & ~n13808 ) ;
  assign n13810 = n13809 ^ n7220 ^ n6988 ;
  assign n13818 = n9496 ^ n7158 ^ n881 ;
  assign n13819 = n13818 ^ n8324 ^ n6751 ;
  assign n13820 = n13819 ^ n4030 ^ n988 ;
  assign n13821 = ( n2670 & n6484 ) | ( n2670 & n13820 ) | ( n6484 & n13820 ) ;
  assign n13822 = n13821 ^ n13211 ^ n12511 ;
  assign n13817 = ( n6075 & n6410 ) | ( n6075 & ~n11726 ) | ( n6410 & ~n11726 ) ;
  assign n13823 = n13822 ^ n13817 ^ n10408 ;
  assign n13811 = n3536 ^ n3515 ^ n2354 ;
  assign n13812 = n13811 ^ n8395 ^ n1442 ;
  assign n13813 = ( n1147 & n2070 ) | ( n1147 & ~n13812 ) | ( n2070 & ~n13812 ) ;
  assign n13814 = n5055 ^ n2855 ^ n1710 ;
  assign n13815 = n13814 ^ n7787 ^ n387 ;
  assign n13816 = ( ~n4570 & n13813 ) | ( ~n4570 & n13815 ) | ( n13813 & n13815 ) ;
  assign n13824 = n13823 ^ n13816 ^ n8087 ;
  assign n13825 = n8050 ^ n6672 ^ n1225 ;
  assign n13826 = ( n1666 & ~n3785 ) | ( n1666 & n9985 ) | ( ~n3785 & n9985 ) ;
  assign n13827 = ( n468 & n4200 ) | ( n468 & ~n13826 ) | ( n4200 & ~n13826 ) ;
  assign n13828 = n13827 ^ n5686 ^ n4414 ;
  assign n13829 = ( n12197 & n13825 ) | ( n12197 & ~n13828 ) | ( n13825 & ~n13828 ) ;
  assign n13830 = n13829 ^ n10813 ^ n1670 ;
  assign n13831 = ( n2399 & n3792 ) | ( n2399 & ~n4048 ) | ( n3792 & ~n4048 ) ;
  assign n13832 = n13831 ^ n13521 ^ n2187 ;
  assign n13833 = n9436 ^ n6618 ^ n1649 ;
  assign n13834 = n13833 ^ n10028 ^ n5171 ;
  assign n13835 = n13834 ^ n10731 ^ n5100 ;
  assign n13836 = ( x65 & n13832 ) | ( x65 & ~n13835 ) | ( n13832 & ~n13835 ) ;
  assign n13837 = ( n4278 & n13592 ) | ( n4278 & n13836 ) | ( n13592 & n13836 ) ;
  assign n13838 = n9737 ^ n7381 ^ n1076 ;
  assign n13839 = n13838 ^ n11823 ^ n9676 ;
  assign n13840 = n13839 ^ n6431 ^ n268 ;
  assign n13841 = ( n3119 & n6038 ) | ( n3119 & ~n9117 ) | ( n6038 & ~n9117 ) ;
  assign n13842 = n2204 ^ n1026 ^ x0 ;
  assign n13843 = ( n5804 & n9855 ) | ( n5804 & ~n13842 ) | ( n9855 & ~n13842 ) ;
  assign n13844 = ( n11637 & ~n13841 ) | ( n11637 & n13843 ) | ( ~n13841 & n13843 ) ;
  assign n13845 = ( n8295 & ~n8974 ) | ( n8295 & n13844 ) | ( ~n8974 & n13844 ) ;
  assign n13846 = n3043 ^ n2301 ^ x20 ;
  assign n13847 = n13846 ^ n1487 ^ n555 ;
  assign n13848 = n11995 ^ n7365 ^ x117 ;
  assign n13849 = ( n5128 & ~n5202 ) | ( n5128 & n13848 ) | ( ~n5202 & n13848 ) ;
  assign n13853 = n3592 ^ n2482 ^ n718 ;
  assign n13851 = n4024 ^ n3120 ^ n3082 ;
  assign n13852 = n13851 ^ n11607 ^ n987 ;
  assign n13850 = n6160 ^ n3479 ^ n585 ;
  assign n13854 = n13853 ^ n13852 ^ n13850 ;
  assign n13855 = ( n349 & ~n3735 ) | ( n349 & n12882 ) | ( ~n3735 & n12882 ) ;
  assign n13856 = n13855 ^ n10890 ^ n10418 ;
  assign n13857 = ( n1605 & ~n1898 ) | ( n1605 & n11304 ) | ( ~n1898 & n11304 ) ;
  assign n13858 = ( n1748 & n11921 ) | ( n1748 & n13857 ) | ( n11921 & n13857 ) ;
  assign n13859 = n6011 ^ n4384 ^ n3078 ;
  assign n13860 = ( n2588 & n2882 ) | ( n2588 & ~n13859 ) | ( n2882 & ~n13859 ) ;
  assign n13861 = ( n3607 & n6862 ) | ( n3607 & n12011 ) | ( n6862 & n12011 ) ;
  assign n13862 = n7338 ^ n3229 ^ n1749 ;
  assign n13863 = n11278 ^ n3076 ^ n394 ;
  assign n13864 = ( ~n2561 & n13862 ) | ( ~n2561 & n13863 ) | ( n13862 & n13863 ) ;
  assign n13865 = ( ~n10369 & n13861 ) | ( ~n10369 & n13864 ) | ( n13861 & n13864 ) ;
  assign n13868 = n12763 ^ n1910 ^ n334 ;
  assign n13867 = ( ~n1056 & n3380 ) | ( ~n1056 & n6222 ) | ( n3380 & n6222 ) ;
  assign n13866 = ( n923 & n1529 ) | ( n923 & ~n7261 ) | ( n1529 & ~n7261 ) ;
  assign n13869 = n13868 ^ n13867 ^ n13866 ;
  assign n13870 = n13869 ^ n12507 ^ n10851 ;
  assign n13871 = ( n3228 & n3957 ) | ( n3228 & ~n6649 ) | ( n3957 & ~n6649 ) ;
  assign n13872 = n13871 ^ n1570 ^ n130 ;
  assign n13873 = ( x112 & n10092 ) | ( x112 & n13872 ) | ( n10092 & n13872 ) ;
  assign n13874 = ( n3559 & n7727 ) | ( n3559 & n10395 ) | ( n7727 & n10395 ) ;
  assign n13875 = ( n4313 & ~n5589 ) | ( n4313 & n10392 ) | ( ~n5589 & n10392 ) ;
  assign n13876 = ( n2505 & n13874 ) | ( n2505 & ~n13875 ) | ( n13874 & ~n13875 ) ;
  assign n13877 = ( ~n13870 & n13873 ) | ( ~n13870 & n13876 ) | ( n13873 & n13876 ) ;
  assign n13878 = n11300 ^ n11166 ^ n10165 ;
  assign n13879 = n7057 ^ n1709 ^ n928 ;
  assign n13881 = ( n615 & n2558 ) | ( n615 & n9117 ) | ( n2558 & n9117 ) ;
  assign n13882 = ( ~n5792 & n10286 ) | ( ~n5792 & n13881 ) | ( n10286 & n13881 ) ;
  assign n13880 = ( n1865 & n4843 ) | ( n1865 & n12516 ) | ( n4843 & n12516 ) ;
  assign n13883 = n13882 ^ n13880 ^ n9976 ;
  assign n13884 = ( n4834 & n6965 ) | ( n4834 & n10375 ) | ( n6965 & n10375 ) ;
  assign n13885 = n13884 ^ n2304 ^ n558 ;
  assign n13886 = ( ~n7240 & n12883 ) | ( ~n7240 & n13885 ) | ( n12883 & n13885 ) ;
  assign n13888 = n3973 ^ n2819 ^ n809 ;
  assign n13887 = n6409 ^ n5004 ^ n4242 ;
  assign n13889 = n13888 ^ n13887 ^ n3993 ;
  assign n13890 = ( ~n10346 & n13886 ) | ( ~n10346 & n13889 ) | ( n13886 & n13889 ) ;
  assign n13891 = n13540 ^ n12309 ^ n4648 ;
  assign n13892 = ( n282 & ~n3502 ) | ( n282 & n13891 ) | ( ~n3502 & n13891 ) ;
  assign n13893 = n766 ^ n391 ^ n356 ;
  assign n13894 = n13893 ^ n9357 ^ n2398 ;
  assign n13895 = n13894 ^ n10732 ^ n9383 ;
  assign n13897 = n3347 ^ n2523 ^ n1706 ;
  assign n13896 = n12397 ^ n6839 ^ n2440 ;
  assign n13898 = n13897 ^ n13896 ^ n3906 ;
  assign n13899 = ( n4289 & n5869 ) | ( n4289 & n13898 ) | ( n5869 & n13898 ) ;
  assign n13904 = ( n1425 & n1735 ) | ( n1425 & n3698 ) | ( n1735 & n3698 ) ;
  assign n13903 = ( n1784 & ~n8474 ) | ( n1784 & n9778 ) | ( ~n8474 & n9778 ) ;
  assign n13900 = ( n182 & n2437 ) | ( n182 & n6357 ) | ( n2437 & n6357 ) ;
  assign n13901 = ( n3135 & n5969 ) | ( n3135 & ~n13900 ) | ( n5969 & ~n13900 ) ;
  assign n13902 = ( n3896 & ~n7265 ) | ( n3896 & n13901 ) | ( ~n7265 & n13901 ) ;
  assign n13905 = n13904 ^ n13903 ^ n13902 ;
  assign n13906 = ( ~n1286 & n2346 ) | ( ~n1286 & n9975 ) | ( n2346 & n9975 ) ;
  assign n13907 = n8842 ^ n7851 ^ n6690 ;
  assign n13910 = n2721 ^ n1333 ^ n1089 ;
  assign n13909 = ( x50 & n2302 ) | ( x50 & ~n9793 ) | ( n2302 & ~n9793 ) ;
  assign n13908 = n11648 ^ n11291 ^ n7952 ;
  assign n13911 = n13910 ^ n13909 ^ n13908 ;
  assign n13918 = ( ~n3755 & n5600 ) | ( ~n3755 & n12184 ) | ( n5600 & n12184 ) ;
  assign n13912 = ( n7833 & n8370 ) | ( n7833 & n10293 ) | ( n8370 & n10293 ) ;
  assign n13913 = ( ~n381 & n1043 ) | ( ~n381 & n2574 ) | ( n1043 & n2574 ) ;
  assign n13914 = n13913 ^ n6303 ^ n4868 ;
  assign n13915 = n5625 ^ n1129 ^ n645 ;
  assign n13916 = ( ~n9690 & n13914 ) | ( ~n9690 & n13915 ) | ( n13914 & n13915 ) ;
  assign n13917 = ( ~n13658 & n13912 ) | ( ~n13658 & n13916 ) | ( n13912 & n13916 ) ;
  assign n13919 = n13918 ^ n13917 ^ n8551 ;
  assign n13920 = ( n1974 & n2997 ) | ( n1974 & n8460 ) | ( n2997 & n8460 ) ;
  assign n13921 = n13920 ^ n11069 ^ n4515 ;
  assign n13922 = n7990 ^ n5384 ^ n1996 ;
  assign n13923 = n13922 ^ n4421 ^ n3956 ;
  assign n13924 = n13923 ^ n11607 ^ n2387 ;
  assign n13925 = n6209 ^ n1290 ^ n251 ;
  assign n13926 = ( n709 & ~n6034 ) | ( n709 & n7912 ) | ( ~n6034 & n7912 ) ;
  assign n13927 = ( ~n3292 & n13571 ) | ( ~n3292 & n13926 ) | ( n13571 & n13926 ) ;
  assign n13928 = ( n8689 & n8880 ) | ( n8689 & n13927 ) | ( n8880 & n13927 ) ;
  assign n13929 = ( ~n1046 & n13925 ) | ( ~n1046 & n13928 ) | ( n13925 & n13928 ) ;
  assign n13930 = n10832 ^ n7874 ^ n4107 ;
  assign n13931 = n12293 ^ n1960 ^ n1344 ;
  assign n13932 = ( n2537 & ~n4504 ) | ( n2537 & n6135 ) | ( ~n4504 & n6135 ) ;
  assign n13933 = n13932 ^ n10913 ^ n7229 ;
  assign n13934 = ( n138 & n13931 ) | ( n138 & ~n13933 ) | ( n13931 & ~n13933 ) ;
  assign n13935 = n13934 ^ n13039 ^ n725 ;
  assign n13936 = ( n11770 & n13930 ) | ( n11770 & ~n13935 ) | ( n13930 & ~n13935 ) ;
  assign n13937 = n6316 ^ n3676 ^ n2780 ;
  assign n13938 = ( ~n312 & n529 ) | ( ~n312 & n5005 ) | ( n529 & n5005 ) ;
  assign n13939 = n13938 ^ n2745 ^ n2436 ;
  assign n13940 = ( ~n478 & n8560 ) | ( ~n478 & n13939 ) | ( n8560 & n13939 ) ;
  assign n13941 = n13940 ^ n970 ^ n718 ;
  assign n13942 = n9924 ^ n3227 ^ n3058 ;
  assign n13943 = ( n10278 & n13941 ) | ( n10278 & n13942 ) | ( n13941 & n13942 ) ;
  assign n13945 = ( n1229 & n5274 ) | ( n1229 & n6294 ) | ( n5274 & n6294 ) ;
  assign n13946 = n13945 ^ n7854 ^ n4101 ;
  assign n13944 = n5804 ^ n5674 ^ n3635 ;
  assign n13947 = n13946 ^ n13944 ^ n12966 ;
  assign n13948 = ( n13937 & n13943 ) | ( n13937 & ~n13947 ) | ( n13943 & ~n13947 ) ;
  assign n13949 = n13948 ^ n9114 ^ n794 ;
  assign n13950 = n4855 ^ n4801 ^ n902 ;
  assign n13951 = ( n942 & n2427 ) | ( n942 & n8747 ) | ( n2427 & n8747 ) ;
  assign n13952 = ( ~n2840 & n3622 ) | ( ~n2840 & n9569 ) | ( n3622 & n9569 ) ;
  assign n13953 = ( n1611 & ~n13951 ) | ( n1611 & n13952 ) | ( ~n13951 & n13952 ) ;
  assign n13954 = n13953 ^ n13250 ^ n187 ;
  assign n13956 = ( n1958 & n5715 ) | ( n1958 & n12133 ) | ( n5715 & n12133 ) ;
  assign n13955 = ( n1045 & ~n1346 ) | ( n1045 & n9362 ) | ( ~n1346 & n9362 ) ;
  assign n13957 = n13956 ^ n13955 ^ n3503 ;
  assign n13958 = n8972 ^ n8216 ^ n3101 ;
  assign n13959 = ( n1663 & n2901 ) | ( n1663 & ~n4932 ) | ( n2901 & ~n4932 ) ;
  assign n13960 = ( ~n2806 & n11664 ) | ( ~n2806 & n13959 ) | ( n11664 & n13959 ) ;
  assign n13961 = n3912 ^ n947 ^ n861 ;
  assign n13962 = ( ~n5869 & n12944 ) | ( ~n5869 & n13961 ) | ( n12944 & n13961 ) ;
  assign n13963 = ( n266 & n13960 ) | ( n266 & n13962 ) | ( n13960 & n13962 ) ;
  assign n13964 = ( n539 & ~n11091 ) | ( n539 & n13455 ) | ( ~n11091 & n13455 ) ;
  assign n13965 = ( x2 & n6454 ) | ( x2 & n11032 ) | ( n6454 & n11032 ) ;
  assign n13966 = ( ~x114 & n9418 ) | ( ~x114 & n13965 ) | ( n9418 & n13965 ) ;
  assign n13967 = ( ~n754 & n6832 ) | ( ~n754 & n13966 ) | ( n6832 & n13966 ) ;
  assign n13968 = n11956 ^ n7221 ^ n3087 ;
  assign n13969 = n12659 ^ n1716 ^ n1592 ;
  assign n13970 = ( x3 & ~n11717 ) | ( x3 & n13969 ) | ( ~n11717 & n13969 ) ;
  assign n13971 = n13390 ^ n9335 ^ n6338 ;
  assign n13972 = ( ~x86 & n786 ) | ( ~x86 & n11577 ) | ( n786 & n11577 ) ;
  assign n13973 = ( x70 & n4901 ) | ( x70 & n13972 ) | ( n4901 & n13972 ) ;
  assign n13974 = ( ~n8075 & n12158 ) | ( ~n8075 & n13973 ) | ( n12158 & n13973 ) ;
  assign n13976 = ( n2641 & ~n3747 ) | ( n2641 & n6818 ) | ( ~n3747 & n6818 ) ;
  assign n13975 = n7247 ^ n3245 ^ n1570 ;
  assign n13977 = n13976 ^ n13975 ^ n11910 ;
  assign n13978 = n13977 ^ n6397 ^ n5197 ;
  assign n13979 = ( ~n6936 & n13974 ) | ( ~n6936 & n13978 ) | ( n13974 & n13978 ) ;
  assign n13980 = ( n7611 & ~n9493 ) | ( n7611 & n13314 ) | ( ~n9493 & n13314 ) ;
  assign n13981 = n13980 ^ n3984 ^ n1898 ;
  assign n13982 = ( ~n511 & n4082 ) | ( ~n511 & n10201 ) | ( n4082 & n10201 ) ;
  assign n13983 = ( ~n382 & n4871 ) | ( ~n382 & n13982 ) | ( n4871 & n13982 ) ;
  assign n13984 = n6642 ^ n5075 ^ n3441 ;
  assign n13985 = ( n8329 & ~n13983 ) | ( n8329 & n13984 ) | ( ~n13983 & n13984 ) ;
  assign n13986 = ( n1714 & n2915 ) | ( n1714 & n3640 ) | ( n2915 & n3640 ) ;
  assign n13987 = ( ~n2853 & n9230 ) | ( ~n2853 & n13986 ) | ( n9230 & n13986 ) ;
  assign n13988 = ( ~n8237 & n13985 ) | ( ~n8237 & n13987 ) | ( n13985 & n13987 ) ;
  assign n13989 = n7479 ^ n5883 ^ n4463 ;
  assign n13990 = ( n698 & ~n4530 ) | ( n698 & n9108 ) | ( ~n4530 & n9108 ) ;
  assign n13991 = ( n5782 & n13989 ) | ( n5782 & n13990 ) | ( n13989 & n13990 ) ;
  assign n13992 = n13991 ^ n6943 ^ n3809 ;
  assign n13993 = ( n264 & n278 ) | ( n264 & n7813 ) | ( n278 & n7813 ) ;
  assign n13994 = n13993 ^ n5262 ^ n4214 ;
  assign n13995 = ( n1563 & ~n3977 ) | ( n1563 & n13994 ) | ( ~n3977 & n13994 ) ;
  assign n13996 = ( n2093 & ~n6917 ) | ( n2093 & n7801 ) | ( ~n6917 & n7801 ) ;
  assign n13997 = ( n4459 & n5376 ) | ( n4459 & ~n13996 ) | ( n5376 & ~n13996 ) ;
  assign n14007 = ( n2070 & n6149 ) | ( n2070 & n7382 ) | ( n6149 & n7382 ) ;
  assign n14004 = ( ~n543 & n4949 ) | ( ~n543 & n9982 ) | ( n4949 & n9982 ) ;
  assign n14005 = n8746 ^ n8008 ^ n566 ;
  assign n14006 = ( ~n9738 & n14004 ) | ( ~n9738 & n14005 ) | ( n14004 & n14005 ) ;
  assign n14002 = ( n6245 & n7953 ) | ( n6245 & n13868 ) | ( n7953 & n13868 ) ;
  assign n13998 = n2656 ^ n2333 ^ n676 ;
  assign n13999 = n13998 ^ n5174 ^ n944 ;
  assign n14000 = n13999 ^ n1961 ^ n1764 ;
  assign n14001 = ( ~n559 & n12919 ) | ( ~n559 & n14000 ) | ( n12919 & n14000 ) ;
  assign n14003 = n14002 ^ n14001 ^ n8567 ;
  assign n14008 = n14007 ^ n14006 ^ n14003 ;
  assign n14009 = ( n10911 & ~n13997 ) | ( n10911 & n14008 ) | ( ~n13997 & n14008 ) ;
  assign n14010 = ( n2438 & n4055 ) | ( n2438 & ~n14009 ) | ( n4055 & ~n14009 ) ;
  assign n14011 = n4731 ^ n3700 ^ n2540 ;
  assign n14012 = ( n660 & n1478 ) | ( n660 & n14011 ) | ( n1478 & n14011 ) ;
  assign n14013 = ( n11552 & n11867 ) | ( n11552 & n14012 ) | ( n11867 & n14012 ) ;
  assign n14014 = n13541 ^ n13212 ^ n4686 ;
  assign n14016 = ( n2649 & ~n4380 ) | ( n2649 & n8857 ) | ( ~n4380 & n8857 ) ;
  assign n14015 = n6245 ^ n5254 ^ n2753 ;
  assign n14017 = n14016 ^ n14015 ^ n11987 ;
  assign n14024 = ( n1298 & ~n2511 ) | ( n1298 & n9112 ) | ( ~n2511 & n9112 ) ;
  assign n14025 = ( ~n4879 & n5189 ) | ( ~n4879 & n14024 ) | ( n5189 & n14024 ) ;
  assign n14026 = ( ~n5391 & n11339 ) | ( ~n5391 & n14025 ) | ( n11339 & n14025 ) ;
  assign n14027 = ( n1663 & n4081 ) | ( n1663 & ~n14026 ) | ( n4081 & ~n14026 ) ;
  assign n14028 = ( n4634 & ~n10383 ) | ( n4634 & n14027 ) | ( ~n10383 & n14027 ) ;
  assign n14022 = ( n1690 & n5730 ) | ( n1690 & ~n6375 ) | ( n5730 & ~n6375 ) ;
  assign n14018 = ( n6245 & n9908 ) | ( n6245 & n12833 ) | ( n9908 & n12833 ) ;
  assign n14019 = n6836 ^ n6253 ^ n2821 ;
  assign n14020 = n14019 ^ n5748 ^ n1957 ;
  assign n14021 = ( n1513 & n14018 ) | ( n1513 & n14020 ) | ( n14018 & n14020 ) ;
  assign n14023 = n14022 ^ n14021 ^ n7011 ;
  assign n14029 = n14028 ^ n14023 ^ n4870 ;
  assign n14030 = n14029 ^ n3645 ^ x102 ;
  assign n14031 = n13016 ^ n10882 ^ n190 ;
  assign n14032 = ( ~n4474 & n8073 ) | ( ~n4474 & n14031 ) | ( n8073 & n14031 ) ;
  assign n14033 = n13634 ^ n8379 ^ n5415 ;
  assign n14034 = n2273 ^ n1862 ^ n1769 ;
  assign n14035 = n4818 ^ n2743 ^ n2537 ;
  assign n14036 = ( n4949 & ~n14034 ) | ( n4949 & n14035 ) | ( ~n14034 & n14035 ) ;
  assign n14037 = ( n5682 & n14033 ) | ( n5682 & ~n14036 ) | ( n14033 & ~n14036 ) ;
  assign n14038 = n14037 ^ n2910 ^ n1827 ;
  assign n14039 = ( n3132 & n13151 ) | ( n3132 & ~n13983 ) | ( n13151 & ~n13983 ) ;
  assign n14040 = ( n6105 & ~n11834 ) | ( n6105 & n14039 ) | ( ~n11834 & n14039 ) ;
  assign n14041 = ( n1923 & n3200 ) | ( n1923 & ~n3956 ) | ( n3200 & ~n3956 ) ;
  assign n14042 = ( n3649 & n10247 ) | ( n3649 & ~n11050 ) | ( n10247 & ~n11050 ) ;
  assign n14043 = ( n1080 & n3299 ) | ( n1080 & ~n7463 ) | ( n3299 & ~n7463 ) ;
  assign n14044 = ( ~n1814 & n11697 ) | ( ~n1814 & n14043 ) | ( n11697 & n14043 ) ;
  assign n14045 = ( n2954 & n9464 ) | ( n2954 & ~n14044 ) | ( n9464 & ~n14044 ) ;
  assign n14046 = ( n14041 & ~n14042 ) | ( n14041 & n14045 ) | ( ~n14042 & n14045 ) ;
  assign n14047 = ( n3274 & n6282 ) | ( n3274 & ~n6594 ) | ( n6282 & ~n6594 ) ;
  assign n14048 = n14047 ^ n11838 ^ n7171 ;
  assign n14054 = ( n1237 & n3991 ) | ( n1237 & n6732 ) | ( n3991 & n6732 ) ;
  assign n14049 = n4377 ^ n2053 ^ n1220 ;
  assign n14050 = n4556 ^ n4238 ^ n1117 ;
  assign n14051 = ( n6524 & ~n10763 ) | ( n6524 & n14050 ) | ( ~n10763 & n14050 ) ;
  assign n14052 = ( n12352 & n14049 ) | ( n12352 & n14051 ) | ( n14049 & n14051 ) ;
  assign n14053 = n14052 ^ n13823 ^ n1698 ;
  assign n14055 = n14054 ^ n14053 ^ n1156 ;
  assign n14056 = n14055 ^ n3359 ^ n2819 ;
  assign n14057 = n5721 ^ n1114 ^ n1087 ;
  assign n14059 = ( n2177 & n3261 ) | ( n2177 & ~n5049 ) | ( n3261 & ~n5049 ) ;
  assign n14058 = n12942 ^ n2575 ^ n1359 ;
  assign n14060 = n14059 ^ n14058 ^ n13270 ;
  assign n14062 = ( n577 & ~n4326 ) | ( n577 & n10886 ) | ( ~n4326 & n10886 ) ;
  assign n14063 = n12477 ^ n6965 ^ n5840 ;
  assign n14064 = ( n9720 & n14062 ) | ( n9720 & ~n14063 ) | ( n14062 & ~n14063 ) ;
  assign n14061 = n6802 ^ n3768 ^ x57 ;
  assign n14065 = n14064 ^ n14061 ^ n11031 ;
  assign n14066 = n11437 ^ n8631 ^ n1204 ;
  assign n14067 = n12087 ^ n2374 ^ n249 ;
  assign n14068 = ( n1949 & ~n3215 ) | ( n1949 & n8171 ) | ( ~n3215 & n8171 ) ;
  assign n14069 = ( n6360 & n10944 ) | ( n6360 & ~n14068 ) | ( n10944 & ~n14068 ) ;
  assign n14070 = ( ~n1700 & n14067 ) | ( ~n1700 & n14069 ) | ( n14067 & n14069 ) ;
  assign n14071 = ( ~n3452 & n14066 ) | ( ~n3452 & n14070 ) | ( n14066 & n14070 ) ;
  assign n14072 = n14071 ^ n8164 ^ n3351 ;
  assign n14075 = n3846 ^ n192 ^ x52 ;
  assign n14073 = ( n4161 & n10491 ) | ( n4161 & n12241 ) | ( n10491 & n12241 ) ;
  assign n14074 = ( n2442 & n7461 ) | ( n2442 & ~n14073 ) | ( n7461 & ~n14073 ) ;
  assign n14076 = n14075 ^ n14074 ^ n7311 ;
  assign n14077 = n7509 ^ n5402 ^ n617 ;
  assign n14078 = ( ~n12062 & n13646 ) | ( ~n12062 & n14077 ) | ( n13646 & n14077 ) ;
  assign n14079 = n12444 ^ n9339 ^ n3187 ;
  assign n14080 = n14079 ^ n13214 ^ n1088 ;
  assign n14081 = ( n4000 & ~n6333 ) | ( n4000 & n8667 ) | ( ~n6333 & n8667 ) ;
  assign n14082 = ( n5946 & ~n10139 ) | ( n5946 & n14081 ) | ( ~n10139 & n14081 ) ;
  assign n14083 = n13165 ^ n12795 ^ n245 ;
  assign n14084 = n4732 ^ n1894 ^ n1437 ;
  assign n14086 = ( ~n2780 & n3723 ) | ( ~n2780 & n6732 ) | ( n3723 & n6732 ) ;
  assign n14087 = ( ~n8155 & n10368 ) | ( ~n8155 & n14086 ) | ( n10368 & n14086 ) ;
  assign n14085 = ( ~n4130 & n5308 ) | ( ~n4130 & n6200 ) | ( n5308 & n6200 ) ;
  assign n14088 = n14087 ^ n14085 ^ n11288 ;
  assign n14089 = n9636 ^ n8320 ^ n1972 ;
  assign n14090 = ( n2784 & ~n6128 ) | ( n2784 & n14089 ) | ( ~n6128 & n14089 ) ;
  assign n14091 = ( n5004 & n5029 ) | ( n5004 & n9599 ) | ( n5029 & n9599 ) ;
  assign n14092 = ( n631 & n7999 ) | ( n631 & n14091 ) | ( n7999 & n14091 ) ;
  assign n14093 = ( n496 & n14090 ) | ( n496 & n14092 ) | ( n14090 & n14092 ) ;
  assign n14094 = n3713 ^ n2831 ^ n2413 ;
  assign n14095 = ( n3760 & n13419 ) | ( n3760 & ~n14094 ) | ( n13419 & ~n14094 ) ;
  assign n14096 = ( n5139 & n11202 ) | ( n5139 & ~n13952 ) | ( n11202 & ~n13952 ) ;
  assign n14097 = ( n3076 & n7031 ) | ( n3076 & ~n14096 ) | ( n7031 & ~n14096 ) ;
  assign n14098 = ( n508 & n8848 ) | ( n508 & ~n14097 ) | ( n8848 & ~n14097 ) ;
  assign n14099 = ( n12919 & ~n14095 ) | ( n12919 & n14098 ) | ( ~n14095 & n14098 ) ;
  assign n14100 = n14099 ^ n1455 ^ n926 ;
  assign n14101 = n9867 ^ n3683 ^ n436 ;
  assign n14102 = n7787 ^ n7250 ^ n1801 ;
  assign n14109 = n9847 ^ n3358 ^ n546 ;
  assign n14110 = ( n4544 & n12750 ) | ( n4544 & ~n14109 ) | ( n12750 & ~n14109 ) ;
  assign n14106 = ( n6338 & ~n7650 ) | ( n6338 & n9370 ) | ( ~n7650 & n9370 ) ;
  assign n14107 = n14106 ^ n7068 ^ n403 ;
  assign n14103 = ( n8258 & n8963 ) | ( n8258 & n9014 ) | ( n8963 & n9014 ) ;
  assign n14104 = n14103 ^ n10695 ^ n359 ;
  assign n14105 = ( n2212 & n8563 ) | ( n2212 & n14104 ) | ( n8563 & n14104 ) ;
  assign n14108 = n14107 ^ n14105 ^ n758 ;
  assign n14111 = n14110 ^ n14108 ^ n1114 ;
  assign n14112 = ( ~n14101 & n14102 ) | ( ~n14101 & n14111 ) | ( n14102 & n14111 ) ;
  assign n14114 = n10359 ^ n9561 ^ n1174 ;
  assign n14113 = n5367 ^ n3768 ^ n3406 ;
  assign n14115 = n14114 ^ n14113 ^ n13811 ;
  assign n14118 = n4443 ^ n2660 ^ n1021 ;
  assign n14119 = n14118 ^ n4193 ^ n1745 ;
  assign n14116 = n9889 ^ n7782 ^ n5244 ;
  assign n14117 = n14116 ^ n8418 ^ n5708 ;
  assign n14120 = n14119 ^ n14117 ^ n14049 ;
  assign n14121 = ( n2356 & n8694 ) | ( n2356 & n11605 ) | ( n8694 & n11605 ) ;
  assign n14122 = ( n4859 & ~n8725 ) | ( n4859 & n14121 ) | ( ~n8725 & n14121 ) ;
  assign n14123 = n14122 ^ n14079 ^ n1663 ;
  assign n14124 = ( ~n1278 & n1733 ) | ( ~n1278 & n3213 ) | ( n1733 & n3213 ) ;
  assign n14125 = ( n251 & n8617 ) | ( n251 & ~n14124 ) | ( n8617 & ~n14124 ) ;
  assign n14128 = n3886 ^ n2214 ^ n1316 ;
  assign n14126 = n4565 ^ n4515 ^ n3124 ;
  assign n14127 = n14126 ^ n2902 ^ n2516 ;
  assign n14129 = n14128 ^ n14127 ^ n3953 ;
  assign n14130 = ( ~n10842 & n11452 ) | ( ~n10842 & n14129 ) | ( n11452 & n14129 ) ;
  assign n14132 = n4371 ^ n3788 ^ n2038 ;
  assign n14131 = ( n3533 & n12181 ) | ( n3533 & n13516 ) | ( n12181 & n13516 ) ;
  assign n14133 = n14132 ^ n14131 ^ n1922 ;
  assign n14134 = ( n1783 & ~n3143 ) | ( n1783 & n14133 ) | ( ~n3143 & n14133 ) ;
  assign n14135 = ( n4081 & n12662 ) | ( n4081 & ~n14134 ) | ( n12662 & ~n14134 ) ;
  assign n14136 = n11369 ^ n3037 ^ n721 ;
  assign n14139 = ( n1261 & ~n2105 ) | ( n1261 & n7177 ) | ( ~n2105 & n7177 ) ;
  assign n14137 = ( n2813 & ~n6567 ) | ( n2813 & n10886 ) | ( ~n6567 & n10886 ) ;
  assign n14138 = n14137 ^ n4847 ^ n1270 ;
  assign n14140 = n14139 ^ n14138 ^ n8274 ;
  assign n14141 = ( n13243 & n14136 ) | ( n13243 & ~n14140 ) | ( n14136 & ~n14140 ) ;
  assign n14142 = ( n2124 & n2211 ) | ( n2124 & ~n4123 ) | ( n2211 & ~n4123 ) ;
  assign n14143 = ( n406 & n2688 ) | ( n406 & ~n14142 ) | ( n2688 & ~n14142 ) ;
  assign n14144 = ( n597 & n12026 ) | ( n597 & n14143 ) | ( n12026 & n14143 ) ;
  assign n14145 = ( n5034 & n14141 ) | ( n5034 & n14144 ) | ( n14141 & n14144 ) ;
  assign n14146 = ( n1021 & n5047 ) | ( n1021 & ~n8055 ) | ( n5047 & ~n8055 ) ;
  assign n14147 = ( n1193 & ~n4040 ) | ( n1193 & n6174 ) | ( ~n4040 & n6174 ) ;
  assign n14148 = n2126 ^ n763 ^ x83 ;
  assign n14149 = ( n1148 & n8310 ) | ( n1148 & ~n9954 ) | ( n8310 & ~n9954 ) ;
  assign n14150 = ( ~n1315 & n8341 ) | ( ~n1315 & n13663 ) | ( n8341 & n13663 ) ;
  assign n14151 = n14150 ^ n6053 ^ n901 ;
  assign n14152 = ( ~n4980 & n5504 ) | ( ~n4980 & n14151 ) | ( n5504 & n14151 ) ;
  assign n14153 = ( ~n7938 & n14149 ) | ( ~n7938 & n14152 ) | ( n14149 & n14152 ) ;
  assign n14154 = ( n8695 & n14148 ) | ( n8695 & n14153 ) | ( n14148 & n14153 ) ;
  assign n14155 = ( ~n14146 & n14147 ) | ( ~n14146 & n14154 ) | ( n14147 & n14154 ) ;
  assign n14156 = n8243 ^ n2458 ^ n2207 ;
  assign n14157 = n14156 ^ n7455 ^ n2539 ;
  assign n14158 = n10659 ^ n10099 ^ n2353 ;
  assign n14161 = ( n6328 & ~n7053 ) | ( n6328 & n9141 ) | ( ~n7053 & n9141 ) ;
  assign n14159 = ( ~n7728 & n10090 ) | ( ~n7728 & n13943 ) | ( n10090 & n13943 ) ;
  assign n14160 = n14159 ^ n3801 ^ n2017 ;
  assign n14162 = n14161 ^ n14160 ^ n1179 ;
  assign n14165 = ( n2370 & ~n3717 ) | ( n2370 & n8883 ) | ( ~n3717 & n8883 ) ;
  assign n14166 = ( n6573 & n10650 ) | ( n6573 & ~n11364 ) | ( n10650 & ~n11364 ) ;
  assign n14167 = ( n5208 & ~n7106 ) | ( n5208 & n14166 ) | ( ~n7106 & n14166 ) ;
  assign n14168 = n13168 ^ n5420 ^ n2781 ;
  assign n14169 = ( n14165 & n14167 ) | ( n14165 & n14168 ) | ( n14167 & n14168 ) ;
  assign n14163 = ( n2574 & n6239 ) | ( n2574 & n10141 ) | ( n6239 & n10141 ) ;
  assign n14164 = n14163 ^ n9854 ^ n2997 ;
  assign n14170 = n14169 ^ n14164 ^ n9133 ;
  assign n14171 = ( n3799 & n4516 ) | ( n3799 & ~n13212 ) | ( n4516 & ~n13212 ) ;
  assign n14172 = ( ~n7005 & n13844 ) | ( ~n7005 & n14171 ) | ( n13844 & n14171 ) ;
  assign n14173 = ( ~n6108 & n6992 ) | ( ~n6108 & n7776 ) | ( n6992 & n7776 ) ;
  assign n14174 = ( n1483 & ~n1582 ) | ( n1483 & n14173 ) | ( ~n1582 & n14173 ) ;
  assign n14175 = n14174 ^ n5150 ^ n4551 ;
  assign n14176 = n14175 ^ n9283 ^ n7885 ;
  assign n14177 = n8356 ^ n5422 ^ n670 ;
  assign n14178 = ( n5468 & n12746 ) | ( n5468 & ~n14177 ) | ( n12746 & ~n14177 ) ;
  assign n14179 = n8324 ^ n6350 ^ n2069 ;
  assign n14180 = ( n1877 & ~n7752 ) | ( n1877 & n9405 ) | ( ~n7752 & n9405 ) ;
  assign n14181 = ( n10649 & n12371 ) | ( n10649 & n14180 ) | ( n12371 & n14180 ) ;
  assign n14182 = ( ~n12797 & n14179 ) | ( ~n12797 & n14181 ) | ( n14179 & n14181 ) ;
  assign n14183 = n7728 ^ n2683 ^ n1464 ;
  assign n14184 = ( n2634 & n7952 ) | ( n2634 & ~n14183 ) | ( n7952 & ~n14183 ) ;
  assign n14185 = n14184 ^ n12883 ^ n2822 ;
  assign n14190 = ( ~n1542 & n2193 ) | ( ~n1542 & n2707 ) | ( n2193 & n2707 ) ;
  assign n14191 = n14190 ^ n6030 ^ n3617 ;
  assign n14188 = ( n1948 & n7498 ) | ( n1948 & ~n11040 ) | ( n7498 & ~n11040 ) ;
  assign n14187 = ( ~n2649 & n5206 ) | ( ~n2649 & n7200 ) | ( n5206 & n7200 ) ;
  assign n14189 = n14188 ^ n14187 ^ n9892 ;
  assign n14186 = ( n1981 & n10194 ) | ( n1981 & ~n10417 ) | ( n10194 & ~n10417 ) ;
  assign n14192 = n14191 ^ n14189 ^ n14186 ;
  assign n14193 = ( n6167 & ~n6534 ) | ( n6167 & n9988 ) | ( ~n6534 & n9988 ) ;
  assign n14194 = ( n8525 & ~n9773 ) | ( n8525 & n11308 ) | ( ~n9773 & n11308 ) ;
  assign n14206 = ( n2621 & n6540 ) | ( n2621 & ~n10882 ) | ( n6540 & ~n10882 ) ;
  assign n14204 = n4365 ^ n4107 ^ x76 ;
  assign n14202 = n12133 ^ n3400 ^ n751 ;
  assign n14199 = ( n3288 & n5310 ) | ( n3288 & ~n7364 ) | ( n5310 & ~n7364 ) ;
  assign n14200 = ( n9430 & n11618 ) | ( n9430 & ~n14199 ) | ( n11618 & ~n14199 ) ;
  assign n14201 = n14200 ^ n5397 ^ n2493 ;
  assign n14203 = n14202 ^ n14201 ^ n3243 ;
  assign n14195 = n12011 ^ n5494 ^ n4026 ;
  assign n14196 = n14195 ^ n10169 ^ n2151 ;
  assign n14197 = n14196 ^ n4901 ^ n4041 ;
  assign n14198 = ( n3976 & ~n6577 ) | ( n3976 & n14197 ) | ( ~n6577 & n14197 ) ;
  assign n14205 = n14204 ^ n14203 ^ n14198 ;
  assign n14207 = n14206 ^ n14205 ^ n9846 ;
  assign n14208 = n13146 ^ n8476 ^ n5106 ;
  assign n14212 = n9735 ^ n2167 ^ x0 ;
  assign n14209 = n8324 ^ n5926 ^ n4811 ;
  assign n14210 = ( n1617 & n2843 ) | ( n1617 & n14209 ) | ( n2843 & n14209 ) ;
  assign n14211 = ( n9849 & ~n13454 ) | ( n9849 & n14210 ) | ( ~n13454 & n14210 ) ;
  assign n14213 = n14212 ^ n14211 ^ n2722 ;
  assign n14218 = n10278 ^ n1550 ^ n952 ;
  assign n14216 = ( ~n209 & n7019 ) | ( ~n209 & n8248 ) | ( n7019 & n8248 ) ;
  assign n14214 = ( n4781 & ~n8344 ) | ( n4781 & n8936 ) | ( ~n8344 & n8936 ) ;
  assign n14215 = ( n6963 & n10470 ) | ( n6963 & n14214 ) | ( n10470 & n14214 ) ;
  assign n14217 = n14216 ^ n14215 ^ n10556 ;
  assign n14219 = n14218 ^ n14217 ^ n2513 ;
  assign n14220 = n13627 ^ n6702 ^ n1966 ;
  assign n14221 = ( n1848 & n7544 ) | ( n1848 & ~n14220 ) | ( n7544 & ~n14220 ) ;
  assign n14222 = ( n939 & ~n2398 ) | ( n939 & n2553 ) | ( ~n2398 & n2553 ) ;
  assign n14223 = n9882 ^ n8557 ^ n8215 ;
  assign n14224 = ( n905 & ~n2358 ) | ( n905 & n8221 ) | ( ~n2358 & n8221 ) ;
  assign n14225 = n14224 ^ n10348 ^ n1623 ;
  assign n14226 = n9034 ^ n4679 ^ n2008 ;
  assign n14227 = ( ~n4298 & n7333 ) | ( ~n4298 & n14226 ) | ( n7333 & n14226 ) ;
  assign n14228 = n14227 ^ n13654 ^ n5511 ;
  assign n14229 = n1492 ^ x30 ^ x1 ;
  assign n14230 = n11114 ^ n5870 ^ n1033 ;
  assign n14231 = n14230 ^ n10255 ^ n6622 ;
  assign n14232 = n11003 ^ n4023 ^ n1291 ;
  assign n14233 = ( ~n3695 & n10976 ) | ( ~n3695 & n14232 ) | ( n10976 & n14232 ) ;
  assign n14235 = ( ~n6747 & n6881 ) | ( ~n6747 & n9149 ) | ( n6881 & n9149 ) ;
  assign n14234 = ( n236 & ~n7865 ) | ( n236 & n8880 ) | ( ~n7865 & n8880 ) ;
  assign n14236 = n14235 ^ n14234 ^ n278 ;
  assign n14237 = n3133 ^ n2236 ^ n170 ;
  assign n14238 = n14237 ^ n5137 ^ n1123 ;
  assign n14239 = ( n6125 & n11247 ) | ( n6125 & n12824 ) | ( n11247 & n12824 ) ;
  assign n14240 = ( n10000 & n12692 ) | ( n10000 & n14239 ) | ( n12692 & n14239 ) ;
  assign n14241 = n14240 ^ n8795 ^ n2311 ;
  assign n14242 = n10047 ^ n3071 ^ n2166 ;
  assign n14243 = n14242 ^ n12482 ^ n6738 ;
  assign n14244 = ( n5947 & n11990 ) | ( n5947 & ~n14243 ) | ( n11990 & ~n14243 ) ;
  assign n14245 = n14244 ^ n13293 ^ n10238 ;
  assign n14246 = n5002 ^ n1185 ^ n340 ;
  assign n14247 = n14246 ^ n8759 ^ n7668 ;
  assign n14248 = ( n3504 & n5621 ) | ( n3504 & n11250 ) | ( n5621 & n11250 ) ;
  assign n14249 = ( n837 & ~n5399 ) | ( n837 & n14248 ) | ( ~n5399 & n14248 ) ;
  assign n14250 = ( n1237 & ~n5435 ) | ( n1237 & n9384 ) | ( ~n5435 & n9384 ) ;
  assign n14251 = n14250 ^ n5923 ^ n3024 ;
  assign n14252 = n11535 ^ n6302 ^ n1897 ;
  assign n14253 = ( n10848 & n14251 ) | ( n10848 & ~n14252 ) | ( n14251 & ~n14252 ) ;
  assign n14255 = ( n313 & n2723 ) | ( n313 & n9026 ) | ( n2723 & n9026 ) ;
  assign n14254 = n12943 ^ n2984 ^ n2858 ;
  assign n14256 = n14255 ^ n14254 ^ n9565 ;
  assign n14257 = ( n7597 & n8108 ) | ( n7597 & n10429 ) | ( n8108 & n10429 ) ;
  assign n14258 = n14257 ^ n9336 ^ n3243 ;
  assign n14259 = n9467 ^ n5922 ^ n1535 ;
  assign n14260 = n11432 ^ n9424 ^ n5753 ;
  assign n14261 = ( n3035 & ~n6110 ) | ( n3035 & n11424 ) | ( ~n6110 & n11424 ) ;
  assign n14268 = n13021 ^ n6121 ^ n4382 ;
  assign n14269 = n14268 ^ n8270 ^ n4369 ;
  assign n14266 = n6852 ^ n6120 ^ n475 ;
  assign n14264 = ( n218 & n392 ) | ( n218 & ~n1244 ) | ( n392 & ~n1244 ) ;
  assign n14263 = ( x34 & n729 ) | ( x34 & n1385 ) | ( n729 & n1385 ) ;
  assign n14262 = n10531 ^ n6680 ^ n6095 ;
  assign n14265 = n14264 ^ n14263 ^ n14262 ;
  assign n14267 = n14266 ^ n14265 ^ n9192 ;
  assign n14270 = n14269 ^ n14267 ^ n3048 ;
  assign n14271 = n11858 ^ n10984 ^ n3808 ;
  assign n14272 = n14271 ^ n10827 ^ n2046 ;
  assign n14273 = n11847 ^ n3457 ^ n293 ;
  assign n14274 = ( n4456 & n6607 ) | ( n4456 & ~n14273 ) | ( n6607 & ~n14273 ) ;
  assign n14275 = ( ~n8543 & n11527 ) | ( ~n8543 & n14274 ) | ( n11527 & n14274 ) ;
  assign n14276 = ( n1008 & ~n4666 ) | ( n1008 & n5980 ) | ( ~n4666 & n5980 ) ;
  assign n14277 = ( n1400 & ~n2498 ) | ( n1400 & n14276 ) | ( ~n2498 & n14276 ) ;
  assign n14278 = ( n2745 & ~n3736 ) | ( n2745 & n7033 ) | ( ~n3736 & n7033 ) ;
  assign n14279 = ( n13074 & n14277 ) | ( n13074 & n14278 ) | ( n14277 & n14278 ) ;
  assign n14280 = ( n1477 & n12012 ) | ( n1477 & ~n14279 ) | ( n12012 & ~n14279 ) ;
  assign n14281 = n14280 ^ n5682 ^ n1822 ;
  assign n14284 = ( n607 & n5160 ) | ( n607 & n5214 ) | ( n5160 & n5214 ) ;
  assign n14285 = ( n3464 & n3942 ) | ( n3464 & n14284 ) | ( n3942 & n14284 ) ;
  assign n14286 = ( n3212 & n4444 ) | ( n3212 & n14285 ) | ( n4444 & n14285 ) ;
  assign n14282 = n1778 ^ n1301 ^ n463 ;
  assign n14283 = ( ~n1263 & n9774 ) | ( ~n1263 & n14282 ) | ( n9774 & n14282 ) ;
  assign n14287 = n14286 ^ n14283 ^ n3922 ;
  assign n14288 = ( n2581 & ~n2876 ) | ( n2581 & n10138 ) | ( ~n2876 & n10138 ) ;
  assign n14289 = ( ~n8298 & n8404 ) | ( ~n8298 & n14288 ) | ( n8404 & n14288 ) ;
  assign n14290 = n14289 ^ n7283 ^ n2617 ;
  assign n14291 = n14290 ^ n11525 ^ n6632 ;
  assign n14292 = ( ~n4426 & n4653 ) | ( ~n4426 & n7452 ) | ( n4653 & n7452 ) ;
  assign n14293 = n5384 ^ n3338 ^ n2814 ;
  assign n14294 = n14293 ^ n8868 ^ n6085 ;
  assign n14295 = ( n2920 & n14292 ) | ( n2920 & n14294 ) | ( n14292 & n14294 ) ;
  assign n14297 = ( ~n2808 & n4771 ) | ( ~n2808 & n5709 ) | ( n4771 & n5709 ) ;
  assign n14298 = n14297 ^ n12275 ^ n1696 ;
  assign n14296 = ( n2476 & ~n2985 ) | ( n2476 & n4012 ) | ( ~n2985 & n4012 ) ;
  assign n14299 = n14298 ^ n14296 ^ n6625 ;
  assign n14300 = n5159 ^ n4114 ^ n1898 ;
  assign n14301 = ( n8682 & ~n13881 ) | ( n8682 & n14300 ) | ( ~n13881 & n14300 ) ;
  assign n14302 = ( n247 & ~n10662 ) | ( n247 & n14301 ) | ( ~n10662 & n14301 ) ;
  assign n14303 = ( n4321 & n9793 ) | ( n4321 & ~n9987 ) | ( n9793 & ~n9987 ) ;
  assign n14308 = ( n1134 & ~n6979 ) | ( n1134 & n8747 ) | ( ~n6979 & n8747 ) ;
  assign n14304 = ( n735 & n4674 ) | ( n735 & n6048 ) | ( n4674 & n6048 ) ;
  assign n14305 = ( n686 & ~n3107 ) | ( n686 & n14304 ) | ( ~n3107 & n14304 ) ;
  assign n14306 = ( n525 & n5774 ) | ( n525 & n14305 ) | ( n5774 & n14305 ) ;
  assign n14307 = n14306 ^ n10927 ^ n2859 ;
  assign n14309 = n14308 ^ n14307 ^ n560 ;
  assign n14313 = ( n4565 & ~n5605 ) | ( n4565 & n7663 ) | ( ~n5605 & n7663 ) ;
  assign n14311 = n7143 ^ n5278 ^ n2731 ;
  assign n14312 = ( n1312 & ~n10286 ) | ( n1312 & n14311 ) | ( ~n10286 & n14311 ) ;
  assign n14310 = ( n6857 & ~n10126 ) | ( n6857 & n13913 ) | ( ~n10126 & n13913 ) ;
  assign n14314 = n14313 ^ n14312 ^ n14310 ;
  assign n14315 = ( n612 & ~n2907 ) | ( n612 & n14314 ) | ( ~n2907 & n14314 ) ;
  assign n14316 = n14045 ^ n8830 ^ n2693 ;
  assign n14317 = n10723 ^ n1119 ^ n419 ;
  assign n14318 = ( ~n4859 & n5799 ) | ( ~n4859 & n7024 ) | ( n5799 & n7024 ) ;
  assign n14319 = ( x64 & ~n4629 ) | ( x64 & n14126 ) | ( ~n4629 & n14126 ) ;
  assign n14320 = ( ~n6927 & n10337 ) | ( ~n6927 & n14319 ) | ( n10337 & n14319 ) ;
  assign n14321 = n14320 ^ n10550 ^ n7990 ;
  assign n14338 = n3953 ^ n3217 ^ n959 ;
  assign n14336 = ( n3100 & ~n3695 ) | ( n3100 & n10200 ) | ( ~n3695 & n10200 ) ;
  assign n14337 = ( n2767 & n7562 ) | ( n2767 & n14336 ) | ( n7562 & n14336 ) ;
  assign n14339 = n14338 ^ n14337 ^ n5645 ;
  assign n14340 = ( n4288 & n5747 ) | ( n4288 & n14339 ) | ( n5747 & n14339 ) ;
  assign n14334 = n12523 ^ n4375 ^ n3460 ;
  assign n14332 = n5858 ^ n5546 ^ n521 ;
  assign n14328 = n9756 ^ n4885 ^ n674 ;
  assign n14329 = ( n1262 & n1763 ) | ( n1262 & ~n9344 ) | ( n1763 & ~n9344 ) ;
  assign n14330 = n6690 ^ n4369 ^ n920 ;
  assign n14331 = ( n14328 & n14329 ) | ( n14328 & ~n14330 ) | ( n14329 & ~n14330 ) ;
  assign n14333 = n14332 ^ n14331 ^ n9991 ;
  assign n14335 = n14334 ^ n14333 ^ n10044 ;
  assign n14322 = ( n2762 & ~n3888 ) | ( n2762 & n9556 ) | ( ~n3888 & n9556 ) ;
  assign n14323 = n8520 ^ n4028 ^ n1427 ;
  assign n14324 = ( n8177 & n10515 ) | ( n8177 & n14323 ) | ( n10515 & n14323 ) ;
  assign n14325 = ( ~n2456 & n6032 ) | ( ~n2456 & n11069 ) | ( n6032 & n11069 ) ;
  assign n14326 = ( ~n4421 & n14324 ) | ( ~n4421 & n14325 ) | ( n14324 & n14325 ) ;
  assign n14327 = ( n5173 & n14322 ) | ( n5173 & ~n14326 ) | ( n14322 & ~n14326 ) ;
  assign n14341 = n14340 ^ n14335 ^ n14327 ;
  assign n14342 = n10498 ^ n5247 ^ n5030 ;
  assign n14343 = n4432 ^ n4134 ^ n1243 ;
  assign n14344 = ( n4087 & n11838 ) | ( n4087 & ~n14343 ) | ( n11838 & ~n14343 ) ;
  assign n14345 = ( ~n7498 & n7709 ) | ( ~n7498 & n14344 ) | ( n7709 & n14344 ) ;
  assign n14346 = n8565 ^ n7300 ^ n2514 ;
  assign n14347 = n7165 ^ n6498 ^ n2247 ;
  assign n14348 = n10954 ^ n688 ^ n621 ;
  assign n14350 = n10182 ^ n5215 ^ n1689 ;
  assign n14349 = n12665 ^ n5077 ^ x48 ;
  assign n14351 = n14350 ^ n14349 ^ n4659 ;
  assign n14352 = ( ~n5434 & n13081 ) | ( ~n5434 & n14351 ) | ( n13081 & n14351 ) ;
  assign n14353 = n7618 ^ n6889 ^ n4539 ;
  assign n14354 = ( n7975 & n12507 ) | ( n7975 & n14353 ) | ( n12507 & n14353 ) ;
  assign n14355 = ( n6048 & ~n14066 ) | ( n6048 & n14354 ) | ( ~n14066 & n14354 ) ;
  assign n14356 = ( n3044 & n6757 ) | ( n3044 & n10338 ) | ( n6757 & n10338 ) ;
  assign n14357 = n3042 ^ n852 ^ n653 ;
  assign n14358 = n14357 ^ n2952 ^ n318 ;
  assign n14359 = n6288 ^ n2624 ^ n202 ;
  assign n14360 = ( n2450 & n14358 ) | ( n2450 & ~n14359 ) | ( n14358 & ~n14359 ) ;
  assign n14361 = ( n3579 & n14356 ) | ( n3579 & ~n14360 ) | ( n14356 & ~n14360 ) ;
  assign n14369 = ( n5412 & ~n9658 ) | ( n5412 & n9908 ) | ( ~n9658 & n9908 ) ;
  assign n14367 = n7463 ^ n6188 ^ n3865 ;
  assign n14368 = ( n1317 & n9212 ) | ( n1317 & n14367 ) | ( n9212 & n14367 ) ;
  assign n14365 = ( n2144 & n9666 ) | ( n2144 & ~n11840 ) | ( n9666 & ~n11840 ) ;
  assign n14366 = ( n4692 & ~n5957 ) | ( n4692 & n14365 ) | ( ~n5957 & n14365 ) ;
  assign n14370 = n14369 ^ n14368 ^ n14366 ;
  assign n14362 = n10518 ^ n1669 ^ n269 ;
  assign n14363 = ( n4703 & ~n10095 ) | ( n4703 & n14362 ) | ( ~n10095 & n14362 ) ;
  assign n14364 = ( n904 & n5610 ) | ( n904 & ~n14363 ) | ( n5610 & ~n14363 ) ;
  assign n14371 = n14370 ^ n14364 ^ n11793 ;
  assign n14372 = n14371 ^ n10429 ^ n5178 ;
  assign n14373 = ( n3962 & ~n8780 ) | ( n3962 & n11293 ) | ( ~n8780 & n11293 ) ;
  assign n14374 = n14373 ^ n3421 ^ n3327 ;
  assign n14375 = ( n7422 & ~n13561 ) | ( n7422 & n14374 ) | ( ~n13561 & n14374 ) ;
  assign n14376 = n2933 ^ n1221 ^ n1013 ;
  assign n14378 = ( n585 & ~n1014 ) | ( n585 & n5968 ) | ( ~n1014 & n5968 ) ;
  assign n14379 = n14378 ^ n3600 ^ n3185 ;
  assign n14380 = ( n1319 & n7172 ) | ( n1319 & ~n14379 ) | ( n7172 & ~n14379 ) ;
  assign n14381 = n14380 ^ n6703 ^ n244 ;
  assign n14382 = n14381 ^ n13418 ^ n527 ;
  assign n14377 = ( n3692 & ~n9510 ) | ( n3692 & n9704 ) | ( ~n9510 & n9704 ) ;
  assign n14383 = n14382 ^ n14377 ^ x108 ;
  assign n14384 = n11661 ^ n6441 ^ n584 ;
  assign n14385 = ( n4540 & ~n9469 ) | ( n4540 & n14384 ) | ( ~n9469 & n14384 ) ;
  assign n14386 = n5057 ^ n3198 ^ n3048 ;
  assign n14387 = n9962 ^ n6805 ^ n1910 ;
  assign n14388 = ( ~n14114 & n14386 ) | ( ~n14114 & n14387 ) | ( n14386 & n14387 ) ;
  assign n14390 = ( ~n651 & n993 ) | ( ~n651 & n3107 ) | ( n993 & n3107 ) ;
  assign n14391 = n14390 ^ n6525 ^ n2722 ;
  assign n14392 = n14391 ^ n6855 ^ n2117 ;
  assign n14389 = n12660 ^ n6189 ^ n508 ;
  assign n14393 = n14392 ^ n14389 ^ n1011 ;
  assign n14394 = ( n941 & n12316 ) | ( n941 & ~n13012 ) | ( n12316 & ~n13012 ) ;
  assign n14395 = ( n3113 & n5937 ) | ( n3113 & ~n14133 ) | ( n5937 & ~n14133 ) ;
  assign n14399 = ( n5278 & ~n6802 ) | ( n5278 & n9449 ) | ( ~n6802 & n9449 ) ;
  assign n14400 = ( x77 & ~n1060 ) | ( x77 & n8290 ) | ( ~n1060 & n8290 ) ;
  assign n14401 = ( n5530 & n14399 ) | ( n5530 & ~n14400 ) | ( n14399 & ~n14400 ) ;
  assign n14396 = ( n2759 & n5383 ) | ( n2759 & n8807 ) | ( n5383 & n8807 ) ;
  assign n14397 = n14396 ^ n14206 ^ n5149 ;
  assign n14398 = ( ~n9476 & n11773 ) | ( ~n9476 & n14397 ) | ( n11773 & n14397 ) ;
  assign n14402 = n14401 ^ n14398 ^ n4868 ;
  assign n14403 = n9345 ^ n3242 ^ n284 ;
  assign n14405 = n8836 ^ n3241 ^ n729 ;
  assign n14404 = ( ~n560 & n998 ) | ( ~n560 & n8306 ) | ( n998 & n8306 ) ;
  assign n14406 = n14405 ^ n14404 ^ n657 ;
  assign n14407 = n9665 ^ n8603 ^ n336 ;
  assign n14408 = n14407 ^ n13119 ^ n3132 ;
  assign n14409 = ( n5437 & n14116 ) | ( n5437 & ~n14408 ) | ( n14116 & ~n14408 ) ;
  assign n14410 = ( n1789 & n11156 ) | ( n1789 & n13787 ) | ( n11156 & n13787 ) ;
  assign n14414 = n13587 ^ n5799 ^ n621 ;
  assign n14411 = ( n1445 & ~n4816 ) | ( n1445 & n12642 ) | ( ~n4816 & n12642 ) ;
  assign n14412 = ( n5646 & n5842 ) | ( n5646 & n14411 ) | ( n5842 & n14411 ) ;
  assign n14413 = ( ~n173 & n10977 ) | ( ~n173 & n14412 ) | ( n10977 & n14412 ) ;
  assign n14415 = n14414 ^ n14413 ^ n10845 ;
  assign n14416 = n12426 ^ n2289 ^ n737 ;
  assign n14417 = n14416 ^ n7838 ^ n1995 ;
  assign n14418 = ( ~n8432 & n8747 ) | ( ~n8432 & n11525 ) | ( n8747 & n11525 ) ;
  assign n14419 = n5785 ^ n1100 ^ n860 ;
  assign n14420 = n14419 ^ n6107 ^ n3509 ;
  assign n14421 = ( n1075 & n13505 ) | ( n1075 & n14420 ) | ( n13505 & n14420 ) ;
  assign n14422 = ( n5143 & n5356 ) | ( n5143 & ~n10545 ) | ( n5356 & ~n10545 ) ;
  assign n14423 = n14422 ^ n9829 ^ n1842 ;
  assign n14424 = n14423 ^ n10265 ^ n5219 ;
  assign n14425 = ( ~n1383 & n13000 ) | ( ~n1383 & n13466 ) | ( n13000 & n13466 ) ;
  assign n14426 = ( n13896 & n14424 ) | ( n13896 & n14425 ) | ( n14424 & n14425 ) ;
  assign n14427 = ( n8987 & n13811 ) | ( n8987 & n14426 ) | ( n13811 & n14426 ) ;
  assign n14428 = n7396 ^ n6697 ^ n1214 ;
  assign n14429 = n3837 ^ n2792 ^ n274 ;
  assign n14430 = ( n4564 & n8860 ) | ( n4564 & n14429 ) | ( n8860 & n14429 ) ;
  assign n14432 = ( n1609 & n2532 ) | ( n1609 & n5106 ) | ( n2532 & n5106 ) ;
  assign n14433 = n14432 ^ n7308 ^ x45 ;
  assign n14431 = n5946 ^ n4227 ^ n1466 ;
  assign n14434 = n14433 ^ n14431 ^ n2555 ;
  assign n14435 = n13976 ^ n12963 ^ n9889 ;
  assign n14436 = ( ~n1276 & n2463 ) | ( ~n1276 & n6820 ) | ( n2463 & n6820 ) ;
  assign n14437 = ( n3321 & ~n10196 ) | ( n3321 & n14436 ) | ( ~n10196 & n14436 ) ;
  assign n14438 = ( n9000 & n9490 ) | ( n9000 & n14437 ) | ( n9490 & n14437 ) ;
  assign n14439 = ( n693 & ~n3230 ) | ( n693 & n14438 ) | ( ~n3230 & n14438 ) ;
  assign n14440 = ( n5480 & ~n11282 ) | ( n5480 & n14439 ) | ( ~n11282 & n14439 ) ;
  assign n14441 = n11099 ^ n8329 ^ n167 ;
  assign n14442 = ( n14435 & ~n14440 ) | ( n14435 & n14441 ) | ( ~n14440 & n14441 ) ;
  assign n14443 = n9040 ^ n8898 ^ n5004 ;
  assign n14444 = ( n5795 & n12588 ) | ( n5795 & ~n14443 ) | ( n12588 & ~n14443 ) ;
  assign n14445 = n5283 ^ n4679 ^ n324 ;
  assign n14446 = n14445 ^ n10405 ^ n672 ;
  assign n14447 = ( ~n5387 & n12000 ) | ( ~n5387 & n14446 ) | ( n12000 & n14446 ) ;
  assign n14448 = n8572 ^ n3237 ^ x127 ;
  assign n14449 = ( n6826 & n7669 ) | ( n6826 & n14448 ) | ( n7669 & n14448 ) ;
  assign n14450 = ( n352 & n5556 ) | ( n352 & n14449 ) | ( n5556 & n14449 ) ;
  assign n14451 = n4711 ^ n3544 ^ n295 ;
  assign n14452 = ( n7416 & ~n8097 ) | ( n7416 & n13322 ) | ( ~n8097 & n13322 ) ;
  assign n14453 = ( n887 & n14451 ) | ( n887 & n14452 ) | ( n14451 & n14452 ) ;
  assign n14454 = n8951 ^ n4517 ^ n1368 ;
  assign n14455 = ( n5456 & ~n8597 ) | ( n5456 & n10241 ) | ( ~n8597 & n10241 ) ;
  assign n14456 = n14455 ^ n12261 ^ n3708 ;
  assign n14457 = ( n13655 & n14454 ) | ( n13655 & ~n14456 ) | ( n14454 & ~n14456 ) ;
  assign n14458 = n5897 ^ n3374 ^ n1434 ;
  assign n14459 = ( n4998 & n9986 ) | ( n4998 & n11602 ) | ( n9986 & n11602 ) ;
  assign n14460 = ( ~n2470 & n8555 ) | ( ~n2470 & n14459 ) | ( n8555 & n14459 ) ;
  assign n14461 = n14460 ^ n13370 ^ n8347 ;
  assign n14462 = n12046 ^ n8360 ^ n1066 ;
  assign n14463 = ( n733 & n1675 ) | ( n733 & ~n4622 ) | ( n1675 & ~n4622 ) ;
  assign n14464 = n14463 ^ n12516 ^ n5942 ;
  assign n14465 = ( n957 & ~n11251 ) | ( n957 & n14464 ) | ( ~n11251 & n14464 ) ;
  assign n14466 = ( n2177 & n3454 ) | ( n2177 & n11908 ) | ( n3454 & n11908 ) ;
  assign n14467 = n6555 ^ n4681 ^ n3309 ;
  assign n14468 = ( n6040 & ~n10157 ) | ( n6040 & n14467 ) | ( ~n10157 & n14467 ) ;
  assign n14469 = ( n1346 & n4473 ) | ( n1346 & ~n12756 ) | ( n4473 & ~n12756 ) ;
  assign n14470 = ( n3118 & n13261 ) | ( n3118 & ~n14469 ) | ( n13261 & ~n14469 ) ;
  assign n14472 = ( ~n858 & n3936 ) | ( ~n858 & n11057 ) | ( n3936 & n11057 ) ;
  assign n14471 = ( ~n1018 & n1289 ) | ( ~n1018 & n4126 ) | ( n1289 & n4126 ) ;
  assign n14473 = n14472 ^ n14471 ^ n319 ;
  assign n14476 = n7076 ^ n5915 ^ n3448 ;
  assign n14474 = ( n832 & n5205 ) | ( n832 & n11623 ) | ( n5205 & n11623 ) ;
  assign n14475 = ( ~n5566 & n7323 ) | ( ~n5566 & n14474 ) | ( n7323 & n14474 ) ;
  assign n14477 = n14476 ^ n14475 ^ n5671 ;
  assign n14478 = n14477 ^ n12026 ^ n5493 ;
  assign n14479 = n14478 ^ n5920 ^ n1520 ;
  assign n14480 = ( n7241 & n7304 ) | ( n7241 & ~n7989 ) | ( n7304 & ~n7989 ) ;
  assign n14481 = ( n5247 & ~n6874 ) | ( n5247 & n14480 ) | ( ~n6874 & n14480 ) ;
  assign n14482 = ( ~n2978 & n6049 ) | ( ~n2978 & n6615 ) | ( n6049 & n6615 ) ;
  assign n14483 = n14482 ^ n13094 ^ n3270 ;
  assign n14484 = ( ~n585 & n1114 ) | ( ~n585 & n2036 ) | ( n1114 & n2036 ) ;
  assign n14485 = ( n2961 & n11351 ) | ( n2961 & ~n14484 ) | ( n11351 & ~n14484 ) ;
  assign n14486 = ( n3087 & n3483 ) | ( n3087 & ~n14485 ) | ( n3483 & ~n14485 ) ;
  assign n14487 = n4870 ^ n954 ^ n714 ;
  assign n14488 = ( n2163 & n7761 ) | ( n2163 & ~n14487 ) | ( n7761 & ~n14487 ) ;
  assign n14489 = ( n4839 & n9085 ) | ( n4839 & n14488 ) | ( n9085 & n14488 ) ;
  assign n14490 = n14489 ^ n10224 ^ n7086 ;
  assign n14491 = n13822 ^ n4266 ^ n961 ;
  assign n14492 = n14387 ^ n5945 ^ n2569 ;
  assign n14493 = ( n11409 & ~n14491 ) | ( n11409 & n14492 ) | ( ~n14491 & n14492 ) ;
  assign n14494 = n9008 ^ n8632 ^ n695 ;
  assign n14495 = ( n1047 & n1573 ) | ( n1047 & n14494 ) | ( n1573 & n14494 ) ;
  assign n14496 = ( ~n1015 & n5117 ) | ( ~n1015 & n14495 ) | ( n5117 & n14495 ) ;
  assign n14497 = ( n7024 & n9522 ) | ( n7024 & n14496 ) | ( n9522 & n14496 ) ;
  assign n14498 = n8191 ^ n5297 ^ n1147 ;
  assign n14499 = n14498 ^ n6410 ^ n4440 ;
  assign n14500 = n14499 ^ n10779 ^ n9332 ;
  assign n14508 = n8414 ^ n3061 ^ n1303 ;
  assign n14509 = n14508 ^ n4184 ^ n2791 ;
  assign n14504 = n4621 ^ n816 ^ n705 ;
  assign n14505 = n5122 ^ n1362 ^ n316 ;
  assign n14506 = ( ~n3000 & n7666 ) | ( ~n3000 & n14505 ) | ( n7666 & n14505 ) ;
  assign n14507 = ( n12661 & n14504 ) | ( n12661 & ~n14506 ) | ( n14504 & ~n14506 ) ;
  assign n14510 = n14509 ^ n14507 ^ n6542 ;
  assign n14501 = n5603 ^ n2277 ^ n540 ;
  assign n14502 = ( ~n3449 & n4670 ) | ( ~n3449 & n14323 ) | ( n4670 & n14323 ) ;
  assign n14503 = ( n12342 & ~n14501 ) | ( n12342 & n14502 ) | ( ~n14501 & n14502 ) ;
  assign n14511 = n14510 ^ n14503 ^ n2033 ;
  assign n14512 = n14511 ^ n4486 ^ n4100 ;
  assign n14513 = n3850 ^ n3208 ^ n1733 ;
  assign n14514 = n14513 ^ n9074 ^ n2855 ;
  assign n14515 = n14514 ^ n13468 ^ n7254 ;
  assign n14520 = ( ~n2893 & n7999 ) | ( ~n2893 & n9726 ) | ( n7999 & n9726 ) ;
  assign n14519 = n12860 ^ n8636 ^ n1237 ;
  assign n14516 = ( ~n792 & n3814 ) | ( ~n792 & n4055 ) | ( n3814 & n4055 ) ;
  assign n14517 = n14516 ^ n4977 ^ n2177 ;
  assign n14518 = ( ~n925 & n3245 ) | ( ~n925 & n14517 ) | ( n3245 & n14517 ) ;
  assign n14521 = n14520 ^ n14519 ^ n14518 ;
  assign n14522 = n11914 ^ n2514 ^ n1680 ;
  assign n14523 = ( ~n2088 & n2575 ) | ( ~n2088 & n14522 ) | ( n2575 & n14522 ) ;
  assign n14524 = ( ~n9524 & n14220 ) | ( ~n9524 & n14523 ) | ( n14220 & n14523 ) ;
  assign n14525 = ( n1372 & ~n11853 ) | ( n1372 & n14524 ) | ( ~n11853 & n14524 ) ;
  assign n14527 = ( n2761 & n7165 ) | ( n2761 & ~n9402 ) | ( n7165 & ~n9402 ) ;
  assign n14528 = ( n6245 & n6635 ) | ( n6245 & n14527 ) | ( n6635 & n14527 ) ;
  assign n14529 = n3828 ^ n2839 ^ n1423 ;
  assign n14530 = ( n6482 & n14528 ) | ( n6482 & n14529 ) | ( n14528 & n14529 ) ;
  assign n14526 = ( n3661 & ~n4503 ) | ( n3661 & n12978 ) | ( ~n4503 & n12978 ) ;
  assign n14531 = n14530 ^ n14526 ^ n1552 ;
  assign n14532 = ( n3289 & ~n5415 ) | ( n3289 & n9391 ) | ( ~n5415 & n9391 ) ;
  assign n14533 = n14532 ^ n13087 ^ n3499 ;
  assign n14534 = n1822 ^ n317 ^ x5 ;
  assign n14535 = n8650 ^ n4783 ^ n326 ;
  assign n14536 = n14535 ^ n12490 ^ n7425 ;
  assign n14537 = n14536 ^ n3199 ^ n1028 ;
  assign n14538 = ( n1490 & ~n4699 ) | ( n1490 & n14537 ) | ( ~n4699 & n14537 ) ;
  assign n14539 = n14538 ^ n3286 ^ n1835 ;
  assign n14540 = ( n6892 & ~n14534 ) | ( n6892 & n14539 ) | ( ~n14534 & n14539 ) ;
  assign n14541 = n8977 ^ n4514 ^ n979 ;
  assign n14542 = ( n2977 & n3738 ) | ( n2977 & ~n8500 ) | ( n3738 & ~n8500 ) ;
  assign n14543 = n11990 ^ n6188 ^ n2864 ;
  assign n14544 = ( ~n3948 & n14542 ) | ( ~n3948 & n14543 ) | ( n14542 & n14543 ) ;
  assign n14545 = ( ~n437 & n14541 ) | ( ~n437 & n14544 ) | ( n14541 & n14544 ) ;
  assign n14546 = ( ~n8590 & n9364 ) | ( ~n8590 & n14545 ) | ( n9364 & n14545 ) ;
  assign n14547 = ( n187 & n2731 ) | ( n187 & ~n7953 ) | ( n2731 & ~n7953 ) ;
  assign n14548 = ( n1425 & n10553 ) | ( n1425 & ~n11320 ) | ( n10553 & ~n11320 ) ;
  assign n14549 = n14548 ^ n11610 ^ n9102 ;
  assign n14550 = ( n2276 & n14042 ) | ( n2276 & n14549 ) | ( n14042 & n14549 ) ;
  assign n14551 = ( n1957 & ~n14547 ) | ( n1957 & n14550 ) | ( ~n14547 & n14550 ) ;
  assign n14552 = n8778 ^ n3605 ^ n201 ;
  assign n14553 = ( n3156 & n3368 ) | ( n3156 & n4378 ) | ( n3368 & n4378 ) ;
  assign n14554 = ( n867 & n8090 ) | ( n867 & n14313 ) | ( n8090 & n14313 ) ;
  assign n14555 = ( n6604 & n14553 ) | ( n6604 & ~n14554 ) | ( n14553 & ~n14554 ) ;
  assign n14556 = n14555 ^ n12450 ^ n7257 ;
  assign n14557 = ( n5857 & n14552 ) | ( n5857 & ~n14556 ) | ( n14552 & ~n14556 ) ;
  assign n14559 = ( n3499 & n6961 ) | ( n3499 & ~n8010 ) | ( n6961 & ~n8010 ) ;
  assign n14558 = ( n4080 & n7761 ) | ( n4080 & n8904 ) | ( n7761 & n8904 ) ;
  assign n14560 = n14559 ^ n14558 ^ n1459 ;
  assign n14561 = ( n2814 & n2906 ) | ( n2814 & ~n7323 ) | ( n2906 & ~n7323 ) ;
  assign n14562 = n14561 ^ n9907 ^ n869 ;
  assign n14563 = n14562 ^ n13591 ^ n9181 ;
  assign n14564 = n14563 ^ n7048 ^ n4373 ;
  assign n14568 = ( n193 & n3743 ) | ( n193 & ~n3863 ) | ( n3743 & ~n3863 ) ;
  assign n14565 = n7253 ^ n4793 ^ n1326 ;
  assign n14566 = n9264 ^ n1352 ^ n805 ;
  assign n14567 = ( n10111 & n14565 ) | ( n10111 & ~n14566 ) | ( n14565 & ~n14566 ) ;
  assign n14569 = n14568 ^ n14567 ^ n10280 ;
  assign n14570 = n10096 ^ n7007 ^ n6856 ;
  assign n14571 = ( n1677 & ~n2008 ) | ( n1677 & n14570 ) | ( ~n2008 & n14570 ) ;
  assign n14572 = n14571 ^ n6435 ^ n6293 ;
  assign n14573 = ( n705 & n3658 ) | ( n705 & n6019 ) | ( n3658 & n6019 ) ;
  assign n14574 = n14573 ^ n7923 ^ n645 ;
  assign n14575 = n7226 ^ n4600 ^ n2238 ;
  assign n14576 = ( n6124 & n6593 ) | ( n6124 & n14575 ) | ( n6593 & n14575 ) ;
  assign n14581 = ( ~n6222 & n7957 ) | ( ~n6222 & n11866 ) | ( n7957 & n11866 ) ;
  assign n14579 = ( n5179 & n7173 ) | ( n5179 & n11696 ) | ( n7173 & n11696 ) ;
  assign n14577 = n10809 ^ n2451 ^ n641 ;
  assign n14578 = ( n642 & n11101 ) | ( n642 & n14577 ) | ( n11101 & n14577 ) ;
  assign n14580 = n14579 ^ n14578 ^ n6266 ;
  assign n14582 = n14581 ^ n14580 ^ n2597 ;
  assign n14583 = n6140 ^ n5455 ^ n1040 ;
  assign n14584 = n14583 ^ n1407 ^ n1393 ;
  assign n14585 = ( n2406 & n3164 ) | ( n2406 & n6745 ) | ( n3164 & n6745 ) ;
  assign n14586 = ( n8852 & n14584 ) | ( n8852 & n14585 ) | ( n14584 & n14585 ) ;
  assign n14587 = ( n1357 & ~n7959 ) | ( n1357 & n9576 ) | ( ~n7959 & n9576 ) ;
  assign n14588 = ( ~n377 & n9833 ) | ( ~n377 & n14587 ) | ( n9833 & n14587 ) ;
  assign n14589 = ( ~n521 & n2105 ) | ( ~n521 & n2812 ) | ( n2105 & n2812 ) ;
  assign n14590 = n14589 ^ n5480 ^ n3865 ;
  assign n14591 = n14590 ^ n7709 ^ n7314 ;
  assign n14592 = n14591 ^ n13379 ^ n8767 ;
  assign n14593 = ( ~n3282 & n3708 ) | ( ~n3282 & n8677 ) | ( n3708 & n8677 ) ;
  assign n14594 = n14593 ^ n11813 ^ n2413 ;
  assign n14596 = n631 ^ n217 ^ x22 ;
  assign n14595 = ( n1597 & n2481 ) | ( n1597 & ~n7410 ) | ( n2481 & ~n7410 ) ;
  assign n14597 = n14596 ^ n14595 ^ n3179 ;
  assign n14598 = ( ~n9833 & n14594 ) | ( ~n9833 & n14597 ) | ( n14594 & n14597 ) ;
  assign n14599 = n12221 ^ n10912 ^ n4695 ;
  assign n14600 = ( n981 & n11645 ) | ( n981 & n13903 ) | ( n11645 & n13903 ) ;
  assign n14601 = ( ~n886 & n14599 ) | ( ~n886 & n14600 ) | ( n14599 & n14600 ) ;
  assign n14602 = n9136 ^ n4249 ^ n257 ;
  assign n14603 = ( n10249 & n11866 ) | ( n10249 & n14602 ) | ( n11866 & n14602 ) ;
  assign n14606 = n6959 ^ n3033 ^ n303 ;
  assign n14604 = n7683 ^ n7390 ^ n2966 ;
  assign n14605 = n14604 ^ n7020 ^ n3212 ;
  assign n14607 = n14606 ^ n14605 ^ n13160 ;
  assign n14608 = ( ~n9811 & n14264 ) | ( ~n9811 & n14607 ) | ( n14264 & n14607 ) ;
  assign n14609 = ( n558 & n4763 ) | ( n558 & n5464 ) | ( n4763 & n5464 ) ;
  assign n14610 = n4842 ^ n1480 ^ n1005 ;
  assign n14611 = n14610 ^ n4910 ^ n700 ;
  assign n14613 = ( n3976 & n4170 ) | ( n3976 & n7900 ) | ( n4170 & n7900 ) ;
  assign n14614 = ( n1722 & n2462 ) | ( n1722 & n14613 ) | ( n2462 & n14613 ) ;
  assign n14612 = n12235 ^ n5750 ^ n614 ;
  assign n14615 = n14614 ^ n14612 ^ n5213 ;
  assign n14619 = ( ~n6524 & n7922 ) | ( ~n6524 & n10905 ) | ( n7922 & n10905 ) ;
  assign n14620 = n14619 ^ n5141 ^ n2800 ;
  assign n14621 = ( ~n3021 & n5800 ) | ( ~n3021 & n14620 ) | ( n5800 & n14620 ) ;
  assign n14617 = n12300 ^ n3260 ^ n216 ;
  assign n14616 = ( n5347 & n8110 ) | ( n5347 & ~n10198 ) | ( n8110 & ~n10198 ) ;
  assign n14618 = n14617 ^ n14616 ^ n6812 ;
  assign n14622 = n14621 ^ n14618 ^ n13102 ;
  assign n14624 = ( ~n8295 & n9828 ) | ( ~n8295 & n12660 ) | ( n9828 & n12660 ) ;
  assign n14623 = n8200 ^ n4985 ^ n4183 ;
  assign n14625 = n14624 ^ n14623 ^ n6582 ;
  assign n14626 = ( n1417 & n3661 ) | ( n1417 & n13886 ) | ( n3661 & n13886 ) ;
  assign n14627 = ( ~n190 & n1388 ) | ( ~n190 & n4378 ) | ( n1388 & n4378 ) ;
  assign n14628 = n10781 ^ n7220 ^ n3364 ;
  assign n14629 = ( n3257 & ~n14627 ) | ( n3257 & n14628 ) | ( ~n14627 & n14628 ) ;
  assign n14630 = ( n3423 & n5734 ) | ( n3423 & n11300 ) | ( n5734 & n11300 ) ;
  assign n14631 = ( n2872 & n11369 ) | ( n2872 & ~n14630 ) | ( n11369 & ~n14630 ) ;
  assign n14632 = ( n443 & ~n3206 ) | ( n443 & n3821 ) | ( ~n3206 & n3821 ) ;
  assign n14633 = n14632 ^ n8345 ^ n3243 ;
  assign n14639 = ( n935 & n5725 ) | ( n935 & n6208 ) | ( n5725 & n6208 ) ;
  assign n14636 = n11303 ^ n9828 ^ n7621 ;
  assign n14637 = ( n3442 & n4703 ) | ( n3442 & ~n14636 ) | ( n4703 & ~n14636 ) ;
  assign n14634 = ( n586 & n3023 ) | ( n586 & n10215 ) | ( n3023 & n10215 ) ;
  assign n14635 = n14634 ^ n14436 ^ n7528 ;
  assign n14638 = n14637 ^ n14635 ^ n2911 ;
  assign n14640 = n14639 ^ n14638 ^ n2249 ;
  assign n14641 = n14640 ^ n13253 ^ n6420 ;
  assign n14642 = ( n14631 & n14633 ) | ( n14631 & ~n14641 ) | ( n14633 & ~n14641 ) ;
  assign n14643 = ( n326 & n569 ) | ( n326 & ~n3811 ) | ( n569 & ~n3811 ) ;
  assign n14644 = n9847 ^ n7571 ^ n4670 ;
  assign n14645 = n5679 ^ n1945 ^ n1729 ;
  assign n14646 = ( n14643 & n14644 ) | ( n14643 & n14645 ) | ( n14644 & n14645 ) ;
  assign n14647 = ( n5847 & n12179 ) | ( n5847 & n14646 ) | ( n12179 & n14646 ) ;
  assign n14649 = ( x109 & n938 ) | ( x109 & n4202 ) | ( n938 & n4202 ) ;
  assign n14650 = ( n7198 & n9134 ) | ( n7198 & n14649 ) | ( n9134 & n14649 ) ;
  assign n14651 = ( n1185 & n4251 ) | ( n1185 & n14650 ) | ( n4251 & n14650 ) ;
  assign n14648 = n2383 ^ n1771 ^ x93 ;
  assign n14652 = n14651 ^ n14648 ^ n9249 ;
  assign n14662 = n6319 ^ n5109 ^ n2501 ;
  assign n14663 = n14662 ^ n14536 ^ n3381 ;
  assign n14664 = ( n3234 & n3637 ) | ( n3234 & ~n14663 ) | ( n3637 & ~n14663 ) ;
  assign n14659 = n4510 ^ n1461 ^ n1279 ;
  assign n14655 = ( x49 & n2178 ) | ( x49 & n2657 ) | ( n2178 & n2657 ) ;
  assign n14656 = n14655 ^ n5859 ^ n3416 ;
  assign n14657 = n14656 ^ n2870 ^ n1057 ;
  assign n14658 = n14657 ^ n9028 ^ n4870 ;
  assign n14653 = ( n1137 & n3570 ) | ( n1137 & ~n7215 ) | ( n3570 & ~n7215 ) ;
  assign n14654 = n14653 ^ n3280 ^ n2209 ;
  assign n14660 = n14659 ^ n14658 ^ n14654 ;
  assign n14661 = n14660 ^ n8033 ^ n5592 ;
  assign n14665 = n14664 ^ n14661 ^ n11120 ;
  assign n14666 = ( n3938 & n7570 ) | ( n3938 & n7969 ) | ( n7570 & n7969 ) ;
  assign n14674 = n13072 ^ n4820 ^ n4422 ;
  assign n14675 = ( ~n1076 & n8747 ) | ( ~n1076 & n14674 ) | ( n8747 & n14674 ) ;
  assign n14676 = ( n5527 & ~n12067 ) | ( n5527 & n14675 ) | ( ~n12067 & n14675 ) ;
  assign n14667 = n12974 ^ n4554 ^ n4433 ;
  assign n14670 = n9287 ^ n7187 ^ n1563 ;
  assign n14668 = n11941 ^ n3484 ^ n2568 ;
  assign n14669 = ( ~n4064 & n13195 ) | ( ~n4064 & n14668 ) | ( n13195 & n14668 ) ;
  assign n14671 = n14670 ^ n14669 ^ n10282 ;
  assign n14672 = ( n2804 & ~n14667 ) | ( n2804 & n14671 ) | ( ~n14667 & n14671 ) ;
  assign n14673 = ( n5019 & n14627 ) | ( n5019 & n14672 ) | ( n14627 & n14672 ) ;
  assign n14677 = n14676 ^ n14673 ^ n12637 ;
  assign n14678 = ( n5291 & n14666 ) | ( n5291 & n14677 ) | ( n14666 & n14677 ) ;
  assign n14679 = ( n1609 & n2746 ) | ( n1609 & ~n14092 ) | ( n2746 & ~n14092 ) ;
  assign n14680 = n9853 ^ n4063 ^ n1520 ;
  assign n14681 = n14680 ^ n3103 ^ x12 ;
  assign n14688 = n12620 ^ n9779 ^ n9003 ;
  assign n14685 = ( n990 & n4013 ) | ( n990 & n9851 ) | ( n4013 & n9851 ) ;
  assign n14686 = n14685 ^ n9264 ^ n7590 ;
  assign n14683 = ( n193 & n251 ) | ( n193 & ~n6747 ) | ( n251 & ~n6747 ) ;
  assign n14684 = n14683 ^ n2616 ^ n497 ;
  assign n14682 = ( n688 & n4750 ) | ( n688 & n10153 ) | ( n4750 & n10153 ) ;
  assign n14687 = n14686 ^ n14684 ^ n14682 ;
  assign n14689 = n14688 ^ n14687 ^ n8010 ;
  assign n14690 = ( n13572 & ~n14681 ) | ( n13572 & n14689 ) | ( ~n14681 & n14689 ) ;
  assign n14691 = ( ~n1114 & n6428 ) | ( ~n1114 & n14537 ) | ( n6428 & n14537 ) ;
  assign n14692 = n3593 ^ n3451 ^ n3108 ;
  assign n14693 = n11820 ^ n5918 ^ n367 ;
  assign n14694 = ( ~n6612 & n10814 ) | ( ~n6612 & n14693 ) | ( n10814 & n14693 ) ;
  assign n14695 = ( n2840 & n7832 ) | ( n2840 & ~n14694 ) | ( n7832 & ~n14694 ) ;
  assign n14696 = ( n13312 & n14692 ) | ( n13312 & ~n14695 ) | ( n14692 & ~n14695 ) ;
  assign n14697 = n14696 ^ n8484 ^ n4482 ;
  assign n14699 = n10715 ^ n4557 ^ n1648 ;
  assign n14698 = n11193 ^ n7847 ^ n4786 ;
  assign n14700 = n14699 ^ n14698 ^ n13490 ;
  assign n14701 = n9570 ^ n7375 ^ n3380 ;
  assign n14702 = n13687 ^ n11845 ^ n1578 ;
  assign n14703 = ( ~x56 & n14701 ) | ( ~x56 & n14702 ) | ( n14701 & n14702 ) ;
  assign n14704 = ( n3170 & n5197 ) | ( n3170 & ~n14703 ) | ( n5197 & ~n14703 ) ;
  assign n14705 = n10842 ^ n8546 ^ n6384 ;
  assign n14706 = ( n7689 & n14587 ) | ( n7689 & ~n14705 ) | ( n14587 & ~n14705 ) ;
  assign n14707 = ( ~n2463 & n3376 ) | ( ~n2463 & n7862 ) | ( n3376 & n7862 ) ;
  assign n14708 = n14707 ^ n8634 ^ n8140 ;
  assign n14709 = ( n295 & n2131 ) | ( n295 & ~n14708 ) | ( n2131 & ~n14708 ) ;
  assign n14710 = ( n3318 & ~n10970 ) | ( n3318 & n11211 ) | ( ~n10970 & n11211 ) ;
  assign n14711 = n14710 ^ n12959 ^ n604 ;
  assign n14712 = ( n1461 & ~n9438 ) | ( n1461 & n10736 ) | ( ~n9438 & n10736 ) ;
  assign n14713 = n14712 ^ n6353 ^ n4002 ;
  assign n14714 = n14713 ^ n6974 ^ n2076 ;
  assign n14715 = ( n4049 & ~n8095 ) | ( n4049 & n14714 ) | ( ~n8095 & n14714 ) ;
  assign n14718 = n6828 ^ n5862 ^ n1748 ;
  assign n14719 = n14718 ^ n10319 ^ n5724 ;
  assign n14716 = n14365 ^ n7666 ^ n3546 ;
  assign n14717 = n14716 ^ n8684 ^ n3763 ;
  assign n14720 = n14719 ^ n14717 ^ n5866 ;
  assign n14721 = ( x69 & ~n10596 ) | ( x69 & n14720 ) | ( ~n10596 & n14720 ) ;
  assign n14722 = ( ~n6123 & n9521 ) | ( ~n6123 & n14721 ) | ( n9521 & n14721 ) ;
  assign n14723 = ( n1787 & n5519 ) | ( n1787 & ~n14722 ) | ( n5519 & ~n14722 ) ;
  assign n14724 = n4928 ^ n3292 ^ n658 ;
  assign n14725 = n14724 ^ n7497 ^ n6878 ;
  assign n14726 = n14725 ^ n13993 ^ n3690 ;
  assign n14727 = ( n1895 & ~n2931 ) | ( n1895 & n11268 ) | ( ~n2931 & n11268 ) ;
  assign n14728 = n14727 ^ n7087 ^ n4099 ;
  assign n14729 = ( n9405 & n11468 ) | ( n9405 & n13704 ) | ( n11468 & n13704 ) ;
  assign n14730 = ( ~n4052 & n7559 ) | ( ~n4052 & n10687 ) | ( n7559 & n10687 ) ;
  assign n14731 = ( n10906 & n11784 ) | ( n10906 & ~n14730 ) | ( n11784 & ~n14730 ) ;
  assign n14732 = ( ~n242 & n7243 ) | ( ~n242 & n13592 ) | ( n7243 & n13592 ) ;
  assign n14733 = n14732 ^ n13169 ^ n6929 ;
  assign n14734 = ( n6940 & n7257 ) | ( n6940 & n14733 ) | ( n7257 & n14733 ) ;
  assign n14735 = ( n6183 & n14731 ) | ( n6183 & n14734 ) | ( n14731 & n14734 ) ;
  assign n14736 = ( ~n12740 & n14729 ) | ( ~n12740 & n14735 ) | ( n14729 & n14735 ) ;
  assign n14737 = n12004 ^ n5776 ^ n1755 ;
  assign n14738 = n14737 ^ n10961 ^ n7107 ;
  assign n14740 = ( n314 & n6064 ) | ( n314 & n10659 ) | ( n6064 & n10659 ) ;
  assign n14739 = n11504 ^ n7403 ^ n5548 ;
  assign n14741 = n14740 ^ n14739 ^ n2262 ;
  assign n14742 = ( n657 & ~n1824 ) | ( n657 & n9192 ) | ( ~n1824 & n9192 ) ;
  assign n14743 = n14742 ^ n10003 ^ n1730 ;
  assign n14744 = ( n10723 & n12800 ) | ( n10723 & n14743 ) | ( n12800 & n14743 ) ;
  assign n14745 = ( ~n350 & n1689 ) | ( ~n350 & n14744 ) | ( n1689 & n14744 ) ;
  assign n14746 = ( n2379 & n7338 ) | ( n2379 & ~n10976 ) | ( n7338 & ~n10976 ) ;
  assign n14747 = ( n2435 & ~n13901 ) | ( n2435 & n14746 ) | ( ~n13901 & n14746 ) ;
  assign n14749 = n2422 ^ n1738 ^ n1088 ;
  assign n14748 = n9766 ^ n9043 ^ n4163 ;
  assign n14750 = n14749 ^ n14748 ^ n2175 ;
  assign n14751 = ( n4790 & n11514 ) | ( n4790 & n14750 ) | ( n11514 & n14750 ) ;
  assign n14753 = n13807 ^ n8306 ^ n8220 ;
  assign n14754 = n4994 ^ n4541 ^ n1051 ;
  assign n14755 = ( n6828 & ~n14753 ) | ( n6828 & n14754 ) | ( ~n14753 & n14754 ) ;
  assign n14752 = ( n10639 & n11891 ) | ( n10639 & ~n13769 ) | ( n11891 & ~n13769 ) ;
  assign n14756 = n14755 ^ n14752 ^ n12830 ;
  assign n14757 = ( n1845 & n3789 ) | ( n1845 & n10561 ) | ( n3789 & n10561 ) ;
  assign n14758 = ( ~n3963 & n10723 ) | ( ~n3963 & n14757 ) | ( n10723 & n14757 ) ;
  assign n14759 = n14758 ^ n3055 ^ n1316 ;
  assign n14762 = ( ~n1706 & n2188 ) | ( ~n1706 & n9589 ) | ( n2188 & n9589 ) ;
  assign n14760 = ( n431 & ~n1984 ) | ( n431 & n5818 ) | ( ~n1984 & n5818 ) ;
  assign n14761 = ( ~n359 & n10089 ) | ( ~n359 & n14760 ) | ( n10089 & n14760 ) ;
  assign n14763 = n14762 ^ n14761 ^ n5800 ;
  assign n14764 = ( n14019 & n14759 ) | ( n14019 & n14763 ) | ( n14759 & n14763 ) ;
  assign n14765 = n13550 ^ n11666 ^ n7867 ;
  assign n14766 = ( ~n1794 & n1893 ) | ( ~n1794 & n3035 ) | ( n1893 & n3035 ) ;
  assign n14767 = ( n2604 & ~n10879 ) | ( n2604 & n14766 ) | ( ~n10879 & n14766 ) ;
  assign n14768 = n13059 ^ n11068 ^ n3131 ;
  assign n14769 = n14768 ^ n14132 ^ n483 ;
  assign n14770 = ( n4681 & n14767 ) | ( n4681 & ~n14769 ) | ( n14767 & ~n14769 ) ;
  assign n14771 = n14066 ^ n10082 ^ n9269 ;
  assign n14773 = ( ~n1531 & n2237 ) | ( ~n1531 & n2796 ) | ( n2237 & n2796 ) ;
  assign n14774 = ( ~n6241 & n6785 ) | ( ~n6241 & n14773 ) | ( n6785 & n14773 ) ;
  assign n14772 = n14562 ^ n13926 ^ n1143 ;
  assign n14775 = n14774 ^ n14772 ^ n2518 ;
  assign n14776 = ( n3658 & n14771 ) | ( n3658 & ~n14775 ) | ( n14771 & ~n14775 ) ;
  assign n14777 = n12318 ^ n7481 ^ n7056 ;
  assign n14778 = ( n2167 & n8702 ) | ( n2167 & n14777 ) | ( n8702 & n14777 ) ;
  assign n14779 = n10650 ^ n8902 ^ n3422 ;
  assign n14780 = ( n1450 & ~n4517 ) | ( n1450 & n4527 ) | ( ~n4517 & n4527 ) ;
  assign n14781 = n14780 ^ n5281 ^ n2612 ;
  assign n14782 = ( n7323 & n7602 ) | ( n7323 & ~n14781 ) | ( n7602 & ~n14781 ) ;
  assign n14783 = ( ~n6238 & n14779 ) | ( ~n6238 & n14782 ) | ( n14779 & n14782 ) ;
  assign n14784 = ( n6595 & ~n8798 ) | ( n6595 & n11263 ) | ( ~n8798 & n11263 ) ;
  assign n14785 = ( n4366 & n9629 ) | ( n4366 & ~n11862 ) | ( n9629 & ~n11862 ) ;
  assign n14786 = ( n14114 & ~n14784 ) | ( n14114 & n14785 ) | ( ~n14784 & n14785 ) ;
  assign n14787 = n12300 ^ n6680 ^ n4083 ;
  assign n14788 = n14787 ^ n2711 ^ n1377 ;
  assign n14793 = n5761 ^ n3466 ^ n271 ;
  assign n14794 = ( n4951 & ~n7377 ) | ( n4951 & n14793 ) | ( ~n7377 & n14793 ) ;
  assign n14795 = ( ~n1567 & n3291 ) | ( ~n1567 & n14794 ) | ( n3291 & n14794 ) ;
  assign n14789 = ( n1346 & ~n4482 ) | ( n1346 & n6357 ) | ( ~n4482 & n6357 ) ;
  assign n14790 = n14789 ^ n8614 ^ n254 ;
  assign n14791 = n14790 ^ n5516 ^ n725 ;
  assign n14792 = n14791 ^ n10619 ^ x16 ;
  assign n14796 = n14795 ^ n14792 ^ n3951 ;
  assign n14797 = ( n12333 & n14788 ) | ( n12333 & n14796 ) | ( n14788 & n14796 ) ;
  assign n14798 = ( n3276 & ~n12644 ) | ( n3276 & n14505 ) | ( ~n12644 & n14505 ) ;
  assign n14801 = n13256 ^ n7934 ^ n6300 ;
  assign n14799 = ( n4241 & n6179 ) | ( n4241 & n7677 ) | ( n6179 & n7677 ) ;
  assign n14800 = n14799 ^ n5440 ^ n3260 ;
  assign n14802 = n14801 ^ n14800 ^ n6265 ;
  assign n14804 = n5101 ^ n2978 ^ n1385 ;
  assign n14803 = ( n3777 & n4225 ) | ( n3777 & n4574 ) | ( n4225 & n4574 ) ;
  assign n14805 = n14804 ^ n14803 ^ n3124 ;
  assign n14811 = ( n3041 & n12238 ) | ( n3041 & ~n12915 ) | ( n12238 & ~n12915 ) ;
  assign n14812 = ( n3231 & n11618 ) | ( n3231 & ~n14811 ) | ( n11618 & ~n14811 ) ;
  assign n14813 = n14812 ^ n6689 ^ n5334 ;
  assign n14814 = n14813 ^ n9377 ^ n6089 ;
  assign n14815 = ( n2092 & ~n3519 ) | ( n2092 & n8782 ) | ( ~n3519 & n8782 ) ;
  assign n14816 = ( ~n2526 & n11718 ) | ( ~n2526 & n14815 ) | ( n11718 & n14815 ) ;
  assign n14817 = ( ~n7235 & n14814 ) | ( ~n7235 & n14816 ) | ( n14814 & n14816 ) ;
  assign n14809 = ( n3776 & n5504 ) | ( n3776 & ~n10306 ) | ( n5504 & ~n10306 ) ;
  assign n14806 = ( n3667 & n4870 ) | ( n3667 & ~n5099 ) | ( n4870 & ~n5099 ) ;
  assign n14807 = n14806 ^ n4036 ^ n941 ;
  assign n14808 = ( ~n8681 & n13379 ) | ( ~n8681 & n14807 ) | ( n13379 & n14807 ) ;
  assign n14810 = n14809 ^ n14808 ^ n1727 ;
  assign n14818 = n14817 ^ n14810 ^ n3414 ;
  assign n14819 = ( n3250 & n10602 ) | ( n3250 & ~n12970 ) | ( n10602 & ~n12970 ) ;
  assign n14820 = ( ~n2398 & n10354 ) | ( ~n2398 & n14819 ) | ( n10354 & n14819 ) ;
  assign n14821 = ( n9788 & n12078 ) | ( n9788 & n14820 ) | ( n12078 & n14820 ) ;
  assign n14822 = ( n1320 & n7125 ) | ( n1320 & ~n14821 ) | ( n7125 & ~n14821 ) ;
  assign n14823 = n9100 ^ n5100 ^ n764 ;
  assign n14824 = n14823 ^ n14429 ^ n8741 ;
  assign n14825 = ( ~x6 & n764 ) | ( ~x6 & n1905 ) | ( n764 & n1905 ) ;
  assign n14826 = n14825 ^ n11415 ^ n5855 ;
  assign n14827 = n14826 ^ n11050 ^ n1031 ;
  assign n14828 = ( ~n808 & n11099 ) | ( ~n808 & n14827 ) | ( n11099 & n14827 ) ;
  assign n14831 = n9698 ^ n5590 ^ n373 ;
  assign n14829 = n11852 ^ n4984 ^ n611 ;
  assign n14830 = ( ~n1266 & n7961 ) | ( ~n1266 & n14829 ) | ( n7961 & n14829 ) ;
  assign n14832 = n14831 ^ n14830 ^ n2424 ;
  assign n14833 = n8586 ^ n7473 ^ n5196 ;
  assign n14834 = ( n2488 & n13073 ) | ( n2488 & n14833 ) | ( n13073 & n14833 ) ;
  assign n14835 = n14834 ^ n10281 ^ n7734 ;
  assign n14841 = n3701 ^ n2357 ^ n1493 ;
  assign n14840 = ( ~n3385 & n5830 ) | ( ~n3385 & n7358 ) | ( n5830 & n7358 ) ;
  assign n14842 = n14841 ^ n14840 ^ n10482 ;
  assign n14837 = n8881 ^ n7168 ^ n5029 ;
  assign n14836 = ( n2111 & ~n9550 ) | ( n2111 & n10774 ) | ( ~n9550 & n10774 ) ;
  assign n14838 = n14837 ^ n14836 ^ n9026 ;
  assign n14839 = ( n9234 & n10006 ) | ( n9234 & ~n14838 ) | ( n10006 & ~n14838 ) ;
  assign n14843 = n14842 ^ n14839 ^ n5838 ;
  assign n14844 = ( ~n3554 & n14835 ) | ( ~n3554 & n14843 ) | ( n14835 & n14843 ) ;
  assign n14845 = ( n2177 & n2482 ) | ( n2177 & n3367 ) | ( n2482 & n3367 ) ;
  assign n14846 = ( n9525 & n12089 ) | ( n9525 & n14845 ) | ( n12089 & n14845 ) ;
  assign n14847 = ( n749 & ~n8921 ) | ( n749 & n14846 ) | ( ~n8921 & n14846 ) ;
  assign n14848 = ( n1065 & n3004 ) | ( n1065 & ~n3312 ) | ( n3004 & ~n3312 ) ;
  assign n14849 = ( n4665 & ~n11110 ) | ( n4665 & n14848 ) | ( ~n11110 & n14848 ) ;
  assign n14850 = n6869 ^ n5152 ^ n568 ;
  assign n14851 = ( ~n793 & n9431 ) | ( ~n793 & n14850 ) | ( n9431 & n14850 ) ;
  assign n14852 = ( n10936 & n14195 ) | ( n10936 & n14851 ) | ( n14195 & n14851 ) ;
  assign n14853 = ( n14847 & n14849 ) | ( n14847 & n14852 ) | ( n14849 & n14852 ) ;
  assign n14857 = ( ~n4812 & n8372 ) | ( ~n4812 & n10497 ) | ( n8372 & n10497 ) ;
  assign n14858 = n14857 ^ n13931 ^ n7756 ;
  assign n14854 = n10997 ^ n5450 ^ n5103 ;
  assign n14855 = ( n736 & n2128 ) | ( n736 & ~n7042 ) | ( n2128 & ~n7042 ) ;
  assign n14856 = ( n14274 & n14854 ) | ( n14274 & n14855 ) | ( n14854 & n14855 ) ;
  assign n14859 = n14858 ^ n14856 ^ n2323 ;
  assign n14860 = n6725 ^ n5297 ^ n2164 ;
  assign n14861 = ( n3633 & n3941 ) | ( n3633 & n5068 ) | ( n3941 & n5068 ) ;
  assign n14862 = n14861 ^ n4901 ^ n1880 ;
  assign n14863 = ( ~n7495 & n14860 ) | ( ~n7495 & n14862 ) | ( n14860 & n14862 ) ;
  assign n14865 = n8827 ^ n2055 ^ n1562 ;
  assign n14864 = ( n3262 & n6177 ) | ( n3262 & ~n14118 ) | ( n6177 & ~n14118 ) ;
  assign n14866 = n14865 ^ n14864 ^ n8272 ;
  assign n14867 = ( n3087 & ~n5765 ) | ( n3087 & n13160 ) | ( ~n5765 & n13160 ) ;
  assign n14868 = ( n590 & ~n14866 ) | ( n590 & n14867 ) | ( ~n14866 & n14867 ) ;
  assign n14869 = n7326 ^ n5870 ^ n3844 ;
  assign n14870 = ( n7654 & ~n8347 ) | ( n7654 & n9151 ) | ( ~n8347 & n9151 ) ;
  assign n14871 = ( n6532 & n14869 ) | ( n6532 & ~n14870 ) | ( n14869 & ~n14870 ) ;
  assign n14872 = ( n1655 & ~n5549 ) | ( n1655 & n14350 ) | ( ~n5549 & n14350 ) ;
  assign n14873 = ( n5545 & n8234 ) | ( n5545 & n9510 ) | ( n8234 & n9510 ) ;
  assign n14874 = n14873 ^ n7912 ^ n4359 ;
  assign n14875 = ( n2188 & n7226 ) | ( n2188 & n14874 ) | ( n7226 & n14874 ) ;
  assign n14876 = ( n9575 & n14872 ) | ( n9575 & n14875 ) | ( n14872 & n14875 ) ;
  assign n14877 = ( n14732 & ~n14871 ) | ( n14732 & n14876 ) | ( ~n14871 & n14876 ) ;
  assign n14884 = n12602 ^ n3768 ^ n1140 ;
  assign n14878 = n12278 ^ n2986 ^ n1372 ;
  assign n14880 = n5564 ^ n3690 ^ n2786 ;
  assign n14879 = n13748 ^ n12545 ^ n821 ;
  assign n14881 = n14880 ^ n14879 ^ n3517 ;
  assign n14882 = n14881 ^ n11099 ^ n3684 ;
  assign n14883 = ( n2548 & n14878 ) | ( n2548 & ~n14882 ) | ( n14878 & ~n14882 ) ;
  assign n14885 = n14884 ^ n14883 ^ n1441 ;
  assign n14887 = n5993 ^ n2093 ^ n2015 ;
  assign n14888 = ( n1817 & n5476 ) | ( n1817 & n14887 ) | ( n5476 & n14887 ) ;
  assign n14886 = ( n818 & n4941 ) | ( n818 & n8005 ) | ( n4941 & n8005 ) ;
  assign n14889 = n14888 ^ n14886 ^ n6409 ;
  assign n14890 = n12136 ^ n6150 ^ n1983 ;
  assign n14891 = n14890 ^ n6501 ^ n6259 ;
  assign n14892 = ( n434 & n14889 ) | ( n434 & n14891 ) | ( n14889 & n14891 ) ;
  assign n14893 = ( ~n3168 & n11960 ) | ( ~n3168 & n12012 ) | ( n11960 & n12012 ) ;
  assign n14894 = ( ~n4092 & n13923 ) | ( ~n4092 & n14893 ) | ( n13923 & n14893 ) ;
  assign n14895 = n7403 ^ n2846 ^ n2485 ;
  assign n14896 = ( n6953 & n11416 ) | ( n6953 & ~n13881 ) | ( n11416 & ~n13881 ) ;
  assign n14897 = ( n220 & n8807 ) | ( n220 & ~n14849 ) | ( n8807 & ~n14849 ) ;
  assign n14898 = ( n748 & n2944 ) | ( n748 & ~n10305 ) | ( n2944 & ~n10305 ) ;
  assign n14899 = ( n10644 & ~n14897 ) | ( n10644 & n14898 ) | ( ~n14897 & n14898 ) ;
  assign n14900 = ( ~n12517 & n14896 ) | ( ~n12517 & n14899 ) | ( n14896 & n14899 ) ;
  assign n14901 = n9579 ^ n7411 ^ x94 ;
  assign n14902 = ( ~n575 & n923 ) | ( ~n575 & n14901 ) | ( n923 & n14901 ) ;
  assign n14903 = n14902 ^ n12225 ^ n8930 ;
  assign n14904 = ( n1501 & n2287 ) | ( n1501 & n10743 ) | ( n2287 & n10743 ) ;
  assign n14905 = n6237 ^ n5352 ^ n2990 ;
  assign n14906 = ( ~n7311 & n7483 ) | ( ~n7311 & n14905 ) | ( n7483 & n14905 ) ;
  assign n14907 = ( n1863 & n14904 ) | ( n1863 & ~n14906 ) | ( n14904 & ~n14906 ) ;
  assign n14908 = ( n2892 & n9527 ) | ( n2892 & n12307 ) | ( n9527 & n12307 ) ;
  assign n14909 = ( n5038 & n5908 ) | ( n5038 & ~n6709 ) | ( n5908 & ~n6709 ) ;
  assign n14910 = ( ~n2741 & n8142 ) | ( ~n2741 & n14909 ) | ( n8142 & n14909 ) ;
  assign n14911 = ( n2077 & n2358 ) | ( n2077 & n2998 ) | ( n2358 & n2998 ) ;
  assign n14914 = n8360 ^ n8099 ^ n7590 ;
  assign n14915 = ( x30 & ~n4141 ) | ( x30 & n14914 ) | ( ~n4141 & n14914 ) ;
  assign n14912 = ( ~n1103 & n4825 ) | ( ~n1103 & n11207 ) | ( n4825 & n11207 ) ;
  assign n14913 = n14912 ^ n9810 ^ n9096 ;
  assign n14916 = n14915 ^ n14913 ^ n13859 ;
  assign n14917 = ( ~n13355 & n14911 ) | ( ~n13355 & n14916 ) | ( n14911 & n14916 ) ;
  assign n14918 = n14917 ^ n9997 ^ n5147 ;
  assign n14919 = ( n2755 & n8865 ) | ( n2755 & ~n10116 ) | ( n8865 & ~n10116 ) ;
  assign n14923 = n11763 ^ n9478 ^ n1552 ;
  assign n14924 = ( n5699 & ~n6316 ) | ( n5699 & n14923 ) | ( ~n6316 & n14923 ) ;
  assign n14921 = n9270 ^ n8448 ^ n5913 ;
  assign n14920 = n11567 ^ n8765 ^ n6456 ;
  assign n14922 = n14921 ^ n14920 ^ n13234 ;
  assign n14925 = n14924 ^ n14922 ^ n6312 ;
  assign n14926 = ( n3291 & n5494 ) | ( n3291 & n5880 ) | ( n5494 & n5880 ) ;
  assign n14927 = n14926 ^ n6460 ^ n5446 ;
  assign n14928 = n14927 ^ n14350 ^ n762 ;
  assign n14929 = ( n5206 & ~n8142 ) | ( n5206 & n14928 ) | ( ~n8142 & n14928 ) ;
  assign n14930 = n3719 ^ n1686 ^ n660 ;
  assign n14931 = n9587 ^ n5175 ^ n441 ;
  assign n14932 = n8088 ^ n7140 ^ n3431 ;
  assign n14933 = n14932 ^ n8477 ^ n4054 ;
  assign n14934 = ( n14930 & n14931 ) | ( n14930 & n14933 ) | ( n14931 & n14933 ) ;
  assign n14935 = ( n1246 & ~n6562 ) | ( n1246 & n14934 ) | ( ~n6562 & n14934 ) ;
  assign n14936 = ( n2261 & n11965 ) | ( n2261 & ~n14935 ) | ( n11965 & ~n14935 ) ;
  assign n14937 = ( n2609 & n2634 ) | ( n2609 & n14936 ) | ( n2634 & n14936 ) ;
  assign n14940 = n10594 ^ n6298 ^ n1134 ;
  assign n14941 = n14940 ^ n7124 ^ n841 ;
  assign n14942 = ( n1261 & ~n1904 ) | ( n1261 & n14941 ) | ( ~n1904 & n14941 ) ;
  assign n14943 = ( n4117 & n8113 ) | ( n4117 & n14942 ) | ( n8113 & n14942 ) ;
  assign n14938 = ( n585 & ~n1032 ) | ( n585 & n12621 ) | ( ~n1032 & n12621 ) ;
  assign n14939 = ( n8484 & ~n11722 ) | ( n8484 & n14938 ) | ( ~n11722 & n14938 ) ;
  assign n14944 = n14943 ^ n14939 ^ n8175 ;
  assign n14945 = n6559 ^ n2884 ^ n1742 ;
  assign n14946 = ( ~n3749 & n9548 ) | ( ~n3749 & n14945 ) | ( n9548 & n14945 ) ;
  assign n14947 = n9488 ^ n3848 ^ n970 ;
  assign n14948 = n13671 ^ n7006 ^ n2204 ;
  assign n14949 = n4638 ^ n1509 ^ n457 ;
  assign n14950 = ( n852 & n14948 ) | ( n852 & n14949 ) | ( n14948 & n14949 ) ;
  assign n14951 = ( n11852 & n14653 ) | ( n11852 & ~n14950 ) | ( n14653 & ~n14950 ) ;
  assign n14953 = n7914 ^ n5690 ^ n2914 ;
  assign n14954 = ( ~n1476 & n5505 ) | ( ~n1476 & n14953 ) | ( n5505 & n14953 ) ;
  assign n14952 = ( n708 & n1381 ) | ( n708 & ~n2588 ) | ( n1381 & ~n2588 ) ;
  assign n14955 = n14954 ^ n14952 ^ n3988 ;
  assign n14956 = n14955 ^ n11089 ^ n8866 ;
  assign n14957 = ( n5368 & n9479 ) | ( n5368 & n14956 ) | ( n9479 & n14956 ) ;
  assign n14958 = ( n5122 & n5367 ) | ( n5122 & ~n11984 ) | ( n5367 & ~n11984 ) ;
  assign n14960 = n3951 ^ n3209 ^ n2530 ;
  assign n14959 = ( n10545 & ~n11070 ) | ( n10545 & n12022 ) | ( ~n11070 & n12022 ) ;
  assign n14961 = n14960 ^ n14959 ^ n14851 ;
  assign n14962 = ( n490 & n1527 ) | ( n490 & n4841 ) | ( n1527 & n4841 ) ;
  assign n14963 = ( ~n2292 & n9369 ) | ( ~n2292 & n14962 ) | ( n9369 & n14962 ) ;
  assign n14964 = ( n732 & n3830 ) | ( n732 & ~n13008 ) | ( n3830 & ~n13008 ) ;
  assign n14969 = ( n3634 & n5912 ) | ( n3634 & ~n11089 ) | ( n5912 & ~n11089 ) ;
  assign n14965 = n2385 ^ n1224 ^ x50 ;
  assign n14966 = ( ~x71 & n1585 ) | ( ~x71 & n4762 ) | ( n1585 & n4762 ) ;
  assign n14967 = ( n11088 & n14965 ) | ( n11088 & ~n14966 ) | ( n14965 & ~n14966 ) ;
  assign n14968 = ( n8808 & n12090 ) | ( n8808 & ~n14967 ) | ( n12090 & ~n14967 ) ;
  assign n14970 = n14969 ^ n14968 ^ n13440 ;
  assign n14974 = ( n1986 & n4204 ) | ( n1986 & n6338 ) | ( n4204 & n6338 ) ;
  assign n14975 = n12767 ^ n10116 ^ n1984 ;
  assign n14976 = ( n1363 & n5772 ) | ( n1363 & n6669 ) | ( n5772 & n6669 ) ;
  assign n14977 = n14976 ^ n12019 ^ n8464 ;
  assign n14978 = ( n13943 & ~n14975 ) | ( n13943 & n14977 ) | ( ~n14975 & n14977 ) ;
  assign n14979 = ( n8782 & ~n14974 ) | ( n8782 & n14978 ) | ( ~n14974 & n14978 ) ;
  assign n14971 = ( n3509 & n7134 ) | ( n3509 & ~n8727 ) | ( n7134 & ~n8727 ) ;
  assign n14972 = ( n7922 & n10622 ) | ( n7922 & n14971 ) | ( n10622 & n14971 ) ;
  assign n14973 = n14972 ^ n10856 ^ n7050 ;
  assign n14980 = n14979 ^ n14973 ^ n4708 ;
  assign n14986 = n5136 ^ n594 ^ n249 ;
  assign n14984 = n13998 ^ n6696 ^ n1808 ;
  assign n14985 = ( ~n1752 & n5935 ) | ( ~n1752 & n14984 ) | ( n5935 & n14984 ) ;
  assign n14981 = n3731 ^ n2621 ^ n1138 ;
  assign n14982 = ( n1642 & ~n7585 ) | ( n1642 & n14981 ) | ( ~n7585 & n14981 ) ;
  assign n14983 = ( n669 & n12390 ) | ( n669 & ~n14982 ) | ( n12390 & ~n14982 ) ;
  assign n14987 = n14986 ^ n14985 ^ n14983 ;
  assign n14988 = ( ~n2686 & n13707 ) | ( ~n2686 & n14817 ) | ( n13707 & n14817 ) ;
  assign n14989 = n4953 ^ n3840 ^ n2225 ;
  assign n14990 = ( n558 & n9052 ) | ( n558 & ~n14989 ) | ( n9052 & ~n14989 ) ;
  assign n14991 = n5406 ^ n4359 ^ x24 ;
  assign n14992 = ( n2492 & n5902 ) | ( n2492 & ~n14991 ) | ( n5902 & ~n14991 ) ;
  assign n14993 = n8058 ^ n6568 ^ n637 ;
  assign n14994 = n14993 ^ n6988 ^ n2892 ;
  assign n14995 = ( n11571 & n14992 ) | ( n11571 & ~n14994 ) | ( n14992 & ~n14994 ) ;
  assign n14996 = ( n6977 & n14990 ) | ( n6977 & n14995 ) | ( n14990 & n14995 ) ;
  assign n14997 = n14996 ^ n8573 ^ n372 ;
  assign n14998 = ( n7501 & n10569 ) | ( n7501 & ~n14997 ) | ( n10569 & ~n14997 ) ;
  assign n14999 = ( n2102 & n5382 ) | ( n2102 & n5654 ) | ( n5382 & n5654 ) ;
  assign n15000 = ( n1511 & n2604 ) | ( n1511 & n4729 ) | ( n2604 & n4729 ) ;
  assign n15001 = ( n5421 & n7986 ) | ( n5421 & ~n15000 ) | ( n7986 & ~n15000 ) ;
  assign n15003 = n9068 ^ n8036 ^ n7094 ;
  assign n15002 = n10725 ^ n10511 ^ n939 ;
  assign n15004 = n15003 ^ n15002 ^ n4903 ;
  assign n15005 = n15004 ^ n12883 ^ n5509 ;
  assign n15007 = n2814 ^ n1377 ^ n724 ;
  assign n15006 = n4812 ^ n3288 ^ x99 ;
  assign n15008 = n15007 ^ n15006 ^ n9482 ;
  assign n15009 = n6711 ^ n4188 ^ n1327 ;
  assign n15010 = ( n14344 & n15008 ) | ( n14344 & n15009 ) | ( n15008 & n15009 ) ;
  assign n15020 = n10571 ^ n6691 ^ n5327 ;
  assign n15019 = n13045 ^ n4445 ^ n4267 ;
  assign n15021 = n15020 ^ n15019 ^ n1943 ;
  assign n15016 = n7683 ^ n6981 ^ n3556 ;
  assign n15014 = ( ~n291 & n1314 ) | ( ~n291 & n4463 ) | ( n1314 & n4463 ) ;
  assign n15015 = n15014 ^ n7811 ^ n5147 ;
  assign n15012 = ( n3624 & ~n9026 ) | ( n3624 & n11263 ) | ( ~n9026 & n11263 ) ;
  assign n15013 = n15012 ^ n6215 ^ n5589 ;
  assign n15017 = n15016 ^ n15015 ^ n15013 ;
  assign n15011 = n9846 ^ n5267 ^ n4238 ;
  assign n15018 = n15017 ^ n15011 ^ n3929 ;
  assign n15022 = n15021 ^ n15018 ^ n9487 ;
  assign n15027 = n7479 ^ n7311 ^ n884 ;
  assign n15028 = ( ~n6285 & n11847 ) | ( ~n6285 & n15027 ) | ( n11847 & n15027 ) ;
  assign n15025 = ( n6092 & n8865 ) | ( n6092 & n10848 ) | ( n8865 & n10848 ) ;
  assign n15026 = ( n6751 & n9188 ) | ( n6751 & ~n15025 ) | ( n9188 & ~n15025 ) ;
  assign n15023 = ( n1984 & n6524 ) | ( n1984 & n9045 ) | ( n6524 & n9045 ) ;
  assign n15024 = ( ~n10473 & n11064 ) | ( ~n10473 & n15023 ) | ( n11064 & n15023 ) ;
  assign n15029 = n15028 ^ n15026 ^ n15024 ;
  assign n15030 = n12903 ^ n7763 ^ n3873 ;
  assign n15031 = n11572 ^ n5530 ^ n3529 ;
  assign n15032 = ( n9764 & n13675 ) | ( n9764 & n15031 ) | ( n13675 & n15031 ) ;
  assign n15033 = ( n1676 & ~n11657 ) | ( n1676 & n13042 ) | ( ~n11657 & n13042 ) ;
  assign n15034 = ( n6488 & n7416 ) | ( n6488 & n13059 ) | ( n7416 & n13059 ) ;
  assign n15035 = n15034 ^ n3945 ^ n994 ;
  assign n15036 = ( n8542 & n15033 ) | ( n8542 & n15035 ) | ( n15033 & n15035 ) ;
  assign n15037 = n11927 ^ n10971 ^ n136 ;
  assign n15038 = n15037 ^ n12492 ^ n6682 ;
  assign n15040 = ( n2499 & ~n5029 ) | ( n2499 & n10199 ) | ( ~n5029 & n10199 ) ;
  assign n15039 = ( n3510 & n3569 ) | ( n3510 & ~n11667 ) | ( n3569 & ~n11667 ) ;
  assign n15041 = n15040 ^ n15039 ^ n5044 ;
  assign n15042 = n7322 ^ n2255 ^ n763 ;
  assign n15043 = n15042 ^ n9082 ^ n251 ;
  assign n15044 = n3397 ^ n3018 ^ n1916 ;
  assign n15045 = n15044 ^ n14264 ^ n5618 ;
  assign n15046 = ( n6008 & ~n12932 ) | ( n6008 & n15045 ) | ( ~n12932 & n15045 ) ;
  assign n15047 = ( n3492 & ~n10943 ) | ( n3492 & n15046 ) | ( ~n10943 & n15046 ) ;
  assign n15048 = n4744 ^ n3768 ^ n2732 ;
  assign n15049 = ( ~n12808 & n13917 ) | ( ~n12808 & n15048 ) | ( n13917 & n15048 ) ;
  assign n15050 = n14381 ^ n5296 ^ n1336 ;
  assign n15051 = ( n2565 & n11513 ) | ( n2565 & ~n14242 ) | ( n11513 & ~n14242 ) ;
  assign n15052 = n15051 ^ n10228 ^ n1775 ;
  assign n15053 = ( n2548 & n7222 ) | ( n2548 & n15052 ) | ( n7222 & n15052 ) ;
  assign n15054 = ( n2673 & n4745 ) | ( n2673 & ~n7992 ) | ( n4745 & ~n7992 ) ;
  assign n15055 = n10963 ^ n2773 ^ n284 ;
  assign n15056 = ( n2745 & n15054 ) | ( n2745 & n15055 ) | ( n15054 & n15055 ) ;
  assign n15057 = n11941 ^ n6157 ^ n2997 ;
  assign n15058 = n15057 ^ n12752 ^ n10868 ;
  assign n15059 = n15058 ^ n11767 ^ n10176 ;
  assign n15060 = ( n841 & n6978 ) | ( n841 & n8768 ) | ( n6978 & n8768 ) ;
  assign n15061 = n1938 ^ n1591 ^ n175 ;
  assign n15062 = ( n1488 & n3029 ) | ( n1488 & n15061 ) | ( n3029 & n15061 ) ;
  assign n15066 = n11426 ^ n6308 ^ n4343 ;
  assign n15067 = n15066 ^ n10532 ^ n3125 ;
  assign n15065 = ( ~x18 & n5620 ) | ( ~x18 & n13020 ) | ( n5620 & n13020 ) ;
  assign n15063 = ( n1275 & n1683 ) | ( n1275 & n3885 ) | ( n1683 & n3885 ) ;
  assign n15064 = ( n11318 & n13368 ) | ( n11318 & n15063 ) | ( n13368 & n15063 ) ;
  assign n15068 = n15067 ^ n15065 ^ n15064 ;
  assign n15069 = ( n3876 & n6387 ) | ( n3876 & n10673 ) | ( n6387 & n10673 ) ;
  assign n15070 = ( n15062 & n15068 ) | ( n15062 & ~n15069 ) | ( n15068 & ~n15069 ) ;
  assign n15071 = n7794 ^ n5297 ^ n2517 ;
  assign n15072 = ( ~n191 & n14005 ) | ( ~n191 & n15071 ) | ( n14005 & n15071 ) ;
  assign n15083 = ( n1623 & n3592 ) | ( n1623 & ~n4604 ) | ( n3592 & ~n4604 ) ;
  assign n15084 = ( n787 & ~n10964 ) | ( n787 & n15083 ) | ( ~n10964 & n15083 ) ;
  assign n15073 = ( x18 & ~n2028 ) | ( x18 & n6525 ) | ( ~n2028 & n6525 ) ;
  assign n15074 = ( n1151 & ~n14494 ) | ( n1151 & n15073 ) | ( ~n14494 & n15073 ) ;
  assign n15075 = ( n3673 & n6416 ) | ( n3673 & ~n7449 ) | ( n6416 & ~n7449 ) ;
  assign n15076 = n15075 ^ n14780 ^ n4745 ;
  assign n15077 = n8037 ^ n7518 ^ n7381 ;
  assign n15078 = n5162 ^ n1007 ^ n893 ;
  assign n15079 = n15078 ^ n13389 ^ n6799 ;
  assign n15080 = ( n6018 & ~n11059 ) | ( n6018 & n15079 ) | ( ~n11059 & n15079 ) ;
  assign n15081 = ( n15076 & n15077 ) | ( n15076 & n15080 ) | ( n15077 & n15080 ) ;
  assign n15082 = ( ~n5323 & n15074 ) | ( ~n5323 & n15081 ) | ( n15074 & n15081 ) ;
  assign n15085 = n15084 ^ n15082 ^ n7515 ;
  assign n15086 = n10771 ^ n9785 ^ n3740 ;
  assign n15087 = ( n2978 & n10023 ) | ( n2978 & n12067 ) | ( n10023 & n12067 ) ;
  assign n15088 = ( ~n9245 & n15086 ) | ( ~n9245 & n15087 ) | ( n15086 & n15087 ) ;
  assign n15090 = n13784 ^ n5553 ^ n1241 ;
  assign n15089 = n11343 ^ n7620 ^ n1733 ;
  assign n15091 = n15090 ^ n15089 ^ n3203 ;
  assign n15092 = ( ~n7277 & n9856 ) | ( ~n7277 & n9966 ) | ( n9856 & n9966 ) ;
  assign n15093 = ( ~n788 & n3399 ) | ( ~n788 & n12904 ) | ( n3399 & n12904 ) ;
  assign n15097 = ( x8 & n1881 ) | ( x8 & n10054 ) | ( n1881 & n10054 ) ;
  assign n15094 = ( n1920 & n5722 ) | ( n1920 & n7884 ) | ( n5722 & n7884 ) ;
  assign n15095 = n15094 ^ n10744 ^ n2845 ;
  assign n15096 = n15095 ^ n12215 ^ n5068 ;
  assign n15098 = n15097 ^ n15096 ^ n4689 ;
  assign n15099 = ( n5074 & n11016 ) | ( n5074 & n15098 ) | ( n11016 & n15098 ) ;
  assign n15100 = ( ~n3384 & n7144 ) | ( ~n3384 & n12046 ) | ( n7144 & n12046 ) ;
  assign n15101 = n15100 ^ n14289 ^ n6133 ;
  assign n15102 = n8432 ^ n3625 ^ n1002 ;
  assign n15103 = ( n405 & n2995 ) | ( n405 & n7180 ) | ( n2995 & n7180 ) ;
  assign n15104 = ( n5900 & n15102 ) | ( n5900 & n15103 ) | ( n15102 & n15103 ) ;
  assign n15105 = n15104 ^ n7426 ^ n1041 ;
  assign n15106 = n11371 ^ n9791 ^ n5685 ;
  assign n15107 = n15106 ^ n13152 ^ n11443 ;
  assign n15108 = n15107 ^ n11866 ^ n5841 ;
  assign n15109 = ( ~n3416 & n6274 ) | ( ~n3416 & n7517 ) | ( n6274 & n7517 ) ;
  assign n15110 = n4993 ^ n3448 ^ n645 ;
  assign n15111 = ( n8328 & n14285 ) | ( n8328 & n15110 ) | ( n14285 & n15110 ) ;
  assign n15112 = ( n1845 & n2032 ) | ( n1845 & n3425 ) | ( n2032 & n3425 ) ;
  assign n15113 = n15112 ^ n1142 ^ n895 ;
  assign n15114 = n15113 ^ n2303 ^ n697 ;
  assign n15118 = ( n2488 & n10126 ) | ( n2488 & ~n13807 ) | ( n10126 & ~n13807 ) ;
  assign n15119 = ( n4431 & ~n11092 ) | ( n4431 & n15118 ) | ( ~n11092 & n15118 ) ;
  assign n15120 = n15119 ^ n7008 ^ n5346 ;
  assign n15117 = n8837 ^ n4011 ^ n934 ;
  assign n15115 = ( n3928 & ~n8634 ) | ( n3928 & n11290 ) | ( ~n8634 & n11290 ) ;
  assign n15116 = n15115 ^ n12542 ^ n11191 ;
  assign n15121 = n15120 ^ n15117 ^ n15116 ;
  assign n15122 = ( n5401 & n15114 ) | ( n5401 & ~n15121 ) | ( n15114 & ~n15121 ) ;
  assign n15123 = n13265 ^ n6463 ^ n4996 ;
  assign n15124 = n15123 ^ n6766 ^ n3774 ;
  assign n15125 = ( ~n7979 & n8361 ) | ( ~n7979 & n11823 ) | ( n8361 & n11823 ) ;
  assign n15126 = n15125 ^ n8427 ^ n6997 ;
  assign n15127 = n15126 ^ n7799 ^ n3297 ;
  assign n15128 = n9539 ^ n2887 ^ n1747 ;
  assign n15129 = ( ~n1940 & n12833 ) | ( ~n1940 & n15128 ) | ( n12833 & n15128 ) ;
  assign n15134 = n6032 ^ n3715 ^ n400 ;
  assign n15135 = n15134 ^ n12058 ^ n3249 ;
  assign n15130 = n6483 ^ n2009 ^ n1931 ;
  assign n15131 = n15130 ^ n6150 ^ n4413 ;
  assign n15132 = n15131 ^ n6141 ^ n1123 ;
  assign n15133 = n15132 ^ n6431 ^ n3706 ;
  assign n15136 = n15135 ^ n15133 ^ n9067 ;
  assign n15137 = n11648 ^ n7544 ^ n3263 ;
  assign n15138 = ( n278 & ~n8972 ) | ( n278 & n15137 ) | ( ~n8972 & n15137 ) ;
  assign n15139 = ( n5725 & n6396 ) | ( n5725 & ~n13741 ) | ( n6396 & ~n13741 ) ;
  assign n15140 = ( n180 & n11720 ) | ( n180 & n15139 ) | ( n11720 & n15139 ) ;
  assign n15143 = ( n1312 & n1505 ) | ( n1312 & ~n7174 ) | ( n1505 & ~n7174 ) ;
  assign n15141 = ( n3430 & n3840 ) | ( n3430 & ~n6880 ) | ( n3840 & ~n6880 ) ;
  assign n15142 = n15141 ^ n3041 ^ n1481 ;
  assign n15144 = n15143 ^ n15142 ^ n2865 ;
  assign n15145 = n15144 ^ n10276 ^ n3932 ;
  assign n15146 = n7940 ^ n4259 ^ n3632 ;
  assign n15149 = ( n6995 & n7199 ) | ( n6995 & n10291 ) | ( n7199 & n10291 ) ;
  assign n15148 = n7475 ^ n4758 ^ n2076 ;
  assign n15147 = n8098 ^ n6069 ^ n4641 ;
  assign n15150 = n15149 ^ n15148 ^ n15147 ;
  assign n15157 = ( n389 & ~n4233 ) | ( n389 & n9174 ) | ( ~n4233 & n9174 ) ;
  assign n15151 = ( n548 & n1407 ) | ( n548 & ~n2872 ) | ( n1407 & ~n2872 ) ;
  assign n15154 = n7811 ^ n7529 ^ n4644 ;
  assign n15152 = ( n493 & n6715 ) | ( n493 & n10605 ) | ( n6715 & n10605 ) ;
  assign n15153 = ( n2842 & n5718 ) | ( n2842 & ~n15152 ) | ( n5718 & ~n15152 ) ;
  assign n15155 = n15154 ^ n15153 ^ n4119 ;
  assign n15156 = ( ~n3906 & n15151 ) | ( ~n3906 & n15155 ) | ( n15151 & n15155 ) ;
  assign n15158 = n15157 ^ n15156 ^ n387 ;
  assign n15159 = ( n569 & ~n1087 ) | ( n569 & n7250 ) | ( ~n1087 & n7250 ) ;
  assign n15160 = n15159 ^ n10778 ^ n592 ;
  assign n15161 = n10809 ^ n7426 ^ n416 ;
  assign n15162 = ( ~n3421 & n10063 ) | ( ~n3421 & n15161 ) | ( n10063 & n15161 ) ;
  assign n15163 = n15162 ^ n12187 ^ n7040 ;
  assign n15164 = ( n1267 & n3909 ) | ( n1267 & ~n6263 ) | ( n3909 & ~n6263 ) ;
  assign n15165 = n15164 ^ n1512 ^ n1113 ;
  assign n15166 = ( n7401 & n10908 ) | ( n7401 & ~n12682 ) | ( n10908 & ~n12682 ) ;
  assign n15167 = ( n6111 & ~n10731 ) | ( n6111 & n15166 ) | ( ~n10731 & n15166 ) ;
  assign n15168 = n15167 ^ n4832 ^ n383 ;
  assign n15169 = ( ~n1788 & n3501 ) | ( ~n1788 & n15168 ) | ( n3501 & n15168 ) ;
  assign n15170 = n15169 ^ n7287 ^ n3756 ;
  assign n15171 = ( n6834 & n14559 ) | ( n6834 & n14995 ) | ( n14559 & n14995 ) ;
  assign n15172 = ( n1309 & n2193 ) | ( n1309 & ~n4218 ) | ( n2193 & ~n4218 ) ;
  assign n15173 = n15172 ^ n10287 ^ n1695 ;
  assign n15174 = ( ~n9195 & n12768 ) | ( ~n9195 & n14232 ) | ( n12768 & n14232 ) ;
  assign n15175 = ( n4605 & ~n15173 ) | ( n4605 & n15174 ) | ( ~n15173 & n15174 ) ;
  assign n15176 = n15175 ^ n1565 ^ n1347 ;
  assign n15177 = n7359 ^ n4228 ^ n286 ;
  assign n15178 = ( ~n419 & n11439 ) | ( ~n419 & n15177 ) | ( n11439 & n15177 ) ;
  assign n15179 = n8290 ^ n585 ^ n479 ;
  assign n15180 = ( n6584 & ~n14976 ) | ( n6584 & n15179 ) | ( ~n14976 & n15179 ) ;
  assign n15181 = n15180 ^ n2152 ^ n1957 ;
  assign n15182 = ( n4588 & n6516 ) | ( n4588 & ~n8959 ) | ( n6516 & ~n8959 ) ;
  assign n15183 = ( n336 & n2991 ) | ( n336 & n6657 ) | ( n2991 & n6657 ) ;
  assign n15184 = ( ~n2610 & n14042 ) | ( ~n2610 & n15183 ) | ( n14042 & n15183 ) ;
  assign n15185 = ( n601 & n15182 ) | ( n601 & ~n15184 ) | ( n15182 & ~n15184 ) ;
  assign n15186 = ( ~x102 & n1877 ) | ( ~x102 & n6657 ) | ( n1877 & n6657 ) ;
  assign n15193 = ( n564 & n726 ) | ( n564 & ~n10087 ) | ( n726 & ~n10087 ) ;
  assign n15190 = n11876 ^ n7574 ^ n332 ;
  assign n15191 = ( n1562 & n1931 ) | ( n1562 & n5592 ) | ( n1931 & n5592 ) ;
  assign n15192 = ( n5217 & n15190 ) | ( n5217 & ~n15191 ) | ( n15190 & ~n15191 ) ;
  assign n15187 = ( n8574 & n12680 ) | ( n8574 & ~n12968 ) | ( n12680 & ~n12968 ) ;
  assign n15188 = ( ~n5176 & n11546 ) | ( ~n5176 & n15187 ) | ( n11546 & n15187 ) ;
  assign n15189 = ( ~n10986 & n11382 ) | ( ~n10986 & n15188 ) | ( n11382 & n15188 ) ;
  assign n15194 = n15193 ^ n15192 ^ n15189 ;
  assign n15195 = ( n1349 & n15186 ) | ( n1349 & ~n15194 ) | ( n15186 & ~n15194 ) ;
  assign n15196 = n15195 ^ n7726 ^ n1887 ;
  assign n15206 = ( n889 & n3432 ) | ( n889 & ~n10578 ) | ( n3432 & ~n10578 ) ;
  assign n15207 = n7688 ^ n815 ^ n571 ;
  assign n15208 = ( n8831 & n13939 ) | ( n8831 & ~n15207 ) | ( n13939 & ~n15207 ) ;
  assign n15209 = ( ~n8878 & n15206 ) | ( ~n8878 & n15208 ) | ( n15206 & n15208 ) ;
  assign n15203 = ( ~n920 & n3857 ) | ( ~n920 & n9725 ) | ( n3857 & n9725 ) ;
  assign n15201 = n5432 ^ n362 ^ x98 ;
  assign n15202 = n15201 ^ n10875 ^ n9476 ;
  assign n15204 = n15203 ^ n15202 ^ n13690 ;
  assign n15197 = n6648 ^ n5549 ^ n3372 ;
  assign n15198 = n15197 ^ n8008 ^ n138 ;
  assign n15199 = n15198 ^ n10808 ^ n7301 ;
  assign n15200 = ( n698 & ~n3069 ) | ( n698 & n15199 ) | ( ~n3069 & n15199 ) ;
  assign n15205 = n15204 ^ n15200 ^ n6846 ;
  assign n15210 = n15209 ^ n15205 ^ n2839 ;
  assign n15216 = n10668 ^ n5462 ^ n2927 ;
  assign n15211 = ( n2342 & n2449 ) | ( n2342 & ~n11153 ) | ( n2449 & ~n11153 ) ;
  assign n15212 = ( n3543 & n9567 ) | ( n3543 & n14451 ) | ( n9567 & n14451 ) ;
  assign n15213 = ( n995 & n4660 ) | ( n995 & n15212 ) | ( n4660 & n15212 ) ;
  assign n15214 = ( n3670 & ~n14917 ) | ( n3670 & n15213 ) | ( ~n14917 & n15213 ) ;
  assign n15215 = ( n13171 & n15211 ) | ( n13171 & ~n15214 ) | ( n15211 & ~n15214 ) ;
  assign n15217 = n15216 ^ n15215 ^ n347 ;
  assign n15219 = ( n5260 & ~n11740 ) | ( n5260 & n13818 ) | ( ~n11740 & n13818 ) ;
  assign n15220 = n15219 ^ n11498 ^ n239 ;
  assign n15218 = ( ~n6814 & n7618 ) | ( ~n6814 & n14460 ) | ( n7618 & n14460 ) ;
  assign n15221 = n15220 ^ n15218 ^ n15137 ;
  assign n15222 = ( n308 & n1486 ) | ( n308 & n3154 ) | ( n1486 & n3154 ) ;
  assign n15223 = ( ~n4480 & n14522 ) | ( ~n4480 & n15222 ) | ( n14522 & n15222 ) ;
  assign n15224 = n15223 ^ n11283 ^ n8465 ;
  assign n15225 = ( n2603 & ~n9130 ) | ( n2603 & n9629 ) | ( ~n9130 & n9629 ) ;
  assign n15226 = n10739 ^ n9930 ^ n8351 ;
  assign n15227 = n15226 ^ n10063 ^ n1196 ;
  assign n15228 = n6147 ^ n4215 ^ x119 ;
  assign n15229 = ( n270 & n7577 ) | ( n270 & n7868 ) | ( n7577 & n7868 ) ;
  assign n15230 = ( n12326 & n15228 ) | ( n12326 & ~n15229 ) | ( n15228 & ~n15229 ) ;
  assign n15231 = ( n1276 & n14334 ) | ( n1276 & n15230 ) | ( n14334 & n15230 ) ;
  assign n15232 = ( n3265 & n3555 ) | ( n3265 & ~n11423 ) | ( n3555 & ~n11423 ) ;
  assign n15233 = ( ~n3600 & n4266 ) | ( ~n3600 & n15232 ) | ( n4266 & n15232 ) ;
  assign n15234 = ( n4795 & ~n10680 ) | ( n4795 & n15233 ) | ( ~n10680 & n15233 ) ;
  assign n15235 = ( n5510 & n10478 ) | ( n5510 & ~n15234 ) | ( n10478 & ~n15234 ) ;
  assign n15236 = n361 ^ n258 ^ n190 ;
  assign n15237 = n15236 ^ n7289 ^ n7231 ;
  assign n15238 = ( ~n1044 & n7607 ) | ( ~n1044 & n9387 ) | ( n7607 & n9387 ) ;
  assign n15239 = n15238 ^ n5701 ^ n2658 ;
  assign n15240 = n2894 ^ n2226 ^ n866 ;
  assign n15241 = n15240 ^ n11945 ^ n9791 ;
  assign n15242 = n15241 ^ n11828 ^ n3187 ;
  assign n15243 = ( ~n14508 & n15239 ) | ( ~n14508 & n15242 ) | ( n15239 & n15242 ) ;
  assign n15244 = ( n1965 & ~n4966 ) | ( n1965 & n7174 ) | ( ~n4966 & n7174 ) ;
  assign n15245 = ( n8118 & n14995 ) | ( n8118 & ~n15244 ) | ( n14995 & ~n15244 ) ;
  assign n15246 = ( n9282 & n12447 ) | ( n9282 & ~n15245 ) | ( n12447 & ~n15245 ) ;
  assign n15247 = n15246 ^ n12568 ^ n10887 ;
  assign n15248 = n9141 ^ n4419 ^ n3547 ;
  assign n15249 = ( n2648 & ~n5113 ) | ( n2648 & n8795 ) | ( ~n5113 & n8795 ) ;
  assign n15250 = ( n7769 & n15248 ) | ( n7769 & ~n15249 ) | ( n15248 & ~n15249 ) ;
  assign n15251 = n15250 ^ n10247 ^ n4492 ;
  assign n15252 = n15251 ^ n13962 ^ n7378 ;
  assign n15253 = n5881 ^ n4506 ^ n3699 ;
  assign n15254 = ( n6622 & n8208 ) | ( n6622 & ~n11789 ) | ( n8208 & ~n11789 ) ;
  assign n15255 = n15254 ^ n13667 ^ n7874 ;
  assign n15256 = n15255 ^ n11720 ^ n7781 ;
  assign n15257 = ( n4663 & n15253 ) | ( n4663 & n15256 ) | ( n15253 & n15256 ) ;
  assign n15258 = ( n1837 & n4251 ) | ( n1837 & n11887 ) | ( n4251 & n11887 ) ;
  assign n15260 = ( n1063 & ~n1623 ) | ( n1063 & n2357 ) | ( ~n1623 & n2357 ) ;
  assign n15261 = n15260 ^ n6338 ^ n6055 ;
  assign n15259 = ( ~n3165 & n4063 ) | ( ~n3165 & n8298 ) | ( n4063 & n8298 ) ;
  assign n15262 = n15261 ^ n15259 ^ n6397 ;
  assign n15264 = n3649 ^ n2819 ^ n1698 ;
  assign n15265 = n15264 ^ n6918 ^ n2614 ;
  assign n15266 = n15265 ^ n9795 ^ n1001 ;
  assign n15263 = n4059 ^ n3503 ^ n2736 ;
  assign n15267 = n15266 ^ n15263 ^ n4919 ;
  assign n15268 = ( n2747 & n4741 ) | ( n2747 & ~n8842 ) | ( n4741 & ~n8842 ) ;
  assign n15269 = n15268 ^ n7801 ^ n1012 ;
  assign n15270 = n15269 ^ n2236 ^ n588 ;
  assign n15271 = n12544 ^ n4255 ^ n3841 ;
  assign n15272 = ( ~n5943 & n6262 ) | ( ~n5943 & n15271 ) | ( n6262 & n15271 ) ;
  assign n15273 = n15272 ^ n10662 ^ n3324 ;
  assign n15274 = n15273 ^ n6694 ^ n1489 ;
  assign n15275 = ( n1245 & ~n6704 ) | ( n1245 & n15274 ) | ( ~n6704 & n15274 ) ;
  assign n15276 = ( x45 & n1677 ) | ( x45 & ~n15275 ) | ( n1677 & ~n15275 ) ;
  assign n15278 = ( ~n1425 & n2108 ) | ( ~n1425 & n11501 ) | ( n2108 & n11501 ) ;
  assign n15277 = n8727 ^ n5883 ^ n2958 ;
  assign n15279 = n15278 ^ n15277 ^ n12457 ;
  assign n15280 = ( n9204 & ~n9514 ) | ( n9204 & n15279 ) | ( ~n9514 & n15279 ) ;
  assign n15282 = ( ~n694 & n10800 ) | ( ~n694 & n12942 ) | ( n10800 & n12942 ) ;
  assign n15283 = n7831 ^ n4447 ^ n1576 ;
  assign n15284 = n15283 ^ x88 ^ x76 ;
  assign n15285 = ( n14197 & ~n15282 ) | ( n14197 & n15284 ) | ( ~n15282 & n15284 ) ;
  assign n15281 = n13138 ^ n8743 ^ n7717 ;
  assign n15286 = n15285 ^ n15281 ^ n7488 ;
  assign n15289 = ( n585 & n5903 ) | ( n585 & n10065 ) | ( n5903 & n10065 ) ;
  assign n15287 = ( n4064 & n5476 ) | ( n4064 & ~n15260 ) | ( n5476 & ~n15260 ) ;
  assign n15288 = ( n4742 & n5126 ) | ( n4742 & ~n15287 ) | ( n5126 & ~n15287 ) ;
  assign n15290 = n15289 ^ n15288 ^ n1521 ;
  assign n15296 = n6801 ^ n1401 ^ n315 ;
  assign n15294 = n2798 ^ n1653 ^ x36 ;
  assign n15295 = n15294 ^ n1981 ^ n1271 ;
  assign n15291 = n7666 ^ n4121 ^ n815 ;
  assign n15292 = ( n2151 & ~n8690 ) | ( n2151 & n14298 ) | ( ~n8690 & n14298 ) ;
  assign n15293 = ( n11653 & ~n15291 ) | ( n11653 & n15292 ) | ( ~n15291 & n15292 ) ;
  assign n15297 = n15296 ^ n15295 ^ n15293 ;
  assign n15298 = n15297 ^ n2660 ^ n575 ;
  assign n15299 = n15298 ^ n11248 ^ n2575 ;
  assign n15300 = n9789 ^ n6165 ^ n3968 ;
  assign n15301 = n15300 ^ n3950 ^ n3813 ;
  assign n15302 = ( n2731 & n3119 ) | ( n2731 & n15301 ) | ( n3119 & n15301 ) ;
  assign n15308 = n5116 ^ n3022 ^ n658 ;
  assign n15303 = n8410 ^ n6417 ^ n4300 ;
  assign n15304 = ( n4664 & n6563 ) | ( n4664 & n15303 ) | ( n6563 & n15303 ) ;
  assign n15305 = ( ~n11919 & n13670 ) | ( ~n11919 & n13927 ) | ( n13670 & n13927 ) ;
  assign n15306 = n15305 ^ n9102 ^ n5006 ;
  assign n15307 = ( n11572 & ~n15304 ) | ( n11572 & n15306 ) | ( ~n15304 & n15306 ) ;
  assign n15309 = n15308 ^ n15307 ^ n10676 ;
  assign n15310 = ( n3025 & n3873 ) | ( n3025 & n6244 ) | ( n3873 & n6244 ) ;
  assign n15311 = n15310 ^ n14613 ^ n14264 ;
  assign n15313 = n14981 ^ n1293 ^ n1226 ;
  assign n15312 = ( n1334 & n1379 ) | ( n1334 & n10874 ) | ( n1379 & n10874 ) ;
  assign n15314 = n15313 ^ n15312 ^ n5106 ;
  assign n15315 = ( ~n2521 & n5951 ) | ( ~n2521 & n11769 ) | ( n5951 & n11769 ) ;
  assign n15316 = n9754 ^ n7384 ^ n2194 ;
  assign n15317 = ( ~n2442 & n3943 ) | ( ~n2442 & n14460 ) | ( n3943 & n14460 ) ;
  assign n15318 = n15317 ^ n11681 ^ n6720 ;
  assign n15319 = ( n5644 & n15316 ) | ( n5644 & n15318 ) | ( n15316 & n15318 ) ;
  assign n15321 = ( ~x68 & n1661 ) | ( ~x68 & n10326 ) | ( n1661 & n10326 ) ;
  assign n15322 = n15321 ^ n10259 ^ n6809 ;
  assign n15320 = n9833 ^ n3700 ^ n3670 ;
  assign n15323 = n15322 ^ n15320 ^ n275 ;
  assign n15324 = n15323 ^ n6546 ^ n4624 ;
  assign n15325 = ( n4357 & ~n12182 ) | ( n4357 & n13069 ) | ( ~n12182 & n13069 ) ;
  assign n15326 = n2686 ^ n1509 ^ n504 ;
  assign n15327 = ( n714 & n5345 ) | ( n714 & ~n15326 ) | ( n5345 & ~n15326 ) ;
  assign n15328 = n12959 ^ n4678 ^ n1853 ;
  assign n15329 = ( n1799 & ~n2497 ) | ( n1799 & n15328 ) | ( ~n2497 & n15328 ) ;
  assign n15330 = ( n6275 & n11384 ) | ( n6275 & ~n15137 ) | ( n11384 & ~n15137 ) ;
  assign n15331 = ( n5740 & n7646 ) | ( n5740 & n8972 ) | ( n7646 & n8972 ) ;
  assign n15332 = ( n5644 & n5737 ) | ( n5644 & n6868 ) | ( n5737 & n6868 ) ;
  assign n15333 = ( ~n807 & n3605 ) | ( ~n807 & n12581 ) | ( n3605 & n12581 ) ;
  assign n15334 = n15333 ^ n4554 ^ n1182 ;
  assign n15335 = ( n440 & n4150 ) | ( n440 & n15334 ) | ( n4150 & n15334 ) ;
  assign n15336 = n13634 ^ n1898 ^ n486 ;
  assign n15337 = ( n3561 & ~n7318 ) | ( n3561 & n15336 ) | ( ~n7318 & n15336 ) ;
  assign n15338 = n13710 ^ n1547 ^ x93 ;
  assign n15339 = ( n7004 & n7986 ) | ( n7004 & n15338 ) | ( n7986 & n15338 ) ;
  assign n15340 = ( n6645 & n15337 ) | ( n6645 & ~n15339 ) | ( n15337 & ~n15339 ) ;
  assign n15341 = n13045 ^ n12728 ^ n6986 ;
  assign n15342 = n15341 ^ n6901 ^ n1286 ;
  assign n15343 = n15342 ^ n9811 ^ n1225 ;
  assign n15344 = n15343 ^ n12340 ^ n1614 ;
  assign n15347 = ( n461 & n1624 ) | ( n461 & ~n9710 ) | ( n1624 & ~n9710 ) ;
  assign n15345 = n15154 ^ n9073 ^ n2837 ;
  assign n15346 = ( n1756 & n11993 ) | ( n1756 & ~n15345 ) | ( n11993 & ~n15345 ) ;
  assign n15348 = n15347 ^ n15346 ^ n14058 ;
  assign n15349 = ( n6862 & n9436 ) | ( n6862 & n15348 ) | ( n9436 & n15348 ) ;
  assign n15350 = ( n8610 & ~n12089 ) | ( n8610 & n14006 ) | ( ~n12089 & n14006 ) ;
  assign n15351 = ( ~n9778 & n12350 ) | ( ~n9778 & n15350 ) | ( n12350 & n15350 ) ;
  assign n15352 = ( n1332 & n11196 ) | ( n1332 & n15351 ) | ( n11196 & n15351 ) ;
  assign n15353 = ( n6553 & n7382 ) | ( n6553 & n8194 ) | ( n7382 & n8194 ) ;
  assign n15354 = ( n6669 & n7919 ) | ( n6669 & ~n15353 ) | ( n7919 & ~n15353 ) ;
  assign n15355 = n9176 ^ n5030 ^ x104 ;
  assign n15356 = n15355 ^ n5010 ^ n2428 ;
  assign n15357 = n15356 ^ n9304 ^ n573 ;
  assign n15362 = n12121 ^ n7569 ^ n4037 ;
  assign n15358 = n5343 ^ n4931 ^ n2606 ;
  assign n15359 = n15358 ^ n4806 ^ n1843 ;
  assign n15360 = ( ~n13301 & n15316 ) | ( ~n13301 & n15359 ) | ( n15316 & n15359 ) ;
  assign n15361 = n15360 ^ n3131 ^ n2519 ;
  assign n15363 = n15362 ^ n15361 ^ n14288 ;
  assign n15365 = n8898 ^ n5975 ^ n2093 ;
  assign n15364 = ( ~n2637 & n3463 ) | ( ~n2637 & n5278 ) | ( n3463 & n5278 ) ;
  assign n15366 = n15365 ^ n15364 ^ n3944 ;
  assign n15368 = n15236 ^ n14562 ^ n399 ;
  assign n15367 = n12004 ^ n6254 ^ n991 ;
  assign n15369 = n15368 ^ n15367 ^ n8860 ;
  assign n15370 = ( n4799 & n6601 ) | ( n4799 & n11161 ) | ( n6601 & n11161 ) ;
  assign n15371 = ( n6581 & n7211 ) | ( n6581 & ~n11758 ) | ( n7211 & ~n11758 ) ;
  assign n15372 = n15371 ^ n7596 ^ n2518 ;
  assign n15373 = ( ~n463 & n1417 ) | ( ~n463 & n15372 ) | ( n1417 & n15372 ) ;
  assign n15374 = ( ~x10 & n9833 ) | ( ~x10 & n15373 ) | ( n9833 & n15373 ) ;
  assign n15379 = n4743 ^ n4202 ^ n2154 ;
  assign n15376 = ( n6703 & n7577 ) | ( n6703 & ~n13831 ) | ( n7577 & ~n13831 ) ;
  assign n15377 = n15376 ^ n4061 ^ n869 ;
  assign n15378 = ( n9720 & n12444 ) | ( n9720 & ~n15377 ) | ( n12444 & ~n15377 ) ;
  assign n15375 = n4949 ^ n4407 ^ n3943 ;
  assign n15380 = n15379 ^ n15378 ^ n15375 ;
  assign n15381 = ( n784 & n2955 ) | ( n784 & ~n7493 ) | ( n2955 & ~n7493 ) ;
  assign n15382 = n15381 ^ n14820 ^ n3674 ;
  assign n15383 = ( ~n4861 & n8488 ) | ( ~n4861 & n8749 ) | ( n8488 & n8749 ) ;
  assign n15384 = ( n3878 & ~n5743 ) | ( n3878 & n15383 ) | ( ~n5743 & n15383 ) ;
  assign n15385 = n15384 ^ n11513 ^ n600 ;
  assign n15386 = ( n11152 & ~n15382 ) | ( n11152 & n15385 ) | ( ~n15382 & n15385 ) ;
  assign n15388 = n15207 ^ n1372 ^ n1065 ;
  assign n15387 = ( n2106 & n5504 ) | ( n2106 & ~n7132 ) | ( n5504 & ~n7132 ) ;
  assign n15389 = n15388 ^ n15387 ^ n1884 ;
  assign n15390 = n10212 ^ n4608 ^ n3883 ;
  assign n15391 = ( n384 & n9610 ) | ( n384 & n15390 ) | ( n9610 & n15390 ) ;
  assign n15392 = ( n411 & n1992 ) | ( n411 & n11570 ) | ( n1992 & n11570 ) ;
  assign n15393 = ( n14353 & ~n15391 ) | ( n14353 & n15392 ) | ( ~n15391 & n15392 ) ;
  assign n15394 = n15393 ^ n9862 ^ n166 ;
  assign n15398 = ( n679 & n2882 ) | ( n679 & ~n6547 ) | ( n2882 & ~n6547 ) ;
  assign n15395 = n11479 ^ n7272 ^ n6256 ;
  assign n15396 = ( n9651 & n12274 ) | ( n9651 & ~n15395 ) | ( n12274 & ~n15395 ) ;
  assign n15397 = n15396 ^ n14034 ^ n1660 ;
  assign n15399 = n15398 ^ n15397 ^ n8288 ;
  assign n15400 = n15399 ^ n8347 ^ n1278 ;
  assign n15401 = n9190 ^ n723 ^ x50 ;
  assign n15402 = n15401 ^ n5320 ^ n2294 ;
  assign n15403 = n15402 ^ n11586 ^ n3281 ;
  assign n15404 = n15360 ^ n14324 ^ n3416 ;
  assign n15405 = n2244 ^ n1380 ^ x27 ;
  assign n15406 = n15405 ^ n8064 ^ n2694 ;
  assign n15407 = ( n4583 & n7743 ) | ( n4583 & ~n15406 ) | ( n7743 & ~n15406 ) ;
  assign n15408 = n15407 ^ n12491 ^ n3675 ;
  assign n15409 = n14009 ^ n6617 ^ n3964 ;
  assign n15410 = ( n5832 & ~n10911 ) | ( n5832 & n14581 ) | ( ~n10911 & n14581 ) ;
  assign n15413 = ( n2874 & n4217 ) | ( n2874 & ~n4958 ) | ( n4217 & ~n4958 ) ;
  assign n15411 = n9115 ^ n6609 ^ n1967 ;
  assign n15412 = ( n10031 & n11538 ) | ( n10031 & ~n15411 ) | ( n11538 & ~n15411 ) ;
  assign n15414 = n15413 ^ n15412 ^ n3321 ;
  assign n15415 = n5285 ^ n4812 ^ n3494 ;
  assign n15416 = n11195 ^ n7770 ^ n532 ;
  assign n15417 = ( n3632 & n6522 ) | ( n3632 & n15416 ) | ( n6522 & n15416 ) ;
  assign n15418 = ( n4561 & n8195 ) | ( n4561 & ~n15417 ) | ( n8195 & ~n15417 ) ;
  assign n15419 = n15418 ^ n10254 ^ x121 ;
  assign n15420 = n11049 ^ n7375 ^ n6131 ;
  assign n15421 = ( n8267 & ~n8544 ) | ( n8267 & n9775 ) | ( ~n8544 & n9775 ) ;
  assign n15422 = ( ~n3957 & n10266 ) | ( ~n3957 & n15421 ) | ( n10266 & n15421 ) ;
  assign n15423 = n15422 ^ n13566 ^ n1727 ;
  assign n15424 = ( n6701 & ~n15420 ) | ( n6701 & n15423 ) | ( ~n15420 & n15423 ) ;
  assign n15425 = ( n15415 & ~n15419 ) | ( n15415 & n15424 ) | ( ~n15419 & n15424 ) ;
  assign n15426 = ( n9602 & ~n10202 ) | ( n9602 & n10966 ) | ( ~n10202 & n10966 ) ;
  assign n15427 = n14627 ^ n4327 ^ n2045 ;
  assign n15428 = n12826 ^ n5424 ^ n1063 ;
  assign n15429 = ( ~n2861 & n9786 ) | ( ~n2861 & n10278 ) | ( n9786 & n10278 ) ;
  assign n15430 = ( n9332 & n10298 ) | ( n9332 & ~n15429 ) | ( n10298 & ~n15429 ) ;
  assign n15431 = ( n3913 & n7764 ) | ( n3913 & ~n11764 ) | ( n7764 & ~n11764 ) ;
  assign n15432 = ( x2 & n11570 ) | ( x2 & n15431 ) | ( n11570 & n15431 ) ;
  assign n15433 = ( ~n9087 & n12920 ) | ( ~n9087 & n15432 ) | ( n12920 & n15432 ) ;
  assign n15434 = n15433 ^ n7303 ^ n5275 ;
  assign n15444 = n13850 ^ n7678 ^ n4426 ;
  assign n15437 = n9198 ^ n3413 ^ n3401 ;
  assign n15438 = ( n8734 & ~n8836 ) | ( n8734 & n15437 ) | ( ~n8836 & n15437 ) ;
  assign n15439 = n3026 ^ n1471 ^ n1022 ;
  assign n15440 = ( n4530 & n10058 ) | ( n4530 & n15439 ) | ( n10058 & n15439 ) ;
  assign n15441 = n15440 ^ n6072 ^ n2278 ;
  assign n15442 = ( n6247 & n9003 ) | ( n6247 & ~n15441 ) | ( n9003 & ~n15441 ) ;
  assign n15443 = ( n4151 & n15438 ) | ( n4151 & ~n15442 ) | ( n15438 & ~n15442 ) ;
  assign n15445 = n15444 ^ n15443 ^ n4499 ;
  assign n15435 = ( n3910 & n4612 ) | ( n3910 & ~n5417 ) | ( n4612 & ~n5417 ) ;
  assign n15436 = n15435 ^ n15368 ^ n13536 ;
  assign n15446 = n15445 ^ n15436 ^ n3108 ;
  assign n15447 = ( n4067 & ~n5427 ) | ( n4067 & n14062 ) | ( ~n5427 & n14062 ) ;
  assign n15448 = n15447 ^ x85 ^ x16 ;
  assign n15451 = ( n2905 & ~n3395 ) | ( n2905 & n11371 ) | ( ~n3395 & n11371 ) ;
  assign n15452 = n12728 ^ n3703 ^ n3424 ;
  assign n15453 = ( n15266 & ~n15451 ) | ( n15266 & n15452 ) | ( ~n15451 & n15452 ) ;
  assign n15449 = n12986 ^ n10578 ^ n7912 ;
  assign n15450 = ( ~n10590 & n14069 ) | ( ~n10590 & n15449 ) | ( n14069 & n15449 ) ;
  assign n15454 = n15453 ^ n15450 ^ n11098 ;
  assign n15455 = n8045 ^ n6631 ^ n4555 ;
  assign n15456 = ( n2898 & n3345 ) | ( n2898 & ~n4269 ) | ( n3345 & ~n4269 ) ;
  assign n15457 = n15456 ^ n5552 ^ n2249 ;
  assign n15458 = ( n1465 & ~n4461 ) | ( n1465 & n5329 ) | ( ~n4461 & n5329 ) ;
  assign n15459 = n13232 ^ n4804 ^ n1002 ;
  assign n15460 = n10970 ^ n10699 ^ n9960 ;
  assign n15461 = ( n2019 & n11347 ) | ( n2019 & ~n15460 ) | ( n11347 & ~n15460 ) ;
  assign n15462 = ( ~n9069 & n15459 ) | ( ~n9069 & n15461 ) | ( n15459 & n15461 ) ;
  assign n15463 = n11355 ^ n10421 ^ n6088 ;
  assign n15464 = n11050 ^ n9988 ^ n2896 ;
  assign n15465 = n11587 ^ n5362 ^ n2348 ;
  assign n15466 = n15465 ^ n15381 ^ n6861 ;
  assign n15467 = ( ~n332 & n1033 ) | ( ~n332 & n9091 ) | ( n1033 & n9091 ) ;
  assign n15468 = ( n1185 & n8008 ) | ( n1185 & n14516 ) | ( n8008 & n14516 ) ;
  assign n15469 = ( ~n1565 & n1645 ) | ( ~n1565 & n15468 ) | ( n1645 & n15468 ) ;
  assign n15470 = n10852 ^ n4627 ^ n1140 ;
  assign n15471 = n15470 ^ n8075 ^ n2113 ;
  assign n15473 = ( n3219 & n6577 ) | ( n3219 & n8763 ) | ( n6577 & n8763 ) ;
  assign n15474 = ( n2627 & n13983 ) | ( n2627 & ~n15473 ) | ( n13983 & ~n15473 ) ;
  assign n15472 = ( ~n5482 & n6184 ) | ( ~n5482 & n7621 ) | ( n6184 & n7621 ) ;
  assign n15475 = n15474 ^ n15472 ^ n1655 ;
  assign n15478 = n7884 ^ n7549 ^ n2859 ;
  assign n15476 = ( ~n4618 & n9849 ) | ( ~n4618 & n10837 ) | ( n9849 & n10837 ) ;
  assign n15477 = n15476 ^ n4921 ^ n589 ;
  assign n15479 = n15478 ^ n15477 ^ n3284 ;
  assign n15480 = ( n256 & n2290 ) | ( n256 & ~n11634 ) | ( n2290 & ~n11634 ) ;
  assign n15481 = ( n2661 & n7162 ) | ( n2661 & ~n15480 ) | ( n7162 & ~n15480 ) ;
  assign n15482 = n15481 ^ n11785 ^ n2650 ;
  assign n15483 = ( n486 & ~n3001 ) | ( n486 & n9540 ) | ( ~n3001 & n9540 ) ;
  assign n15484 = ( ~n650 & n12601 ) | ( ~n650 & n15483 ) | ( n12601 & n15483 ) ;
  assign n15485 = n15484 ^ n9750 ^ n5950 ;
  assign n15486 = n8749 ^ n7016 ^ n6295 ;
  assign n15487 = ( n1411 & ~n2748 ) | ( n1411 & n15486 ) | ( ~n2748 & n15486 ) ;
  assign n15488 = n15487 ^ n9816 ^ n5662 ;
  assign n15489 = n14268 ^ n9223 ^ n616 ;
  assign n15490 = ( n2904 & n15159 ) | ( n2904 & n15489 ) | ( n15159 & n15489 ) ;
  assign n15491 = n15490 ^ n2455 ^ n2298 ;
  assign n15492 = ( n10912 & ~n12354 ) | ( n10912 & n15491 ) | ( ~n12354 & n15491 ) ;
  assign n15493 = ( n6239 & n15488 ) | ( n6239 & ~n15492 ) | ( n15488 & ~n15492 ) ;
  assign n15495 = n2182 ^ n863 ^ x101 ;
  assign n15494 = n3731 ^ n1740 ^ n1085 ;
  assign n15496 = n15495 ^ n15494 ^ n7336 ;
  assign n15497 = ( n8798 & ~n10025 ) | ( n8798 & n15496 ) | ( ~n10025 & n15496 ) ;
  assign n15505 = ( ~n1908 & n4853 ) | ( ~n1908 & n8008 ) | ( n4853 & n8008 ) ;
  assign n15506 = n15505 ^ n2399 ^ n1807 ;
  assign n15501 = n6713 ^ n4500 ^ n2559 ;
  assign n15499 = n1350 ^ n921 ^ n141 ;
  assign n15500 = ( n2185 & ~n10339 ) | ( n2185 & n15499 ) | ( ~n10339 & n15499 ) ;
  assign n15498 = ( ~n2636 & n3358 ) | ( ~n2636 & n11330 ) | ( n3358 & n11330 ) ;
  assign n15502 = n15501 ^ n15500 ^ n15498 ;
  assign n15503 = ( n4386 & ~n12716 ) | ( n4386 & n15502 ) | ( ~n12716 & n15502 ) ;
  assign n15504 = ( n442 & n10723 ) | ( n442 & n15503 ) | ( n10723 & n15503 ) ;
  assign n15507 = n15506 ^ n15504 ^ n1896 ;
  assign n15508 = ( n6686 & n9985 ) | ( n6686 & n12164 ) | ( n9985 & n12164 ) ;
  assign n15510 = n12352 ^ n5153 ^ n1178 ;
  assign n15509 = n5826 ^ n3995 ^ n2390 ;
  assign n15511 = n15510 ^ n15509 ^ n3630 ;
  assign n15512 = ( n1877 & ~n15508 ) | ( n1877 & n15511 ) | ( ~n15508 & n15511 ) ;
  assign n15513 = ( n264 & ~n7641 ) | ( n264 & n13008 ) | ( ~n7641 & n13008 ) ;
  assign n15514 = n15513 ^ n14063 ^ n1049 ;
  assign n15515 = ( n884 & ~n2797 ) | ( n884 & n11461 ) | ( ~n2797 & n11461 ) ;
  assign n15516 = n15515 ^ n6795 ^ x125 ;
  assign n15517 = ( n12405 & n15514 ) | ( n12405 & ~n15516 ) | ( n15514 & ~n15516 ) ;
  assign n15520 = n9564 ^ n7414 ^ n6646 ;
  assign n15519 = ( ~n2449 & n5683 ) | ( ~n2449 & n14391 ) | ( n5683 & n14391 ) ;
  assign n15521 = n15520 ^ n15519 ^ n11264 ;
  assign n15518 = n7184 ^ n6576 ^ n213 ;
  assign n15522 = n15521 ^ n15518 ^ n14801 ;
  assign n15523 = n8183 ^ n4406 ^ n1028 ;
  assign n15526 = ( n2673 & ~n6120 ) | ( n2673 & n10872 ) | ( ~n6120 & n10872 ) ;
  assign n15525 = n5889 ^ n4515 ^ n1191 ;
  assign n15524 = n14286 ^ n4860 ^ n3846 ;
  assign n15527 = n15526 ^ n15525 ^ n15524 ;
  assign n15528 = ( n558 & n3635 ) | ( n558 & n7394 ) | ( n3635 & n7394 ) ;
  assign n15529 = n10596 ^ n5303 ^ n2276 ;
  assign n15530 = n15529 ^ n8000 ^ x84 ;
  assign n15531 = n15530 ^ n10305 ^ n4785 ;
  assign n15532 = ( n1358 & n15528 ) | ( n1358 & ~n15531 ) | ( n15528 & ~n15531 ) ;
  assign n15533 = n6524 ^ n5974 ^ n3346 ;
  assign n15534 = n15533 ^ n11621 ^ n4976 ;
  assign n15535 = ( ~n2310 & n5671 ) | ( ~n2310 & n15534 ) | ( n5671 & n15534 ) ;
  assign n15536 = ( ~n15063 & n15277 ) | ( ~n15063 & n15535 ) | ( n15277 & n15535 ) ;
  assign n15537 = n9169 ^ n5103 ^ n3597 ;
  assign n15538 = n15537 ^ n15526 ^ n2108 ;
  assign n15539 = ( ~n6983 & n8936 ) | ( ~n6983 & n13592 ) | ( n8936 & n13592 ) ;
  assign n15541 = n12814 ^ n5313 ^ n1827 ;
  assign n15540 = ( ~n2115 & n9917 ) | ( ~n2115 & n10094 ) | ( n9917 & n10094 ) ;
  assign n15542 = n15541 ^ n15540 ^ n1572 ;
  assign n15543 = ( ~n9658 & n15539 ) | ( ~n9658 & n15542 ) | ( n15539 & n15542 ) ;
  assign n15544 = n12941 ^ n3139 ^ x2 ;
  assign n15545 = n15544 ^ n9668 ^ n5436 ;
  assign n15546 = n10697 ^ n7939 ^ n3496 ;
  assign n15547 = n15546 ^ n6016 ^ n3894 ;
  assign n15548 = n10923 ^ n10085 ^ n5482 ;
  assign n15549 = ( n1433 & n5411 ) | ( n1433 & ~n15179 ) | ( n5411 & ~n15179 ) ;
  assign n15550 = ( n6999 & n13564 ) | ( n6999 & n15549 ) | ( n13564 & n15549 ) ;
  assign n15551 = ( ~n12496 & n15548 ) | ( ~n12496 & n15550 ) | ( n15548 & n15550 ) ;
  assign n15552 = ( n11152 & n13036 ) | ( n11152 & ~n15379 ) | ( n13036 & ~n15379 ) ;
  assign n15553 = n7302 ^ n4631 ^ n1985 ;
  assign n15554 = n15553 ^ n9963 ^ n5122 ;
  assign n15555 = ( n5896 & n15552 ) | ( n5896 & ~n15554 ) | ( n15552 & ~n15554 ) ;
  assign n15556 = ( n2301 & ~n15551 ) | ( n2301 & n15555 ) | ( ~n15551 & n15555 ) ;
  assign n15557 = n7490 ^ n1273 ^ n853 ;
  assign n15558 = n8836 ^ n7449 ^ n226 ;
  assign n15559 = ( ~n1880 & n8703 ) | ( ~n1880 & n14542 ) | ( n8703 & n14542 ) ;
  assign n15560 = ( n951 & ~n6717 ) | ( n951 & n15559 ) | ( ~n6717 & n15559 ) ;
  assign n15561 = ( n5243 & n15558 ) | ( n5243 & n15560 ) | ( n15558 & n15560 ) ;
  assign n15562 = n15541 ^ n6322 ^ n6058 ;
  assign n15563 = n4417 ^ n2368 ^ n615 ;
  assign n15564 = ( ~n1793 & n8025 ) | ( ~n1793 & n15563 ) | ( n8025 & n15563 ) ;
  assign n15565 = n9993 ^ n9873 ^ n2634 ;
  assign n15566 = ( n3753 & n8747 ) | ( n3753 & ~n15565 ) | ( n8747 & ~n15565 ) ;
  assign n15567 = ( n370 & n2257 ) | ( n370 & n3687 ) | ( n2257 & n3687 ) ;
  assign n15568 = n15567 ^ n10735 ^ n4629 ;
  assign n15569 = ( ~x50 & n3754 ) | ( ~x50 & n15568 ) | ( n3754 & n15568 ) ;
  assign n15570 = ( n223 & n994 ) | ( n223 & ~n5798 ) | ( n994 & ~n5798 ) ;
  assign n15571 = ( n3464 & n4548 ) | ( n3464 & n15570 ) | ( n4548 & n15570 ) ;
  assign n15572 = n15571 ^ n6053 ^ n1214 ;
  assign n15575 = n13287 ^ n9259 ^ n608 ;
  assign n15573 = n1449 ^ n1399 ^ n691 ;
  assign n15574 = n15573 ^ n5174 ^ n4379 ;
  assign n15576 = n15575 ^ n15574 ^ n3063 ;
  assign n15577 = n15576 ^ n9519 ^ n329 ;
  assign n15578 = ( ~n3229 & n5445 ) | ( ~n3229 & n12774 ) | ( n5445 & n12774 ) ;
  assign n15579 = ( ~n3974 & n5607 ) | ( ~n3974 & n7829 ) | ( n5607 & n7829 ) ;
  assign n15580 = n15579 ^ n9785 ^ n9183 ;
  assign n15581 = ( n2886 & n15578 ) | ( n2886 & n15580 ) | ( n15578 & n15580 ) ;
  assign n15582 = n4577 ^ n2566 ^ n1166 ;
  assign n15583 = ( n2546 & n6711 ) | ( n2546 & n15582 ) | ( n6711 & n15582 ) ;
  assign n15584 = ( n834 & ~n5309 ) | ( n834 & n15583 ) | ( ~n5309 & n15583 ) ;
  assign n15587 = n4119 ^ n3416 ^ n1108 ;
  assign n15586 = ( n6786 & n7543 ) | ( n6786 & ~n7993 ) | ( n7543 & ~n7993 ) ;
  assign n15585 = n10804 ^ n8216 ^ n909 ;
  assign n15588 = n15587 ^ n15586 ^ n15585 ;
  assign n15589 = n11621 ^ n8817 ^ n4256 ;
  assign n15590 = n12583 ^ n5704 ^ n1433 ;
  assign n15591 = ( ~n10541 & n14930 ) | ( ~n10541 & n15590 ) | ( n14930 & n15590 ) ;
  assign n15592 = n9193 ^ n5699 ^ n188 ;
  assign n15593 = ( n1853 & n8618 ) | ( n1853 & ~n15592 ) | ( n8618 & ~n15592 ) ;
  assign n15595 = ( n2455 & n5001 ) | ( n2455 & n15023 ) | ( n5001 & n15023 ) ;
  assign n15594 = ( n1683 & ~n7118 ) | ( n1683 & n13039 ) | ( ~n7118 & n13039 ) ;
  assign n15596 = n15595 ^ n15594 ^ n6806 ;
  assign n15597 = n15413 ^ n9662 ^ n3276 ;
  assign n15598 = ( n2580 & n5439 ) | ( n2580 & ~n5700 ) | ( n5439 & ~n5700 ) ;
  assign n15599 = ( ~n6558 & n15597 ) | ( ~n6558 & n15598 ) | ( n15597 & n15598 ) ;
  assign n15600 = ( n1662 & n3570 ) | ( n1662 & ~n8814 ) | ( n3570 & ~n8814 ) ;
  assign n15601 = ( n246 & ~n2205 ) | ( n246 & n8464 ) | ( ~n2205 & n8464 ) ;
  assign n15602 = n15601 ^ n7884 ^ n4026 ;
  assign n15603 = ( n258 & n3289 ) | ( n258 & n11468 ) | ( n3289 & n11468 ) ;
  assign n15604 = ( ~n2864 & n8892 ) | ( ~n2864 & n15603 ) | ( n8892 & n15603 ) ;
  assign n15605 = ( n2801 & n9056 ) | ( n2801 & n15604 ) | ( n9056 & n15604 ) ;
  assign n15606 = n15605 ^ n11783 ^ n3856 ;
  assign n15607 = n15046 ^ n12639 ^ n9004 ;
  assign n15608 = ( ~n15602 & n15606 ) | ( ~n15602 & n15607 ) | ( n15606 & n15607 ) ;
  assign n15609 = n13722 ^ n8980 ^ n6586 ;
  assign n15610 = ( ~n1684 & n6703 ) | ( ~n1684 & n15609 ) | ( n6703 & n15609 ) ;
  assign n15611 = n14285 ^ n5687 ^ n854 ;
  assign n15613 = n8963 ^ n7642 ^ n5594 ;
  assign n15612 = ( n848 & n5048 ) | ( n848 & ~n5235 ) | ( n5048 & ~n5235 ) ;
  assign n15614 = n15613 ^ n15612 ^ n8225 ;
  assign n15615 = n15614 ^ n10167 ^ n7059 ;
  assign n15616 = n14595 ^ n6342 ^ n3518 ;
  assign n15617 = ( n1170 & n13797 ) | ( n1170 & ~n15616 ) | ( n13797 & ~n15616 ) ;
  assign n15618 = n15617 ^ n5477 ^ n1187 ;
  assign n15619 = ( n443 & n2296 ) | ( n443 & n15618 ) | ( n2296 & n15618 ) ;
  assign n15620 = ( ~n15611 & n15615 ) | ( ~n15611 & n15619 ) | ( n15615 & n15619 ) ;
  assign n15621 = n9063 ^ n5194 ^ n4770 ;
  assign n15622 = n15621 ^ n14966 ^ n8947 ;
  assign n15629 = n8896 ^ n7131 ^ n229 ;
  assign n15625 = n14667 ^ n6011 ^ n5070 ;
  assign n15626 = n15625 ^ n11038 ^ n2972 ;
  assign n15627 = n15626 ^ n10492 ^ n9403 ;
  assign n15624 = ( n1039 & n4894 ) | ( n1039 & n5027 ) | ( n4894 & n5027 ) ;
  assign n15628 = n15627 ^ n15624 ^ n8596 ;
  assign n15623 = n11805 ^ n5640 ^ n283 ;
  assign n15630 = n15629 ^ n15628 ^ n15623 ;
  assign n15631 = n15630 ^ n12754 ^ n12236 ;
  assign n15632 = n13379 ^ n11735 ^ n1974 ;
  assign n15633 = n8818 ^ n4324 ^ n2634 ;
  assign n15635 = ( n1762 & ~n2278 ) | ( n1762 & n11200 ) | ( ~n2278 & n11200 ) ;
  assign n15634 = ( ~n3937 & n6319 ) | ( ~n3937 & n11002 ) | ( n6319 & n11002 ) ;
  assign n15636 = n15635 ^ n15634 ^ n9957 ;
  assign n15637 = ( n4525 & ~n9731 ) | ( n4525 & n15636 ) | ( ~n9731 & n15636 ) ;
  assign n15641 = ( n1708 & n7312 ) | ( n1708 & ~n12998 ) | ( n7312 & ~n12998 ) ;
  assign n15638 = ( n3654 & n8327 ) | ( n3654 & n12784 ) | ( n8327 & n12784 ) ;
  assign n15639 = ( n7444 & n15510 ) | ( n7444 & n15638 ) | ( n15510 & n15638 ) ;
  assign n15640 = n15639 ^ n12371 ^ n654 ;
  assign n15642 = n15641 ^ n15640 ^ n9918 ;
  assign n15643 = n15642 ^ n15318 ^ n12350 ;
  assign n15644 = n6036 ^ n3715 ^ n817 ;
  assign n15645 = ( n2799 & n10606 ) | ( n2799 & n15644 ) | ( n10606 & n15644 ) ;
  assign n15646 = n15645 ^ n11432 ^ n4361 ;
  assign n15647 = n15646 ^ n5219 ^ n1152 ;
  assign n15648 = n14639 ^ n7396 ^ n226 ;
  assign n15649 = n15648 ^ n8884 ^ n6705 ;
  assign n15650 = ( ~n6309 & n13479 ) | ( ~n6309 & n15333 ) | ( n13479 & n15333 ) ;
  assign n15651 = n15650 ^ n14938 ^ n7454 ;
  assign n15652 = n819 ^ n742 ^ n254 ;
  assign n15653 = ( ~n4018 & n15253 ) | ( ~n4018 & n15652 ) | ( n15253 & n15652 ) ;
  assign n15654 = ( n5087 & n7942 ) | ( n5087 & ~n15653 ) | ( n7942 & ~n15653 ) ;
  assign n15657 = n10478 ^ n10287 ^ n8977 ;
  assign n15655 = ( ~n1510 & n4555 ) | ( ~n1510 & n6660 ) | ( n4555 & n6660 ) ;
  assign n15656 = ( ~n708 & n9556 ) | ( ~n708 & n15655 ) | ( n9556 & n15655 ) ;
  assign n15658 = n15657 ^ n15656 ^ n2091 ;
  assign n15671 = ( ~n1504 & n5335 ) | ( ~n1504 & n7557 ) | ( n5335 & n7557 ) ;
  assign n15672 = n15671 ^ n14020 ^ n5457 ;
  assign n15673 = ( n7263 & n10465 ) | ( n7263 & ~n15672 ) | ( n10465 & ~n15672 ) ;
  assign n15674 = n14959 ^ n14114 ^ n1857 ;
  assign n15675 = ( n7406 & n15673 ) | ( n7406 & n15674 ) | ( n15673 & n15674 ) ;
  assign n15661 = n3155 ^ n1924 ^ n828 ;
  assign n15659 = ( n2284 & n3821 ) | ( n2284 & ~n6410 ) | ( n3821 & ~n6410 ) ;
  assign n15660 = ( n7473 & ~n8922 ) | ( n7473 & n15659 ) | ( ~n8922 & n15659 ) ;
  assign n15662 = n15661 ^ n15660 ^ n423 ;
  assign n15663 = n14268 ^ n6340 ^ n4994 ;
  assign n15664 = n15663 ^ n4636 ^ n4117 ;
  assign n15665 = ( x57 & n4213 ) | ( x57 & n15664 ) | ( n4213 & n15664 ) ;
  assign n15666 = ( ~x9 & n3497 ) | ( ~x9 & n8378 ) | ( n3497 & n8378 ) ;
  assign n15667 = ( n777 & n5625 ) | ( n777 & ~n15666 ) | ( n5625 & ~n15666 ) ;
  assign n15668 = ( n15662 & n15665 ) | ( n15662 & ~n15667 ) | ( n15665 & ~n15667 ) ;
  assign n15669 = ( n5160 & n14924 ) | ( n5160 & ~n15668 ) | ( n14924 & ~n15668 ) ;
  assign n15670 = ( n2845 & n11061 ) | ( n2845 & n15669 ) | ( n11061 & n15669 ) ;
  assign n15676 = n15675 ^ n15670 ^ n3678 ;
  assign n15678 = n12733 ^ n11468 ^ n8107 ;
  assign n15677 = ( n3549 & ~n6593 ) | ( n3549 & n8556 ) | ( ~n6593 & n8556 ) ;
  assign n15679 = n15678 ^ n15677 ^ n9620 ;
  assign n15680 = ( ~x111 & n4566 ) | ( ~x111 & n9265 ) | ( n4566 & n9265 ) ;
  assign n15681 = n15680 ^ n13749 ^ n5301 ;
  assign n15682 = n15017 ^ n7993 ^ n4037 ;
  assign n15683 = ( ~n1477 & n2722 ) | ( ~n1477 & n15682 ) | ( n2722 & n15682 ) ;
  assign n15684 = ( n6173 & n14785 ) | ( n6173 & ~n15683 ) | ( n14785 & ~n15683 ) ;
  assign n15685 = n9407 ^ n9310 ^ n2327 ;
  assign n15686 = n4669 ^ n4449 ^ n2168 ;
  assign n15687 = ( n3245 & ~n10486 ) | ( n3245 & n15686 ) | ( ~n10486 & n15686 ) ;
  assign n15688 = n15687 ^ n11641 ^ n1555 ;
  assign n15689 = ( ~n683 & n15685 ) | ( ~n683 & n15688 ) | ( n15685 & n15688 ) ;
  assign n15695 = ( n265 & n1172 ) | ( n265 & n5169 ) | ( n1172 & n5169 ) ;
  assign n15696 = ( n3226 & ~n10471 ) | ( n3226 & n15695 ) | ( ~n10471 & n15695 ) ;
  assign n15697 = n15696 ^ n7334 ^ n3857 ;
  assign n15698 = n15697 ^ n9578 ^ n3497 ;
  assign n15690 = ( n1648 & n2645 ) | ( n1648 & ~n6603 ) | ( n2645 & ~n6603 ) ;
  assign n15691 = ( n4377 & ~n4811 ) | ( n4377 & n8367 ) | ( ~n4811 & n8367 ) ;
  assign n15692 = ( n8215 & ~n15690 ) | ( n8215 & n15691 ) | ( ~n15690 & n15691 ) ;
  assign n15693 = ( n768 & ~n5429 ) | ( n768 & n14426 ) | ( ~n5429 & n14426 ) ;
  assign n15694 = ( n7248 & ~n15692 ) | ( n7248 & n15693 ) | ( ~n15692 & n15693 ) ;
  assign n15699 = n15698 ^ n15694 ^ n793 ;
  assign n15700 = n7763 ^ n5102 ^ n3935 ;
  assign n15701 = ( n3137 & ~n14846 ) | ( n3137 & n15700 ) | ( ~n14846 & n15700 ) ;
  assign n15702 = n15701 ^ n3167 ^ n2092 ;
  assign n15703 = n7231 ^ n5720 ^ n1034 ;
  assign n15708 = n5950 ^ n4207 ^ n2258 ;
  assign n15709 = ( n773 & n9442 ) | ( n773 & n15708 ) | ( n9442 & n15708 ) ;
  assign n15710 = n15709 ^ n9141 ^ n4856 ;
  assign n15706 = n14034 ^ n2342 ^ n1802 ;
  assign n15705 = n10629 ^ n5105 ^ n3450 ;
  assign n15704 = ( n3240 & ~n5286 ) | ( n3240 & n14443 ) | ( ~n5286 & n14443 ) ;
  assign n15707 = n15706 ^ n15705 ^ n15704 ;
  assign n15711 = n15710 ^ n15707 ^ n4853 ;
  assign n15714 = n7358 ^ n6554 ^ n585 ;
  assign n15715 = n572 ^ n552 ^ n188 ;
  assign n15716 = n15715 ^ n3454 ^ n1152 ;
  assign n15717 = ( ~n2397 & n12846 ) | ( ~n2397 & n15716 ) | ( n12846 & n15716 ) ;
  assign n15718 = ( n13398 & n15714 ) | ( n13398 & ~n15717 ) | ( n15714 & ~n15717 ) ;
  assign n15719 = n15718 ^ n11770 ^ n975 ;
  assign n15712 = n11498 ^ n9875 ^ n8054 ;
  assign n15713 = ( ~n8845 & n11329 ) | ( ~n8845 & n15712 ) | ( n11329 & n15712 ) ;
  assign n15720 = n15719 ^ n15713 ^ n13250 ;
  assign n15730 = ( n385 & ~n4076 ) | ( n385 & n13910 ) | ( ~n4076 & n13910 ) ;
  assign n15721 = n7182 ^ n2162 ^ n1232 ;
  assign n15722 = ( ~n6484 & n11735 ) | ( ~n6484 & n15721 ) | ( n11735 & n15721 ) ;
  assign n15723 = ( n4554 & ~n14152 ) | ( n4554 & n15722 ) | ( ~n14152 & n15722 ) ;
  assign n15725 = n12053 ^ n9059 ^ n4741 ;
  assign n15724 = ( n1801 & ~n2702 ) | ( n1801 & n6297 ) | ( ~n2702 & n6297 ) ;
  assign n15726 = n15725 ^ n15724 ^ n7536 ;
  assign n15727 = n15726 ^ n10525 ^ n4550 ;
  assign n15728 = n15727 ^ n7058 ^ n3655 ;
  assign n15729 = ( n11934 & n15723 ) | ( n11934 & ~n15728 ) | ( n15723 & ~n15728 ) ;
  assign n15731 = n15730 ^ n15729 ^ n11978 ;
  assign n15733 = ( n1373 & n1916 ) | ( n1373 & ~n8800 ) | ( n1916 & ~n8800 ) ;
  assign n15732 = ( ~n425 & n5480 ) | ( ~n425 & n14794 ) | ( n5480 & n14794 ) ;
  assign n15734 = n15733 ^ n15732 ^ n4298 ;
  assign n15735 = ( n4154 & ~n13620 ) | ( n4154 & n15734 ) | ( ~n13620 & n15734 ) ;
  assign n15740 = ( n1287 & n3535 ) | ( n1287 & n11612 ) | ( n3535 & n11612 ) ;
  assign n15737 = n14226 ^ n11569 ^ n2319 ;
  assign n15738 = ( n2003 & ~n3222 ) | ( n2003 & n15737 ) | ( ~n3222 & n15737 ) ;
  assign n15739 = n15738 ^ n7312 ^ n5031 ;
  assign n15736 = ( n2355 & n6569 ) | ( n2355 & n7145 ) | ( n6569 & n7145 ) ;
  assign n15741 = n15740 ^ n15739 ^ n15736 ;
  assign n15744 = ( n8014 & n9740 ) | ( n8014 & n12795 ) | ( n9740 & n12795 ) ;
  assign n15742 = n13931 ^ n5976 ^ n3134 ;
  assign n15743 = n15742 ^ n13301 ^ n11336 ;
  assign n15745 = n15744 ^ n15743 ^ n9122 ;
  assign n15746 = n13220 ^ n1751 ^ n823 ;
  assign n15747 = ( n2952 & n9813 ) | ( n2952 & ~n15746 ) | ( n9813 & ~n15746 ) ;
  assign n15748 = ( n507 & ~n6228 ) | ( n507 & n15747 ) | ( ~n6228 & n15747 ) ;
  assign n15749 = ( n9271 & ~n14378 ) | ( n9271 & n14561 ) | ( ~n14378 & n14561 ) ;
  assign n15750 = ( ~n1950 & n6886 ) | ( ~n1950 & n15749 ) | ( n6886 & n15749 ) ;
  assign n15751 = ( n1375 & ~n4437 ) | ( n1375 & n5955 ) | ( ~n4437 & n5955 ) ;
  assign n15752 = ( ~n7109 & n7567 ) | ( ~n7109 & n15751 ) | ( n7567 & n15751 ) ;
  assign n15753 = n6801 ^ n5293 ^ n4953 ;
  assign n15754 = ( n7918 & n9291 ) | ( n7918 & ~n15753 ) | ( n9291 & ~n15753 ) ;
  assign n15759 = n15161 ^ n9298 ^ n1798 ;
  assign n15758 = n9558 ^ n7087 ^ n5814 ;
  assign n15756 = ( n896 & ~n7893 ) | ( n896 & n10309 ) | ( ~n7893 & n10309 ) ;
  assign n15755 = ( n2772 & n8369 ) | ( n2772 & ~n12784 ) | ( n8369 & ~n12784 ) ;
  assign n15757 = n15756 ^ n15755 ^ n2117 ;
  assign n15760 = n15759 ^ n15758 ^ n15757 ;
  assign n15761 = ( n3829 & n15754 ) | ( n3829 & ~n15760 ) | ( n15754 & ~n15760 ) ;
  assign n15762 = n15761 ^ n8512 ^ n7808 ;
  assign n15763 = ( x118 & ~n2473 ) | ( x118 & n6270 ) | ( ~n2473 & n6270 ) ;
  assign n15764 = ( n12115 & n12699 ) | ( n12115 & ~n15763 ) | ( n12699 & ~n15763 ) ;
  assign n15765 = ( ~n236 & n2892 ) | ( ~n236 & n6012 ) | ( n2892 & n6012 ) ;
  assign n15766 = ( n7196 & n14737 ) | ( n7196 & ~n15765 ) | ( n14737 & ~n15765 ) ;
  assign n15768 = ( ~n2776 & n3652 ) | ( ~n2776 & n5343 ) | ( n3652 & n5343 ) ;
  assign n15769 = ( n5200 & ~n8906 ) | ( n5200 & n15768 ) | ( ~n8906 & n15768 ) ;
  assign n15767 = n5248 ^ n3946 ^ n1721 ;
  assign n15770 = n15769 ^ n15767 ^ n14695 ;
  assign n15771 = n15770 ^ n9048 ^ n8446 ;
  assign n15772 = ( n4133 & n8091 ) | ( n4133 & n13310 ) | ( n8091 & n13310 ) ;
  assign n15773 = n15772 ^ n8539 ^ n4749 ;
  assign n15774 = n15773 ^ n5280 ^ n1408 ;
  assign n15775 = ( n2490 & ~n4940 ) | ( n2490 & n9978 ) | ( ~n4940 & n9978 ) ;
  assign n15776 = n15775 ^ n15693 ^ n4212 ;
  assign n15779 = n13249 ^ n7991 ^ n511 ;
  assign n15780 = ( n2706 & n2805 ) | ( n2706 & ~n8526 ) | ( n2805 & ~n8526 ) ;
  assign n15781 = ( ~n13692 & n15779 ) | ( ~n13692 & n15780 ) | ( n15779 & n15780 ) ;
  assign n15777 = n7880 ^ n6733 ^ n6446 ;
  assign n15778 = ( n3374 & n14579 ) | ( n3374 & n15777 ) | ( n14579 & n15777 ) ;
  assign n15782 = n15781 ^ n15778 ^ n11997 ;
  assign n15783 = ( n415 & n3030 ) | ( n415 & n9523 ) | ( n3030 & n9523 ) ;
  assign n15784 = ( ~n229 & n5795 ) | ( ~n229 & n6808 ) | ( n5795 & n6808 ) ;
  assign n15785 = n9924 ^ n8139 ^ n3467 ;
  assign n15786 = ( n2006 & ~n9489 ) | ( n2006 & n15785 ) | ( ~n9489 & n15785 ) ;
  assign n15787 = n11955 ^ n11439 ^ n6717 ;
  assign n15788 = ( n10512 & n14620 ) | ( n10512 & ~n15787 ) | ( n14620 & ~n15787 ) ;
  assign n15789 = n11778 ^ n4039 ^ n918 ;
  assign n15790 = n15789 ^ n12136 ^ n5375 ;
  assign n15791 = ( n5520 & ~n8131 ) | ( n5520 & n8488 ) | ( ~n8131 & n8488 ) ;
  assign n15792 = n13082 ^ n10096 ^ n2241 ;
  assign n15793 = ( n1121 & n5976 ) | ( n1121 & ~n15792 ) | ( n5976 & ~n15792 ) ;
  assign n15794 = ( ~n15790 & n15791 ) | ( ~n15790 & n15793 ) | ( n15791 & n15793 ) ;
  assign n15795 = n9541 ^ n4679 ^ n4142 ;
  assign n15796 = n15795 ^ n15515 ^ n10011 ;
  assign n15797 = ( ~n3656 & n4629 ) | ( ~n3656 & n10519 ) | ( n4629 & n10519 ) ;
  assign n15798 = ( n2941 & n11990 ) | ( n2941 & n15797 ) | ( n11990 & n15797 ) ;
  assign n15799 = ( n2479 & n15796 ) | ( n2479 & n15798 ) | ( n15796 & n15798 ) ;
  assign n15800 = n12480 ^ n4881 ^ n2339 ;
  assign n15801 = ( ~n329 & n6886 ) | ( ~n329 & n12125 ) | ( n6886 & n12125 ) ;
  assign n15802 = ( n7119 & n9482 ) | ( n7119 & ~n15801 ) | ( n9482 & ~n15801 ) ;
  assign n15803 = ( n1876 & n15800 ) | ( n1876 & n15802 ) | ( n15800 & n15802 ) ;
  assign n15804 = ( n2730 & ~n11733 ) | ( n2730 & n14390 ) | ( ~n11733 & n14390 ) ;
  assign n15805 = ( ~n1748 & n4633 ) | ( ~n1748 & n12760 ) | ( n4633 & n12760 ) ;
  assign n15806 = ( n1382 & n12823 ) | ( n1382 & ~n14297 ) | ( n12823 & ~n14297 ) ;
  assign n15807 = ( n2227 & ~n2483 ) | ( n2227 & n3613 ) | ( ~n2483 & n3613 ) ;
  assign n15808 = ( n4210 & n8918 ) | ( n4210 & ~n12508 ) | ( n8918 & ~n12508 ) ;
  assign n15809 = ( n208 & n15807 ) | ( n208 & ~n15808 ) | ( n15807 & ~n15808 ) ;
  assign n15810 = ( n7609 & n15806 ) | ( n7609 & n15809 ) | ( n15806 & n15809 ) ;
  assign n15811 = n7327 ^ n3831 ^ x119 ;
  assign n15812 = n10350 ^ n9100 ^ n8489 ;
  assign n15813 = ( n8694 & n15811 ) | ( n8694 & ~n15812 ) | ( n15811 & ~n15812 ) ;
  assign n15814 = n12575 ^ n12167 ^ n11598 ;
  assign n15815 = n15814 ^ n11773 ^ n130 ;
  assign n15816 = ( ~n901 & n1185 ) | ( ~n901 & n2538 ) | ( n1185 & n2538 ) ;
  assign n15817 = ( n6204 & n13942 ) | ( n6204 & n15816 ) | ( n13942 & n15816 ) ;
  assign n15818 = n15817 ^ n7922 ^ n3335 ;
  assign n15819 = ( n15813 & n15815 ) | ( n15813 & ~n15818 ) | ( n15815 & ~n15818 ) ;
  assign n15820 = ( ~n3374 & n3399 ) | ( ~n3374 & n7315 ) | ( n3399 & n7315 ) ;
  assign n15821 = ( n3461 & n6171 ) | ( n3461 & ~n8181 ) | ( n6171 & ~n8181 ) ;
  assign n15822 = n15821 ^ n10119 ^ n3889 ;
  assign n15823 = ( n3482 & n6690 ) | ( n3482 & n15822 ) | ( n6690 & n15822 ) ;
  assign n15824 = ( n15067 & n15820 ) | ( n15067 & n15823 ) | ( n15820 & n15823 ) ;
  assign n15827 = n11057 ^ n4078 ^ x8 ;
  assign n15828 = ( ~n730 & n4864 ) | ( ~n730 & n15827 ) | ( n4864 & n15827 ) ;
  assign n15825 = n12908 ^ n8397 ^ n2956 ;
  assign n15826 = n15825 ^ n12044 ^ n2786 ;
  assign n15829 = n15828 ^ n15826 ^ n8914 ;
  assign n15834 = ( n6719 & n6914 ) | ( n6719 & n10886 ) | ( n6914 & n10886 ) ;
  assign n15835 = n15834 ^ n14300 ^ n1669 ;
  assign n15836 = n15835 ^ n9383 ^ n1488 ;
  assign n15830 = n3999 ^ n3618 ^ n549 ;
  assign n15831 = n15551 ^ n12951 ^ n4639 ;
  assign n15832 = ( n1765 & ~n2527 ) | ( n1765 & n15831 ) | ( ~n2527 & n15831 ) ;
  assign n15833 = ( n10537 & n15830 ) | ( n10537 & ~n15832 ) | ( n15830 & ~n15832 ) ;
  assign n15837 = n15836 ^ n15833 ^ n4519 ;
  assign n15839 = n5236 ^ n2075 ^ n585 ;
  assign n15838 = ( ~n462 & n5773 ) | ( ~n462 & n7000 ) | ( n5773 & n7000 ) ;
  assign n15840 = n15839 ^ n15838 ^ n8296 ;
  assign n15841 = n15840 ^ n12868 ^ n8022 ;
  assign n15842 = ( n2236 & ~n3836 ) | ( n2236 & n7224 ) | ( ~n3836 & n7224 ) ;
  assign n15843 = n6984 ^ n5010 ^ n2503 ;
  assign n15844 = ( n3724 & n9143 ) | ( n3724 & n15843 ) | ( n9143 & n15843 ) ;
  assign n15845 = ( ~n5154 & n8222 ) | ( ~n5154 & n15844 ) | ( n8222 & n15844 ) ;
  assign n15846 = n15845 ^ n8477 ^ n2398 ;
  assign n15847 = ( n15841 & n15842 ) | ( n15841 & ~n15846 ) | ( n15842 & ~n15846 ) ;
  assign n15854 = n5260 ^ n4985 ^ n2010 ;
  assign n15851 = n7158 ^ n741 ^ n169 ;
  assign n15852 = ( n2341 & n6221 ) | ( n2341 & n15851 ) | ( n6221 & n15851 ) ;
  assign n15853 = ( n7124 & ~n7987 ) | ( n7124 & n15852 ) | ( ~n7987 & n15852 ) ;
  assign n15855 = n15854 ^ n15853 ^ n430 ;
  assign n15848 = n5312 ^ n2930 ^ n1930 ;
  assign n15849 = n15848 ^ n12045 ^ n675 ;
  assign n15850 = ( n7360 & n8702 ) | ( n7360 & ~n15849 ) | ( n8702 & ~n15849 ) ;
  assign n15856 = n15855 ^ n15850 ^ n2879 ;
  assign n15857 = n14237 ^ n3223 ^ n1183 ;
  assign n15858 = ( n3803 & n15856 ) | ( n3803 & ~n15857 ) | ( n15856 & ~n15857 ) ;
  assign n15859 = ( n1869 & n10293 ) | ( n1869 & ~n13817 ) | ( n10293 & ~n13817 ) ;
  assign n15860 = n15859 ^ n5610 ^ n2884 ;
  assign n15865 = ( n131 & n1338 ) | ( n131 & ~n2261 ) | ( n1338 & ~n2261 ) ;
  assign n15863 = ( n1074 & n4492 ) | ( n1074 & n7624 ) | ( n4492 & n7624 ) ;
  assign n15864 = n15863 ^ n6757 ^ n1335 ;
  assign n15861 = n15848 ^ n5806 ^ n350 ;
  assign n15862 = n15861 ^ n12068 ^ n11712 ;
  assign n15866 = n15865 ^ n15864 ^ n15862 ;
  assign n15867 = n9092 ^ n7329 ^ n7004 ;
  assign n15868 = n12275 ^ n8564 ^ n3748 ;
  assign n15869 = n15278 ^ n10700 ^ n10221 ;
  assign n15870 = ( n2521 & n15868 ) | ( n2521 & ~n15869 ) | ( n15868 & ~n15869 ) ;
  assign n15871 = ( n8095 & n15867 ) | ( n8095 & n15870 ) | ( n15867 & n15870 ) ;
  assign n15876 = n10651 ^ n1693 ^ n549 ;
  assign n15872 = n8849 ^ n8757 ^ n3472 ;
  assign n15873 = ( n576 & n5044 ) | ( n576 & ~n6810 ) | ( n5044 & ~n6810 ) ;
  assign n15874 = ( n11173 & ~n13045 ) | ( n11173 & n15873 ) | ( ~n13045 & n15873 ) ;
  assign n15875 = ( ~n10710 & n15872 ) | ( ~n10710 & n15874 ) | ( n15872 & n15874 ) ;
  assign n15877 = n15876 ^ n15875 ^ n12609 ;
  assign n15878 = n7450 ^ n4963 ^ n4592 ;
  assign n15879 = n15878 ^ n14762 ^ n9312 ;
  assign n15880 = ( n9106 & n10723 ) | ( n9106 & ~n15879 ) | ( n10723 & ~n15879 ) ;
  assign n15881 = n15880 ^ n8884 ^ n4905 ;
  assign n15882 = ( n10758 & ~n15877 ) | ( n10758 & n15881 ) | ( ~n15877 & n15881 ) ;
  assign n15884 = ( n1792 & n3981 ) | ( n1792 & n8620 ) | ( n3981 & n8620 ) ;
  assign n15883 = ( n933 & ~n3421 ) | ( n933 & n9163 ) | ( ~n3421 & n9163 ) ;
  assign n15885 = n15884 ^ n15883 ^ n1127 ;
  assign n15886 = ( n1231 & n2023 ) | ( n1231 & ~n15885 ) | ( n2023 & ~n15885 ) ;
  assign n15887 = ( n6794 & ~n14132 ) | ( n6794 & n14990 ) | ( ~n14132 & n14990 ) ;
  assign n15888 = ( n4449 & ~n15886 ) | ( n4449 & n15887 ) | ( ~n15886 & n15887 ) ;
  assign n15889 = ( n2405 & ~n8722 ) | ( n2405 & n15888 ) | ( ~n8722 & n15888 ) ;
  assign n15890 = n5429 ^ n5342 ^ n3258 ;
  assign n15891 = n15890 ^ n13291 ^ n6262 ;
  assign n15892 = n13834 ^ n9728 ^ n2222 ;
  assign n15896 = n4270 ^ n3767 ^ n1027 ;
  assign n15897 = n15896 ^ n7598 ^ n1372 ;
  assign n15898 = n15897 ^ n1008 ^ n539 ;
  assign n15899 = n15898 ^ n4679 ^ n1828 ;
  assign n15900 = n15899 ^ n12078 ^ n7162 ;
  assign n15893 = ( n3281 & ~n6046 ) | ( n3281 & n10116 ) | ( ~n6046 & n10116 ) ;
  assign n15894 = ( ~n5243 & n9880 ) | ( ~n5243 & n15893 ) | ( n9880 & n15893 ) ;
  assign n15895 = n15894 ^ n15827 ^ n643 ;
  assign n15901 = n15900 ^ n15895 ^ n12004 ;
  assign n15902 = n15901 ^ n6547 ^ n4521 ;
  assign n15903 = n8298 ^ n1956 ^ n1287 ;
  assign n15904 = ( ~n601 & n4870 ) | ( ~n601 & n15903 ) | ( n4870 & n15903 ) ;
  assign n15905 = n15904 ^ n5311 ^ n4929 ;
  assign n15906 = n15905 ^ n8560 ^ n7025 ;
  assign n15907 = ( n1056 & n3051 ) | ( n1056 & n15906 ) | ( n3051 & n15906 ) ;
  assign n15908 = n6984 ^ n2353 ^ x23 ;
  assign n15909 = ( ~n1988 & n4488 ) | ( ~n1988 & n15908 ) | ( n4488 & n15908 ) ;
  assign n15910 = ( n167 & n5254 ) | ( n167 & n15909 ) | ( n5254 & n15909 ) ;
  assign n15911 = n15910 ^ n6689 ^ n1940 ;
  assign n15915 = n8603 ^ n6471 ^ n3145 ;
  assign n15914 = n7229 ^ n6835 ^ x23 ;
  assign n15912 = n7410 ^ n2927 ^ n1838 ;
  assign n15913 = n15912 ^ n3977 ^ n3253 ;
  assign n15916 = n15915 ^ n15914 ^ n15913 ;
  assign n15917 = ( ~n4330 & n7266 ) | ( ~n4330 & n8325 ) | ( n7266 & n8325 ) ;
  assign n15918 = ( n10167 & n10551 ) | ( n10167 & ~n15917 ) | ( n10551 & ~n15917 ) ;
  assign n15919 = n13484 ^ n7039 ^ n2955 ;
  assign n15920 = ( n10426 & n11910 ) | ( n10426 & ~n15919 ) | ( n11910 & ~n15919 ) ;
  assign n15921 = ( n4009 & n5474 ) | ( n4009 & ~n15920 ) | ( n5474 & ~n15920 ) ;
  assign n15922 = n15921 ^ n4083 ^ n1724 ;
  assign n15926 = n5327 ^ n3306 ^ n2760 ;
  assign n15928 = ( n1562 & n13456 ) | ( n1562 & ~n15020 ) | ( n13456 & ~n15020 ) ;
  assign n15927 = ( n2289 & ~n5324 ) | ( n2289 & n8051 ) | ( ~n5324 & n8051 ) ;
  assign n15929 = n15928 ^ n15927 ^ n893 ;
  assign n15930 = n15929 ^ n5538 ^ n584 ;
  assign n15931 = ( n15172 & ~n15926 ) | ( n15172 & n15930 ) | ( ~n15926 & n15930 ) ;
  assign n15923 = ( n2494 & n13914 ) | ( n2494 & ~n14649 ) | ( n13914 & ~n14649 ) ;
  assign n15924 = n12667 ^ n5006 ^ n2124 ;
  assign n15925 = ( ~n1323 & n15923 ) | ( ~n1323 & n15924 ) | ( n15923 & n15924 ) ;
  assign n15932 = n15931 ^ n15925 ^ n11464 ;
  assign n15933 = n4492 ^ n3792 ^ n467 ;
  assign n15934 = n15933 ^ n8073 ^ n2675 ;
  assign n15935 = n15934 ^ n9441 ^ n8437 ;
  assign n15936 = ( n2185 & n9443 ) | ( n2185 & ~n13429 ) | ( n9443 & ~n13429 ) ;
  assign n15937 = n15936 ^ n3216 ^ n1596 ;
  assign n15938 = n1907 ^ n591 ^ x2 ;
  assign n15939 = n15938 ^ n12648 ^ n2108 ;
  assign n15940 = n11834 ^ n6427 ^ n5829 ;
  assign n15941 = ( ~n1077 & n9138 ) | ( ~n1077 & n15940 ) | ( n9138 & n15940 ) ;
  assign n15943 = ( ~n2418 & n3086 ) | ( ~n2418 & n6444 ) | ( n3086 & n6444 ) ;
  assign n15942 = n7476 ^ n4437 ^ n670 ;
  assign n15944 = n15943 ^ n15942 ^ n8041 ;
  assign n15945 = ( n2779 & n5420 ) | ( n2779 & n14437 ) | ( n5420 & n14437 ) ;
  assign n15946 = ( n2075 & n3642 ) | ( n2075 & n13893 ) | ( n3642 & n13893 ) ;
  assign n15947 = ( n5438 & ~n15405 ) | ( n5438 & n15946 ) | ( ~n15405 & n15946 ) ;
  assign n15948 = ( ~n2742 & n15945 ) | ( ~n2742 & n15947 ) | ( n15945 & n15947 ) ;
  assign n15949 = n6912 ^ n5361 ^ n1198 ;
  assign n15950 = ( n11187 & n13548 ) | ( n11187 & ~n15949 ) | ( n13548 & ~n15949 ) ;
  assign n15957 = ( ~n8925 & n10313 ) | ( ~n8925 & n13255 ) | ( n10313 & n13255 ) ;
  assign n15956 = n9122 ^ n2064 ^ n1933 ;
  assign n15951 = ( ~n3626 & n5117 ) | ( ~n3626 & n11449 ) | ( n5117 & n11449 ) ;
  assign n15952 = ( x113 & n3360 ) | ( x113 & ~n5122 ) | ( n3360 & ~n5122 ) ;
  assign n15953 = n15952 ^ n3178 ^ n2603 ;
  assign n15954 = ( n5916 & n8382 ) | ( n5916 & n15953 ) | ( n8382 & n15953 ) ;
  assign n15955 = ( n2495 & n15951 ) | ( n2495 & ~n15954 ) | ( n15951 & ~n15954 ) ;
  assign n15958 = n15957 ^ n15956 ^ n15955 ;
  assign n15959 = n12370 ^ n8705 ^ n5901 ;
  assign n15960 = n15959 ^ n15516 ^ n10244 ;
  assign n15961 = ( ~n3310 & n10142 ) | ( ~n3310 & n15204 ) | ( n10142 & n15204 ) ;
  assign n15962 = n9009 ^ n3603 ^ n2022 ;
  assign n15963 = n12701 ^ n5861 ^ n754 ;
  assign n15964 = ( ~n1041 & n7394 ) | ( ~n1041 & n9081 ) | ( n7394 & n9081 ) ;
  assign n15965 = ( n12660 & n12895 ) | ( n12660 & n15800 ) | ( n12895 & n15800 ) ;
  assign n15966 = ( n3417 & n15964 ) | ( n3417 & n15965 ) | ( n15964 & n15965 ) ;
  assign n15967 = n15625 ^ n8095 ^ n7365 ;
  assign n15968 = ( n8523 & ~n10194 ) | ( n8523 & n15967 ) | ( ~n10194 & n15967 ) ;
  assign n15971 = ( n206 & n5645 ) | ( n206 & ~n8250 ) | ( n5645 & ~n8250 ) ;
  assign n15970 = ( ~n2991 & n7022 ) | ( ~n2991 & n14491 ) | ( n7022 & n14491 ) ;
  assign n15969 = ( n3259 & ~n9462 ) | ( n3259 & n9519 ) | ( ~n9462 & n9519 ) ;
  assign n15972 = n15971 ^ n15970 ^ n15969 ;
  assign n15975 = n7382 ^ n6312 ^ n407 ;
  assign n15974 = ( n10329 & n11044 ) | ( n10329 & ~n12205 ) | ( n11044 & ~n12205 ) ;
  assign n15973 = n13809 ^ n8484 ^ n4042 ;
  assign n15976 = n15975 ^ n15974 ^ n15973 ;
  assign n15977 = ( n15968 & n15972 ) | ( n15968 & n15976 ) | ( n15972 & n15976 ) ;
  assign n15978 = n9469 ^ n6566 ^ x104 ;
  assign n15979 = n15978 ^ n10808 ^ n1197 ;
  assign n15980 = ( n4522 & ~n11711 ) | ( n4522 & n15979 ) | ( ~n11711 & n15979 ) ;
  assign n15981 = ( ~n10320 & n10331 ) | ( ~n10320 & n15245 ) | ( n10331 & n15245 ) ;
  assign n15982 = n6155 ^ n3401 ^ n3025 ;
  assign n15983 = ( n10014 & n10974 ) | ( n10014 & n15982 ) | ( n10974 & n15982 ) ;
  assign n15984 = n15983 ^ n13806 ^ n7847 ;
  assign n15985 = n13187 ^ n3898 ^ n2950 ;
  assign n15986 = ( n1063 & ~n13348 ) | ( n1063 & n14719 ) | ( ~n13348 & n14719 ) ;
  assign n15987 = ( n8269 & ~n14333 ) | ( n8269 & n15986 ) | ( ~n14333 & n15986 ) ;
  assign n15991 = ( n3199 & n11797 ) | ( n3199 & n14886 ) | ( n11797 & n14886 ) ;
  assign n15988 = ( n5832 & n9774 ) | ( n5832 & n13529 ) | ( n9774 & n13529 ) ;
  assign n15989 = n15988 ^ n4778 ^ n1669 ;
  assign n15990 = ( ~n4218 & n12823 ) | ( ~n4218 & n15989 ) | ( n12823 & n15989 ) ;
  assign n15992 = n15991 ^ n15990 ^ n3210 ;
  assign n15994 = n5170 ^ n2042 ^ n1668 ;
  assign n15993 = n14152 ^ n12975 ^ n8164 ;
  assign n15995 = n15994 ^ n15993 ^ n7990 ;
  assign n15996 = n14613 ^ n4014 ^ n802 ;
  assign n15997 = ( n2284 & ~n7997 ) | ( n2284 & n12725 ) | ( ~n7997 & n12725 ) ;
  assign n15998 = n15997 ^ n9579 ^ n7059 ;
  assign n15999 = n15998 ^ n12186 ^ n11677 ;
  assign n16000 = ( n6790 & n15996 ) | ( n6790 & n15999 ) | ( n15996 & n15999 ) ;
  assign n16001 = n12576 ^ n12549 ^ n3918 ;
  assign n16003 = ( n1713 & n2375 ) | ( n1713 & n5968 ) | ( n2375 & n5968 ) ;
  assign n16002 = ( ~n1154 & n5151 ) | ( ~n1154 & n14575 ) | ( n5151 & n14575 ) ;
  assign n16004 = n16003 ^ n16002 ^ n15518 ;
  assign n16005 = n9178 ^ n6383 ^ n2564 ;
  assign n16006 = n3871 ^ n681 ^ n610 ;
  assign n16007 = ( ~n3539 & n6280 ) | ( ~n3539 & n13866 ) | ( n6280 & n13866 ) ;
  assign n16008 = ( n3133 & n16006 ) | ( n3133 & ~n16007 ) | ( n16006 & ~n16007 ) ;
  assign n16009 = ( n9582 & n9666 ) | ( n9582 & ~n16008 ) | ( n9666 & ~n16008 ) ;
  assign n16010 = n9306 ^ n8801 ^ n3016 ;
  assign n16011 = n6534 ^ n1968 ^ n1307 ;
  assign n16012 = ( n1073 & n1467 ) | ( n1073 & n3101 ) | ( n1467 & n3101 ) ;
  assign n16013 = ( ~n10713 & n10870 ) | ( ~n10713 & n16012 ) | ( n10870 & n16012 ) ;
  assign n16015 = n14583 ^ n5709 ^ n1744 ;
  assign n16016 = ( n476 & n10053 ) | ( n476 & n16015 ) | ( n10053 & n16015 ) ;
  assign n16014 = n3630 ^ n3471 ^ n165 ;
  assign n16017 = n16016 ^ n16014 ^ n6686 ;
  assign n16018 = n15621 ^ n11077 ^ n5169 ;
  assign n16019 = ( ~n3054 & n14138 ) | ( ~n3054 & n16018 ) | ( n14138 & n16018 ) ;
  assign n16020 = n14941 ^ n6107 ^ n377 ;
  assign n16021 = n16020 ^ n10488 ^ n515 ;
  assign n16026 = ( n3556 & n4165 ) | ( n3556 & n7720 ) | ( n4165 & n7720 ) ;
  assign n16024 = n6361 ^ n3835 ^ n1525 ;
  assign n16022 = n10825 ^ n9236 ^ n156 ;
  assign n16023 = ( n6042 & ~n9572 ) | ( n6042 & n16022 ) | ( ~n9572 & n16022 ) ;
  assign n16025 = n16024 ^ n16023 ^ n8143 ;
  assign n16027 = n16026 ^ n16025 ^ n7362 ;
  assign n16029 = n8228 ^ n4870 ^ n3468 ;
  assign n16028 = n7153 ^ n5106 ^ n4910 ;
  assign n16030 = n16029 ^ n16028 ^ n2647 ;
  assign n16032 = n4879 ^ n1299 ^ n382 ;
  assign n16033 = n16032 ^ n9383 ^ n1126 ;
  assign n16031 = n5540 ^ n2864 ^ n2458 ;
  assign n16034 = n16033 ^ n16031 ^ n1599 ;
  assign n16035 = n11255 ^ n9128 ^ n972 ;
  assign n16036 = n10159 ^ n8890 ^ n1814 ;
  assign n16037 = ( n811 & n16035 ) | ( n811 & n16036 ) | ( n16035 & n16036 ) ;
  assign n16038 = ( ~n5855 & n14927 ) | ( ~n5855 & n15236 ) | ( n14927 & n15236 ) ;
  assign n16039 = ( ~n3452 & n8116 ) | ( ~n3452 & n13171 ) | ( n8116 & n13171 ) ;
  assign n16047 = ( ~n674 & n1968 ) | ( ~n674 & n10019 ) | ( n1968 & n10019 ) ;
  assign n16048 = ( n4952 & ~n8214 ) | ( n4952 & n16047 ) | ( ~n8214 & n16047 ) ;
  assign n16040 = n4640 ^ n4551 ^ n1933 ;
  assign n16044 = ( n2431 & n8428 ) | ( n2431 & ~n11582 ) | ( n8428 & ~n11582 ) ;
  assign n16041 = ( n4137 & n7163 ) | ( n4137 & n10553 ) | ( n7163 & n10553 ) ;
  assign n16042 = n16041 ^ n6403 ^ n2824 ;
  assign n16043 = ( n6080 & ~n8010 ) | ( n6080 & n16042 ) | ( ~n8010 & n16042 ) ;
  assign n16045 = n16044 ^ n16043 ^ n4845 ;
  assign n16046 = ( n519 & n16040 ) | ( n519 & n16045 ) | ( n16040 & n16045 ) ;
  assign n16049 = n16048 ^ n16046 ^ n5617 ;
  assign n16050 = ( ~n1290 & n7030 ) | ( ~n1290 & n12764 ) | ( n7030 & n12764 ) ;
  assign n16051 = n16050 ^ n15867 ^ n1530 ;
  assign n16052 = n15377 ^ n7159 ^ n3207 ;
  assign n16053 = ( n2278 & n8844 ) | ( n2278 & ~n9802 ) | ( n8844 & ~n9802 ) ;
  assign n16054 = n16053 ^ n496 ^ n482 ;
  assign n16055 = n15872 ^ n12522 ^ n4069 ;
  assign n16056 = n16055 ^ n9003 ^ n1592 ;
  assign n16057 = n16056 ^ n6690 ^ n6264 ;
  assign n16058 = ( ~n6471 & n7774 ) | ( ~n6471 & n9561 ) | ( n7774 & n9561 ) ;
  assign n16059 = n4256 ^ n3807 ^ n3119 ;
  assign n16060 = ( ~n4558 & n16058 ) | ( ~n4558 & n16059 ) | ( n16058 & n16059 ) ;
  assign n16061 = ( n3190 & n3448 ) | ( n3190 & ~n8252 ) | ( n3448 & ~n8252 ) ;
  assign n16062 = ( n4526 & ~n16060 ) | ( n4526 & n16061 ) | ( ~n16060 & n16061 ) ;
  assign n16069 = n10135 ^ n5843 ^ n4437 ;
  assign n16068 = ( n7114 & n12017 ) | ( n7114 & n12170 ) | ( n12017 & n12170 ) ;
  assign n16063 = n8773 ^ n1821 ^ n1462 ;
  assign n16064 = n12379 ^ n8508 ^ n1144 ;
  assign n16065 = n16064 ^ n13996 ^ n5902 ;
  assign n16066 = n16065 ^ n12215 ^ n7821 ;
  assign n16067 = ( n6394 & ~n16063 ) | ( n6394 & n16066 ) | ( ~n16063 & n16066 ) ;
  assign n16070 = n16069 ^ n16068 ^ n16067 ;
  assign n16073 = ( n2534 & n3847 ) | ( n2534 & n14129 ) | ( n3847 & n14129 ) ;
  assign n16071 = ( n3826 & n8511 ) | ( n3826 & ~n13601 ) | ( n8511 & ~n13601 ) ;
  assign n16072 = ( n8768 & ~n9865 ) | ( n8768 & n16071 ) | ( ~n9865 & n16071 ) ;
  assign n16074 = n16073 ^ n16072 ^ n142 ;
  assign n16078 = n13478 ^ n5721 ^ n4666 ;
  assign n16076 = n9479 ^ n5218 ^ n943 ;
  assign n16077 = ( ~n3050 & n9403 ) | ( ~n3050 & n16076 ) | ( n9403 & n16076 ) ;
  assign n16075 = ( x46 & n2088 ) | ( x46 & n6297 ) | ( n2088 & n6297 ) ;
  assign n16079 = n16078 ^ n16077 ^ n16075 ;
  assign n16080 = ( n1762 & ~n3190 ) | ( n1762 & n11228 ) | ( ~n3190 & n11228 ) ;
  assign n16081 = ( n202 & n3380 ) | ( n202 & ~n4852 ) | ( n3380 & ~n4852 ) ;
  assign n16082 = n16081 ^ n11602 ^ n4531 ;
  assign n16083 = n8422 ^ n2617 ^ n550 ;
  assign n16084 = ( n1877 & ~n16082 ) | ( n1877 & n16083 ) | ( ~n16082 & n16083 ) ;
  assign n16085 = ( n1315 & n9572 ) | ( n1315 & n13138 ) | ( n9572 & n13138 ) ;
  assign n16086 = n16085 ^ n10505 ^ n8754 ;
  assign n16087 = n16086 ^ n5335 ^ n2935 ;
  assign n16089 = ( ~n193 & n5081 ) | ( ~n193 & n6542 ) | ( n5081 & n6542 ) ;
  assign n16090 = n16089 ^ n6128 ^ n2457 ;
  assign n16091 = ( n1383 & ~n8125 ) | ( n1383 & n16090 ) | ( ~n8125 & n16090 ) ;
  assign n16088 = n10290 ^ n8858 ^ x2 ;
  assign n16092 = n16091 ^ n16088 ^ n14140 ;
  assign n16093 = n13261 ^ n12932 ^ n5654 ;
  assign n16094 = ( n8966 & n12231 ) | ( n8966 & n16093 ) | ( n12231 & n16093 ) ;
  assign n16095 = ( n6929 & n15112 ) | ( n6929 & n15549 ) | ( n15112 & n15549 ) ;
  assign n16096 = n16095 ^ n15293 ^ n465 ;
  assign n16097 = n14920 ^ n4768 ^ n4071 ;
  assign n16100 = n9424 ^ n3574 ^ n933 ;
  assign n16101 = n16100 ^ n13564 ^ n5194 ;
  assign n16102 = ( n7974 & n14766 ) | ( n7974 & ~n16101 ) | ( n14766 & ~n16101 ) ;
  assign n16098 = n7769 ^ n5128 ^ n1684 ;
  assign n16099 = n16098 ^ n6164 ^ n1245 ;
  assign n16103 = n16102 ^ n16099 ^ n1676 ;
  assign n16107 = ( n4018 & n7356 ) | ( n4018 & ~n9136 ) | ( n7356 & ~n9136 ) ;
  assign n16105 = ( n1324 & n4114 ) | ( n1324 & ~n10665 ) | ( n4114 & ~n10665 ) ;
  assign n16106 = ( n4936 & ~n11933 ) | ( n4936 & n16105 ) | ( ~n11933 & n16105 ) ;
  assign n16104 = n15751 ^ n13468 ^ n5377 ;
  assign n16108 = n16107 ^ n16106 ^ n16104 ;
  assign n16109 = n7314 ^ n5191 ^ n3691 ;
  assign n16110 = ( n5748 & n14714 ) | ( n5748 & n16109 ) | ( n14714 & n16109 ) ;
  assign n16111 = n16110 ^ n12390 ^ n3767 ;
  assign n16113 = n7035 ^ n4637 ^ n1172 ;
  assign n16112 = n13208 ^ n5171 ^ n833 ;
  assign n16114 = n16113 ^ n16112 ^ n9041 ;
  assign n16115 = ( n1283 & n6235 ) | ( n1283 & n11154 ) | ( n6235 & n11154 ) ;
  assign n16116 = n16115 ^ n10391 ^ n2664 ;
  assign n16117 = n8435 ^ n4433 ^ n3493 ;
  assign n16118 = n16117 ^ n10794 ^ n6248 ;
  assign n16119 = n14292 ^ n5859 ^ n1512 ;
  assign n16120 = n7567 ^ n1807 ^ n1173 ;
  assign n16121 = ( n13983 & n16119 ) | ( n13983 & ~n16120 ) | ( n16119 & ~n16120 ) ;
  assign n16122 = ( ~n1779 & n5524 ) | ( ~n1779 & n5771 ) | ( n5524 & n5771 ) ;
  assign n16123 = n16122 ^ n14471 ^ n247 ;
  assign n16124 = ( n4731 & ~n10062 ) | ( n4731 & n12294 ) | ( ~n10062 & n12294 ) ;
  assign n16125 = n11842 ^ n4437 ^ n1718 ;
  assign n16126 = ( ~n2815 & n5010 ) | ( ~n2815 & n16125 ) | ( n5010 & n16125 ) ;
  assign n16127 = n10212 ^ n9847 ^ n7920 ;
  assign n16128 = n16127 ^ n6332 ^ n2628 ;
  assign n16129 = ( n16124 & n16126 ) | ( n16124 & ~n16128 ) | ( n16126 & ~n16128 ) ;
  assign n16130 = n11470 ^ n10370 ^ n515 ;
  assign n16131 = n8843 ^ n4191 ^ n2530 ;
  assign n16132 = n16131 ^ n14513 ^ n10920 ;
  assign n16133 = ( n434 & n16130 ) | ( n434 & ~n16132 ) | ( n16130 & ~n16132 ) ;
  assign n16134 = ( n6319 & n16129 ) | ( n6319 & n16133 ) | ( n16129 & n16133 ) ;
  assign n16135 = ( n796 & n6578 ) | ( n796 & n7701 ) | ( n6578 & n7701 ) ;
  assign n16136 = ( n3585 & n7326 ) | ( n3585 & ~n16135 ) | ( n7326 & ~n16135 ) ;
  assign n16137 = n11784 ^ n10557 ^ n3520 ;
  assign n16138 = ( n3106 & n16136 ) | ( n3106 & ~n16137 ) | ( n16136 & ~n16137 ) ;
  assign n16139 = ( ~n1517 & n5585 ) | ( ~n1517 & n14694 ) | ( n5585 & n14694 ) ;
  assign n16140 = ( x72 & n509 ) | ( x72 & ~n9966 ) | ( n509 & ~n9966 ) ;
  assign n16141 = ( ~n2122 & n7762 ) | ( ~n2122 & n15806 ) | ( n7762 & n15806 ) ;
  assign n16142 = n7621 ^ n5304 ^ n3112 ;
  assign n16143 = ( n765 & n4777 ) | ( n765 & ~n16142 ) | ( n4777 & ~n16142 ) ;
  assign n16144 = ( n11736 & n15575 ) | ( n11736 & n16143 ) | ( n15575 & n16143 ) ;
  assign n16145 = ( ~n11218 & n16141 ) | ( ~n11218 & n16144 ) | ( n16141 & n16144 ) ;
  assign n16146 = ( n2431 & n5630 ) | ( n2431 & ~n16145 ) | ( n5630 & ~n16145 ) ;
  assign n16147 = ( n16139 & ~n16140 ) | ( n16139 & n16146 ) | ( ~n16140 & n16146 ) ;
  assign n16151 = n3731 ^ n2050 ^ n2042 ;
  assign n16148 = ( n478 & ~n5450 ) | ( n478 & n12429 ) | ( ~n5450 & n12429 ) ;
  assign n16149 = n16148 ^ n8560 ^ n5450 ;
  assign n16150 = ( n5194 & n6468 ) | ( n5194 & n16149 ) | ( n6468 & n16149 ) ;
  assign n16152 = n16151 ^ n16150 ^ n2981 ;
  assign n16153 = n16152 ^ n7536 ^ n644 ;
  assign n16154 = n7349 ^ n6193 ^ n3693 ;
  assign n16155 = ( ~n6727 & n14476 ) | ( ~n6727 & n16154 ) | ( n14476 & n16154 ) ;
  assign n16156 = n16155 ^ n10012 ^ n4890 ;
  assign n16157 = ( n14186 & ~n16153 ) | ( n14186 & n16156 ) | ( ~n16153 & n16156 ) ;
  assign n16160 = n13276 ^ n8773 ^ n8427 ;
  assign n16161 = ( n8430 & n15304 ) | ( n8430 & ~n16160 ) | ( n15304 & ~n16160 ) ;
  assign n16158 = ( ~n3431 & n7198 ) | ( ~n3431 & n13795 ) | ( n7198 & n13795 ) ;
  assign n16159 = n16158 ^ n3254 ^ n3208 ;
  assign n16162 = n16161 ^ n16159 ^ n12999 ;
  assign n16163 = ( ~n7526 & n10387 ) | ( ~n7526 & n10965 ) | ( n10387 & n10965 ) ;
  assign n16164 = ( ~n1917 & n16015 ) | ( ~n1917 & n16163 ) | ( n16015 & n16163 ) ;
  assign n16165 = ( n11596 & n14329 ) | ( n11596 & n16164 ) | ( n14329 & n16164 ) ;
  assign n16166 = n16165 ^ n5731 ^ n5349 ;
  assign n16167 = n12182 ^ n5048 ^ n4044 ;
  assign n16168 = ( n275 & n2498 ) | ( n275 & ~n13064 ) | ( n2498 & ~n13064 ) ;
  assign n16169 = ( n13784 & ~n16167 ) | ( n13784 & n16168 ) | ( ~n16167 & n16168 ) ;
  assign n16170 = n16169 ^ n5194 ^ n3245 ;
  assign n16171 = n11331 ^ n9640 ^ n4795 ;
  assign n16172 = n16171 ^ n13488 ^ n1177 ;
  assign n16173 = n12312 ^ n4647 ^ n4025 ;
  assign n16174 = n5230 ^ n4114 ^ n2422 ;
  assign n16175 = n16174 ^ n3391 ^ n2117 ;
  assign n16176 = n16175 ^ n13000 ^ n4329 ;
  assign n16177 = n6167 ^ n4856 ^ n1735 ;
  assign n16178 = ( n255 & ~n1843 ) | ( n255 & n5023 ) | ( ~n1843 & n5023 ) ;
  assign n16179 = n16178 ^ n4637 ^ n1485 ;
  assign n16180 = ( n320 & ~n16177 ) | ( n320 & n16179 ) | ( ~n16177 & n16179 ) ;
  assign n16181 = n6057 ^ n3441 ^ n438 ;
  assign n16182 = ( n1666 & ~n11820 ) | ( n1666 & n16181 ) | ( ~n11820 & n16181 ) ;
  assign n16183 = ( n5312 & n5827 ) | ( n5312 & n13774 ) | ( n5827 & n13774 ) ;
  assign n16184 = ( n14613 & ~n16182 ) | ( n14613 & n16183 ) | ( ~n16182 & n16183 ) ;
  assign n16185 = n16184 ^ n15609 ^ n1165 ;
  assign n16188 = n4316 ^ n3336 ^ n193 ;
  assign n16187 = n15715 ^ n3770 ^ n3006 ;
  assign n16186 = ( n1367 & n5407 ) | ( n1367 & n8789 ) | ( n5407 & n8789 ) ;
  assign n16189 = n16188 ^ n16187 ^ n16186 ;
  assign n16190 = n16189 ^ n1996 ^ n1176 ;
  assign n16191 = n16190 ^ n14020 ^ n585 ;
  assign n16192 = ( ~n797 & n12130 ) | ( ~n797 & n13067 ) | ( n12130 & n13067 ) ;
  assign n16193 = ( n2956 & n5848 ) | ( n2956 & n15202 ) | ( n5848 & n15202 ) ;
  assign n16194 = n11456 ^ n3378 ^ n1015 ;
  assign n16195 = ( n9474 & n16193 ) | ( n9474 & ~n16194 ) | ( n16193 & ~n16194 ) ;
  assign n16196 = n14445 ^ n8334 ^ n1133 ;
  assign n16197 = n5840 ^ n5210 ^ n1025 ;
  assign n16198 = n14283 ^ n5069 ^ n3136 ;
  assign n16199 = ( n2599 & ~n16197 ) | ( n2599 & n16198 ) | ( ~n16197 & n16198 ) ;
  assign n16200 = n10650 ^ n10533 ^ n9764 ;
  assign n16201 = n6901 ^ n3997 ^ n1390 ;
  assign n16202 = n15834 ^ n9401 ^ n158 ;
  assign n16203 = ( n2921 & n11162 ) | ( n2921 & ~n16202 ) | ( n11162 & ~n16202 ) ;
  assign n16204 = n4487 ^ n4264 ^ n2953 ;
  assign n16205 = ( ~n1122 & n4603 ) | ( ~n1122 & n16204 ) | ( n4603 & n16204 ) ;
  assign n16206 = ( n726 & n3304 ) | ( n726 & n3645 ) | ( n3304 & n3645 ) ;
  assign n16207 = ( n3791 & n6660 ) | ( n3791 & ~n16206 ) | ( n6660 & ~n16206 ) ;
  assign n16208 = ( n12860 & n16205 ) | ( n12860 & ~n16207 ) | ( n16205 & ~n16207 ) ;
  assign n16209 = n16208 ^ n5876 ^ n3928 ;
  assign n16210 = ( n3103 & n6760 ) | ( n3103 & n13280 ) | ( n6760 & n13280 ) ;
  assign n16211 = ( n389 & n1997 ) | ( n389 & ~n15843 ) | ( n1997 & ~n15843 ) ;
  assign n16212 = ( n733 & ~n9104 ) | ( n733 & n16211 ) | ( ~n9104 & n16211 ) ;
  assign n16213 = n10614 ^ n2229 ^ n2167 ;
  assign n16214 = n16213 ^ n12205 ^ n8805 ;
  assign n16215 = n16214 ^ n11062 ^ n2210 ;
  assign n16218 = ( n3142 & ~n4380 ) | ( n3142 & n11318 ) | ( ~n4380 & n11318 ) ;
  assign n16219 = n16218 ^ n8038 ^ n7012 ;
  assign n16220 = n16219 ^ n14091 ^ n3627 ;
  assign n16216 = ( n8892 & n9612 ) | ( n8892 & n14506 ) | ( n9612 & n14506 ) ;
  assign n16217 = n16216 ^ n6898 ^ n5782 ;
  assign n16221 = n16220 ^ n16217 ^ n6443 ;
  assign n16232 = n7896 ^ n3957 ^ n1006 ;
  assign n16231 = n4579 ^ n1230 ^ n196 ;
  assign n16229 = ( n2228 & n5099 ) | ( n2228 & n7481 ) | ( n5099 & n7481 ) ;
  assign n16227 = ( n992 & ~n2928 ) | ( n992 & n3678 ) | ( ~n2928 & n3678 ) ;
  assign n16228 = ( n2422 & n4746 ) | ( n2422 & ~n16227 ) | ( n4746 & ~n16227 ) ;
  assign n16225 = ( n589 & n1880 ) | ( n589 & n12278 ) | ( n1880 & n12278 ) ;
  assign n16226 = n16225 ^ n11668 ^ n6702 ;
  assign n16230 = n16229 ^ n16228 ^ n16226 ;
  assign n16233 = n16232 ^ n16231 ^ n16230 ;
  assign n16222 = n12485 ^ n11544 ^ n4579 ;
  assign n16223 = ( n2295 & n4229 ) | ( n2295 & n16222 ) | ( n4229 & n16222 ) ;
  assign n16224 = ( ~n6039 & n7245 ) | ( ~n6039 & n16223 ) | ( n7245 & n16223 ) ;
  assign n16234 = n16233 ^ n16224 ^ n9831 ;
  assign n16235 = ( n3722 & n3912 ) | ( n3722 & ~n5818 ) | ( n3912 & ~n5818 ) ;
  assign n16239 = ( ~x37 & n3484 ) | ( ~x37 & n12676 ) | ( n3484 & n12676 ) ;
  assign n16240 = ( n1596 & ~n2130 ) | ( n1596 & n16239 ) | ( ~n2130 & n16239 ) ;
  assign n16236 = ( ~n2638 & n6819 ) | ( ~n2638 & n9357 ) | ( n6819 & n9357 ) ;
  assign n16237 = ( n1915 & ~n6512 ) | ( n1915 & n16236 ) | ( ~n6512 & n16236 ) ;
  assign n16238 = ( ~n8892 & n12701 ) | ( ~n8892 & n16237 ) | ( n12701 & n16237 ) ;
  assign n16241 = n16240 ^ n16238 ^ n10153 ;
  assign n16242 = ( n7449 & n16235 ) | ( n7449 & n16241 ) | ( n16235 & n16241 ) ;
  assign n16243 = ( n894 & n11378 ) | ( n894 & ~n11765 ) | ( n11378 & ~n11765 ) ;
  assign n16244 = n16243 ^ n12233 ^ n1496 ;
  assign n16245 = ( n3424 & n7648 ) | ( n3424 & n16244 ) | ( n7648 & n16244 ) ;
  assign n16246 = n7214 ^ n1338 ^ n262 ;
  assign n16248 = ( ~n428 & n3650 ) | ( ~n428 & n4646 ) | ( n3650 & n4646 ) ;
  assign n16249 = ( n5830 & ~n7178 ) | ( n5830 & n16248 ) | ( ~n7178 & n16248 ) ;
  assign n16247 = ( ~n5375 & n8209 ) | ( ~n5375 & n15204 ) | ( n8209 & n15204 ) ;
  assign n16250 = n16249 ^ n16247 ^ n1701 ;
  assign n16251 = ( n1185 & n4161 ) | ( n1185 & ~n16143 ) | ( n4161 & ~n16143 ) ;
  assign n16255 = n11594 ^ n8828 ^ n616 ;
  assign n16256 = n16255 ^ n11504 ^ n8566 ;
  assign n16254 = ( ~n3134 & n12900 ) | ( ~n3134 & n14269 ) | ( n12900 & n14269 ) ;
  assign n16252 = ( ~n5811 & n6698 ) | ( ~n5811 & n10219 ) | ( n6698 & n10219 ) ;
  assign n16253 = ( n8026 & n12544 ) | ( n8026 & ~n16252 ) | ( n12544 & ~n16252 ) ;
  assign n16257 = n16256 ^ n16254 ^ n16253 ;
  assign n16258 = n6561 ^ n4166 ^ n1002 ;
  assign n16259 = ( n3663 & n8534 ) | ( n3663 & ~n16258 ) | ( n8534 & ~n16258 ) ;
  assign n16260 = ( n15114 & n16257 ) | ( n15114 & n16259 ) | ( n16257 & n16259 ) ;
  assign n16261 = n9972 ^ n5759 ^ n1605 ;
  assign n16262 = n16261 ^ n13735 ^ n10555 ;
  assign n16263 = ( n2369 & ~n4110 ) | ( n2369 & n7340 ) | ( ~n4110 & n7340 ) ;
  assign n16264 = ( ~n2966 & n4185 ) | ( ~n2966 & n4462 ) | ( n4185 & n4462 ) ;
  assign n16265 = ( n1366 & ~n1428 ) | ( n1366 & n16264 ) | ( ~n1428 & n16264 ) ;
  assign n16266 = ( x54 & n472 ) | ( x54 & n4651 ) | ( n472 & n4651 ) ;
  assign n16267 = ( n4035 & n7767 ) | ( n4035 & n16266 ) | ( n7767 & n16266 ) ;
  assign n16268 = n6702 ^ n6506 ^ n5297 ;
  assign n16269 = ( ~n2589 & n4542 ) | ( ~n2589 & n16268 ) | ( n4542 & n16268 ) ;
  assign n16270 = ( ~n1814 & n3165 ) | ( ~n1814 & n9915 ) | ( n3165 & n9915 ) ;
  assign n16271 = n16270 ^ n7578 ^ n3344 ;
  assign n16272 = ( ~n3669 & n15767 ) | ( ~n3669 & n16271 ) | ( n15767 & n16271 ) ;
  assign n16273 = ( n2038 & ~n4599 ) | ( n2038 & n16272 ) | ( ~n4599 & n16272 ) ;
  assign n16275 = n8222 ^ n1181 ^ n764 ;
  assign n16274 = ( n1357 & ~n7821 ) | ( n1357 & n9988 ) | ( ~n7821 & n9988 ) ;
  assign n16276 = n16275 ^ n16274 ^ n986 ;
  assign n16277 = n16276 ^ n14890 ^ n2934 ;
  assign n16278 = ( n3622 & n12834 ) | ( n3622 & ~n13146 ) | ( n12834 & ~n13146 ) ;
  assign n16279 = n16278 ^ n15826 ^ n9776 ;
  assign n16280 = ( ~n665 & n1719 ) | ( ~n665 & n3816 ) | ( n1719 & n3816 ) ;
  assign n16281 = n16280 ^ n5206 ^ n3327 ;
  assign n16282 = n16281 ^ n2269 ^ n1607 ;
  assign n16283 = ( ~n1730 & n6652 ) | ( ~n1730 & n16282 ) | ( n6652 & n16282 ) ;
  assign n16293 = ( ~n444 & n2829 ) | ( ~n444 & n10031 ) | ( n2829 & n10031 ) ;
  assign n16294 = n16293 ^ n8775 ^ n5691 ;
  assign n16291 = n12908 ^ n4589 ^ n1446 ;
  assign n16286 = n7187 ^ n5357 ^ n1027 ;
  assign n16287 = ( n301 & n11052 ) | ( n301 & n16286 ) | ( n11052 & n16286 ) ;
  assign n16288 = ( n3577 & n5464 ) | ( n3577 & ~n16287 ) | ( n5464 & ~n16287 ) ;
  assign n16284 = n12862 ^ n7688 ^ n6387 ;
  assign n16285 = n16284 ^ n8042 ^ n2765 ;
  assign n16289 = n16288 ^ n16285 ^ n7094 ;
  assign n16290 = ( n7534 & n9298 ) | ( n7534 & ~n16289 ) | ( n9298 & ~n16289 ) ;
  assign n16292 = n16291 ^ n16290 ^ n1274 ;
  assign n16295 = n16294 ^ n16292 ^ n15234 ;
  assign n16297 = n6302 ^ n5448 ^ n4504 ;
  assign n16296 = ( n3758 & n6424 ) | ( n3758 & ~n12301 ) | ( n6424 & ~n12301 ) ;
  assign n16298 = n16297 ^ n16296 ^ n15220 ;
  assign n16303 = n6309 ^ n3640 ^ n1378 ;
  assign n16304 = ( n6830 & n15883 ) | ( n6830 & ~n16303 ) | ( n15883 & ~n16303 ) ;
  assign n16299 = ( n592 & n1557 ) | ( n592 & ~n13375 ) | ( n1557 & ~n13375 ) ;
  assign n16300 = ( n1067 & n1796 ) | ( n1067 & n8453 ) | ( n1796 & n8453 ) ;
  assign n16301 = ( n13191 & n16299 ) | ( n13191 & ~n16300 ) | ( n16299 & ~n16300 ) ;
  assign n16302 = ( n3051 & n5436 ) | ( n3051 & n16301 ) | ( n5436 & n16301 ) ;
  assign n16305 = n16304 ^ n16302 ^ n10790 ;
  assign n16306 = n14548 ^ n10708 ^ n7078 ;
  assign n16307 = ( n1321 & ~n6865 ) | ( n1321 & n16306 ) | ( ~n6865 & n16306 ) ;
  assign n16308 = n10843 ^ n4510 ^ n1627 ;
  assign n16309 = n16308 ^ n11542 ^ n3369 ;
  assign n16314 = n7669 ^ n3739 ^ n1972 ;
  assign n16312 = n6148 ^ n5684 ^ n3154 ;
  assign n16310 = ( n797 & ~n2725 ) | ( n797 & n4804 ) | ( ~n2725 & n4804 ) ;
  assign n16311 = ( n7532 & ~n10737 ) | ( n7532 & n16310 ) | ( ~n10737 & n16310 ) ;
  assign n16313 = n16312 ^ n16311 ^ n1417 ;
  assign n16315 = n16314 ^ n16313 ^ n9203 ;
  assign n16316 = ( n2351 & ~n4683 ) | ( n2351 & n13555 ) | ( ~n4683 & n13555 ) ;
  assign n16317 = ( ~x70 & n7077 ) | ( ~x70 & n16316 ) | ( n7077 & n16316 ) ;
  assign n16318 = ( n8214 & n9267 ) | ( n8214 & ~n11011 ) | ( n9267 & ~n11011 ) ;
  assign n16319 = ( n6177 & n12239 ) | ( n6177 & n16318 ) | ( n12239 & n16318 ) ;
  assign n16320 = ( n1708 & n6688 ) | ( n1708 & n16319 ) | ( n6688 & n16319 ) ;
  assign n16321 = ( ~n2876 & n3964 ) | ( ~n2876 & n10200 ) | ( n3964 & n10200 ) ;
  assign n16322 = ( ~n3611 & n7056 ) | ( ~n3611 & n10131 ) | ( n7056 & n10131 ) ;
  assign n16323 = n3509 ^ n732 ^ n473 ;
  assign n16324 = ( ~n10311 & n12667 ) | ( ~n10311 & n16323 ) | ( n12667 & n16323 ) ;
  assign n16340 = n7370 ^ n5567 ^ n218 ;
  assign n16341 = n16340 ^ n7509 ^ n6642 ;
  assign n16339 = n14384 ^ n11355 ^ n3720 ;
  assign n16337 = n13501 ^ n2724 ^ n282 ;
  assign n16335 = n9006 ^ n3627 ^ n2058 ;
  assign n16336 = ( n1088 & n1236 ) | ( n1088 & ~n16335 ) | ( n1236 & ~n16335 ) ;
  assign n16325 = n15526 ^ n5409 ^ n1397 ;
  assign n16326 = ( ~n3314 & n5843 ) | ( ~n3314 & n16325 ) | ( n5843 & n16325 ) ;
  assign n16327 = n9316 ^ n6499 ^ n3041 ;
  assign n16328 = ( ~n2861 & n16326 ) | ( ~n2861 & n16327 ) | ( n16326 & n16327 ) ;
  assign n16331 = n6049 ^ n2633 ^ n986 ;
  assign n16332 = ( n717 & ~n9006 ) | ( n717 & n16331 ) | ( ~n9006 & n16331 ) ;
  assign n16329 = n10346 ^ n8506 ^ n6681 ;
  assign n16330 = ( n6216 & n12473 ) | ( n6216 & n16329 ) | ( n12473 & n16329 ) ;
  assign n16333 = n16332 ^ n16330 ^ n3723 ;
  assign n16334 = ( ~n5316 & n16328 ) | ( ~n5316 & n16333 ) | ( n16328 & n16333 ) ;
  assign n16338 = n16337 ^ n16336 ^ n16334 ;
  assign n16342 = n16341 ^ n16339 ^ n16338 ;
  assign n16343 = ( n3238 & ~n7851 ) | ( n3238 & n11023 ) | ( ~n7851 & n11023 ) ;
  assign n16344 = ( n10573 & ~n15917 ) | ( n10573 & n16343 ) | ( ~n15917 & n16343 ) ;
  assign n16346 = ( n1241 & ~n3731 ) | ( n1241 & n14942 ) | ( ~n3731 & n14942 ) ;
  assign n16345 = ( n448 & ~n7856 ) | ( n448 & n7990 ) | ( ~n7856 & n7990 ) ;
  assign n16347 = n16346 ^ n16345 ^ n14264 ;
  assign n16348 = ( n4288 & n9094 ) | ( n4288 & n10442 ) | ( n9094 & n10442 ) ;
  assign n16349 = ( ~n1051 & n4594 ) | ( ~n1051 & n16348 ) | ( n4594 & n16348 ) ;
  assign n16350 = ( n1531 & n13553 ) | ( n1531 & ~n16349 ) | ( n13553 & ~n16349 ) ;
  assign n16351 = ( n1411 & n2285 ) | ( n1411 & n14323 ) | ( n2285 & n14323 ) ;
  assign n16352 = n2930 ^ n2466 ^ n1268 ;
  assign n16355 = ( ~n342 & n3940 ) | ( ~n342 & n5604 ) | ( n3940 & n5604 ) ;
  assign n16353 = n6195 ^ n3483 ^ n2210 ;
  assign n16354 = ( n2160 & n12052 ) | ( n2160 & ~n16353 ) | ( n12052 & ~n16353 ) ;
  assign n16356 = n16355 ^ n16354 ^ n6754 ;
  assign n16357 = ( n1558 & ~n7768 ) | ( n1558 & n16356 ) | ( ~n7768 & n16356 ) ;
  assign n16358 = ( n11481 & ~n16352 ) | ( n11481 & n16357 ) | ( ~n16352 & n16357 ) ;
  assign n16359 = n16358 ^ n6208 ^ n4855 ;
  assign n16360 = ( ~n11632 & n12906 ) | ( ~n11632 & n16359 ) | ( n12906 & n16359 ) ;
  assign n16361 = ( n1397 & n3034 ) | ( n1397 & ~n4368 ) | ( n3034 & ~n4368 ) ;
  assign n16362 = ( n1936 & n4228 ) | ( n1936 & n5415 ) | ( n4228 & n5415 ) ;
  assign n16363 = ( n11723 & n16361 ) | ( n11723 & ~n16362 ) | ( n16361 & ~n16362 ) ;
  assign n16364 = ( n5440 & n10933 ) | ( n5440 & ~n14803 ) | ( n10933 & ~n14803 ) ;
  assign n16365 = ( n808 & n12688 ) | ( n808 & ~n16364 ) | ( n12688 & ~n16364 ) ;
  assign n16366 = ( x110 & n6473 ) | ( x110 & n13422 ) | ( n6473 & n13422 ) ;
  assign n16367 = n16366 ^ n6424 ^ n3120 ;
  assign n16370 = n5548 ^ n3270 ^ n716 ;
  assign n16369 = ( n612 & n4570 ) | ( n612 & ~n9076 ) | ( n4570 & ~n9076 ) ;
  assign n16368 = ( n4886 & n5671 ) | ( n4886 & ~n14419 ) | ( n5671 & ~n14419 ) ;
  assign n16371 = n16370 ^ n16369 ^ n16368 ;
  assign n16372 = ( n134 & n2563 ) | ( n134 & n2924 ) | ( n2563 & n2924 ) ;
  assign n16373 = ( n1219 & n15953 ) | ( n1219 & n16372 ) | ( n15953 & n16372 ) ;
  assign n16374 = n16373 ^ n12732 ^ n9330 ;
  assign n16375 = ( ~n3525 & n16371 ) | ( ~n3525 & n16374 ) | ( n16371 & n16374 ) ;
  assign n16376 = ( ~n4119 & n6030 ) | ( ~n4119 & n10297 ) | ( n6030 & n10297 ) ;
  assign n16377 = n16376 ^ n13023 ^ n10168 ;
  assign n16379 = n3714 ^ n3015 ^ n1549 ;
  assign n16378 = ( x80 & n6384 ) | ( x80 & n15045 ) | ( n6384 & n15045 ) ;
  assign n16380 = n16379 ^ n16378 ^ n15560 ;
  assign n16381 = ( n856 & n6987 ) | ( n856 & n16076 ) | ( n6987 & n16076 ) ;
  assign n16385 = ( x53 & ~n4546 ) | ( x53 & n10962 ) | ( ~n4546 & n10962 ) ;
  assign n16383 = n11429 ^ n1117 ^ x20 ;
  assign n16384 = ( n3326 & ~n3971 ) | ( n3326 & n16383 ) | ( ~n3971 & n16383 ) ;
  assign n16382 = ( n2032 & ~n10972 ) | ( n2032 & n14091 ) | ( ~n10972 & n14091 ) ;
  assign n16386 = n16385 ^ n16384 ^ n16382 ;
  assign n16387 = ( n12046 & ~n16381 ) | ( n12046 & n16386 ) | ( ~n16381 & n16386 ) ;
  assign n16388 = n6864 ^ n3687 ^ n655 ;
  assign n16389 = n13529 ^ n3093 ^ n1954 ;
  assign n16390 = ( n3827 & n16388 ) | ( n3827 & ~n16389 ) | ( n16388 & ~n16389 ) ;
  assign n16391 = ( n12713 & n16387 ) | ( n12713 & n16390 ) | ( n16387 & n16390 ) ;
  assign n16392 = ( ~n850 & n4354 ) | ( ~n850 & n16391 ) | ( n4354 & n16391 ) ;
  assign n16393 = n10017 ^ n9043 ^ n7276 ;
  assign n16394 = n16393 ^ n8919 ^ n1024 ;
  assign n16395 = n16394 ^ n11922 ^ n9432 ;
  assign n16396 = ( n11300 & ~n14338 ) | ( n11300 & n15486 ) | ( ~n14338 & n15486 ) ;
  assign n16397 = ( n1802 & n1916 ) | ( n1802 & ~n2099 ) | ( n1916 & ~n2099 ) ;
  assign n16398 = ( ~n6262 & n13654 ) | ( ~n6262 & n16397 ) | ( n13654 & n16397 ) ;
  assign n16399 = ( ~n6516 & n15367 ) | ( ~n6516 & n16398 ) | ( n15367 & n16398 ) ;
  assign n16400 = n14979 ^ n12102 ^ n11001 ;
  assign n16401 = ( n3271 & ~n3711 ) | ( n3271 & n11040 ) | ( ~n3711 & n11040 ) ;
  assign n16402 = n10276 ^ n9876 ^ n4982 ;
  assign n16403 = n11672 ^ n6387 ^ x29 ;
  assign n16404 = ( n10788 & n15832 ) | ( n10788 & ~n16403 ) | ( n15832 & ~n16403 ) ;
  assign n16405 = ( n16401 & n16402 ) | ( n16401 & n16404 ) | ( n16402 & n16404 ) ;
  assign n16415 = n7153 ^ n5836 ^ n1172 ;
  assign n16416 = ( n3069 & ~n5824 ) | ( n3069 & n16415 ) | ( ~n5824 & n16415 ) ;
  assign n16411 = ( n1819 & n3325 ) | ( n1819 & n12965 ) | ( n3325 & n12965 ) ;
  assign n16412 = ( n2427 & n10127 ) | ( n2427 & n16411 ) | ( n10127 & n16411 ) ;
  assign n16410 = n11326 ^ n10829 ^ n3242 ;
  assign n16413 = n16412 ^ n16410 ^ n12241 ;
  assign n16409 = n14311 ^ n6002 ^ n4622 ;
  assign n16414 = n16413 ^ n16409 ^ n6720 ;
  assign n16417 = n16416 ^ n16414 ^ n2407 ;
  assign n16406 = n12431 ^ n7414 ^ n721 ;
  assign n16407 = ( ~n3452 & n7924 ) | ( ~n3452 & n16406 ) | ( n7924 & n16406 ) ;
  assign n16408 = ( ~n8460 & n8655 ) | ( ~n8460 & n16407 ) | ( n8655 & n16407 ) ;
  assign n16418 = n16417 ^ n16408 ^ n10845 ;
  assign n16421 = n8065 ^ n5572 ^ n3753 ;
  assign n16422 = n16421 ^ n13566 ^ n5594 ;
  assign n16419 = ( n4204 & ~n6513 ) | ( n4204 & n11703 ) | ( ~n6513 & n11703 ) ;
  assign n16420 = n16419 ^ n12022 ^ n10756 ;
  assign n16423 = n16422 ^ n16420 ^ n11061 ;
  assign n16424 = n16423 ^ n13298 ^ n10755 ;
  assign n16428 = n8896 ^ n8486 ^ n1058 ;
  assign n16427 = n9670 ^ n9163 ^ x99 ;
  assign n16429 = n16428 ^ n16427 ^ n10619 ;
  assign n16426 = n11551 ^ n8941 ^ n6386 ;
  assign n16425 = ( n267 & ~n12335 ) | ( n267 & n12682 ) | ( ~n12335 & n12682 ) ;
  assign n16430 = n16429 ^ n16426 ^ n16425 ;
  assign n16439 = n16047 ^ n10374 ^ n1075 ;
  assign n16440 = n16439 ^ n11654 ^ n11240 ;
  assign n16433 = n3678 ^ n2098 ^ n1819 ;
  assign n16434 = ( n5623 & n10525 ) | ( n5623 & ~n16433 ) | ( n10525 & ~n16433 ) ;
  assign n16435 = ( n4321 & n8140 ) | ( n4321 & n8381 ) | ( n8140 & n8381 ) ;
  assign n16436 = ( n5044 & ~n5803 ) | ( n5044 & n16435 ) | ( ~n5803 & n16435 ) ;
  assign n16437 = n16436 ^ n6545 ^ n2197 ;
  assign n16438 = ( n7784 & n16434 ) | ( n7784 & ~n16437 ) | ( n16434 & ~n16437 ) ;
  assign n16431 = n5379 ^ n4947 ^ n684 ;
  assign n16432 = n16431 ^ n14829 ^ n11565 ;
  assign n16441 = n16440 ^ n16438 ^ n16432 ;
  assign n16443 = ( n1515 & n7927 ) | ( n1515 & n9967 ) | ( n7927 & n9967 ) ;
  assign n16444 = n1155 ^ n789 ^ x110 ;
  assign n16445 = n16444 ^ n2550 ^ n937 ;
  assign n16446 = n16445 ^ n10914 ^ n2280 ;
  assign n16447 = n16446 ^ n15560 ^ n9369 ;
  assign n16448 = ( n1436 & n4555 ) | ( n1436 & ~n14044 ) | ( n4555 & ~n14044 ) ;
  assign n16449 = ( n16443 & n16447 ) | ( n16443 & n16448 ) | ( n16447 & n16448 ) ;
  assign n16442 = ( n896 & ~n6145 ) | ( n896 & n8515 ) | ( ~n6145 & n8515 ) ;
  assign n16450 = n16449 ^ n16442 ^ n14864 ;
  assign n16451 = ( n2214 & n8340 ) | ( n2214 & ~n13412 ) | ( n8340 & ~n13412 ) ;
  assign n16452 = ( n12148 & n13463 ) | ( n12148 & n16451 ) | ( n13463 & n16451 ) ;
  assign n16454 = ( ~n4833 & n6486 ) | ( ~n4833 & n15062 ) | ( n6486 & n15062 ) ;
  assign n16453 = n15895 ^ n13168 ^ n6753 ;
  assign n16455 = n16454 ^ n16453 ^ n2726 ;
  assign n16456 = ( n859 & ~n2541 ) | ( n859 & n3523 ) | ( ~n2541 & n3523 ) ;
  assign n16457 = n16456 ^ n4194 ^ n2585 ;
  assign n16460 = n7109 ^ n5408 ^ n1668 ;
  assign n16458 = ( ~n142 & n3722 ) | ( ~n142 & n6883 ) | ( n3722 & n6883 ) ;
  assign n16459 = n16458 ^ n16293 ^ n6216 ;
  assign n16461 = n16460 ^ n16459 ^ n5003 ;
  assign n16462 = n16369 ^ n10419 ^ n1020 ;
  assign n16463 = n16462 ^ n13761 ^ n3626 ;
  assign n16464 = n16463 ^ n11027 ^ n6708 ;
  assign n16465 = n16464 ^ n13322 ^ n887 ;
  assign n16466 = ( n6239 & n7869 ) | ( n6239 & n11283 ) | ( n7869 & n11283 ) ;
  assign n16467 = ( n5474 & ~n11967 ) | ( n5474 & n16466 ) | ( ~n11967 & n16466 ) ;
  assign n16468 = n3444 ^ n1279 ^ n962 ;
  assign n16469 = ( ~n2140 & n11468 ) | ( ~n2140 & n12535 ) | ( n11468 & n12535 ) ;
  assign n16470 = ( n5627 & n16468 ) | ( n5627 & ~n16469 ) | ( n16468 & ~n16469 ) ;
  assign n16481 = n9076 ^ n6432 ^ n4466 ;
  assign n16482 = ( ~n3909 & n11350 ) | ( ~n3909 & n16481 ) | ( n11350 & n16481 ) ;
  assign n16479 = n9058 ^ n5524 ^ n2152 ;
  assign n16480 = ( n5231 & n12780 ) | ( n5231 & n16479 ) | ( n12780 & n16479 ) ;
  assign n16483 = n16482 ^ n16480 ^ n9667 ;
  assign n16477 = ( n720 & n9144 ) | ( n720 & n10831 ) | ( n9144 & n10831 ) ;
  assign n16478 = ( n12846 & ~n14510 ) | ( n12846 & n16477 ) | ( ~n14510 & n16477 ) ;
  assign n16475 = ( n4515 & n5798 ) | ( n4515 & n10622 ) | ( n5798 & n10622 ) ;
  assign n16473 = n7432 ^ n2137 ^ n773 ;
  assign n16471 = n5381 ^ n3529 ^ n1397 ;
  assign n16472 = n16471 ^ n4647 ^ n426 ;
  assign n16474 = n16473 ^ n16472 ^ n10545 ;
  assign n16476 = n16475 ^ n16474 ^ n12311 ;
  assign n16484 = n16483 ^ n16478 ^ n16476 ;
  assign n16492 = n11596 ^ n4919 ^ x105 ;
  assign n16493 = n16492 ^ n10814 ^ n8236 ;
  assign n16485 = n10872 ^ n6550 ^ n2582 ;
  assign n16486 = n16485 ^ n5284 ^ n3479 ;
  assign n16487 = n16228 ^ n11110 ^ n436 ;
  assign n16488 = ( n1138 & n11207 ) | ( n1138 & ~n16487 ) | ( n11207 & ~n16487 ) ;
  assign n16489 = ( ~n922 & n16486 ) | ( ~n922 & n16488 ) | ( n16486 & n16488 ) ;
  assign n16490 = n14940 ^ n11334 ^ n6484 ;
  assign n16491 = ( n5950 & ~n16489 ) | ( n5950 & n16490 ) | ( ~n16489 & n16490 ) ;
  assign n16494 = n16493 ^ n16491 ^ n12450 ;
  assign n16495 = n6786 ^ n2198 ^ n273 ;
  assign n16496 = n16495 ^ n7683 ^ n4016 ;
  assign n16497 = n16496 ^ n10608 ^ n3319 ;
  assign n16502 = ( n3887 & n9943 ) | ( n3887 & n10465 ) | ( n9943 & n10465 ) ;
  assign n16498 = n8327 ^ n5330 ^ n3677 ;
  assign n16499 = ( n961 & n4008 ) | ( n961 & n5830 ) | ( n4008 & n5830 ) ;
  assign n16500 = ( n1223 & n16498 ) | ( n1223 & n16499 ) | ( n16498 & n16499 ) ;
  assign n16501 = n16500 ^ n9330 ^ n6215 ;
  assign n16503 = n16502 ^ n16501 ^ n8566 ;
  assign n16505 = ( ~n3943 & n7937 ) | ( ~n3943 & n12271 ) | ( n7937 & n12271 ) ;
  assign n16504 = n16041 ^ n12784 ^ n298 ;
  assign n16506 = n16505 ^ n16504 ^ n4806 ;
  assign n16507 = n12754 ^ n7422 ^ n4673 ;
  assign n16508 = ( n3582 & n9970 ) | ( n3582 & ~n16507 ) | ( n9970 & ~n16507 ) ;
  assign n16509 = n10670 ^ n7809 ^ n1095 ;
  assign n16510 = ( n221 & n11077 ) | ( n221 & ~n16509 ) | ( n11077 & ~n16509 ) ;
  assign n16511 = n16510 ^ n3748 ^ n1153 ;
  assign n16512 = ( n2780 & ~n4157 ) | ( n2780 & n16511 ) | ( ~n4157 & n16511 ) ;
  assign n16513 = n16512 ^ n11477 ^ n1380 ;
  assign n16514 = ( n3780 & n16366 ) | ( n3780 & ~n16513 ) | ( n16366 & ~n16513 ) ;
  assign n16519 = ( ~n2717 & n5472 ) | ( ~n2717 & n13663 ) | ( n5472 & n13663 ) ;
  assign n16520 = ( ~n4045 & n6217 ) | ( ~n4045 & n16519 ) | ( n6217 & n16519 ) ;
  assign n16521 = ( n8403 & n9789 ) | ( n8403 & n16520 ) | ( n9789 & n16520 ) ;
  assign n16515 = ( n591 & ~n1431 ) | ( n591 & n14436 ) | ( ~n1431 & n14436 ) ;
  assign n16516 = ( n1972 & ~n4777 ) | ( n1972 & n8266 ) | ( ~n4777 & n8266 ) ;
  assign n16517 = ( ~n640 & n16515 ) | ( ~n640 & n16516 ) | ( n16515 & n16516 ) ;
  assign n16518 = ( n2725 & n9134 ) | ( n2725 & ~n16517 ) | ( n9134 & ~n16517 ) ;
  assign n16522 = n16521 ^ n16518 ^ n3447 ;
  assign n16526 = n15264 ^ n12661 ^ n3018 ;
  assign n16527 = ( n3395 & n4816 ) | ( n3395 & n16526 ) | ( n4816 & n16526 ) ;
  assign n16525 = n13341 ^ n9186 ^ n5923 ;
  assign n16523 = n9914 ^ n3423 ^ n3371 ;
  assign n16524 = ( n7277 & ~n7980 ) | ( n7277 & n16523 ) | ( ~n7980 & n16523 ) ;
  assign n16528 = n16527 ^ n16525 ^ n16524 ;
  assign n16529 = n13976 ^ n5128 ^ n1820 ;
  assign n16530 = n8501 ^ n1996 ^ n1053 ;
  assign n16531 = n16530 ^ n4876 ^ n3277 ;
  assign n16532 = ( ~n3530 & n5068 ) | ( ~n3530 & n16531 ) | ( n5068 & n16531 ) ;
  assign n16533 = n4582 ^ n3652 ^ n1298 ;
  assign n16534 = ( n7926 & ~n9612 ) | ( n7926 & n16533 ) | ( ~n9612 & n16533 ) ;
  assign n16535 = ( ~n3917 & n11112 ) | ( ~n3917 & n16534 ) | ( n11112 & n16534 ) ;
  assign n16536 = n16535 ^ n8132 ^ n7019 ;
  assign n16537 = n9226 ^ n7569 ^ n4444 ;
  assign n16538 = ( ~n7374 & n8043 ) | ( ~n7374 & n16537 ) | ( n8043 & n16537 ) ;
  assign n16539 = n14391 ^ n3329 ^ x89 ;
  assign n16540 = n16539 ^ n12667 ^ n10998 ;
  assign n16541 = ( n6728 & n8975 ) | ( n6728 & ~n16540 ) | ( n8975 & ~n16540 ) ;
  assign n16542 = n13998 ^ n7211 ^ n5108 ;
  assign n16543 = n16542 ^ n9986 ^ n1062 ;
  assign n16544 = n13745 ^ n9550 ^ n6728 ;
  assign n16545 = n16544 ^ n12635 ^ n12079 ;
  assign n16546 = ( n4798 & ~n8238 ) | ( n4798 & n16545 ) | ( ~n8238 & n16545 ) ;
  assign n16547 = n16546 ^ n9746 ^ n7898 ;
  assign n16548 = ( ~n905 & n1016 ) | ( ~n905 & n8932 ) | ( n1016 & n8932 ) ;
  assign n16549 = n16548 ^ n6293 ^ n3412 ;
  assign n16550 = ( ~n5356 & n11239 ) | ( ~n5356 & n16549 ) | ( n11239 & n16549 ) ;
  assign n16554 = ( n2835 & n2902 ) | ( n2835 & ~n3600 ) | ( n2902 & ~n3600 ) ;
  assign n16551 = ( ~n8383 & n11003 ) | ( ~n8383 & n12901 ) | ( n11003 & n12901 ) ;
  assign n16552 = ( n5631 & ~n8370 ) | ( n5631 & n16551 ) | ( ~n8370 & n16551 ) ;
  assign n16553 = ( n2073 & ~n8302 ) | ( n2073 & n16552 ) | ( ~n8302 & n16552 ) ;
  assign n16555 = n16554 ^ n16553 ^ n11967 ;
  assign n16556 = n16555 ^ n8673 ^ n4590 ;
  assign n16557 = n5324 ^ n4002 ^ x103 ;
  assign n16558 = ( n1369 & n9937 ) | ( n1369 & ~n16557 ) | ( n9937 & ~n16557 ) ;
  assign n16559 = n16558 ^ n14187 ^ n9033 ;
  assign n16560 = ( n3713 & ~n5782 ) | ( n3713 & n16518 ) | ( ~n5782 & n16518 ) ;
  assign n16565 = ( n3017 & ~n7253 ) | ( n3017 & n15212 ) | ( ~n7253 & n15212 ) ;
  assign n16563 = ( n132 & n2827 ) | ( n132 & ~n3336 ) | ( n2827 & ~n3336 ) ;
  assign n16564 = ( ~n2601 & n4787 ) | ( ~n2601 & n16563 ) | ( n4787 & n16563 ) ;
  assign n16561 = n8288 ^ n6618 ^ n2872 ;
  assign n16562 = ( n4037 & n14405 ) | ( n4037 & n16561 ) | ( n14405 & n16561 ) ;
  assign n16566 = n16565 ^ n16564 ^ n16562 ;
  assign n16567 = ( n8996 & ~n10963 ) | ( n8996 & n13304 ) | ( ~n10963 & n13304 ) ;
  assign n16568 = ( ~n7067 & n13288 ) | ( ~n7067 & n14952 ) | ( n13288 & n14952 ) ;
  assign n16569 = ( ~n1249 & n1530 ) | ( ~n1249 & n16241 ) | ( n1530 & n16241 ) ;
  assign n16570 = n13049 ^ n3219 ^ n2945 ;
  assign n16573 = ( n1165 & n6867 ) | ( n1165 & ~n14788 ) | ( n6867 & ~n14788 ) ;
  assign n16572 = ( ~n1148 & n2279 ) | ( ~n1148 & n2457 ) | ( n2279 & n2457 ) ;
  assign n16574 = n16573 ^ n16572 ^ n10242 ;
  assign n16571 = n9408 ^ n1447 ^ n1019 ;
  assign n16575 = n16574 ^ n16571 ^ n5620 ;
  assign n16576 = ( n1304 & n7349 ) | ( n1304 & ~n16555 ) | ( n7349 & ~n16555 ) ;
  assign n16577 = n13789 ^ n7116 ^ n1933 ;
  assign n16578 = ( ~n5723 & n6170 ) | ( ~n5723 & n16577 ) | ( n6170 & n16577 ) ;
  assign n16579 = ( ~n1022 & n12162 ) | ( ~n1022 & n16578 ) | ( n12162 & n16578 ) ;
  assign n16580 = ( ~n569 & n5811 ) | ( ~n569 & n15879 ) | ( n5811 & n15879 ) ;
  assign n16581 = ( n1497 & ~n4483 ) | ( n1497 & n7135 ) | ( ~n4483 & n7135 ) ;
  assign n16582 = ( n5683 & n11673 ) | ( n5683 & n16581 ) | ( n11673 & n16581 ) ;
  assign n16583 = ( n3234 & ~n3569 ) | ( n3234 & n5247 ) | ( ~n3569 & n5247 ) ;
  assign n16584 = n3168 ^ n2694 ^ n297 ;
  assign n16585 = ( n15159 & n16583 ) | ( n15159 & ~n16584 ) | ( n16583 & ~n16584 ) ;
  assign n16589 = ( ~n2720 & n3821 ) | ( ~n2720 & n15102 ) | ( n3821 & n15102 ) ;
  assign n16586 = ( x96 & n1189 ) | ( x96 & n2240 ) | ( n1189 & n2240 ) ;
  assign n16587 = ( ~n2469 & n7798 ) | ( ~n2469 & n16586 ) | ( n7798 & n16586 ) ;
  assign n16588 = ( n12448 & n13329 ) | ( n12448 & n16587 ) | ( n13329 & n16587 ) ;
  assign n16590 = n16589 ^ n16588 ^ n14126 ;
  assign n16591 = n16590 ^ n9723 ^ n8090 ;
  assign n16592 = ( ~n5046 & n16585 ) | ( ~n5046 & n16591 ) | ( n16585 & n16591 ) ;
  assign n16593 = n13243 ^ n8202 ^ n220 ;
  assign n16594 = ( n886 & n14205 ) | ( n886 & ~n16593 ) | ( n14205 & ~n16593 ) ;
  assign n16596 = ( n6120 & n10107 ) | ( n6120 & n12071 ) | ( n10107 & n12071 ) ;
  assign n16595 = n9234 ^ n8950 ^ n2475 ;
  assign n16597 = n16596 ^ n16595 ^ n14578 ;
  assign n16601 = ( n2226 & n6530 ) | ( n2226 & n13448 ) | ( n6530 & n13448 ) ;
  assign n16598 = ( n938 & n1312 ) | ( n938 & ~n10744 ) | ( n1312 & ~n10744 ) ;
  assign n16599 = ( n1696 & ~n4690 ) | ( n1696 & n16598 ) | ( ~n4690 & n16598 ) ;
  assign n16600 = n16599 ^ n12856 ^ n1338 ;
  assign n16602 = n16601 ^ n16600 ^ n3076 ;
  assign n16604 = n9806 ^ n8295 ^ n5730 ;
  assign n16603 = ( ~n6365 & n7479 ) | ( ~n6365 & n13910 ) | ( n7479 & n13910 ) ;
  assign n16605 = n16604 ^ n16603 ^ n8968 ;
  assign n16606 = ( n2764 & n8419 ) | ( n2764 & n12835 ) | ( n8419 & n12835 ) ;
  assign n16607 = ( n1227 & n13723 ) | ( n1227 & ~n16606 ) | ( n13723 & ~n16606 ) ;
  assign n16608 = ( n3066 & n6757 ) | ( n3066 & ~n7243 ) | ( n6757 & ~n7243 ) ;
  assign n16609 = n13690 ^ n1404 ^ n129 ;
  assign n16610 = ( n4671 & n16608 ) | ( n4671 & ~n16609 ) | ( n16608 & ~n16609 ) ;
  assign n16611 = ( n1621 & n9248 ) | ( n1621 & n16610 ) | ( n9248 & n16610 ) ;
  assign n16612 = ( n5038 & n15284 ) | ( n5038 & n16611 ) | ( n15284 & n16611 ) ;
  assign n16613 = ( n313 & n3062 ) | ( n313 & ~n3234 ) | ( n3062 & ~n3234 ) ;
  assign n16614 = ( ~n4666 & n9856 ) | ( ~n4666 & n14516 ) | ( n9856 & n14516 ) ;
  assign n16615 = ( ~n14053 & n16613 ) | ( ~n14053 & n16614 ) | ( n16613 & n16614 ) ;
  assign n16618 = ( n3092 & ~n4195 ) | ( n3092 & n12104 ) | ( ~n4195 & n12104 ) ;
  assign n16616 = ( n3703 & n7238 ) | ( n3703 & n8402 ) | ( n7238 & n8402 ) ;
  assign n16617 = n16616 ^ n2053 ^ n1085 ;
  assign n16619 = n16618 ^ n16617 ^ n16169 ;
  assign n16620 = ( n4128 & n7060 ) | ( n4128 & n7479 ) | ( n7060 & n7479 ) ;
  assign n16621 = n16620 ^ n7840 ^ n7153 ;
  assign n16622 = ( n1893 & n9780 ) | ( n1893 & n16587 ) | ( n9780 & n16587 ) ;
  assign n16623 = ( n13523 & n16621 ) | ( n13523 & n16622 ) | ( n16621 & n16622 ) ;
  assign n16624 = ( n4709 & ~n13233 ) | ( n4709 & n16623 ) | ( ~n13233 & n16623 ) ;
  assign n16625 = n9587 ^ n7264 ^ n5347 ;
  assign n16628 = n10664 ^ n4472 ^ n570 ;
  assign n16626 = n6785 ^ n6742 ^ n4732 ;
  assign n16627 = ( n884 & n3503 ) | ( n884 & ~n16626 ) | ( n3503 & ~n16626 ) ;
  assign n16629 = n16628 ^ n16627 ^ n2180 ;
  assign n16637 = ( ~n1150 & n2863 ) | ( ~n1150 & n3960 ) | ( n2863 & n3960 ) ;
  assign n16638 = n16637 ^ n1805 ^ n803 ;
  assign n16630 = ( n892 & n931 ) | ( n892 & ~n1073 ) | ( n931 & ~n1073 ) ;
  assign n16631 = n16630 ^ n5054 ^ n1132 ;
  assign n16632 = n16631 ^ n12777 ^ n12274 ;
  assign n16633 = n4845 ^ n884 ^ n311 ;
  assign n16634 = n16633 ^ n3486 ^ n1831 ;
  assign n16635 = n16634 ^ n4156 ^ n3553 ;
  assign n16636 = ( n3372 & ~n16632 ) | ( n3372 & n16635 ) | ( ~n16632 & n16635 ) ;
  assign n16639 = n16638 ^ n16636 ^ n7961 ;
  assign n16642 = ( n541 & ~n4819 ) | ( n541 & n6863 ) | ( ~n4819 & n6863 ) ;
  assign n16643 = ( n1968 & n5822 ) | ( n1968 & n16642 ) | ( n5822 & n16642 ) ;
  assign n16640 = ( n5395 & n6731 ) | ( n5395 & ~n11392 ) | ( n6731 & ~n11392 ) ;
  assign n16641 = ( ~n10291 & n10913 ) | ( ~n10291 & n16640 ) | ( n10913 & n16640 ) ;
  assign n16644 = n16643 ^ n16641 ^ n11908 ;
  assign n16645 = ( ~n5899 & n16639 ) | ( ~n5899 & n16644 ) | ( n16639 & n16644 ) ;
  assign n16648 = n8122 ^ n7769 ^ n557 ;
  assign n16646 = ( n575 & n4229 ) | ( n575 & ~n11728 ) | ( n4229 & ~n11728 ) ;
  assign n16647 = n16646 ^ n14246 ^ n5698 ;
  assign n16649 = n16648 ^ n16647 ^ n2983 ;
  assign n16650 = ( n141 & n343 ) | ( n141 & ~n3442 ) | ( n343 & ~n3442 ) ;
  assign n16651 = ( n4073 & n7177 ) | ( n4073 & ~n16650 ) | ( n7177 & ~n16650 ) ;
  assign n16652 = n5518 ^ n3750 ^ n1655 ;
  assign n16653 = ( ~n5919 & n9082 ) | ( ~n5919 & n16652 ) | ( n9082 & n16652 ) ;
  assign n16654 = n15565 ^ n11844 ^ n2042 ;
  assign n16655 = ( n1792 & n8500 ) | ( n1792 & ~n16654 ) | ( n8500 & ~n16654 ) ;
  assign n16656 = n16655 ^ n6231 ^ n5213 ;
  assign n16658 = ( n2021 & n4919 ) | ( n2021 & n7775 ) | ( n4919 & n7775 ) ;
  assign n16659 = n16658 ^ n8327 ^ n2742 ;
  assign n16657 = ( n1686 & n6614 ) | ( n1686 & n13373 ) | ( n6614 & n13373 ) ;
  assign n16660 = n16659 ^ n16657 ^ n8539 ;
  assign n16661 = ( n2046 & n2306 ) | ( n2046 & ~n7123 ) | ( n2306 & ~n7123 ) ;
  assign n16662 = ( n6107 & n16660 ) | ( n6107 & ~n16661 ) | ( n16660 & ~n16661 ) ;
  assign n16663 = n16662 ^ n16272 ^ x105 ;
  assign n16664 = ( n6324 & n16656 ) | ( n6324 & ~n16663 ) | ( n16656 & ~n16663 ) ;
  assign n16665 = n5824 ^ n1794 ^ n1704 ;
  assign n16666 = ( n5841 & n12846 ) | ( n5841 & ~n16665 ) | ( n12846 & ~n16665 ) ;
  assign n16668 = ( n1708 & ~n6579 ) | ( n1708 & n15034 ) | ( ~n6579 & n15034 ) ;
  assign n16669 = n16668 ^ n15415 ^ n7861 ;
  assign n16670 = ( ~n1148 & n13583 ) | ( ~n1148 & n16669 ) | ( n13583 & n16669 ) ;
  assign n16667 = n6601 ^ n4783 ^ n1019 ;
  assign n16671 = n16670 ^ n16667 ^ n7756 ;
  assign n16672 = ( n2837 & n7072 ) | ( n2837 & ~n11762 ) | ( n7072 & ~n11762 ) ;
  assign n16673 = ( ~n16666 & n16671 ) | ( ~n16666 & n16672 ) | ( n16671 & n16672 ) ;
  assign n16674 = ( n468 & ~n1222 ) | ( n468 & n2485 ) | ( ~n1222 & n2485 ) ;
  assign n16675 = ( n6661 & n7216 ) | ( n6661 & n9692 ) | ( n7216 & n9692 ) ;
  assign n16676 = n13311 ^ n8956 ^ n851 ;
  assign n16677 = ( n5101 & ~n13130 ) | ( n5101 & n16676 ) | ( ~n13130 & n16676 ) ;
  assign n16678 = ( n1029 & n4218 ) | ( n1029 & ~n13836 ) | ( n4218 & ~n13836 ) ;
  assign n16679 = ( n10380 & ~n10856 ) | ( n10380 & n14838 ) | ( ~n10856 & n14838 ) ;
  assign n16680 = ( ~n3156 & n5320 ) | ( ~n3156 & n11778 ) | ( n5320 & n11778 ) ;
  assign n16681 = n3840 ^ n2132 ^ n391 ;
  assign n16682 = n14237 ^ n8185 ^ n6877 ;
  assign n16683 = n16682 ^ n2226 ^ n932 ;
  assign n16684 = ( n5385 & n6075 ) | ( n5385 & n7459 ) | ( n6075 & n7459 ) ;
  assign n16685 = ( ~n2417 & n3918 ) | ( ~n2417 & n16684 ) | ( n3918 & n16684 ) ;
  assign n16687 = n7434 ^ n5863 ^ n2444 ;
  assign n16686 = n13564 ^ n7218 ^ n467 ;
  assign n16688 = n16687 ^ n16686 ^ n15230 ;
  assign n16689 = ( n1246 & n8755 ) | ( n1246 & n10326 ) | ( n8755 & n10326 ) ;
  assign n16690 = n2489 ^ n2055 ^ x18 ;
  assign n16691 = n5963 ^ n4083 ^ n683 ;
  assign n16692 = ( ~n8930 & n16690 ) | ( ~n8930 & n16691 ) | ( n16690 & n16691 ) ;
  assign n16693 = n16692 ^ n6018 ^ n3622 ;
  assign n16694 = ( n5345 & n12353 ) | ( n5345 & ~n15283 ) | ( n12353 & ~n15283 ) ;
  assign n16695 = ( n16689 & n16693 ) | ( n16689 & n16694 ) | ( n16693 & n16694 ) ;
  assign n16696 = ( n848 & n849 ) | ( n848 & n16695 ) | ( n849 & n16695 ) ;
  assign n16697 = n15035 ^ n5140 ^ n3049 ;
  assign n16698 = n6135 ^ n4848 ^ n3935 ;
  assign n16699 = ( ~n3820 & n15769 ) | ( ~n3820 & n16698 ) | ( n15769 & n16698 ) ;
  assign n16700 = ( n1305 & n4564 ) | ( n1305 & n5957 ) | ( n4564 & n5957 ) ;
  assign n16701 = ( n4608 & n13322 ) | ( n4608 & ~n16700 ) | ( n13322 & ~n16700 ) ;
  assign n16702 = ( n2076 & ~n11273 ) | ( n2076 & n11571 ) | ( ~n11273 & n11571 ) ;
  assign n16703 = ( n5489 & n10587 ) | ( n5489 & n16702 ) | ( n10587 & n16702 ) ;
  assign n16706 = ( n734 & n858 ) | ( n734 & ~n6633 ) | ( n858 & ~n6633 ) ;
  assign n16705 = ( n5972 & n10473 ) | ( n5972 & n15360 ) | ( n10473 & n15360 ) ;
  assign n16704 = ( ~n1402 & n7046 ) | ( ~n1402 & n9201 ) | ( n7046 & n9201 ) ;
  assign n16707 = n16706 ^ n16705 ^ n16704 ;
  assign n16708 = ( ~n603 & n1209 ) | ( ~n603 & n4349 ) | ( n1209 & n4349 ) ;
  assign n16709 = ( n4822 & n12108 ) | ( n4822 & n16708 ) | ( n12108 & n16708 ) ;
  assign n16710 = ( x17 & n223 ) | ( x17 & ~n6219 ) | ( n223 & ~n6219 ) ;
  assign n16711 = ( n3956 & n4145 ) | ( n3956 & ~n9314 ) | ( n4145 & ~n9314 ) ;
  assign n16712 = ( n888 & n8697 ) | ( n888 & ~n16711 ) | ( n8697 & ~n16711 ) ;
  assign n16713 = n16712 ^ n15613 ^ n3341 ;
  assign n16714 = ( n10419 & ~n16710 ) | ( n10419 & n16713 ) | ( ~n16710 & n16713 ) ;
  assign n16715 = ( ~n3988 & n14710 ) | ( ~n3988 & n16714 ) | ( n14710 & n16714 ) ;
  assign n16716 = n15130 ^ n9735 ^ n8058 ;
  assign n16720 = n13861 ^ n13039 ^ n12971 ;
  assign n16721 = n16720 ^ n16385 ^ n10710 ;
  assign n16722 = ( n790 & n12732 ) | ( n790 & n16721 ) | ( n12732 & n16721 ) ;
  assign n16718 = ( n6495 & n7336 ) | ( n6495 & ~n13012 ) | ( n7336 & ~n13012 ) ;
  assign n16719 = n16718 ^ n9907 ^ n5371 ;
  assign n16717 = n16669 ^ n9304 ^ n8865 ;
  assign n16723 = n16722 ^ n16719 ^ n16717 ;
  assign n16724 = n11580 ^ n11167 ^ n1223 ;
  assign n16725 = n11736 ^ n4695 ^ n2007 ;
  assign n16726 = ( n1554 & n7092 ) | ( n1554 & n8594 ) | ( n7092 & n8594 ) ;
  assign n16727 = n10377 ^ n9050 ^ n8906 ;
  assign n16728 = ( n269 & ~n16726 ) | ( n269 & n16727 ) | ( ~n16726 & n16727 ) ;
  assign n16729 = n5466 ^ n2995 ^ n2988 ;
  assign n16730 = ( ~n6421 & n8603 ) | ( ~n6421 & n11003 ) | ( n8603 & n11003 ) ;
  assign n16731 = ( ~n7020 & n7271 ) | ( ~n7020 & n10282 ) | ( n7271 & n10282 ) ;
  assign n16732 = ( ~n6991 & n16730 ) | ( ~n6991 & n16731 ) | ( n16730 & n16731 ) ;
  assign n16733 = ( n1661 & n7902 ) | ( n1661 & ~n8685 ) | ( n7902 & ~n8685 ) ;
  assign n16734 = n16733 ^ n6336 ^ n3863 ;
  assign n16735 = ( ~n12288 & n16446 ) | ( ~n12288 & n16734 ) | ( n16446 & n16734 ) ;
  assign n16736 = n15310 ^ n11214 ^ n1060 ;
  assign n16737 = ( n3481 & n16735 ) | ( n3481 & ~n16736 ) | ( n16735 & ~n16736 ) ;
  assign n16739 = ( n2365 & n5204 ) | ( n2365 & n6412 ) | ( n5204 & n6412 ) ;
  assign n16738 = ( n3207 & n3791 ) | ( n3207 & ~n12386 ) | ( n3791 & ~n12386 ) ;
  assign n16740 = n16739 ^ n16738 ^ n1196 ;
  assign n16741 = ( n1910 & n4609 ) | ( n1910 & ~n16740 ) | ( n4609 & ~n16740 ) ;
  assign n16742 = n15533 ^ n14808 ^ n11020 ;
  assign n16743 = ( ~n13580 & n16741 ) | ( ~n13580 & n16742 ) | ( n16741 & n16742 ) ;
  assign n16744 = ( n2884 & n13066 ) | ( n2884 & n13940 ) | ( n13066 & n13940 ) ;
  assign n16745 = ( n10601 & n12496 ) | ( n10601 & n16744 ) | ( n12496 & n16744 ) ;
  assign n16746 = n13501 ^ n12989 ^ n10116 ;
  assign n16747 = ( ~n1737 & n2703 ) | ( ~n1737 & n16746 ) | ( n2703 & n16746 ) ;
  assign n16748 = ( ~n7210 & n10728 ) | ( ~n7210 & n15526 ) | ( n10728 & n15526 ) ;
  assign n16749 = ( ~n617 & n6419 ) | ( ~n617 & n7180 ) | ( n6419 & n7180 ) ;
  assign n16750 = n16749 ^ n1028 ^ n811 ;
  assign n16755 = n8103 ^ n4765 ^ n2502 ;
  assign n16752 = n5528 ^ n4265 ^ n2050 ;
  assign n16751 = n5572 ^ n2796 ^ n500 ;
  assign n16753 = n16752 ^ n16751 ^ n9125 ;
  assign n16754 = n16753 ^ n9038 ^ n5130 ;
  assign n16756 = n16755 ^ n16754 ^ n16429 ;
  assign n16757 = ( ~n7354 & n9782 ) | ( ~n7354 & n13994 ) | ( n9782 & n13994 ) ;
  assign n16758 = n16757 ^ n8055 ^ n4546 ;
  assign n16759 = n12992 ^ n5856 ^ x110 ;
  assign n16760 = ( n949 & ~n3461 ) | ( n949 & n16759 ) | ( ~n3461 & n16759 ) ;
  assign n16761 = ( n504 & n6849 ) | ( n504 & n16760 ) | ( n6849 & n16760 ) ;
  assign n16762 = n16761 ^ n9387 ^ n6132 ;
  assign n16763 = n13236 ^ n11154 ^ n4102 ;
  assign n16764 = ( n2481 & ~n13370 ) | ( n2481 & n16763 ) | ( ~n13370 & n16763 ) ;
  assign n16765 = ( n6704 & ~n9587 ) | ( n6704 & n11845 ) | ( ~n9587 & n11845 ) ;
  assign n16766 = n10297 ^ n5691 ^ n880 ;
  assign n16767 = n16766 ^ n10133 ^ n3721 ;
  assign n16768 = ( n4838 & ~n5497 ) | ( n4838 & n5661 ) | ( ~n5497 & n5661 ) ;
  assign n16769 = ( n5073 & n12240 ) | ( n5073 & n16768 ) | ( n12240 & n16768 ) ;
  assign n16770 = n5435 ^ n4695 ^ x52 ;
  assign n16771 = ( n1517 & n7998 ) | ( n1517 & ~n16770 ) | ( n7998 & ~n16770 ) ;
  assign n16772 = ( n520 & n3681 ) | ( n520 & n4247 ) | ( n3681 & n4247 ) ;
  assign n16773 = ( n311 & n605 ) | ( n311 & ~n6961 ) | ( n605 & ~n6961 ) ;
  assign n16774 = ( n4911 & n16772 ) | ( n4911 & ~n16773 ) | ( n16772 & ~n16773 ) ;
  assign n16775 = n5666 ^ n1823 ^ x59 ;
  assign n16776 = ( n6319 & n16774 ) | ( n6319 & ~n16775 ) | ( n16774 & ~n16775 ) ;
  assign n16779 = n8308 ^ n6625 ^ n2397 ;
  assign n16780 = ( n5745 & n11251 ) | ( n5745 & n16779 ) | ( n11251 & n16779 ) ;
  assign n16777 = ( n730 & ~n3543 ) | ( n730 & n15851 ) | ( ~n3543 & n15851 ) ;
  assign n16778 = ( n3588 & ~n12612 ) | ( n3588 & n16777 ) | ( ~n12612 & n16777 ) ;
  assign n16781 = n16780 ^ n16778 ^ n5924 ;
  assign n16783 = n11150 ^ n2743 ^ n2121 ;
  assign n16782 = n14298 ^ n8409 ^ n7680 ;
  assign n16784 = n16783 ^ n16782 ^ n11395 ;
  assign n16785 = n7322 ^ n5455 ^ n2522 ;
  assign n16786 = ( n1715 & ~n16222 ) | ( n1715 & n16785 ) | ( ~n16222 & n16785 ) ;
  assign n16787 = n8298 ^ n7414 ^ n2468 ;
  assign n16788 = n16787 ^ n11424 ^ n2229 ;
  assign n16789 = ( ~n6095 & n9954 ) | ( ~n6095 & n10129 ) | ( n9954 & n10129 ) ;
  assign n16790 = ( n4226 & n13590 ) | ( n4226 & ~n16789 ) | ( n13590 & ~n16789 ) ;
  assign n16791 = ( n2511 & n6146 ) | ( n2511 & n8612 ) | ( n6146 & n8612 ) ;
  assign n16792 = ( ~n2398 & n3858 ) | ( ~n2398 & n16791 ) | ( n3858 & n16791 ) ;
  assign n16793 = n8525 ^ n8448 ^ n775 ;
  assign n16794 = ( n5742 & n12880 ) | ( n5742 & ~n16793 ) | ( n12880 & ~n16793 ) ;
  assign n16795 = n14147 ^ n2555 ^ n1808 ;
  assign n16799 = ( ~n4399 & n9219 ) | ( ~n4399 & n12823 ) | ( n9219 & n12823 ) ;
  assign n16800 = ( ~n2376 & n14799 ) | ( ~n2376 & n16799 ) | ( n14799 & n16799 ) ;
  assign n16797 = n13757 ^ n12777 ^ n2983 ;
  assign n16796 = ( n5227 & n5303 ) | ( n5227 & ~n11335 ) | ( n5303 & ~n11335 ) ;
  assign n16798 = n16797 ^ n16796 ^ n8064 ;
  assign n16801 = n16800 ^ n16798 ^ n13250 ;
  assign n16802 = ( n396 & ~n1500 ) | ( n396 & n7311 ) | ( ~n1500 & n7311 ) ;
  assign n16803 = n16802 ^ n3318 ^ n1397 ;
  assign n16804 = ( ~n11468 & n15700 ) | ( ~n11468 & n16803 ) | ( n15700 & n16803 ) ;
  assign n16806 = ( n140 & ~n5218 ) | ( n140 & n16089 ) | ( ~n5218 & n16089 ) ;
  assign n16805 = ( n4930 & n11545 ) | ( n4930 & ~n13279 ) | ( n11545 & ~n13279 ) ;
  assign n16807 = n16806 ^ n16805 ^ n15449 ;
  assign n16808 = n4358 ^ n3477 ^ n138 ;
  assign n16809 = n6680 ^ n1598 ^ n407 ;
  assign n16810 = ( n4312 & n7248 ) | ( n4312 & ~n13277 ) | ( n7248 & ~n13277 ) ;
  assign n16811 = ( n3652 & ~n16809 ) | ( n3652 & n16810 ) | ( ~n16809 & n16810 ) ;
  assign n16812 = n16811 ^ n8834 ^ n2263 ;
  assign n16813 = n7955 ^ n4236 ^ n3045 ;
  assign n16814 = n12833 ^ n2667 ^ n978 ;
  assign n16815 = n16814 ^ n6914 ^ n2841 ;
  assign n16816 = n16815 ^ n5921 ^ n1608 ;
  assign n16817 = ( n4812 & n16813 ) | ( n4812 & ~n16816 ) | ( n16813 & ~n16816 ) ;
  assign n16818 = ( n4629 & n6251 ) | ( n4629 & n16817 ) | ( n6251 & n16817 ) ;
  assign n16819 = n7408 ^ n6737 ^ n5427 ;
  assign n16820 = n16819 ^ n6172 ^ n4512 ;
  assign n16821 = n15715 ^ n6181 ^ n2496 ;
  assign n16822 = ( ~n2927 & n6130 ) | ( ~n2927 & n16821 ) | ( n6130 & n16821 ) ;
  assign n16823 = n8591 ^ n7107 ^ n1109 ;
  assign n16824 = ( n1818 & n16822 ) | ( n1818 & ~n16823 ) | ( n16822 & ~n16823 ) ;
  assign n16825 = n16824 ^ n2568 ^ n616 ;
  assign n16826 = ( n359 & n2139 ) | ( n359 & ~n16825 ) | ( n2139 & ~n16825 ) ;
  assign n16829 = ( n2507 & n6008 ) | ( n2507 & ~n6896 ) | ( n6008 & ~n6896 ) ;
  assign n16830 = n5885 ^ n4649 ^ n1812 ;
  assign n16831 = ( n2977 & n16829 ) | ( n2977 & ~n16830 ) | ( n16829 & ~n16830 ) ;
  assign n16832 = n16831 ^ n13386 ^ n8066 ;
  assign n16827 = n9098 ^ n2257 ^ n1237 ;
  assign n16828 = ( n3087 & n15027 ) | ( n3087 & ~n16827 ) | ( n15027 & ~n16827 ) ;
  assign n16833 = n16832 ^ n16828 ^ n11176 ;
  assign n16834 = n6114 ^ n5208 ^ n3647 ;
  assign n16835 = n16834 ^ n16809 ^ n287 ;
  assign n16836 = ( n3738 & n4935 ) | ( n3738 & n15079 ) | ( n4935 & n15079 ) ;
  assign n16837 = n16836 ^ n12804 ^ n12271 ;
  assign n16838 = ( n8376 & n9957 ) | ( n8376 & ~n11657 ) | ( n9957 & ~n11657 ) ;
  assign n16839 = ( n5157 & n13897 ) | ( n5157 & n16838 ) | ( n13897 & n16838 ) ;
  assign n16840 = n14714 ^ n10459 ^ n996 ;
  assign n16841 = ( n4485 & ~n5295 ) | ( n4485 & n16840 ) | ( ~n5295 & n16840 ) ;
  assign n16842 = ( n1132 & n12710 ) | ( n1132 & n13055 ) | ( n12710 & n13055 ) ;
  assign n16843 = ( n5299 & ~n8221 ) | ( n5299 & n16842 ) | ( ~n8221 & n16842 ) ;
  assign n16844 = n14142 ^ n4193 ^ n3484 ;
  assign n16845 = n16844 ^ n16483 ^ n3119 ;
  assign n16846 = n10189 ^ n3065 ^ n2658 ;
  assign n16847 = ( n8449 & n13833 ) | ( n8449 & ~n16846 ) | ( n13833 & ~n16846 ) ;
  assign n16848 = n13531 ^ n8796 ^ n5516 ;
  assign n16849 = n16848 ^ n9545 ^ n6671 ;
  assign n16855 = n6260 ^ n2462 ^ n2280 ;
  assign n16854 = ( ~n290 & n6309 ) | ( ~n290 & n7813 ) | ( n6309 & n7813 ) ;
  assign n16856 = n16855 ^ n16854 ^ n2157 ;
  assign n16850 = n8484 ^ n4663 ^ n1105 ;
  assign n16851 = ( n10911 & ~n13023 ) | ( n10911 & n16850 ) | ( ~n13023 & n16850 ) ;
  assign n16852 = ( n5548 & ~n13255 ) | ( n5548 & n16851 ) | ( ~n13255 & n16851 ) ;
  assign n16853 = ( n3953 & n6217 ) | ( n3953 & n16852 ) | ( n6217 & n16852 ) ;
  assign n16857 = n16856 ^ n16853 ^ n10749 ;
  assign n16858 = n11496 ^ n10250 ^ n2187 ;
  assign n16859 = n14981 ^ n8471 ^ n2718 ;
  assign n16860 = ( n1031 & ~n6230 ) | ( n1031 & n16859 ) | ( ~n6230 & n16859 ) ;
  assign n16861 = ( n1144 & n6877 ) | ( n1144 & n16860 ) | ( n6877 & n16860 ) ;
  assign n16862 = ( n1333 & n6070 ) | ( n1333 & ~n8126 ) | ( n6070 & ~n8126 ) ;
  assign n16863 = ( n2964 & n3763 ) | ( n2964 & n16862 ) | ( n3763 & n16862 ) ;
  assign n16864 = ( n5691 & n6034 ) | ( n5691 & n16863 ) | ( n6034 & n16863 ) ;
  assign n16865 = ( ~n5930 & n16861 ) | ( ~n5930 & n16864 ) | ( n16861 & n16864 ) ;
  assign n16866 = ( ~n16303 & n16858 ) | ( ~n16303 & n16865 ) | ( n16858 & n16865 ) ;
  assign n16870 = ( n4812 & ~n5712 ) | ( n4812 & n7471 ) | ( ~n5712 & n7471 ) ;
  assign n16871 = ( n1097 & n2385 ) | ( n1097 & n16870 ) | ( n2385 & n16870 ) ;
  assign n16868 = n7805 ^ n4914 ^ n2225 ;
  assign n16869 = n16868 ^ n16107 ^ n14524 ;
  assign n16867 = ( n1679 & n1920 ) | ( n1679 & n9281 ) | ( n1920 & n9281 ) ;
  assign n16872 = n16871 ^ n16869 ^ n16867 ;
  assign n16873 = ( n2880 & n10931 ) | ( n2880 & n12011 ) | ( n10931 & n12011 ) ;
  assign n16874 = ( n1071 & n1452 ) | ( n1071 & ~n16873 ) | ( n1452 & ~n16873 ) ;
  assign n16875 = n16874 ^ n13991 ^ n8942 ;
  assign n16876 = ( n9929 & n16058 ) | ( n9929 & ~n16875 ) | ( n16058 & ~n16875 ) ;
  assign n16877 = n16876 ^ n16014 ^ n11172 ;
  assign n16878 = n13495 ^ n11515 ^ n6270 ;
  assign n16879 = ( n10314 & ~n16359 ) | ( n10314 & n16878 ) | ( ~n16359 & n16878 ) ;
  assign n16882 = ( ~n1254 & n5099 ) | ( ~n1254 & n9921 ) | ( n5099 & n9921 ) ;
  assign n16880 = n8612 ^ n7161 ^ n6102 ;
  assign n16881 = ( n13558 & n14429 ) | ( n13558 & ~n16880 ) | ( n14429 & ~n16880 ) ;
  assign n16883 = n16882 ^ n16881 ^ n12480 ;
  assign n16886 = ( n1180 & ~n2762 ) | ( n1180 & n3491 ) | ( ~n2762 & n3491 ) ;
  assign n16884 = ( ~n1469 & n3886 ) | ( ~n1469 & n5553 ) | ( n3886 & n5553 ) ;
  assign n16885 = ( n2439 & ~n11856 ) | ( n2439 & n16884 ) | ( ~n11856 & n16884 ) ;
  assign n16887 = n16886 ^ n16885 ^ n5254 ;
  assign n16888 = ( n1694 & n3480 ) | ( n1694 & ~n9228 ) | ( n3480 & ~n9228 ) ;
  assign n16889 = n16888 ^ n12620 ^ n8491 ;
  assign n16890 = ( n326 & ~n1016 ) | ( n326 & n14190 ) | ( ~n1016 & n14190 ) ;
  assign n16891 = n16890 ^ n4967 ^ n4702 ;
  assign n16892 = ( n6752 & ~n8946 ) | ( n6752 & n16891 ) | ( ~n8946 & n16891 ) ;
  assign n16893 = n16892 ^ n7146 ^ n2393 ;
  assign n16894 = ( ~n1409 & n11637 ) | ( ~n1409 & n16893 ) | ( n11637 & n16893 ) ;
  assign n16895 = ( n6332 & ~n16889 ) | ( n6332 & n16894 ) | ( ~n16889 & n16894 ) ;
  assign n16896 = ( n5457 & ~n13355 ) | ( n5457 & n16895 ) | ( ~n13355 & n16895 ) ;
  assign n16897 = n13389 ^ n3165 ^ n2715 ;
  assign n16898 = ( n7002 & ~n10453 ) | ( n7002 & n16897 ) | ( ~n10453 & n16897 ) ;
  assign n16899 = ( n5584 & n7253 ) | ( n5584 & ~n16898 ) | ( n7253 & ~n16898 ) ;
  assign n16900 = ( n6660 & ~n10546 ) | ( n6660 & n14401 ) | ( ~n10546 & n14401 ) ;
  assign n16901 = n7453 ^ n4403 ^ n639 ;
  assign n16902 = ( ~n7522 & n12663 ) | ( ~n7522 & n16901 ) | ( n12663 & n16901 ) ;
  assign n16903 = ( n2098 & n8312 ) | ( n2098 & n16902 ) | ( n8312 & n16902 ) ;
  assign n16904 = n1828 ^ n1616 ^ n1147 ;
  assign n16907 = ( n2366 & ~n3082 ) | ( n2366 & n6609 ) | ( ~n3082 & n6609 ) ;
  assign n16905 = n10318 ^ n2809 ^ n2456 ;
  assign n16906 = ( n2241 & n11019 ) | ( n2241 & ~n16905 ) | ( n11019 & ~n16905 ) ;
  assign n16908 = n16907 ^ n16906 ^ n3113 ;
  assign n16909 = n16908 ^ n11855 ^ n4015 ;
  assign n16910 = n10958 ^ n2051 ^ n478 ;
  assign n16918 = n8568 ^ n2501 ^ n1318 ;
  assign n16919 = n9978 ^ n9631 ^ n7396 ;
  assign n16920 = ( ~n1946 & n16918 ) | ( ~n1946 & n16919 ) | ( n16918 & n16919 ) ;
  assign n16916 = ( n922 & n1503 ) | ( n922 & ~n4034 ) | ( n1503 & ~n4034 ) ;
  assign n16915 = ( n2156 & ~n9188 ) | ( n2156 & n14107 ) | ( ~n9188 & n14107 ) ;
  assign n16917 = n16916 ^ n16915 ^ n7132 ;
  assign n16921 = n16920 ^ n16917 ^ n1213 ;
  assign n16913 = n15821 ^ n11486 ^ n2714 ;
  assign n16914 = n16913 ^ n4430 ^ n4181 ;
  assign n16911 = ( n3404 & n4809 ) | ( n3404 & ~n11122 ) | ( n4809 & ~n11122 ) ;
  assign n16912 = ( n4604 & ~n11466 ) | ( n4604 & n16911 ) | ( ~n11466 & n16911 ) ;
  assign n16922 = n16921 ^ n16914 ^ n16912 ;
  assign n16923 = n7588 ^ n2292 ^ n2044 ;
  assign n16924 = ( n4821 & ~n5182 ) | ( n4821 & n15704 ) | ( ~n5182 & n15704 ) ;
  assign n16925 = ( ~n10172 & n16923 ) | ( ~n10172 & n16924 ) | ( n16923 & n16924 ) ;
  assign n16926 = ( n2134 & n3141 ) | ( n2134 & n10171 ) | ( n3141 & n10171 ) ;
  assign n16927 = n16926 ^ n15102 ^ n5950 ;
  assign n16928 = ( n1338 & n13776 ) | ( n1338 & n16927 ) | ( n13776 & n16927 ) ;
  assign n16930 = n14565 ^ n5984 ^ n4329 ;
  assign n16929 = n14206 ^ n4010 ^ n2849 ;
  assign n16931 = n16930 ^ n16929 ^ n9591 ;
  assign n16932 = ( n2624 & n8891 ) | ( n2624 & n16931 ) | ( n8891 & n16931 ) ;
  assign n16933 = n14729 ^ n14561 ^ n2055 ;
  assign n16934 = ( n301 & n1067 ) | ( n301 & n3827 ) | ( n1067 & n3827 ) ;
  assign n16935 = ( n237 & ~n16331 ) | ( n237 & n16934 ) | ( ~n16331 & n16934 ) ;
  assign n16936 = ( n2626 & ~n10627 ) | ( n2626 & n13533 ) | ( ~n10627 & n13533 ) ;
  assign n16937 = n16936 ^ n16356 ^ n11097 ;
  assign n16939 = n7313 ^ n6276 ^ n4175 ;
  assign n16938 = n16154 ^ n14043 ^ n13180 ;
  assign n16940 = n16939 ^ n16938 ^ n8008 ;
  assign n16941 = n10786 ^ n5668 ^ n5317 ;
  assign n16942 = n16941 ^ n4437 ^ n2576 ;
  assign n16943 = ( n10253 & n11897 ) | ( n10253 & n15908 ) | ( n11897 & n15908 ) ;
  assign n16944 = n16943 ^ n12919 ^ n12760 ;
  assign n16945 = ( n15666 & ~n16942 ) | ( n15666 & n16944 ) | ( ~n16942 & n16944 ) ;
  assign n16946 = ( n187 & ~n3927 ) | ( n187 & n10633 ) | ( ~n3927 & n10633 ) ;
  assign n16947 = ( n4475 & ~n6692 ) | ( n4475 & n9754 ) | ( ~n6692 & n9754 ) ;
  assign n16948 = n16947 ^ n12058 ^ n9300 ;
  assign n16949 = n15449 ^ n13361 ^ n5817 ;
  assign n16950 = n16949 ^ n7915 ^ n301 ;
  assign n16951 = ( x15 & n173 ) | ( x15 & ~n16950 ) | ( n173 & ~n16950 ) ;
  assign n16952 = ( n12428 & ~n14436 ) | ( n12428 & n16951 ) | ( ~n14436 & n16951 ) ;
  assign n16953 = ( ~n1823 & n2789 ) | ( ~n1823 & n6395 ) | ( n2789 & n6395 ) ;
  assign n16954 = ( n2336 & ~n6044 ) | ( n2336 & n7006 ) | ( ~n6044 & n7006 ) ;
  assign n16955 = n16954 ^ n11897 ^ n8165 ;
  assign n16956 = ( n2066 & n9438 ) | ( n2066 & ~n16955 ) | ( n9438 & ~n16955 ) ;
  assign n16959 = ( n2261 & n3396 ) | ( n2261 & ~n3492 ) | ( n3396 & ~n3492 ) ;
  assign n16957 = n8345 ^ n3036 ^ n2878 ;
  assign n16958 = ( n14966 & n15759 ) | ( n14966 & ~n16957 ) | ( n15759 & ~n16957 ) ;
  assign n16960 = n16959 ^ n16958 ^ n15806 ;
  assign n16961 = n14314 ^ n8837 ^ n1144 ;
  assign n16962 = n15770 ^ n12845 ^ n6968 ;
  assign n16963 = ( ~n1824 & n3169 ) | ( ~n1824 & n11211 ) | ( n3169 & n11211 ) ;
  assign n16964 = n16963 ^ n15700 ^ n14628 ;
  assign n16965 = n16964 ^ n10695 ^ n2104 ;
  assign n16966 = ( ~n9079 & n9256 ) | ( ~n9079 & n16965 ) | ( n9256 & n16965 ) ;
  assign n16967 = n13315 ^ n3174 ^ n949 ;
  assign n16968 = ( x110 & n2674 ) | ( x110 & ~n2697 ) | ( n2674 & ~n2697 ) ;
  assign n16969 = n16968 ^ n4216 ^ n3553 ;
  assign n16970 = ( n4379 & n16967 ) | ( n4379 & ~n16969 ) | ( n16967 & ~n16969 ) ;
  assign n16971 = n16970 ^ n2565 ^ n1932 ;
  assign n16972 = ( n1021 & n6656 ) | ( n1021 & ~n16936 ) | ( n6656 & ~n16936 ) ;
  assign n16973 = n8041 ^ n4503 ^ x25 ;
  assign n16974 = ( n5744 & ~n10887 ) | ( n5744 & n16973 ) | ( ~n10887 & n16973 ) ;
  assign n16975 = ( n8610 & n15272 ) | ( n8610 & ~n15863 ) | ( n15272 & ~n15863 ) ;
  assign n16976 = n16975 ^ n14994 ^ n2520 ;
  assign n16977 = n11560 ^ n9771 ^ n1134 ;
  assign n16978 = n16977 ^ n5851 ^ n5224 ;
  assign n16979 = ( n2024 & ~n3043 ) | ( n2024 & n8281 ) | ( ~n3043 & n8281 ) ;
  assign n16980 = n14855 ^ n2921 ^ x77 ;
  assign n16981 = ( ~n4721 & n15273 ) | ( ~n4721 & n16980 ) | ( n15273 & n16980 ) ;
  assign n16982 = ( n14749 & n16979 ) | ( n14749 & n16981 ) | ( n16979 & n16981 ) ;
  assign n16983 = n12544 ^ n9237 ^ n7126 ;
  assign n16984 = n3067 ^ n1688 ^ n826 ;
  assign n16985 = ( n2691 & n16983 ) | ( n2691 & ~n16984 ) | ( n16983 & ~n16984 ) ;
  assign n16986 = ( n1100 & ~n4072 ) | ( n1100 & n8563 ) | ( ~n4072 & n8563 ) ;
  assign n16991 = ( n4827 & ~n9806 ) | ( n4827 & n14390 ) | ( ~n9806 & n14390 ) ;
  assign n16988 = n7296 ^ n1889 ^ n430 ;
  assign n16989 = ( n13564 & n14407 ) | ( n13564 & ~n16988 ) | ( n14407 & ~n16988 ) ;
  assign n16990 = n16989 ^ n10114 ^ n691 ;
  assign n16987 = n12881 ^ n4768 ^ n1464 ;
  assign n16992 = n16991 ^ n16990 ^ n16987 ;
  assign n16993 = ( n5593 & ~n10074 ) | ( n5593 & n13171 ) | ( ~n10074 & n13171 ) ;
  assign n16994 = n16993 ^ n16741 ^ n4441 ;
  assign n16995 = ( n7700 & n12910 ) | ( n7700 & n16994 ) | ( n12910 & n16994 ) ;
  assign n16999 = n12586 ^ n6835 ^ n382 ;
  assign n16996 = ( n5872 & ~n13910 ) | ( n5872 & n15272 ) | ( ~n13910 & n15272 ) ;
  assign n16997 = n7609 ^ n3635 ^ n1015 ;
  assign n16998 = ( ~n4986 & n16996 ) | ( ~n4986 & n16997 ) | ( n16996 & n16997 ) ;
  assign n17000 = n16999 ^ n16998 ^ n11520 ;
  assign n17003 = n4764 ^ n2580 ^ n1808 ;
  assign n17004 = n17003 ^ n11323 ^ n4457 ;
  assign n17001 = ( ~n1922 & n6447 ) | ( ~n1922 & n12248 ) | ( n6447 & n12248 ) ;
  assign n17002 = ( n1460 & ~n2614 ) | ( n1460 & n17001 ) | ( ~n2614 & n17001 ) ;
  assign n17005 = n17004 ^ n17002 ^ n12538 ;
  assign n17006 = n13496 ^ n12844 ^ n2717 ;
  assign n17007 = n13527 ^ n4760 ^ n4181 ;
  assign n17008 = ( n17005 & n17006 ) | ( n17005 & ~n17007 ) | ( n17006 & ~n17007 ) ;
  assign n17009 = ( n999 & n8583 ) | ( n999 & n17008 ) | ( n8583 & n17008 ) ;
  assign n17010 = n6892 ^ n6465 ^ n2932 ;
  assign n17011 = ( ~n12924 & n16384 ) | ( ~n12924 & n17010 ) | ( n16384 & n17010 ) ;
  assign n17012 = n17011 ^ n12944 ^ n8846 ;
  assign n17015 = n8879 ^ n4455 ^ n3922 ;
  assign n17014 = ( n812 & n3138 ) | ( n812 & n4499 ) | ( n3138 & n4499 ) ;
  assign n17013 = ( n1481 & n6884 ) | ( n1481 & n15199 ) | ( n6884 & n15199 ) ;
  assign n17016 = n17015 ^ n17014 ^ n17013 ;
  assign n17017 = n16243 ^ n5020 ^ n944 ;
  assign n17018 = n15998 ^ n12661 ^ n6227 ;
  assign n17019 = ( n5692 & ~n17017 ) | ( n5692 & n17018 ) | ( ~n17017 & n17018 ) ;
  assign n17020 = n17019 ^ n13989 ^ n12903 ;
  assign n17021 = ( ~n5415 & n13942 ) | ( ~n5415 & n14573 ) | ( n13942 & n14573 ) ;
  assign n17022 = n17021 ^ n4840 ^ n1172 ;
  assign n17023 = ( ~n3919 & n12187 ) | ( ~n3919 & n17022 ) | ( n12187 & n17022 ) ;
  assign n17024 = ( n7468 & n16504 ) | ( n7468 & n17023 ) | ( n16504 & n17023 ) ;
  assign n17025 = ( ~n828 & n4504 ) | ( ~n828 & n15152 ) | ( n4504 & n15152 ) ;
  assign n17026 = ( ~n263 & n6120 ) | ( ~n263 & n17015 ) | ( n6120 & n17015 ) ;
  assign n17027 = ( ~n4252 & n9004 ) | ( ~n4252 & n17026 ) | ( n9004 & n17026 ) ;
  assign n17028 = ( n2155 & n17025 ) | ( n2155 & ~n17027 ) | ( n17025 & ~n17027 ) ;
  assign n17029 = ( n1237 & n3594 ) | ( n1237 & n12514 ) | ( n3594 & n12514 ) ;
  assign n17031 = ( n4441 & n13818 ) | ( n4441 & ~n15003 ) | ( n13818 & ~n15003 ) ;
  assign n17030 = ( x111 & ~n9158 ) | ( x111 & n12826 ) | ( ~n9158 & n12826 ) ;
  assign n17032 = n17031 ^ n17030 ^ n173 ;
  assign n17033 = ( ~n4817 & n8526 ) | ( ~n4817 & n14367 ) | ( n8526 & n14367 ) ;
  assign n17034 = ( n17029 & ~n17032 ) | ( n17029 & n17033 ) | ( ~n17032 & n17033 ) ;
  assign n17035 = n9795 ^ n6698 ^ n530 ;
  assign n17036 = ( ~n3858 & n10818 ) | ( ~n3858 & n17035 ) | ( n10818 & n17035 ) ;
  assign n17037 = n14784 ^ n6518 ^ n4161 ;
  assign n17039 = ( ~n440 & n2633 ) | ( ~n440 & n14214 ) | ( n2633 & n14214 ) ;
  assign n17038 = ( n7563 & ~n7687 ) | ( n7563 & n9314 ) | ( ~n7687 & n9314 ) ;
  assign n17040 = n17039 ^ n17038 ^ n14173 ;
  assign n17041 = ( n7441 & ~n17037 ) | ( n7441 & n17040 ) | ( ~n17037 & n17040 ) ;
  assign n17042 = ( ~x30 & n2418 ) | ( ~x30 & n4603 ) | ( n2418 & n4603 ) ;
  assign n17043 = ( n3036 & ~n6804 ) | ( n3036 & n10489 ) | ( ~n6804 & n10489 ) ;
  assign n17044 = n17043 ^ n6130 ^ n6076 ;
  assign n17045 = ( n3430 & n3831 ) | ( n3430 & ~n8538 ) | ( n3831 & ~n8538 ) ;
  assign n17046 = ( n1938 & ~n3344 ) | ( n1938 & n9182 ) | ( ~n3344 & n9182 ) ;
  assign n17047 = ( n6099 & n7186 ) | ( n6099 & n17046 ) | ( n7186 & n17046 ) ;
  assign n17048 = ( n4339 & n4552 ) | ( n4339 & ~n16106 ) | ( n4552 & ~n16106 ) ;
  assign n17049 = ( n17045 & ~n17047 ) | ( n17045 & n17048 ) | ( ~n17047 & n17048 ) ;
  assign n17050 = ( n5047 & n17044 ) | ( n5047 & n17049 ) | ( n17044 & n17049 ) ;
  assign n17051 = n17050 ^ n13436 ^ n288 ;
  assign n17052 = ( n2009 & n17042 ) | ( n2009 & n17051 ) | ( n17042 & n17051 ) ;
  assign n17053 = n12526 ^ n3956 ^ n537 ;
  assign n17054 = ( n6166 & n6434 ) | ( n6166 & ~n10537 ) | ( n6434 & ~n10537 ) ;
  assign n17055 = ( n357 & n7667 ) | ( n357 & n17054 ) | ( n7667 & n17054 ) ;
  assign n17056 = n6430 ^ n5311 ^ n190 ;
  assign n17057 = ( n11736 & n17055 ) | ( n11736 & ~n17056 ) | ( n17055 & ~n17056 ) ;
  assign n17058 = ( n642 & ~n2785 ) | ( n642 & n5904 ) | ( ~n2785 & n5904 ) ;
  assign n17059 = ( n17053 & n17057 ) | ( n17053 & ~n17058 ) | ( n17057 & ~n17058 ) ;
  assign n17060 = ( ~n4842 & n11882 ) | ( ~n4842 & n13611 ) | ( n11882 & n13611 ) ;
  assign n17061 = n4651 ^ n1536 ^ n1050 ;
  assign n17062 = ( n6334 & ~n7434 ) | ( n6334 & n17061 ) | ( ~n7434 & n17061 ) ;
  assign n17069 = n5668 ^ n3117 ^ n1087 ;
  assign n17063 = n3139 ^ n1573 ^ n1524 ;
  assign n17064 = n17063 ^ n2378 ^ n682 ;
  assign n17065 = ( n327 & n1153 ) | ( n327 & n17064 ) | ( n1153 & n17064 ) ;
  assign n17066 = ( n3323 & n10334 ) | ( n3323 & ~n17065 ) | ( n10334 & ~n17065 ) ;
  assign n17067 = n12440 ^ n11813 ^ n3794 ;
  assign n17068 = ( n10781 & ~n17066 ) | ( n10781 & n17067 ) | ( ~n17066 & n17067 ) ;
  assign n17070 = n17069 ^ n17068 ^ n3127 ;
  assign n17072 = ( n721 & ~n6801 ) | ( n721 & n7428 ) | ( ~n6801 & n7428 ) ;
  assign n17071 = ( n4740 & n6799 ) | ( n4740 & ~n14215 ) | ( n6799 & ~n14215 ) ;
  assign n17073 = n17072 ^ n17071 ^ n16623 ;
  assign n17074 = ( n17062 & n17070 ) | ( n17062 & ~n17073 ) | ( n17070 & ~n17073 ) ;
  assign n17075 = ( n884 & n1448 ) | ( n884 & ~n9761 ) | ( n1448 & ~n9761 ) ;
  assign n17076 = ( n1277 & n5529 ) | ( n1277 & n17075 ) | ( n5529 & n17075 ) ;
  assign n17077 = n17076 ^ n11299 ^ n4686 ;
  assign n17078 = ( ~n4600 & n5196 ) | ( ~n4600 & n17077 ) | ( n5196 & n17077 ) ;
  assign n17079 = n11025 ^ n8730 ^ n7715 ;
  assign n17082 = ( n3512 & ~n4985 ) | ( n3512 & n6338 ) | ( ~n4985 & n6338 ) ;
  assign n17080 = ( n3989 & n6428 ) | ( n3989 & ~n15964 ) | ( n6428 & ~n15964 ) ;
  assign n17081 = ( n14532 & n15613 ) | ( n14532 & n17080 ) | ( n15613 & n17080 ) ;
  assign n17083 = n17082 ^ n17081 ^ n14932 ;
  assign n17084 = ( n9551 & ~n11711 ) | ( n9551 & n17083 ) | ( ~n11711 & n17083 ) ;
  assign n17085 = n17084 ^ n5983 ^ n939 ;
  assign n17086 = n8543 ^ n4982 ^ n3918 ;
  assign n17087 = n15406 ^ n14819 ^ n13993 ;
  assign n17089 = n14718 ^ n7857 ^ n6258 ;
  assign n17088 = n13998 ^ n8337 ^ n3728 ;
  assign n17090 = n17089 ^ n17088 ^ n478 ;
  assign n17091 = ( ~n4993 & n10103 ) | ( ~n4993 & n17090 ) | ( n10103 & n17090 ) ;
  assign n17092 = n15341 ^ n11678 ^ n1983 ;
  assign n17093 = n17092 ^ n11505 ^ n2981 ;
  assign n17094 = n17093 ^ n8737 ^ n1571 ;
  assign n17095 = n17094 ^ n9686 ^ n8763 ;
  assign n17096 = n14983 ^ n13944 ^ n12830 ;
  assign n17097 = ( n5187 & n7432 ) | ( n5187 & n11148 ) | ( n7432 & n11148 ) ;
  assign n17098 = ( n4641 & ~n7640 ) | ( n4641 & n9144 ) | ( ~n7640 & n9144 ) ;
  assign n17099 = n17098 ^ n4929 ^ n3966 ;
  assign n17100 = n11238 ^ n10165 ^ n3922 ;
  assign n17101 = n17100 ^ n16354 ^ n2404 ;
  assign n17102 = ( ~n3403 & n10021 ) | ( ~n3403 & n13931 ) | ( n10021 & n13931 ) ;
  assign n17103 = n17102 ^ n16512 ^ n9152 ;
  assign n17106 = n6391 ^ n4453 ^ n3180 ;
  assign n17107 = n17106 ^ n10438 ^ n8419 ;
  assign n17104 = ( n1835 & n4225 ) | ( n1835 & n8240 ) | ( n4225 & n8240 ) ;
  assign n17105 = ( n2099 & ~n5323 ) | ( n2099 & n17104 ) | ( ~n5323 & n17104 ) ;
  assign n17108 = n17107 ^ n17105 ^ n16381 ;
  assign n17109 = ( ~n5766 & n7583 ) | ( ~n5766 & n17108 ) | ( n7583 & n17108 ) ;
  assign n17110 = n7136 ^ n5251 ^ n220 ;
  assign n17111 = n17110 ^ n5046 ^ n166 ;
  assign n17112 = ( n583 & n5952 ) | ( n583 & ~n17111 ) | ( n5952 & ~n17111 ) ;
  assign n17113 = ( ~n6258 & n7185 ) | ( ~n6258 & n17112 ) | ( n7185 & n17112 ) ;
  assign n17114 = n11717 ^ n5488 ^ n3128 ;
  assign n17115 = ( n2889 & n4345 ) | ( n2889 & ~n17114 ) | ( n4345 & ~n17114 ) ;
  assign n17116 = n17115 ^ n13268 ^ n5902 ;
  assign n17117 = n17116 ^ n8315 ^ n6397 ;
  assign n17118 = ( ~n634 & n1749 ) | ( ~n634 & n13671 ) | ( n1749 & n13671 ) ;
  assign n17119 = n17118 ^ n13941 ^ n3884 ;
  assign n17120 = ( n5359 & n8777 ) | ( n5359 & ~n16371 ) | ( n8777 & ~n16371 ) ;
  assign n17121 = ( ~n485 & n6450 ) | ( ~n485 & n12961 ) | ( n6450 & n12961 ) ;
  assign n17122 = ( ~n8216 & n11351 ) | ( ~n8216 & n17121 ) | ( n11351 & n17121 ) ;
  assign n17123 = ( n8004 & ~n8593 ) | ( n8004 & n17122 ) | ( ~n8593 & n17122 ) ;
  assign n17124 = n1784 ^ n1748 ^ n1666 ;
  assign n17125 = ( n1143 & n1296 ) | ( n1143 & ~n17124 ) | ( n1296 & ~n17124 ) ;
  assign n17126 = n17125 ^ n7165 ^ n526 ;
  assign n17127 = n17126 ^ n7926 ^ n4773 ;
  assign n17128 = n17127 ^ n15721 ^ n7607 ;
  assign n17133 = n15540 ^ n7531 ^ n6456 ;
  assign n17131 = n12947 ^ n10683 ^ n398 ;
  assign n17129 = n16481 ^ n10239 ^ n545 ;
  assign n17130 = ( n4064 & n11297 ) | ( n4064 & ~n17129 ) | ( n11297 & ~n17129 ) ;
  assign n17132 = n17131 ^ n17130 ^ n5339 ;
  assign n17134 = n17133 ^ n17132 ^ n7494 ;
  assign n17140 = n9496 ^ n7590 ^ n2856 ;
  assign n17136 = n12860 ^ n10737 ^ n3803 ;
  assign n17137 = n17136 ^ n10011 ^ n1433 ;
  assign n17138 = n8692 ^ n8065 ^ n3120 ;
  assign n17139 = ( n7714 & ~n17137 ) | ( n7714 & n17138 ) | ( ~n17137 & n17138 ) ;
  assign n17135 = ( n8951 & ~n15441 ) | ( n8951 & n15956 ) | ( ~n15441 & n15956 ) ;
  assign n17141 = n17140 ^ n17139 ^ n17135 ;
  assign n17142 = ( n1841 & n5881 ) | ( n1841 & n9149 ) | ( n5881 & n9149 ) ;
  assign n17144 = n15416 ^ n5461 ^ n1205 ;
  assign n17143 = ( n1979 & n10866 ) | ( n1979 & n12078 ) | ( n10866 & n12078 ) ;
  assign n17145 = n17144 ^ n17143 ^ n4195 ;
  assign n17149 = n10574 ^ n7381 ^ n2057 ;
  assign n17146 = n7108 ^ n5675 ^ n3234 ;
  assign n17147 = n17146 ^ n7755 ^ n5601 ;
  assign n17148 = ( ~n4251 & n16218 ) | ( ~n4251 & n17147 ) | ( n16218 & n17147 ) ;
  assign n17150 = n17149 ^ n17148 ^ n10014 ;
  assign n17151 = n10422 ^ n4483 ^ n3981 ;
  assign n17152 = ( ~n5010 & n10547 ) | ( ~n5010 & n13023 ) | ( n10547 & n13023 ) ;
  assign n17153 = ( ~n3886 & n6172 ) | ( ~n3886 & n17152 ) | ( n6172 & n17152 ) ;
  assign n17154 = n17153 ^ n15277 ^ n12355 ;
  assign n17155 = ( n6966 & n7885 ) | ( n6966 & n17154 ) | ( n7885 & n17154 ) ;
  assign n17156 = ( n9275 & ~n17151 ) | ( n9275 & n17155 ) | ( ~n17151 & n17155 ) ;
  assign n17157 = ( ~n1878 & n4784 ) | ( ~n1878 & n10082 ) | ( n4784 & n10082 ) ;
  assign n17158 = ( n6211 & n6401 ) | ( n6211 & n10300 ) | ( n6401 & n10300 ) ;
  assign n17159 = ( n3053 & ~n3435 ) | ( n3053 & n17158 ) | ( ~n3435 & n17158 ) ;
  assign n17160 = ( n1182 & n6590 ) | ( n1182 & ~n16744 ) | ( n6590 & ~n16744 ) ;
  assign n17161 = ( ~n2038 & n2904 ) | ( ~n2038 & n14022 ) | ( n2904 & n14022 ) ;
  assign n17162 = ( n17159 & n17160 ) | ( n17159 & ~n17161 ) | ( n17160 & ~n17161 ) ;
  assign n17163 = n13503 ^ n8742 ^ n265 ;
  assign n17164 = ( ~n4040 & n9688 ) | ( ~n4040 & n13459 ) | ( n9688 & n13459 ) ;
  assign n17165 = n9428 ^ n4585 ^ n3304 ;
  assign n17166 = n17165 ^ n7085 ^ n3053 ;
  assign n17167 = ( ~n1145 & n11406 ) | ( ~n1145 & n17166 ) | ( n11406 & n17166 ) ;
  assign n17168 = n15726 ^ n6834 ^ n4388 ;
  assign n17169 = n17168 ^ n12767 ^ n1777 ;
  assign n17170 = ( n147 & n17167 ) | ( n147 & ~n17169 ) | ( n17167 & ~n17169 ) ;
  assign n17171 = ( n2089 & ~n17164 ) | ( n2089 & n17170 ) | ( ~n17164 & n17170 ) ;
  assign n17172 = ( n5679 & n7577 ) | ( n5679 & ~n14106 ) | ( n7577 & ~n14106 ) ;
  assign n17173 = ( n6317 & ~n14136 ) | ( n6317 & n17172 ) | ( ~n14136 & n17172 ) ;
  assign n17174 = n10791 ^ n9754 ^ n7959 ;
  assign n17175 = n13446 ^ n6933 ^ n5609 ;
  assign n17176 = n17175 ^ n15186 ^ n1647 ;
  assign n17177 = ( n7489 & n7490 ) | ( n7489 & n17176 ) | ( n7490 & n17176 ) ;
  assign n17178 = ( n332 & ~n17174 ) | ( n332 & n17177 ) | ( ~n17174 & n17177 ) ;
  assign n17179 = n16669 ^ n9349 ^ n318 ;
  assign n17180 = ( n703 & ~n2124 ) | ( n703 & n12131 ) | ( ~n2124 & n12131 ) ;
  assign n17181 = ( ~n10470 & n17179 ) | ( ~n10470 & n17180 ) | ( n17179 & n17180 ) ;
  assign n17182 = ( n4407 & ~n7134 ) | ( n4407 & n10556 ) | ( ~n7134 & n10556 ) ;
  assign n17183 = ( ~n3293 & n9506 ) | ( ~n3293 & n9930 ) | ( n9506 & n9930 ) ;
  assign n17184 = n17183 ^ n14681 ^ n10436 ;
  assign n17185 = n8737 ^ n8370 ^ n3852 ;
  assign n17186 = n13066 ^ n12943 ^ n6352 ;
  assign n17187 = n17186 ^ n10477 ^ n8383 ;
  assign n17188 = ( ~n1241 & n6447 ) | ( ~n1241 & n17187 ) | ( n6447 & n17187 ) ;
  assign n17189 = ( n11527 & n16650 ) | ( n11527 & ~n17188 ) | ( n16650 & ~n17188 ) ;
  assign n17190 = n9437 ^ n7751 ^ n6537 ;
  assign n17191 = ( n7730 & n9435 ) | ( n7730 & n11480 ) | ( n9435 & n11480 ) ;
  assign n17192 = ( n2884 & ~n17190 ) | ( n2884 & n17191 ) | ( ~n17190 & n17191 ) ;
  assign n17194 = ( ~n1101 & n2242 ) | ( ~n1101 & n11411 ) | ( n2242 & n11411 ) ;
  assign n17193 = ( ~n5541 & n9887 ) | ( ~n5541 & n12895 ) | ( n9887 & n12895 ) ;
  assign n17195 = n17194 ^ n17193 ^ n12875 ;
  assign n17196 = n17195 ^ n14732 ^ n5246 ;
  assign n17197 = n8327 ^ n7636 ^ n7014 ;
  assign n17198 = n17197 ^ n7242 ^ n5783 ;
  assign n17199 = ( n3854 & n7863 ) | ( n3854 & ~n14090 ) | ( n7863 & ~n14090 ) ;
  assign n17200 = ( n3327 & n7088 ) | ( n3327 & n7985 ) | ( n7088 & n7985 ) ;
  assign n17201 = ( ~n6251 & n6693 ) | ( ~n6251 & n12659 ) | ( n6693 & n12659 ) ;
  assign n17202 = ( n17199 & n17200 ) | ( n17199 & n17201 ) | ( n17200 & n17201 ) ;
  assign n17204 = ( n2472 & ~n2848 ) | ( n2472 & n6684 ) | ( ~n2848 & n6684 ) ;
  assign n17203 = n16167 ^ n9517 ^ n462 ;
  assign n17205 = n17204 ^ n17203 ^ n16621 ;
  assign n17206 = n14491 ^ n9498 ^ n620 ;
  assign n17207 = n17206 ^ n16980 ^ n233 ;
  assign n17208 = ( n7353 & ~n10063 ) | ( n7353 & n17207 ) | ( ~n10063 & n17207 ) ;
  assign n17209 = ( n7371 & ~n8543 ) | ( n7371 & n17208 ) | ( ~n8543 & n17208 ) ;
  assign n17210 = ( n4580 & ~n9574 ) | ( n4580 & n10858 ) | ( ~n9574 & n10858 ) ;
  assign n17211 = n10441 ^ n9519 ^ n3639 ;
  assign n17212 = n8970 ^ n6410 ^ n6359 ;
  assign n17213 = ( n4121 & n4321 ) | ( n4121 & ~n9755 ) | ( n4321 & ~n9755 ) ;
  assign n17214 = n13484 ^ n5515 ^ n1411 ;
  assign n17215 = ( n2158 & n7650 ) | ( n2158 & ~n17214 ) | ( n7650 & ~n17214 ) ;
  assign n17216 = n17215 ^ n12095 ^ n1375 ;
  assign n17217 = ( ~n4239 & n17213 ) | ( ~n4239 & n17216 ) | ( n17213 & n17216 ) ;
  assign n17219 = n10650 ^ n6964 ^ n6179 ;
  assign n17220 = ( n225 & n2712 ) | ( n225 & ~n17219 ) | ( n2712 & ~n17219 ) ;
  assign n17221 = ( ~n246 & n269 ) | ( ~n246 & n17220 ) | ( n269 & n17220 ) ;
  assign n17218 = ( n3821 & n9334 ) | ( n3821 & ~n11410 ) | ( n9334 & ~n11410 ) ;
  assign n17222 = n17221 ^ n17218 ^ n16682 ;
  assign n17223 = n15119 ^ n7283 ^ n511 ;
  assign n17224 = ( n4343 & ~n10589 ) | ( n4343 & n17223 ) | ( ~n10589 & n17223 ) ;
  assign n17225 = n10692 ^ n7276 ^ n3407 ;
  assign n17226 = ( n1128 & ~n8389 ) | ( n1128 & n10255 ) | ( ~n8389 & n10255 ) ;
  assign n17227 = ( ~n8882 & n12798 ) | ( ~n8882 & n17226 ) | ( n12798 & n17226 ) ;
  assign n17228 = ( ~n2237 & n3908 ) | ( ~n2237 & n12895 ) | ( n3908 & n12895 ) ;
  assign n17229 = ( n15530 & ~n16255 ) | ( n15530 & n17228 ) | ( ~n16255 & n17228 ) ;
  assign n17230 = n14044 ^ n7248 ^ n251 ;
  assign n17231 = ( n4264 & n4884 ) | ( n4264 & ~n8625 ) | ( n4884 & ~n8625 ) ;
  assign n17232 = n17231 ^ n6930 ^ n840 ;
  assign n17233 = n17232 ^ n12763 ^ n12015 ;
  assign n17234 = ( ~n3607 & n4963 ) | ( ~n3607 & n11909 ) | ( n4963 & n11909 ) ;
  assign n17235 = ( x32 & ~n3283 ) | ( x32 & n17234 ) | ( ~n3283 & n17234 ) ;
  assign n17236 = n15565 ^ n13085 ^ n7271 ;
  assign n17237 = ( n1679 & ~n5974 ) | ( n1679 & n11047 ) | ( ~n5974 & n11047 ) ;
  assign n17238 = ( ~n2967 & n7229 ) | ( ~n2967 & n11127 ) | ( n7229 & n11127 ) ;
  assign n17239 = n16169 ^ n15508 ^ n1301 ;
  assign n17240 = ( ~n8785 & n11013 ) | ( ~n8785 & n14165 ) | ( n11013 & n14165 ) ;
  assign n17241 = n12193 ^ n7631 ^ n6352 ;
  assign n17242 = ( n184 & n17240 ) | ( n184 & n17241 ) | ( n17240 & n17241 ) ;
  assign n17243 = ( ~n3335 & n5109 ) | ( ~n3335 & n10121 ) | ( n5109 & n10121 ) ;
  assign n17244 = ( n5131 & n11250 ) | ( n5131 & ~n16564 ) | ( n11250 & ~n16564 ) ;
  assign n17245 = n14906 ^ n3274 ^ n2894 ;
  assign n17246 = ( ~n3289 & n17244 ) | ( ~n3289 & n17245 ) | ( n17244 & n17245 ) ;
  assign n17247 = n14701 ^ n7027 ^ n165 ;
  assign n17248 = n15525 ^ n9058 ^ n5928 ;
  assign n17249 = ( n1366 & n16648 ) | ( n1366 & n17248 ) | ( n16648 & n17248 ) ;
  assign n17250 = n17249 ^ n10645 ^ n975 ;
  assign n17251 = n17250 ^ n13859 ^ n5206 ;
  assign n17252 = ( ~n5483 & n15003 ) | ( ~n5483 & n17251 ) | ( n15003 & n17251 ) ;
  assign n17253 = n17252 ^ n15845 ^ n2325 ;
  assign n17254 = n17253 ^ n13400 ^ n363 ;
  assign n17255 = n11673 ^ n5935 ^ n838 ;
  assign n17256 = ( ~n2313 & n5258 ) | ( ~n2313 & n5700 ) | ( n5258 & n5700 ) ;
  assign n17257 = ( n5161 & n7171 ) | ( n5161 & ~n16239 ) | ( n7171 & ~n16239 ) ;
  assign n17258 = ( n3765 & n17256 ) | ( n3765 & ~n17257 ) | ( n17256 & ~n17257 ) ;
  assign n17259 = n2821 ^ n2378 ^ n1285 ;
  assign n17260 = n17259 ^ n11771 ^ n8890 ;
  assign n17261 = ( n14476 & ~n17258 ) | ( n14476 & n17260 ) | ( ~n17258 & n17260 ) ;
  assign n17262 = ( n439 & n3931 ) | ( n439 & ~n16733 ) | ( n3931 & ~n16733 ) ;
  assign n17263 = n17262 ^ n6473 ^ n3766 ;
  assign n17264 = n7999 ^ n7796 ^ x65 ;
  assign n17265 = ( n3143 & n17116 ) | ( n3143 & ~n17264 ) | ( n17116 & ~n17264 ) ;
  assign n17266 = n10632 ^ n8986 ^ n3177 ;
  assign n17267 = ( ~n4069 & n5280 ) | ( ~n4069 & n10144 ) | ( n5280 & n10144 ) ;
  assign n17268 = ( ~n11944 & n12446 ) | ( ~n11944 & n17267 ) | ( n12446 & n17267 ) ;
  assign n17272 = ( n1763 & n4513 ) | ( n1763 & ~n11487 ) | ( n4513 & ~n11487 ) ;
  assign n17271 = ( x56 & ~n968 ) | ( x56 & n11054 ) | ( ~n968 & n11054 ) ;
  assign n17269 = ( n1830 & ~n2535 ) | ( n1830 & n7109 ) | ( ~n2535 & n7109 ) ;
  assign n17270 = ( n6285 & n14377 ) | ( n6285 & n17269 ) | ( n14377 & n17269 ) ;
  assign n17273 = n17272 ^ n17271 ^ n17270 ;
  assign n17274 = ( n5578 & n17268 ) | ( n5578 & ~n17273 ) | ( n17268 & ~n17273 ) ;
  assign n17275 = ( n2148 & n6793 ) | ( n2148 & n8890 ) | ( n6793 & n8890 ) ;
  assign n17276 = n4784 ^ n4234 ^ n3238 ;
  assign n17277 = n17276 ^ n4661 ^ n2315 ;
  assign n17278 = ( n185 & n350 ) | ( n185 & n9301 ) | ( n350 & n9301 ) ;
  assign n17279 = n17278 ^ n8160 ^ n205 ;
  assign n17280 = ( ~n17275 & n17277 ) | ( ~n17275 & n17279 ) | ( n17277 & n17279 ) ;
  assign n17281 = n11159 ^ n1915 ^ n1185 ;
  assign n17282 = ( ~n1323 & n14760 ) | ( ~n1323 & n17281 ) | ( n14760 & n17281 ) ;
  assign n17283 = ( n5058 & ~n7205 ) | ( n5058 & n17282 ) | ( ~n7205 & n17282 ) ;
  assign n17284 = n14451 ^ n3611 ^ n3315 ;
  assign n17285 = n4757 ^ n965 ^ n740 ;
  assign n17290 = ( ~n3655 & n4342 ) | ( ~n3655 & n5730 ) | ( n4342 & n5730 ) ;
  assign n17289 = ( ~n3196 & n4243 ) | ( ~n3196 & n16411 ) | ( n4243 & n16411 ) ;
  assign n17291 = n17290 ^ n17289 ^ n10345 ;
  assign n17288 = ( n4115 & n14273 ) | ( n4115 & ~n15066 ) | ( n14273 & ~n15066 ) ;
  assign n17286 = n11702 ^ n6598 ^ n473 ;
  assign n17287 = n17286 ^ n15849 ^ n7538 ;
  assign n17292 = n17291 ^ n17288 ^ n17287 ;
  assign n17293 = ( n1140 & n1374 ) | ( n1140 & ~n3517 ) | ( n1374 & ~n3517 ) ;
  assign n17294 = n17293 ^ n15894 ^ n15431 ;
  assign n17295 = n17294 ^ n10698 ^ n9794 ;
  assign n17296 = ( n3058 & n7086 ) | ( n3058 & ~n9579 ) | ( n7086 & ~n9579 ) ;
  assign n17297 = ( n1583 & n5869 ) | ( n1583 & ~n11256 ) | ( n5869 & ~n11256 ) ;
  assign n17298 = ( n2144 & n2663 ) | ( n2144 & ~n17297 ) | ( n2663 & ~n17297 ) ;
  assign n17299 = ( n3686 & n13020 ) | ( n3686 & n17122 ) | ( n13020 & n17122 ) ;
  assign n17300 = ( n2373 & n17298 ) | ( n2373 & n17299 ) | ( n17298 & n17299 ) ;
  assign n17301 = n17083 ^ n13101 ^ n12341 ;
  assign n17302 = ( ~n1372 & n2932 ) | ( ~n1372 & n10031 ) | ( n2932 & n10031 ) ;
  assign n17303 = n17302 ^ n11621 ^ n10856 ;
  assign n17304 = ( n4957 & ~n15183 ) | ( n4957 & n15848 ) | ( ~n15183 & n15848 ) ;
  assign n17305 = n5540 ^ n4372 ^ n3809 ;
  assign n17306 = ( n3530 & n3746 ) | ( n3530 & n17305 ) | ( n3746 & n17305 ) ;
  assign n17307 = ( n8084 & n17304 ) | ( n8084 & ~n17306 ) | ( n17304 & ~n17306 ) ;
  assign n17308 = ( ~n198 & n3555 ) | ( ~n198 & n13972 ) | ( n3555 & n13972 ) ;
  assign n17309 = ( n16773 & ~n17307 ) | ( n16773 & n17308 ) | ( ~n17307 & n17308 ) ;
  assign n17310 = n10574 ^ n5314 ^ n335 ;
  assign n17311 = n17310 ^ n15057 ^ n12704 ;
  assign n17312 = ( n6422 & n12589 ) | ( n6422 & n14753 ) | ( n12589 & n14753 ) ;
  assign n17313 = ( n11703 & ~n13381 ) | ( n11703 & n16181 ) | ( ~n13381 & n16181 ) ;
  assign n17314 = ( n6077 & n6462 ) | ( n6077 & ~n11181 ) | ( n6462 & ~n11181 ) ;
  assign n17315 = ( ~n3597 & n12838 ) | ( ~n3597 & n13241 ) | ( n12838 & n13241 ) ;
  assign n17316 = ( n5794 & n17288 ) | ( n5794 & n17315 ) | ( n17288 & n17315 ) ;
  assign n17317 = ( ~n14055 & n17314 ) | ( ~n14055 & n17316 ) | ( n17314 & n17316 ) ;
  assign n17319 = n11437 ^ n9510 ^ n3088 ;
  assign n17318 = n6405 ^ n5572 ^ n1147 ;
  assign n17320 = n17319 ^ n17318 ^ n6254 ;
  assign n17321 = n11444 ^ n10948 ^ n4421 ;
  assign n17322 = ( n2973 & ~n7850 ) | ( n2973 & n8384 ) | ( ~n7850 & n8384 ) ;
  assign n17323 = n17322 ^ n13203 ^ n12590 ;
  assign n17324 = ( n12267 & ~n16991 ) | ( n12267 & n17323 ) | ( ~n16991 & n17323 ) ;
  assign n17325 = ( ~n5200 & n5485 ) | ( ~n5200 & n7074 ) | ( n5485 & n7074 ) ;
  assign n17326 = ( n9420 & ~n10026 ) | ( n9420 & n17325 ) | ( ~n10026 & n17325 ) ;
  assign n17327 = ( n4745 & n15090 ) | ( n4745 & ~n15166 ) | ( n15090 & ~n15166 ) ;
  assign n17328 = ( n2037 & n17326 ) | ( n2037 & ~n17327 ) | ( n17326 & ~n17327 ) ;
  assign n17329 = n17328 ^ n3837 ^ n911 ;
  assign n17330 = n16420 ^ n10607 ^ n8590 ;
  assign n17332 = ( ~n3152 & n11680 ) | ( ~n3152 & n13022 ) | ( n11680 & n13022 ) ;
  assign n17331 = n13053 ^ n10043 ^ n9354 ;
  assign n17333 = n17332 ^ n17331 ^ n1946 ;
  assign n17334 = ( n3988 & n4354 ) | ( n3988 & n17333 ) | ( n4354 & n17333 ) ;
  assign n17335 = n12385 ^ n10657 ^ n7636 ;
  assign n17336 = ( n2421 & ~n4988 ) | ( n2421 & n17335 ) | ( ~n4988 & n17335 ) ;
  assign n17339 = n15013 ^ n11027 ^ n5226 ;
  assign n17338 = n10500 ^ n7453 ^ n2076 ;
  assign n17337 = n15472 ^ n6013 ^ n5708 ;
  assign n17340 = n17339 ^ n17338 ^ n17337 ;
  assign n17341 = n11501 ^ n8064 ^ n6623 ;
  assign n17342 = n17341 ^ n2322 ^ n1989 ;
  assign n17343 = n10664 ^ n2871 ^ n1812 ;
  assign n17344 = ( n1796 & ~n4044 ) | ( n1796 & n11872 ) | ( ~n4044 & n11872 ) ;
  assign n17345 = ( ~n13039 & n17343 ) | ( ~n13039 & n17344 ) | ( n17343 & n17344 ) ;
  assign n17346 = n17345 ^ n11357 ^ n9282 ;
  assign n17347 = n15953 ^ n3548 ^ n2672 ;
  assign n17348 = ( ~n2435 & n4848 ) | ( ~n2435 & n17347 ) | ( n4848 & n17347 ) ;
  assign n17349 = n17348 ^ n10551 ^ n7457 ;
  assign n17350 = ( n2405 & ~n5329 ) | ( n2405 & n17349 ) | ( ~n5329 & n17349 ) ;
  assign n17351 = n9021 ^ n8438 ^ n6375 ;
  assign n17352 = n17351 ^ n16288 ^ n15551 ;
  assign n17353 = ( ~n2647 & n3232 ) | ( ~n2647 & n17352 ) | ( n3232 & n17352 ) ;
  assign n17354 = ( n315 & n13016 ) | ( n315 & n17353 ) | ( n13016 & n17353 ) ;
  assign n17355 = n12984 ^ n7368 ^ n4485 ;
  assign n17360 = n9099 ^ n1961 ^ n1568 ;
  assign n17361 = n17360 ^ n6464 ^ n1029 ;
  assign n17359 = ( n2474 & n5016 ) | ( n2474 & ~n16044 ) | ( n5016 & ~n16044 ) ;
  assign n17357 = ( ~n7563 & n8511 ) | ( ~n7563 & n13842 ) | ( n8511 & n13842 ) ;
  assign n17356 = ( ~n4983 & n10350 ) | ( ~n4983 & n13536 ) | ( n10350 & n13536 ) ;
  assign n17358 = n17357 ^ n17356 ^ n11976 ;
  assign n17362 = n17361 ^ n17359 ^ n17358 ;
  assign n17366 = ( ~n932 & n1731 ) | ( ~n932 & n2178 ) | ( n1731 & n2178 ) ;
  assign n17363 = n10667 ^ n6602 ^ n4828 ;
  assign n17364 = n17363 ^ n5074 ^ n1260 ;
  assign n17365 = n17364 ^ n11213 ^ n8688 ;
  assign n17367 = n17366 ^ n17365 ^ n11000 ;
  assign n17368 = ( n1240 & n5802 ) | ( n1240 & ~n9929 ) | ( n5802 & ~n9929 ) ;
  assign n17369 = ( ~n1993 & n7427 ) | ( ~n1993 & n17368 ) | ( n7427 & n17368 ) ;
  assign n17370 = n7010 ^ n3401 ^ n1426 ;
  assign n17371 = n8488 ^ n3984 ^ n2358 ;
  assign n17372 = ( n7810 & n15872 ) | ( n7810 & ~n17371 ) | ( n15872 & ~n17371 ) ;
  assign n17373 = ( n3102 & ~n12235 ) | ( n3102 & n17372 ) | ( ~n12235 & n17372 ) ;
  assign n17374 = n17373 ^ n12637 ^ n6762 ;
  assign n17375 = n17374 ^ n15737 ^ n5489 ;
  assign n17376 = ( ~n3741 & n17370 ) | ( ~n3741 & n17375 ) | ( n17370 & n17375 ) ;
  assign n17377 = ( ~n6262 & n7409 ) | ( ~n6262 & n17376 ) | ( n7409 & n17376 ) ;
  assign n17378 = n16014 ^ n1899 ^ x105 ;
  assign n17379 = n6987 ^ n3034 ^ x64 ;
  assign n17380 = n17379 ^ n5903 ^ n481 ;
  assign n17381 = n11412 ^ n5259 ^ n1503 ;
  assign n17382 = ( ~n10572 & n10627 ) | ( ~n10572 & n17381 ) | ( n10627 & n17381 ) ;
  assign n17383 = ( n3475 & n7363 ) | ( n3475 & ~n8475 ) | ( n7363 & ~n8475 ) ;
  assign n17384 = ( n12801 & ~n13096 ) | ( n12801 & n17383 ) | ( ~n13096 & n17383 ) ;
  assign n17385 = n15678 ^ n13726 ^ n7473 ;
  assign n17386 = ( n10624 & n12291 ) | ( n10624 & ~n14927 ) | ( n12291 & ~n14927 ) ;
  assign n17387 = n17386 ^ n11956 ^ n11111 ;
  assign n17388 = ( ~n7195 & n15719 ) | ( ~n7195 & n17387 ) | ( n15719 & n17387 ) ;
  assign n17390 = n5913 ^ n3142 ^ n372 ;
  assign n17391 = ( ~n9852 & n12532 ) | ( ~n9852 & n17390 ) | ( n12532 & n17390 ) ;
  assign n17392 = ( n1668 & ~n12297 ) | ( n1668 & n17391 ) | ( ~n12297 & n17391 ) ;
  assign n17393 = ( ~n2064 & n14042 ) | ( ~n2064 & n17392 ) | ( n14042 & n17392 ) ;
  assign n17389 = n7444 ^ n6660 ^ n4941 ;
  assign n17394 = n17393 ^ n17389 ^ n3374 ;
  assign n17395 = ( ~n3979 & n6570 ) | ( ~n3979 & n7719 ) | ( n6570 & n7719 ) ;
  assign n17396 = ( ~n9297 & n14271 ) | ( ~n9297 & n17395 ) | ( n14271 & n17395 ) ;
  assign n17400 = n4859 ^ n2236 ^ n1840 ;
  assign n17398 = n13510 ^ n12824 ^ n8210 ;
  assign n17399 = n17398 ^ n1754 ^ n208 ;
  assign n17401 = n17400 ^ n17399 ^ n6605 ;
  assign n17397 = ( n3786 & n12444 ) | ( n3786 & ~n14579 ) | ( n12444 & ~n14579 ) ;
  assign n17402 = n17401 ^ n17397 ^ n16086 ;
  assign n17403 = ( n249 & n4974 ) | ( n249 & ~n8036 ) | ( n4974 & ~n8036 ) ;
  assign n17404 = n17403 ^ n11551 ^ n3016 ;
  assign n17405 = n15204 ^ n8154 ^ n130 ;
  assign n17406 = ( n7292 & ~n10983 ) | ( n7292 & n17405 ) | ( ~n10983 & n17405 ) ;
  assign n17411 = ( n499 & n1231 ) | ( n499 & ~n10346 ) | ( n1231 & ~n10346 ) ;
  assign n17412 = ( n1287 & ~n6036 ) | ( n1287 & n17411 ) | ( ~n6036 & n17411 ) ;
  assign n17408 = ( n3237 & n4092 ) | ( n3237 & n8025 ) | ( n4092 & n8025 ) ;
  assign n17409 = ( ~n232 & n4371 ) | ( ~n232 & n17408 ) | ( n4371 & n17408 ) ;
  assign n17410 = ( n8802 & n13825 ) | ( n8802 & n17409 ) | ( n13825 & n17409 ) ;
  assign n17407 = ( n271 & ~n4290 ) | ( n271 & n16586 ) | ( ~n4290 & n16586 ) ;
  assign n17413 = n17412 ^ n17410 ^ n17407 ;
  assign n17414 = n9803 ^ n6502 ^ n6421 ;
  assign n17415 = n17414 ^ n11830 ^ n10875 ;
  assign n17416 = ( n4525 & n6469 ) | ( n4525 & n15495 ) | ( n6469 & n15495 ) ;
  assign n17417 = ( ~n506 & n858 ) | ( ~n506 & n17416 ) | ( n858 & n17416 ) ;
  assign n17418 = ( n1226 & n2139 ) | ( n1226 & n3066 ) | ( n2139 & n3066 ) ;
  assign n17419 = ( n10472 & n11120 ) | ( n10472 & n11283 ) | ( n11120 & n11283 ) ;
  assign n17420 = ( ~n4909 & n7853 ) | ( ~n4909 & n17419 ) | ( n7853 & n17419 ) ;
  assign n17421 = n9050 ^ n8518 ^ n2354 ;
  assign n17422 = n16388 ^ n11193 ^ n1279 ;
  assign n17423 = ( n5921 & n17421 ) | ( n5921 & ~n17422 ) | ( n17421 & ~n17422 ) ;
  assign n17424 = ( ~n729 & n3944 ) | ( ~n729 & n4375 ) | ( n3944 & n4375 ) ;
  assign n17425 = n7059 ^ n5438 ^ n4722 ;
  assign n17426 = n17425 ^ n13481 ^ n12989 ;
  assign n17427 = n17426 ^ n15923 ^ n2450 ;
  assign n17428 = n11485 ^ n7479 ^ n2228 ;
  assign n17429 = ( n1562 & n1779 ) | ( n1562 & n5006 ) | ( n1779 & n5006 ) ;
  assign n17430 = n12569 ^ n10412 ^ n2547 ;
  assign n17431 = ( n2117 & n17429 ) | ( n2117 & n17430 ) | ( n17429 & n17430 ) ;
  assign n17432 = n17431 ^ n2280 ^ n890 ;
  assign n17433 = ( n1760 & n17428 ) | ( n1760 & n17432 ) | ( n17428 & n17432 ) ;
  assign n17434 = ( n2097 & n4602 ) | ( n2097 & n6360 ) | ( n4602 & n6360 ) ;
  assign n17435 = ( n2280 & n7495 ) | ( n2280 & n7554 ) | ( n7495 & n7554 ) ;
  assign n17436 = ( n789 & n3822 ) | ( n789 & n17435 ) | ( n3822 & n17435 ) ;
  assign n17437 = ( n2646 & ~n17434 ) | ( n2646 & n17436 ) | ( ~n17434 & n17436 ) ;
  assign n17438 = n17166 ^ n8994 ^ n8386 ;
  assign n17439 = n13821 ^ n8131 ^ n3218 ;
  assign n17440 = ( ~n1296 & n10346 ) | ( ~n1296 & n17439 ) | ( n10346 & n17439 ) ;
  assign n17444 = ( n637 & n1219 ) | ( n637 & n3228 ) | ( n1219 & n3228 ) ;
  assign n17441 = n3835 ^ n2810 ^ n1532 ;
  assign n17442 = n17441 ^ n6227 ^ n3867 ;
  assign n17443 = ( n5215 & ~n10216 ) | ( n5215 & n17442 ) | ( ~n10216 & n17442 ) ;
  assign n17445 = n17444 ^ n17443 ^ n5073 ;
  assign n17446 = n13684 ^ n9788 ^ n6042 ;
  assign n17449 = n15714 ^ n15065 ^ n7918 ;
  assign n17447 = n6725 ^ n4492 ^ n576 ;
  assign n17448 = ( n3539 & n5313 ) | ( n3539 & ~n17447 ) | ( n5313 & ~n17447 ) ;
  assign n17450 = n17449 ^ n17448 ^ n15216 ;
  assign n17451 = n9334 ^ n6435 ^ n1562 ;
  assign n17452 = ( n1411 & n5168 ) | ( n1411 & ~n10694 ) | ( n5168 & ~n10694 ) ;
  assign n17453 = ( ~n3596 & n10401 ) | ( ~n3596 & n17452 ) | ( n10401 & n17452 ) ;
  assign n17454 = n17453 ^ n11948 ^ n3789 ;
  assign n17455 = ( n9074 & n17451 ) | ( n9074 & ~n17454 ) | ( n17451 & ~n17454 ) ;
  assign n17456 = n16823 ^ n9056 ^ n9051 ;
  assign n17457 = ( n5741 & ~n7638 ) | ( n5741 & n17456 ) | ( ~n7638 & n17456 ) ;
  assign n17462 = n14277 ^ n3407 ^ n2043 ;
  assign n17463 = n17462 ^ n7628 ^ n754 ;
  assign n17464 = n17463 ^ n5283 ^ n1985 ;
  assign n17459 = ( n1154 & n3641 ) | ( n1154 & n11200 ) | ( n3641 & n11200 ) ;
  assign n17460 = ( ~n8366 & n9075 ) | ( ~n8366 & n17459 ) | ( n9075 & n17459 ) ;
  assign n17458 = ( ~n7777 & n11813 ) | ( ~n7777 & n14693 ) | ( n11813 & n14693 ) ;
  assign n17461 = n17460 ^ n17458 ^ n5134 ;
  assign n17465 = n17464 ^ n17461 ^ n13042 ;
  assign n17466 = ( n5587 & ~n9238 ) | ( n5587 & n14128 ) | ( ~n9238 & n14128 ) ;
  assign n17467 = ( n3111 & n8314 ) | ( n3111 & ~n17466 ) | ( n8314 & ~n17466 ) ;
  assign n17468 = n13333 ^ n4293 ^ n670 ;
  assign n17469 = ( n12453 & n17467 ) | ( n12453 & ~n17468 ) | ( n17467 & ~n17468 ) ;
  assign n17470 = ( n3683 & n10950 ) | ( n3683 & n11336 ) | ( n10950 & n11336 ) ;
  assign n17471 = n17470 ^ n6329 ^ n2388 ;
  assign n17472 = ( n6957 & ~n14045 ) | ( n6957 & n17471 ) | ( ~n14045 & n17471 ) ;
  assign n17473 = n13598 ^ n4782 ^ n482 ;
  assign n17474 = n14282 ^ n9709 ^ n1241 ;
  assign n17475 = ( n7522 & ~n9742 ) | ( n7522 & n16659 ) | ( ~n9742 & n16659 ) ;
  assign n17476 = ( n17271 & ~n17474 ) | ( n17271 & n17475 ) | ( ~n17474 & n17475 ) ;
  assign n17477 = ( n12670 & n17473 ) | ( n12670 & ~n17476 ) | ( n17473 & ~n17476 ) ;
  assign n17478 = ( n1674 & n5142 ) | ( n1674 & n11717 ) | ( n5142 & n11717 ) ;
  assign n17479 = ( n6425 & ~n10363 ) | ( n6425 & n12440 ) | ( ~n10363 & n12440 ) ;
  assign n17480 = ( n8881 & n17168 ) | ( n8881 & ~n17479 ) | ( n17168 & ~n17479 ) ;
  assign n17488 = ( n3800 & ~n9554 ) | ( n3800 & n12600 ) | ( ~n9554 & n12600 ) ;
  assign n17489 = n17488 ^ n7635 ^ n4303 ;
  assign n17490 = ( n2112 & n6648 ) | ( n2112 & ~n17489 ) | ( n6648 & ~n17489 ) ;
  assign n17491 = n17490 ^ n10793 ^ n605 ;
  assign n17486 = n6972 ^ n1795 ^ n758 ;
  assign n17487 = ( n753 & n15603 ) | ( n753 & n17486 ) | ( n15603 & n17486 ) ;
  assign n17492 = n17491 ^ n17487 ^ n987 ;
  assign n17481 = n13739 ^ n11408 ^ n10827 ;
  assign n17483 = n2348 ^ n1391 ^ n382 ;
  assign n17482 = n13558 ^ n11142 ^ n5825 ;
  assign n17484 = n17483 ^ n17482 ^ n13686 ;
  assign n17485 = ( n7057 & ~n17481 ) | ( n7057 & n17484 ) | ( ~n17481 & n17484 ) ;
  assign n17493 = n17492 ^ n17485 ^ n3467 ;
  assign n17497 = ( n401 & n7263 ) | ( n401 & ~n11993 ) | ( n7263 & ~n11993 ) ;
  assign n17496 = ( n629 & ~n8159 ) | ( n629 & n16076 ) | ( ~n8159 & n16076 ) ;
  assign n17494 = n8838 ^ n6947 ^ n4218 ;
  assign n17495 = ( n6154 & n9228 ) | ( n6154 & ~n17494 ) | ( n9228 & ~n17494 ) ;
  assign n17498 = n17497 ^ n17496 ^ n17495 ;
  assign n17499 = n17498 ^ n10354 ^ n1841 ;
  assign n17500 = n10837 ^ n1396 ^ n1147 ;
  assign n17501 = ( n4101 & ~n16059 ) | ( n4101 & n17500 ) | ( ~n16059 & n17500 ) ;
  assign n17502 = n17501 ^ n8062 ^ n3535 ;
  assign n17503 = ( n293 & ~n3600 ) | ( n293 & n3620 ) | ( ~n3600 & n3620 ) ;
  assign n17504 = n17503 ^ n11718 ^ n1529 ;
  assign n17505 = n17504 ^ n2395 ^ n2147 ;
  assign n17506 = ( n6106 & n9163 ) | ( n6106 & n16045 ) | ( n9163 & n16045 ) ;
  assign n17507 = n15544 ^ n4873 ^ n3485 ;
  assign n17508 = ( n5390 & n8192 ) | ( n5390 & ~n17507 ) | ( n8192 & ~n17507 ) ;
  assign n17509 = ( n5348 & n16214 ) | ( n5348 & ~n17508 ) | ( n16214 & ~n17508 ) ;
  assign n17510 = ( n823 & n851 ) | ( n823 & n4920 ) | ( n851 & n4920 ) ;
  assign n17511 = n17510 ^ n7709 ^ n7018 ;
  assign n17512 = ( n2208 & n8363 ) | ( n2208 & ~n17511 ) | ( n8363 & ~n17511 ) ;
  assign n17513 = ( ~n2475 & n8016 ) | ( ~n2475 & n12285 ) | ( n8016 & n12285 ) ;
  assign n17514 = n17513 ^ n9069 ^ n4069 ;
  assign n17515 = n15143 ^ n9737 ^ n6645 ;
  assign n17516 = ( ~x5 & n1195 ) | ( ~x5 & n2285 ) | ( n1195 & n2285 ) ;
  assign n17517 = ( ~n1935 & n5406 ) | ( ~n1935 & n16906 ) | ( n5406 & n16906 ) ;
  assign n17518 = ( n4804 & n6045 ) | ( n4804 & n10092 ) | ( n6045 & n10092 ) ;
  assign n17519 = n17518 ^ n16875 ^ n2747 ;
  assign n17520 = n15921 ^ n7507 ^ n5203 ;
  assign n17521 = ( n1278 & n6651 ) | ( n1278 & ~n11197 ) | ( n6651 & ~n11197 ) ;
  assign n17522 = n17521 ^ n10054 ^ n9151 ;
  assign n17523 = ( n2166 & n3744 ) | ( n2166 & ~n4363 ) | ( n3744 & ~n4363 ) ;
  assign n17524 = n17523 ^ n6883 ^ n5360 ;
  assign n17525 = ( n1122 & n1765 ) | ( n1122 & n13766 ) | ( n1765 & n13766 ) ;
  assign n17526 = ( ~n7336 & n17524 ) | ( ~n7336 & n17525 ) | ( n17524 & n17525 ) ;
  assign n17527 = ( n8951 & n17522 ) | ( n8951 & n17526 ) | ( n17522 & n17526 ) ;
  assign n17528 = ( n189 & n946 ) | ( n189 & ~n6852 ) | ( n946 & ~n6852 ) ;
  assign n17529 = ( n4780 & ~n10472 ) | ( n4780 & n12595 ) | ( ~n10472 & n12595 ) ;
  assign n17530 = n17529 ^ n13926 ^ n2445 ;
  assign n17531 = ( n16130 & n17528 ) | ( n16130 & ~n17530 ) | ( n17528 & ~n17530 ) ;
  assign n17537 = n13745 ^ n7049 ^ n5959 ;
  assign n17538 = n16815 ^ n13762 ^ n2376 ;
  assign n17539 = n10495 ^ n7510 ^ n6163 ;
  assign n17540 = n17539 ^ n10043 ^ n4650 ;
  assign n17541 = ( n17537 & ~n17538 ) | ( n17537 & n17540 ) | ( ~n17538 & n17540 ) ;
  assign n17534 = n6855 ^ n5041 ^ n3238 ;
  assign n17535 = n17534 ^ n7447 ^ n1127 ;
  assign n17533 = ( n13607 & n13761 ) | ( n13607 & n14432 ) | ( n13761 & n14432 ) ;
  assign n17532 = n9243 ^ n7918 ^ n3873 ;
  assign n17536 = n17535 ^ n17533 ^ n17532 ;
  assign n17542 = n17541 ^ n17536 ^ n15530 ;
  assign n17544 = n12862 ^ n9204 ^ n1960 ;
  assign n17545 = n17544 ^ n9098 ^ n7311 ;
  assign n17543 = ( n1489 & ~n5424 ) | ( n1489 & n10301 ) | ( ~n5424 & n10301 ) ;
  assign n17546 = n17545 ^ n17543 ^ n466 ;
  assign n17547 = ( ~n674 & n2967 ) | ( ~n674 & n4785 ) | ( n2967 & n4785 ) ;
  assign n17548 = ( n3862 & ~n6443 ) | ( n3862 & n13928 ) | ( ~n6443 & n13928 ) ;
  assign n17549 = ( n5508 & ~n9059 ) | ( n5508 & n17548 ) | ( ~n9059 & n17548 ) ;
  assign n17550 = ( n6299 & ~n17547 ) | ( n6299 & n17549 ) | ( ~n17547 & n17549 ) ;
  assign n17551 = n6584 ^ n1786 ^ n1114 ;
  assign n17552 = ( n594 & ~n1233 ) | ( n594 & n17551 ) | ( ~n1233 & n17551 ) ;
  assign n17554 = ( n1796 & ~n2264 ) | ( n1796 & n4634 ) | ( ~n2264 & n4634 ) ;
  assign n17553 = n16712 ^ n15722 ^ n1165 ;
  assign n17555 = n17554 ^ n17553 ^ n10910 ;
  assign n17556 = ( n16109 & n17552 ) | ( n16109 & ~n17555 ) | ( n17552 & ~n17555 ) ;
  assign n17559 = n12282 ^ n9172 ^ n6294 ;
  assign n17557 = n5221 ^ n4108 ^ n1478 ;
  assign n17558 = n17557 ^ n9222 ^ n1945 ;
  assign n17560 = n17559 ^ n17558 ^ n5506 ;
  assign n17561 = ( ~n4891 & n12305 ) | ( ~n4891 & n16163 ) | ( n12305 & n16163 ) ;
  assign n17562 = ( n8873 & ~n17386 ) | ( n8873 & n17561 ) | ( ~n17386 & n17561 ) ;
  assign n17563 = ( n5817 & ~n11910 ) | ( n5817 & n17562 ) | ( ~n11910 & n17562 ) ;
  assign n17564 = ( n4345 & n5449 ) | ( n4345 & ~n6416 ) | ( n5449 & ~n6416 ) ;
  assign n17565 = n17564 ^ n10482 ^ n5311 ;
  assign n17567 = n14921 ^ n8694 ^ n2342 ;
  assign n17566 = n10922 ^ n8994 ^ n6406 ;
  assign n17568 = n17567 ^ n17566 ^ n16585 ;
  assign n17569 = ( n4796 & n11114 ) | ( n4796 & n15023 ) | ( n11114 & n15023 ) ;
  assign n17570 = n17569 ^ n6028 ^ n6009 ;
  assign n17571 = ( ~n9707 & n13931 ) | ( ~n9707 & n17570 ) | ( n13931 & n17570 ) ;
  assign n17572 = n17571 ^ n11347 ^ n8571 ;
  assign n17575 = ( n832 & n5891 ) | ( n832 & ~n10266 ) | ( n5891 & ~n10266 ) ;
  assign n17573 = n14753 ^ n5173 ^ n1910 ;
  assign n17574 = ( ~n12879 & n16091 ) | ( ~n12879 & n17573 ) | ( n16091 & n17573 ) ;
  assign n17576 = n17575 ^ n17574 ^ n14696 ;
  assign n17584 = ( n2891 & n4504 ) | ( n2891 & n16959 ) | ( n4504 & n16959 ) ;
  assign n17585 = n11854 ^ n11089 ^ n2652 ;
  assign n17586 = ( ~n10908 & n17584 ) | ( ~n10908 & n17585 ) | ( n17584 & n17585 ) ;
  assign n17577 = n7094 ^ n5734 ^ n2889 ;
  assign n17578 = ( n4647 & ~n5522 ) | ( n4647 & n17577 ) | ( ~n5522 & n17577 ) ;
  assign n17579 = n9733 ^ n2137 ^ n1941 ;
  assign n17580 = ( ~n2699 & n5327 ) | ( ~n2699 & n17579 ) | ( n5327 & n17579 ) ;
  assign n17581 = n17580 ^ n15166 ^ n4768 ;
  assign n17582 = n17581 ^ n17401 ^ n17390 ;
  assign n17583 = ( n1078 & n17578 ) | ( n1078 & n17582 ) | ( n17578 & n17582 ) ;
  assign n17587 = n17586 ^ n17583 ^ n16850 ;
  assign n17588 = ( n13417 & n15199 ) | ( n13417 & n17466 ) | ( n15199 & n17466 ) ;
  assign n17589 = ( x35 & ~n1239 ) | ( x35 & n6857 ) | ( ~n1239 & n6857 ) ;
  assign n17590 = ( ~n14607 & n15202 ) | ( ~n14607 & n17589 ) | ( n15202 & n17589 ) ;
  assign n17591 = n10838 ^ n6546 ^ n2557 ;
  assign n17592 = n16222 ^ n8415 ^ n5110 ;
  assign n17593 = ( n10345 & ~n17591 ) | ( n10345 & n17592 ) | ( ~n17591 & n17592 ) ;
  assign n17594 = ( ~n1817 & n16101 ) | ( ~n1817 & n17593 ) | ( n16101 & n17593 ) ;
  assign n17598 = n9623 ^ n3001 ^ n455 ;
  assign n17595 = ( n1069 & n8791 ) | ( n1069 & n9957 ) | ( n8791 & n9957 ) ;
  assign n17596 = ( n4015 & n7912 ) | ( n4015 & ~n17595 ) | ( n7912 & ~n17595 ) ;
  assign n17597 = ( n4340 & ~n16006 ) | ( n4340 & n17596 ) | ( ~n16006 & n17596 ) ;
  assign n17599 = n17598 ^ n17597 ^ n15798 ;
  assign n17600 = n9710 ^ n5935 ^ n4936 ;
  assign n17601 = n17600 ^ n15736 ^ n8507 ;
  assign n17602 = ( n6480 & n8380 ) | ( n6480 & n9383 ) | ( n8380 & n9383 ) ;
  assign n17603 = n15342 ^ n1575 ^ n348 ;
  assign n17604 = ( ~n7253 & n17602 ) | ( ~n7253 & n17603 ) | ( n17602 & n17603 ) ;
  assign n17605 = ( n7865 & ~n13137 ) | ( n7865 & n17604 ) | ( ~n13137 & n17604 ) ;
  assign n17606 = n14870 ^ n8534 ^ n2831 ;
  assign n17607 = ( n6353 & n7525 ) | ( n6353 & ~n17606 ) | ( n7525 & ~n17606 ) ;
  assign n17608 = n13223 ^ n4558 ^ n3737 ;
  assign n17609 = ( n1072 & n1219 ) | ( n1072 & n8688 ) | ( n1219 & n8688 ) ;
  assign n17610 = n17609 ^ n10950 ^ n5058 ;
  assign n17611 = n13451 ^ n2137 ^ n396 ;
  assign n17612 = n17611 ^ n8376 ^ n794 ;
  assign n17613 = n17612 ^ n16229 ^ n11406 ;
  assign n17614 = ( n9539 & n17610 ) | ( n9539 & n17613 ) | ( n17610 & n17613 ) ;
  assign n17615 = ( n1006 & n9054 ) | ( n1006 & ~n17614 ) | ( n9054 & ~n17614 ) ;
  assign n17616 = n9236 ^ n5435 ^ n3740 ;
  assign n17617 = n17616 ^ n14520 ^ n7978 ;
  assign n17618 = ( n800 & ~n5146 ) | ( n800 & n11705 ) | ( ~n5146 & n11705 ) ;
  assign n17619 = n17618 ^ n11068 ^ n4358 ;
  assign n17638 = n13043 ^ n4806 ^ n2564 ;
  assign n17635 = n3533 ^ n1565 ^ n1277 ;
  assign n17636 = ( ~n209 & n2200 ) | ( ~n209 & n17635 ) | ( n2200 & n17635 ) ;
  assign n17631 = n4808 ^ n749 ^ n440 ;
  assign n17632 = n17631 ^ n14535 ^ n4936 ;
  assign n17633 = ( ~n449 & n2409 ) | ( ~n449 & n16799 ) | ( n2409 & n16799 ) ;
  assign n17634 = ( n1679 & n17632 ) | ( n1679 & ~n17633 ) | ( n17632 & ~n17633 ) ;
  assign n17620 = n13722 ^ n11596 ^ n5346 ;
  assign n17627 = n15865 ^ n15066 ^ n13292 ;
  assign n17626 = n17015 ^ n6992 ^ n6799 ;
  assign n17624 = ( n2061 & n5795 ) | ( n2061 & ~n9958 ) | ( n5795 & ~n9958 ) ;
  assign n17621 = n11479 ^ n7693 ^ n3001 ;
  assign n17622 = n17621 ^ n9813 ^ n2792 ;
  assign n17623 = ( n14250 & n17412 ) | ( n14250 & n17622 ) | ( n17412 & n17622 ) ;
  assign n17625 = n17624 ^ n17623 ^ n15742 ;
  assign n17628 = n17627 ^ n17626 ^ n17625 ;
  assign n17629 = n17628 ^ n4796 ^ n1270 ;
  assign n17630 = ( n5209 & n17620 ) | ( n5209 & n17629 ) | ( n17620 & n17629 ) ;
  assign n17637 = n17636 ^ n17634 ^ n17630 ;
  assign n17639 = n17638 ^ n17637 ^ n9108 ;
  assign n17640 = ( n4003 & n10328 ) | ( n4003 & ~n13499 ) | ( n10328 & ~n13499 ) ;
  assign n17641 = n17640 ^ n5190 ^ n2386 ;
  assign n17642 = n14960 ^ n10127 ^ n2512 ;
  assign n17643 = ( n333 & n10410 ) | ( n333 & ~n17642 ) | ( n10410 & ~n17642 ) ;
  assign n17644 = ( ~n5322 & n12548 ) | ( ~n5322 & n17643 ) | ( n12548 & n17643 ) ;
  assign n17645 = n17644 ^ n8518 ^ n4318 ;
  assign n17646 = ( n2451 & n17641 ) | ( n2451 & ~n17645 ) | ( n17641 & ~n17645 ) ;
  assign n17647 = n4838 ^ n2418 ^ n2118 ;
  assign n17648 = n9936 ^ n9292 ^ n2331 ;
  assign n17649 = ( n17521 & n17647 ) | ( n17521 & n17648 ) | ( n17647 & n17648 ) ;
  assign n17650 = n17649 ^ n6235 ^ n4631 ;
  assign n17651 = n8326 ^ n5245 ^ n1930 ;
  assign n17652 = ( n8992 & n17275 ) | ( n8992 & ~n17651 ) | ( n17275 & ~n17651 ) ;
  assign n17653 = ( n7426 & n8643 ) | ( n7426 & n17652 ) | ( n8643 & n17652 ) ;
  assign n17655 = ( n3683 & n8601 ) | ( n3683 & ~n13773 ) | ( n8601 & ~n13773 ) ;
  assign n17654 = ( n1693 & n7169 ) | ( n1693 & ~n8694 ) | ( n7169 & ~n8694 ) ;
  assign n17656 = n17655 ^ n17654 ^ n2996 ;
  assign n17657 = n17656 ^ n2372 ^ n1465 ;
  assign n17662 = n11527 ^ n9425 ^ n9329 ;
  assign n17658 = ( n5363 & n6146 ) | ( n5363 & n13114 ) | ( n6146 & n13114 ) ;
  assign n17659 = ( n3418 & ~n5351 ) | ( n3418 & n17658 ) | ( ~n5351 & n17658 ) ;
  assign n17660 = n9145 ^ n3380 ^ n3200 ;
  assign n17661 = ( ~n1604 & n17659 ) | ( ~n1604 & n17660 ) | ( n17659 & n17660 ) ;
  assign n17663 = n17662 ^ n17661 ^ n17273 ;
  assign n17664 = n5994 ^ n5048 ^ n3760 ;
  assign n17665 = ( ~n12631 & n13793 ) | ( ~n12631 & n17664 ) | ( n13793 & n17664 ) ;
  assign n17666 = ( n1876 & n3942 ) | ( n1876 & ~n3960 ) | ( n3942 & ~n3960 ) ;
  assign n17667 = ( n7677 & n13478 ) | ( n7677 & ~n16551 ) | ( n13478 & ~n16551 ) ;
  assign n17668 = ( n7088 & n11366 ) | ( n7088 & ~n15683 ) | ( n11366 & ~n15683 ) ;
  assign n17669 = n17668 ^ n6095 ^ n1741 ;
  assign n17670 = ( n257 & n12072 ) | ( n257 & ~n12337 ) | ( n12072 & ~n12337 ) ;
  assign n17671 = ( n633 & n1455 ) | ( n633 & ~n13516 ) | ( n1455 & ~n13516 ) ;
  assign n17672 = n17671 ^ n9619 ^ n4193 ;
  assign n17673 = n17672 ^ n6145 ^ n5455 ;
  assign n17674 = n12864 ^ n10028 ^ n6256 ;
  assign n17675 = n17674 ^ n8133 ^ n1535 ;
  assign n17676 = n16390 ^ n4769 ^ n4151 ;
  assign n17677 = ( n2554 & n8481 ) | ( n2554 & ~n9885 ) | ( n8481 & ~n9885 ) ;
  assign n17678 = n14758 ^ n9340 ^ n9082 ;
  assign n17679 = n13578 ^ n9881 ^ n6720 ;
  assign n17680 = ( ~n377 & n3968 ) | ( ~n377 & n17111 ) | ( n3968 & n17111 ) ;
  assign n17681 = ( n8634 & ~n12514 ) | ( n8634 & n17680 ) | ( ~n12514 & n17680 ) ;
  assign n17683 = n17267 ^ n15867 ^ n10269 ;
  assign n17682 = n7867 ^ n6618 ^ n5303 ;
  assign n17684 = n17683 ^ n17682 ^ n15550 ;
  assign n17685 = ( n2011 & n3796 ) | ( n2011 & ~n13797 ) | ( n3796 & ~n13797 ) ;
  assign n17686 = ( ~n12824 & n14254 ) | ( ~n12824 & n17685 ) | ( n14254 & n17685 ) ;
  assign n17687 = n17686 ^ n14976 ^ n907 ;
  assign n17688 = ( ~n3542 & n9467 ) | ( ~n3542 & n14967 ) | ( n9467 & n14967 ) ;
  assign n17689 = n17688 ^ n15613 ^ n11552 ;
  assign n17690 = ( ~n2581 & n10877 ) | ( ~n2581 & n14373 ) | ( n10877 & n14373 ) ;
  assign n17691 = n16870 ^ n10851 ^ n3792 ;
  assign n17692 = n17691 ^ n16081 ^ n2843 ;
  assign n17693 = n15790 ^ n12760 ^ n9786 ;
  assign n17694 = ( n1755 & n11913 ) | ( n1755 & n16643 ) | ( n11913 & n16643 ) ;
  assign n17695 = ( n897 & n6271 ) | ( n897 & n7669 ) | ( n6271 & n7669 ) ;
  assign n17696 = ( n17693 & n17694 ) | ( n17693 & ~n17695 ) | ( n17694 & ~n17695 ) ;
  assign n17697 = ( ~n6102 & n9389 ) | ( ~n6102 & n13654 ) | ( n9389 & n13654 ) ;
  assign n17698 = n17697 ^ n13521 ^ n13483 ;
  assign n17699 = n14422 ^ n14104 ^ n11921 ;
  assign n17700 = ( n4724 & n6907 ) | ( n4724 & n14199 ) | ( n6907 & n14199 ) ;
  assign n17701 = ( n1444 & n7541 ) | ( n1444 & ~n17700 ) | ( n7541 & ~n17700 ) ;
  assign n17702 = n13580 ^ n12150 ^ n6620 ;
  assign n17703 = ( n993 & n3052 ) | ( n993 & n17702 ) | ( n3052 & n17702 ) ;
  assign n17704 = n17703 ^ n11112 ^ n5803 ;
  assign n17705 = n10462 ^ n7827 ^ n6497 ;
  assign n17706 = ( n5408 & n17704 ) | ( n5408 & ~n17705 ) | ( n17704 & ~n17705 ) ;
  assign n17709 = ( ~n3774 & n7643 ) | ( ~n3774 & n12962 ) | ( n7643 & n12962 ) ;
  assign n17708 = n14066 ^ n13160 ^ n1724 ;
  assign n17710 = n17709 ^ n17708 ^ n12688 ;
  assign n17707 = n9660 ^ n6009 ^ n2993 ;
  assign n17711 = n17710 ^ n17707 ^ n9729 ;
  assign n17712 = ( n6686 & n13677 ) | ( n6686 & ~n15840 ) | ( n13677 & ~n15840 ) ;
  assign n17713 = n17695 ^ n6986 ^ n3569 ;
  assign n17714 = ( n1020 & n2841 ) | ( n1020 & n10007 ) | ( n2841 & n10007 ) ;
  assign n17715 = n17714 ^ n3781 ^ n1630 ;
  assign n17716 = ( n6339 & ~n7124 ) | ( n6339 & n7269 ) | ( ~n7124 & n7269 ) ;
  assign n17717 = n11222 ^ n7133 ^ n798 ;
  assign n17718 = ( n7133 & n17318 ) | ( n7133 & ~n17717 ) | ( n17318 & ~n17717 ) ;
  assign n17719 = ( ~n12119 & n17716 ) | ( ~n12119 & n17718 ) | ( n17716 & n17718 ) ;
  assign n17721 = n13486 ^ n6796 ^ n5419 ;
  assign n17722 = ( n467 & n7882 ) | ( n467 & n17721 ) | ( n7882 & n17721 ) ;
  assign n17720 = ( n8972 & ~n10738 ) | ( n8972 & n12511 ) | ( ~n10738 & n12511 ) ;
  assign n17723 = n17722 ^ n17720 ^ n5837 ;
  assign n17724 = n9300 ^ n6467 ^ n3268 ;
  assign n17725 = n17724 ^ n10754 ^ n1316 ;
  assign n17726 = n16519 ^ n2753 ^ n2080 ;
  assign n17727 = n10756 ^ n7156 ^ n5253 ;
  assign n17728 = n17727 ^ n17460 ^ n3587 ;
  assign n17729 = ( n321 & n5936 ) | ( n321 & n9220 ) | ( n5936 & n9220 ) ;
  assign n17730 = ( n4895 & ~n12961 ) | ( n4895 & n17729 ) | ( ~n12961 & n17729 ) ;
  assign n17731 = n14847 ^ n12098 ^ n3556 ;
  assign n17732 = ( n8082 & n10153 ) | ( n8082 & ~n17731 ) | ( n10153 & ~n17731 ) ;
  assign n17733 = ( n9623 & n17730 ) | ( n9623 & n17732 ) | ( n17730 & n17732 ) ;
  assign n17734 = ( n1967 & n4787 ) | ( n1967 & n13590 ) | ( n4787 & n13590 ) ;
  assign n17735 = n17734 ^ n9801 ^ n3555 ;
  assign n17736 = ( n1942 & n2393 ) | ( n1942 & ~n3235 ) | ( n2393 & ~n3235 ) ;
  assign n17737 = n17593 ^ n3045 ^ n2101 ;
  assign n17738 = n12119 ^ n11597 ^ n3385 ;
  assign n17739 = n17738 ^ n16333 ^ n5251 ;
  assign n17740 = ( n3438 & n6080 ) | ( n3438 & ~n11092 ) | ( n6080 & ~n11092 ) ;
  assign n17741 = n13531 ^ n8274 ^ x0 ;
  assign n17742 = ( n2048 & n17740 ) | ( n2048 & n17741 ) | ( n17740 & n17741 ) ;
  assign n17744 = n12766 ^ n6818 ^ n2890 ;
  assign n17743 = n17264 ^ n9108 ^ n5598 ;
  assign n17745 = n17744 ^ n17743 ^ n15888 ;
  assign n17746 = ( n1673 & ~n9441 ) | ( n1673 & n10007 ) | ( ~n9441 & n10007 ) ;
  assign n17747 = ( n1606 & n7254 ) | ( n1606 & ~n17746 ) | ( n7254 & ~n17746 ) ;
  assign n17748 = n17747 ^ n7731 ^ n1546 ;
  assign n17749 = n11758 ^ n1765 ^ n1230 ;
  assign n17750 = n17749 ^ n9052 ^ n2355 ;
  assign n17751 = ( ~n9704 & n13008 ) | ( ~n9704 & n17750 ) | ( n13008 & n17750 ) ;
  assign n17752 = n8434 ^ n2401 ^ n459 ;
  assign n17753 = n11672 ^ n6208 ^ n4097 ;
  assign n17754 = ( n3449 & ~n11359 ) | ( n3449 & n11994 ) | ( ~n11359 & n11994 ) ;
  assign n17755 = n17754 ^ n16650 ^ n8251 ;
  assign n17756 = n11882 ^ n9462 ^ n1019 ;
  assign n17757 = ( n7993 & ~n9740 ) | ( n7993 & n17756 ) | ( ~n9740 & n17756 ) ;
  assign n17758 = ( n6814 & n13897 ) | ( n6814 & n17757 ) | ( n13897 & n17757 ) ;
  assign n17759 = n17758 ^ n5299 ^ n439 ;
  assign n17760 = ( n11840 & n13904 ) | ( n11840 & ~n17759 ) | ( n13904 & ~n17759 ) ;
  assign n17761 = ( n1176 & ~n5460 ) | ( n1176 & n6201 ) | ( ~n5460 & n6201 ) ;
  assign n17762 = ( n6660 & ~n17290 ) | ( n6660 & n17761 ) | ( ~n17290 & n17761 ) ;
  assign n17763 = ( n6722 & n17537 ) | ( n6722 & ~n17762 ) | ( n17537 & ~n17762 ) ;
  assign n17764 = ( ~n1408 & n2536 ) | ( ~n1408 & n11393 ) | ( n2536 & n11393 ) ;
  assign n17765 = n17764 ^ n15582 ^ n5801 ;
  assign n17766 = ( ~n5670 & n9984 ) | ( ~n5670 & n17765 ) | ( n9984 & n17765 ) ;
  assign n17767 = n16187 ^ n14278 ^ n10412 ;
  assign n17768 = n17767 ^ n4153 ^ n398 ;
  assign n17769 = n7028 ^ n3516 ^ n1276 ;
  assign n17770 = n17769 ^ n8114 ^ n502 ;
  assign n17771 = n17770 ^ n16595 ^ n1827 ;
  assign n17772 = ( n5232 & ~n13572 ) | ( n5232 & n17771 ) | ( ~n13572 & n17771 ) ;
  assign n17773 = ( n1496 & n2683 ) | ( n1496 & ~n9230 ) | ( n2683 & ~n9230 ) ;
  assign n17774 = ( n2302 & n13687 ) | ( n2302 & ~n17773 ) | ( n13687 & ~n17773 ) ;
  assign n17782 = n11061 ^ n6952 ^ n940 ;
  assign n17779 = n13959 ^ n13402 ^ n9127 ;
  assign n17778 = ( n1022 & n3900 ) | ( n1022 & ~n6511 ) | ( n3900 & ~n6511 ) ;
  assign n17780 = n17779 ^ n17778 ^ n14211 ;
  assign n17781 = ( ~n5767 & n17137 ) | ( ~n5767 & n17780 ) | ( n17137 & n17780 ) ;
  assign n17775 = n4765 ^ n4533 ^ n441 ;
  assign n17776 = ( n2351 & n2875 ) | ( n2351 & ~n10148 ) | ( n2875 & ~n10148 ) ;
  assign n17777 = ( n14197 & n17775 ) | ( n14197 & n17776 ) | ( n17775 & n17776 ) ;
  assign n17783 = n17782 ^ n17781 ^ n17777 ;
  assign n17787 = ( ~n1901 & n3783 ) | ( ~n1901 & n8262 ) | ( n3783 & n8262 ) ;
  assign n17785 = n9301 ^ n3836 ^ n3437 ;
  assign n17784 = n7177 ^ n6964 ^ n5254 ;
  assign n17786 = n17785 ^ n17784 ^ n4221 ;
  assign n17788 = n17787 ^ n17786 ^ n16731 ;
  assign n17793 = n7685 ^ n6852 ^ n4953 ;
  assign n17794 = n17793 ^ n4061 ^ n1388 ;
  assign n17795 = ( n1843 & ~n10851 ) | ( n1843 & n15686 ) | ( ~n10851 & n15686 ) ;
  assign n17796 = ( n5884 & ~n17794 ) | ( n5884 & n17795 ) | ( ~n17794 & n17795 ) ;
  assign n17789 = n6117 ^ n5022 ^ n1156 ;
  assign n17790 = n17789 ^ n11351 ^ n4483 ;
  assign n17791 = n17790 ^ n17573 ^ n8935 ;
  assign n17792 = ( n1210 & ~n2999 ) | ( n1210 & n17791 ) | ( ~n2999 & n17791 ) ;
  assign n17797 = n17796 ^ n17792 ^ n8048 ;
  assign n17798 = ( n4477 & ~n16832 ) | ( n4477 & n17797 ) | ( ~n16832 & n17797 ) ;
  assign n17799 = ( n249 & n7355 ) | ( n249 & n8739 ) | ( n7355 & n8739 ) ;
  assign n17800 = ( n3155 & ~n4922 ) | ( n3155 & n8257 ) | ( ~n4922 & n8257 ) ;
  assign n17801 = n17800 ^ n8382 ^ n8019 ;
  assign n17802 = n5556 ^ n4530 ^ n3722 ;
  assign n17803 = ( n4555 & n13036 ) | ( n4555 & n17802 ) | ( n13036 & n17802 ) ;
  assign n17804 = n17803 ^ n6417 ^ n1671 ;
  assign n17805 = ( n17799 & n17801 ) | ( n17799 & n17804 ) | ( n17801 & n17804 ) ;
  assign n17806 = ( ~n9264 & n12810 ) | ( ~n9264 & n13324 ) | ( n12810 & n13324 ) ;
  assign n17808 = ( ~n3514 & n4007 ) | ( ~n3514 & n8298 ) | ( n4007 & n8298 ) ;
  assign n17807 = ( n2976 & n12873 ) | ( n2976 & n13246 ) | ( n12873 & n13246 ) ;
  assign n17809 = n17808 ^ n17807 ^ n10286 ;
  assign n17810 = ( n13091 & n13344 ) | ( n13091 & ~n17809 ) | ( n13344 & ~n17809 ) ;
  assign n17811 = ( n6829 & n10626 ) | ( n6829 & ~n12536 ) | ( n10626 & ~n12536 ) ;
  assign n17812 = ( ~n5259 & n7892 ) | ( ~n5259 & n16768 ) | ( n7892 & n16768 ) ;
  assign n17813 = n17812 ^ n741 ^ n355 ;
  assign n17814 = ( n15411 & n17811 ) | ( n15411 & ~n17813 ) | ( n17811 & ~n17813 ) ;
  assign n17815 = ( n997 & n1406 ) | ( n997 & ~n7861 ) | ( n1406 & ~n7861 ) ;
  assign n17816 = n17815 ^ n15978 ^ n14195 ;
  assign n17817 = n9908 ^ n8028 ^ n3163 ;
  assign n17818 = ( n253 & n2890 ) | ( n253 & ~n16637 ) | ( n2890 & ~n16637 ) ;
  assign n17819 = ( n823 & n7318 ) | ( n823 & n17818 ) | ( n7318 & n17818 ) ;
  assign n17820 = ( n12974 & n17817 ) | ( n12974 & ~n17819 ) | ( n17817 & ~n17819 ) ;
  assign n17821 = ( n10405 & n17816 ) | ( n10405 & ~n17820 ) | ( n17816 & ~n17820 ) ;
  assign n17822 = ( n12426 & n12429 ) | ( n12426 & ~n14619 ) | ( n12429 & ~n14619 ) ;
  assign n17823 = n17822 ^ n13391 ^ n4713 ;
  assign n17824 = ( ~x8 & n10782 ) | ( ~x8 & n17823 ) | ( n10782 & n17823 ) ;
  assign n17825 = ( n1686 & n3831 ) | ( n1686 & ~n3873 ) | ( n3831 & ~n3873 ) ;
  assign n17826 = n8788 ^ n3142 ^ n2033 ;
  assign n17827 = n4165 ^ n2025 ^ n852 ;
  assign n17832 = ( n10862 & ~n16229 ) | ( n10862 & n17409 ) | ( ~n16229 & n17409 ) ;
  assign n17830 = n7701 ^ n5563 ^ n4769 ;
  assign n17831 = n17830 ^ n9788 ^ n7263 ;
  assign n17828 = n13537 ^ n8774 ^ n5187 ;
  assign n17829 = n17828 ^ n17738 ^ n4430 ;
  assign n17833 = n17832 ^ n17831 ^ n17829 ;
  assign n17834 = ( n2022 & ~n17827 ) | ( n2022 & n17833 ) | ( ~n17827 & n17833 ) ;
  assign n17835 = n10550 ^ n1242 ^ n235 ;
  assign n17836 = ( n1047 & ~n6015 ) | ( n1047 & n17835 ) | ( ~n6015 & n17835 ) ;
  assign n17837 = n10648 ^ n9016 ^ n266 ;
  assign n17838 = n13654 ^ n10054 ^ n6183 ;
  assign n17839 = n17838 ^ n7132 ^ n5566 ;
  assign n17840 = ( n15883 & n16482 ) | ( n15883 & ~n17839 ) | ( n16482 & ~n17839 ) ;
  assign n17841 = ( ~n1039 & n5731 ) | ( ~n1039 & n8600 ) | ( n5731 & n8600 ) ;
  assign n17842 = n17841 ^ n17717 ^ n16844 ;
  assign n17843 = n17842 ^ n15516 ^ n7100 ;
  assign n17844 = n5800 ^ n5372 ^ n3332 ;
  assign n17845 = ( n1966 & n10146 ) | ( n1966 & n17844 ) | ( n10146 & n17844 ) ;
  assign n17846 = n13598 ^ n5104 ^ n256 ;
  assign n17847 = ( n7103 & n9873 ) | ( n7103 & n17846 ) | ( n9873 & n17846 ) ;
  assign n17848 = n7632 ^ n5106 ^ n3766 ;
  assign n17849 = ( n15406 & n17714 ) | ( n15406 & n17848 ) | ( n17714 & n17848 ) ;
  assign n17851 = n7402 ^ n5670 ^ n3333 ;
  assign n17850 = n7874 ^ n6994 ^ n2893 ;
  assign n17852 = n17851 ^ n17850 ^ n1026 ;
  assign n17853 = ( n1240 & n5631 ) | ( n1240 & ~n14639 ) | ( n5631 & ~n14639 ) ;
  assign n17854 = ( ~n11275 & n13871 ) | ( ~n11275 & n17853 ) | ( n13871 & n17853 ) ;
  assign n17855 = n15991 ^ n7108 ^ n166 ;
  assign n17856 = ( ~n4191 & n4637 ) | ( ~n4191 & n17855 ) | ( n4637 & n17855 ) ;
  assign n17857 = ( n8164 & n8300 ) | ( n8164 & n9054 ) | ( n8300 & n9054 ) ;
  assign n17858 = n17857 ^ n4038 ^ n213 ;
  assign n17861 = ( n3439 & ~n6004 ) | ( n3439 & n8177 ) | ( ~n6004 & n8177 ) ;
  assign n17859 = ( n2526 & ~n12267 ) | ( n2526 & n12678 ) | ( ~n12267 & n12678 ) ;
  assign n17860 = n17859 ^ n16600 ^ n5664 ;
  assign n17862 = n17861 ^ n17860 ^ n11616 ;
  assign n17863 = n13855 ^ n12376 ^ n3127 ;
  assign n17864 = n17863 ^ n17067 ^ n10685 ;
  assign n17865 = ( n423 & n662 ) | ( n423 & n3077 ) | ( n662 & n3077 ) ;
  assign n17866 = n15272 ^ n11890 ^ n8011 ;
  assign n17867 = ( n15580 & n17865 ) | ( n15580 & n17866 ) | ( n17865 & n17866 ) ;
  assign n17868 = n12482 ^ n5749 ^ n4804 ;
  assign n17869 = n7070 ^ n5946 ^ n1714 ;
  assign n17872 = n13745 ^ n7385 ^ n3597 ;
  assign n17870 = ( n1806 & ~n7416 ) | ( n1806 & n15359 ) | ( ~n7416 & n15359 ) ;
  assign n17871 = n17870 ^ n16706 ^ n2219 ;
  assign n17873 = n17872 ^ n17871 ^ n2955 ;
  assign n17874 = n12173 ^ n10244 ^ n9334 ;
  assign n17875 = n17874 ^ n11320 ^ n7056 ;
  assign n17876 = n10106 ^ n1734 ^ n456 ;
  assign n17877 = ( n5575 & ~n8539 ) | ( n5575 & n17876 ) | ( ~n8539 & n17876 ) ;
  assign n17878 = ( n13706 & ~n15388 ) | ( n13706 & n17877 ) | ( ~n15388 & n17877 ) ;
  assign n17879 = ( ~n3125 & n6114 ) | ( ~n3125 & n6990 ) | ( n6114 & n6990 ) ;
  assign n17880 = ( n891 & ~n7215 ) | ( n891 & n8227 ) | ( ~n7215 & n8227 ) ;
  assign n17881 = ( n7853 & n17879 ) | ( n7853 & ~n17880 ) | ( n17879 & ~n17880 ) ;
  assign n17883 = n8960 ^ n7700 ^ n2439 ;
  assign n17882 = ( n904 & ~n3763 ) | ( n904 & n12544 ) | ( ~n3763 & n12544 ) ;
  assign n17884 = n17883 ^ n17882 ^ n2050 ;
  assign n17885 = ( ~n131 & n1016 ) | ( ~n131 & n17884 ) | ( n1016 & n17884 ) ;
  assign n17887 = ( n3088 & n4948 ) | ( n3088 & n16736 ) | ( n4948 & n16736 ) ;
  assign n17886 = n16676 ^ n5501 ^ n1702 ;
  assign n17888 = n17887 ^ n17886 ^ n10501 ;
  assign n17889 = ( n13245 & ~n13253 ) | ( n13245 & n15139 ) | ( ~n13253 & n15139 ) ;
  assign n17890 = ( ~n700 & n5861 ) | ( ~n700 & n8481 ) | ( n5861 & n8481 ) ;
  assign n17891 = ( ~n4857 & n10740 ) | ( ~n4857 & n17890 ) | ( n10740 & n17890 ) ;
  assign n17892 = ( ~n6141 & n6199 ) | ( ~n6141 & n16599 ) | ( n6199 & n16599 ) ;
  assign n17893 = n17892 ^ n5154 ^ n621 ;
  assign n17894 = n16007 ^ n9044 ^ n8889 ;
  assign n17895 = ( n3353 & n3706 ) | ( n3353 & n17894 ) | ( n3706 & n17894 ) ;
  assign n17896 = n17895 ^ n11232 ^ n4428 ;
  assign n17897 = ( n4182 & n10133 ) | ( n4182 & n10204 ) | ( n10133 & n10204 ) ;
  assign n17898 = ( ~n5773 & n7489 ) | ( ~n5773 & n15336 ) | ( n7489 & n15336 ) ;
  assign n17899 = n17898 ^ n4024 ^ n653 ;
  assign n17900 = ( n17644 & n17897 ) | ( n17644 & n17899 ) | ( n17897 & n17899 ) ;
  assign n17901 = n13819 ^ n4538 ^ n2978 ;
  assign n17902 = n17901 ^ n11465 ^ n6291 ;
  assign n17903 = ( n310 & n6174 ) | ( n310 & ~n8248 ) | ( n6174 & ~n8248 ) ;
  assign n17904 = ( n3610 & n12002 ) | ( n3610 & n17903 ) | ( n12002 & n17903 ) ;
  assign n17905 = ( n9482 & n14495 ) | ( n9482 & ~n17539 ) | ( n14495 & ~n17539 ) ;
  assign n17906 = n9164 ^ n1173 ^ n631 ;
  assign n17907 = ( n882 & n7758 ) | ( n882 & ~n9725 ) | ( n7758 & ~n9725 ) ;
  assign n17908 = ( n12658 & n17906 ) | ( n12658 & n17907 ) | ( n17906 & n17907 ) ;
  assign n17909 = n14042 ^ n9591 ^ n7979 ;
  assign n17910 = ( n449 & n3820 ) | ( n449 & ~n17909 ) | ( n3820 & ~n17909 ) ;
  assign n17911 = ( n1901 & n8497 ) | ( n1901 & ~n10964 ) | ( n8497 & ~n10964 ) ;
  assign n17912 = ( ~n2563 & n3139 ) | ( ~n2563 & n17911 ) | ( n3139 & n17911 ) ;
  assign n17913 = ( n6705 & ~n12231 ) | ( n6705 & n17912 ) | ( ~n12231 & n17912 ) ;
  assign n17914 = n8538 ^ n6123 ^ n1003 ;
  assign n17915 = ( n4658 & ~n15405 ) | ( n4658 & n17914 ) | ( ~n15405 & n17914 ) ;
  assign n17916 = ( n1036 & ~n8178 ) | ( n1036 & n17915 ) | ( ~n8178 & n17915 ) ;
  assign n17917 = n17032 ^ n7759 ^ n4840 ;
  assign n17918 = n12513 ^ n9928 ^ n8513 ;
  assign n17919 = ( n8653 & n17299 ) | ( n8653 & n17918 ) | ( n17299 & n17918 ) ;
  assign n17920 = ( ~n1043 & n6215 ) | ( ~n1043 & n15655 ) | ( n6215 & n15655 ) ;
  assign n17921 = n17920 ^ n17428 ^ n4385 ;
  assign n17922 = ( ~n8405 & n9850 ) | ( ~n8405 & n17921 ) | ( n9850 & n17921 ) ;
  assign n17923 = n9937 ^ n9677 ^ n4212 ;
  assign n17924 = n17923 ^ n11339 ^ n3746 ;
  assign n17928 = ( ~n574 & n2577 ) | ( ~n574 & n14807 ) | ( n2577 & n14807 ) ;
  assign n17925 = n4253 ^ n3698 ^ n3276 ;
  assign n17926 = n11763 ^ n4029 ^ n968 ;
  assign n17927 = ( n250 & n17925 ) | ( n250 & n17926 ) | ( n17925 & n17926 ) ;
  assign n17929 = n17928 ^ n17927 ^ n17488 ;
  assign n17935 = ( x51 & n4515 ) | ( x51 & ~n6904 ) | ( n4515 & ~n6904 ) ;
  assign n17930 = n7714 ^ n4475 ^ n3510 ;
  assign n17931 = n10958 ^ n5064 ^ n4645 ;
  assign n17932 = ( n975 & ~n3555 ) | ( n975 & n9050 ) | ( ~n3555 & n9050 ) ;
  assign n17933 = ( ~n8227 & n16179 ) | ( ~n8227 & n17932 ) | ( n16179 & n17932 ) ;
  assign n17934 = ( n17930 & n17931 ) | ( n17930 & n17933 ) | ( n17931 & n17933 ) ;
  assign n17936 = n17935 ^ n17934 ^ n2124 ;
  assign n17937 = ( n2422 & n4368 ) | ( n2422 & ~n5824 ) | ( n4368 & ~n5824 ) ;
  assign n17938 = ( n2284 & ~n16206 ) | ( n2284 & n17937 ) | ( ~n16206 & n17937 ) ;
  assign n17939 = n11475 ^ n6411 ^ n2598 ;
  assign n17940 = n17939 ^ n10388 ^ x124 ;
  assign n17947 = ( n508 & n13116 ) | ( n508 & ~n14216 ) | ( n13116 & ~n14216 ) ;
  assign n17948 = ( n1475 & ~n17482 ) | ( n1475 & n17947 ) | ( ~n17482 & n17947 ) ;
  assign n17941 = n15839 ^ n13383 ^ n11148 ;
  assign n17942 = ( n1561 & n2584 ) | ( n1561 & ~n4443 ) | ( n2584 & ~n4443 ) ;
  assign n17943 = ( n6373 & n8425 ) | ( n6373 & ~n17942 ) | ( n8425 & ~n17942 ) ;
  assign n17944 = n17943 ^ n12683 ^ n8203 ;
  assign n17945 = n17792 ^ n13811 ^ n8089 ;
  assign n17946 = ( n17941 & n17944 ) | ( n17941 & ~n17945 ) | ( n17944 & ~n17945 ) ;
  assign n17949 = n17948 ^ n17946 ^ n16774 ;
  assign n17950 = n13039 ^ n8249 ^ n2911 ;
  assign n17951 = n17950 ^ n10083 ^ n2456 ;
  assign n17952 = n4478 ^ n3638 ^ n882 ;
  assign n17953 = ( n10208 & n17951 ) | ( n10208 & ~n17952 ) | ( n17951 & ~n17952 ) ;
  assign n17957 = ( ~n5994 & n6854 ) | ( ~n5994 & n8080 ) | ( n6854 & n8080 ) ;
  assign n17955 = ( n4184 & ~n4650 ) | ( n4184 & n8295 ) | ( ~n4650 & n8295 ) ;
  assign n17956 = n17955 ^ n4636 ^ n2201 ;
  assign n17958 = n17957 ^ n17956 ^ n5142 ;
  assign n17954 = n17767 ^ n2977 ^ n811 ;
  assign n17959 = n17958 ^ n17954 ^ n13150 ;
  assign n17960 = n17581 ^ n15736 ^ n9438 ;
  assign n17961 = ( ~n11376 & n13944 ) | ( ~n11376 & n17960 ) | ( n13944 & n17960 ) ;
  assign n17962 = n17961 ^ n15177 ^ n11042 ;
  assign n17964 = n13945 ^ n13550 ^ n2849 ;
  assign n17963 = ( n1295 & ~n12900 ) | ( n1295 & n17322 ) | ( ~n12900 & n17322 ) ;
  assign n17965 = n17964 ^ n17963 ^ n10068 ;
  assign n17966 = ( n4392 & n13548 ) | ( n4392 & n17965 ) | ( n13548 & n17965 ) ;
  assign n17967 = ( n7017 & n17962 ) | ( n7017 & ~n17966 ) | ( n17962 & ~n17966 ) ;
  assign n17968 = n13022 ^ n10473 ^ n5124 ;
  assign n17969 = ( n871 & n3971 ) | ( n871 & n7452 ) | ( n3971 & n7452 ) ;
  assign n17970 = ( n3257 & ~n9439 ) | ( n3257 & n17969 ) | ( ~n9439 & n17969 ) ;
  assign n17971 = ( n5763 & ~n15379 ) | ( n5763 & n17970 ) | ( ~n15379 & n17970 ) ;
  assign n17972 = ( n2996 & n17968 ) | ( n2996 & n17971 ) | ( n17968 & n17971 ) ;
  assign n17973 = n13735 ^ n3818 ^ n1362 ;
  assign n17974 = n17973 ^ n14154 ^ n8639 ;
  assign n17975 = n17974 ^ n16316 ^ n12277 ;
  assign n17976 = n16397 ^ n3766 ^ n1063 ;
  assign n17977 = n17976 ^ n14659 ^ n10497 ;
  assign n17979 = n10931 ^ n6287 ^ n3624 ;
  assign n17980 = n9125 ^ n1318 ^ n1279 ;
  assign n17981 = ( ~n192 & n17979 ) | ( ~n192 & n17980 ) | ( n17979 & n17980 ) ;
  assign n17982 = n17981 ^ n2051 ^ n1899 ;
  assign n17978 = ( ~n2516 & n13516 ) | ( ~n2516 & n16964 ) | ( n13516 & n16964 ) ;
  assign n17983 = n17982 ^ n17978 ^ n12477 ;
  assign n17984 = n17534 ^ n7264 ^ n3939 ;
  assign n17989 = ( ~n760 & n3351 ) | ( ~n760 & n9268 ) | ( n3351 & n9268 ) ;
  assign n17990 = n15433 ^ n14737 ^ n2602 ;
  assign n17991 = ( n7308 & ~n17989 ) | ( n7308 & n17990 ) | ( ~n17989 & n17990 ) ;
  assign n17985 = n6408 ^ n6304 ^ n1740 ;
  assign n17986 = n17985 ^ n10206 ^ n4432 ;
  assign n17987 = ( n7325 & n11106 ) | ( n7325 & n17986 ) | ( n11106 & n17986 ) ;
  assign n17988 = n17987 ^ n10724 ^ n9266 ;
  assign n17992 = n17991 ^ n17988 ^ n3963 ;
  assign n17993 = n2692 ^ n2395 ^ n742 ;
  assign n17994 = ( n7310 & ~n8205 ) | ( n7310 & n17993 ) | ( ~n8205 & n17993 ) ;
  assign n17995 = n17994 ^ n17614 ^ n1694 ;
  assign n17996 = ( x68 & ~n2320 ) | ( x68 & n8854 ) | ( ~n2320 & n8854 ) ;
  assign n17997 = n17996 ^ n10313 ^ n5211 ;
  assign n18000 = n7363 ^ n179 ^ x57 ;
  assign n17999 = n13175 ^ n11110 ^ n7631 ;
  assign n17998 = n13817 ^ n11701 ^ n10719 ;
  assign n18001 = n18000 ^ n17999 ^ n17998 ;
  assign n18002 = ( n4407 & n7899 ) | ( n4407 & n10583 ) | ( n7899 & n10583 ) ;
  assign n18003 = n18002 ^ n15026 ^ n10739 ;
  assign n18004 = n4152 ^ n3876 ^ n2749 ;
  assign n18005 = n16229 ^ n8483 ^ n6446 ;
  assign n18006 = n18005 ^ n8269 ^ n6246 ;
  assign n18007 = ( n297 & n13838 ) | ( n297 & n18006 ) | ( n13838 & n18006 ) ;
  assign n18008 = ( x105 & ~n18004 ) | ( x105 & n18007 ) | ( ~n18004 & n18007 ) ;
  assign n18009 = ( n1526 & n7630 ) | ( n1526 & n12024 ) | ( n7630 & n12024 ) ;
  assign n18011 = n16665 ^ n9196 ^ n4254 ;
  assign n18010 = ( n2850 & ~n10328 ) | ( n2850 & n12134 ) | ( ~n10328 & n12134 ) ;
  assign n18012 = n18011 ^ n18010 ^ n16632 ;
  assign n18013 = ( ~n16710 & n16917 ) | ( ~n16710 & n18012 ) | ( n16917 & n18012 ) ;
  assign n18014 = n13506 ^ n9929 ^ n1536 ;
  assign n18015 = ( n6012 & n12303 ) | ( n6012 & ~n18014 ) | ( n12303 & ~n18014 ) ;
  assign n18016 = n12422 ^ n7658 ^ n4481 ;
  assign n18017 = ( n7212 & ~n12797 ) | ( n7212 & n18016 ) | ( ~n12797 & n18016 ) ;
  assign n18018 = n18017 ^ n15849 ^ n4515 ;
  assign n18019 = ( n1472 & n5973 ) | ( n1472 & ~n11763 ) | ( n5973 & ~n11763 ) ;
  assign n18020 = ( ~n8500 & n14886 ) | ( ~n8500 & n18019 ) | ( n14886 & n18019 ) ;
  assign n18021 = ( n17792 & n18018 ) | ( n17792 & n18020 ) | ( n18018 & n18020 ) ;
  assign n18022 = n18021 ^ n16109 ^ n1498 ;
  assign n18024 = ( n1288 & ~n5383 ) | ( n1288 & n15974 ) | ( ~n5383 & n15974 ) ;
  assign n18023 = ( x112 & ~n6659 ) | ( x112 & n7925 ) | ( ~n6659 & n7925 ) ;
  assign n18025 = n18024 ^ n18023 ^ n17456 ;
  assign n18026 = ( ~n5732 & n7867 ) | ( ~n5732 & n8509 ) | ( n7867 & n8509 ) ;
  assign n18027 = n18026 ^ n15230 ^ n6357 ;
  assign n18028 = ( n4084 & ~n7513 ) | ( n4084 & n13991 ) | ( ~n7513 & n13991 ) ;
  assign n18032 = n13781 ^ n7923 ^ n3293 ;
  assign n18029 = ( n854 & ~n6366 ) | ( n854 & n15040 ) | ( ~n6366 & n15040 ) ;
  assign n18030 = ( ~n4211 & n8767 ) | ( ~n4211 & n18029 ) | ( n8767 & n18029 ) ;
  assign n18031 = n18030 ^ n13938 ^ n6871 ;
  assign n18033 = n18032 ^ n18031 ^ n11904 ;
  assign n18034 = ( n3554 & n4221 ) | ( n3554 & n8032 ) | ( n4221 & n8032 ) ;
  assign n18035 = ( ~n3679 & n5874 ) | ( ~n3679 & n18034 ) | ( n5874 & n18034 ) ;
  assign n18036 = ( ~n3160 & n5491 ) | ( ~n3160 & n9958 ) | ( n5491 & n9958 ) ;
  assign n18037 = ( n1699 & n2617 ) | ( n1699 & n18036 ) | ( n2617 & n18036 ) ;
  assign n18038 = ( n218 & n1858 ) | ( n218 & n3509 ) | ( n1858 & n3509 ) ;
  assign n18039 = ( n8904 & n18037 ) | ( n8904 & n18038 ) | ( n18037 & n18038 ) ;
  assign n18040 = n14561 ^ n4569 ^ n656 ;
  assign n18041 = ( n2012 & ~n5274 ) | ( n2012 & n18040 ) | ( ~n5274 & n18040 ) ;
  assign n18042 = ( n11881 & n13484 ) | ( n11881 & n18041 ) | ( n13484 & n18041 ) ;
  assign n18043 = n4149 ^ n3790 ^ n1487 ;
  assign n18044 = n18043 ^ n12823 ^ n11189 ;
  assign n18045 = n16280 ^ n10405 ^ n1536 ;
  assign n18049 = n13595 ^ n9542 ^ n6635 ;
  assign n18050 = ( n9974 & ~n13004 ) | ( n9974 & n18049 ) | ( ~n13004 & n18049 ) ;
  assign n18046 = n8154 ^ n6499 ^ n1679 ;
  assign n18047 = n4816 ^ n2111 ^ n547 ;
  assign n18048 = ( n5768 & n18046 ) | ( n5768 & ~n18047 ) | ( n18046 & ~n18047 ) ;
  assign n18051 = n18050 ^ n18048 ^ n7068 ;
  assign n18056 = n14873 ^ n5392 ^ n4726 ;
  assign n18052 = n8773 ^ n8320 ^ n1303 ;
  assign n18053 = ( n1009 & ~n3434 ) | ( n1009 & n12966 ) | ( ~n3434 & n12966 ) ;
  assign n18054 = ( n7511 & n18052 ) | ( n7511 & n18053 ) | ( n18052 & n18053 ) ;
  assign n18055 = ( n3354 & ~n5097 ) | ( n3354 & n18054 ) | ( ~n5097 & n18054 ) ;
  assign n18057 = n18056 ^ n18055 ^ n13580 ;
  assign n18058 = n9496 ^ n8331 ^ n2083 ;
  assign n18059 = n9658 ^ n9009 ^ n4905 ;
  assign n18060 = n18059 ^ n12672 ^ n1316 ;
  assign n18061 = ( ~n7403 & n18058 ) | ( ~n7403 & n18060 ) | ( n18058 & n18060 ) ;
  assign n18062 = n13807 ^ n7689 ^ n6926 ;
  assign n18063 = ( n1651 & ~n18061 ) | ( n1651 & n18062 ) | ( ~n18061 & n18062 ) ;
  assign n18064 = n11443 ^ n10003 ^ n5623 ;
  assign n18065 = ( n1083 & ~n11610 ) | ( n1083 & n18064 ) | ( ~n11610 & n18064 ) ;
  assign n18066 = n14911 ^ n2691 ^ n385 ;
  assign n18067 = n18066 ^ n13021 ^ n7262 ;
  assign n18068 = n18067 ^ n7849 ^ n1683 ;
  assign n18069 = ( n3650 & ~n5046 ) | ( n3650 & n6181 ) | ( ~n5046 & n6181 ) ;
  assign n18070 = n18069 ^ n6894 ^ n3689 ;
  assign n18071 = ( ~n2150 & n14819 ) | ( ~n2150 & n18070 ) | ( n14819 & n18070 ) ;
  assign n18073 = n5766 ^ n1007 ^ n736 ;
  assign n18072 = ( n794 & ~n1576 ) | ( n794 & n4775 ) | ( ~n1576 & n4775 ) ;
  assign n18074 = n18073 ^ n18072 ^ n5119 ;
  assign n18075 = n18074 ^ n6437 ^ n1378 ;
  assign n18076 = ( n1985 & n6873 ) | ( n1985 & ~n18075 ) | ( n6873 & ~n18075 ) ;
  assign n18077 = ( ~n9684 & n11129 ) | ( ~n9684 & n11338 ) | ( n11129 & n11338 ) ;
  assign n18078 = ( ~x30 & n2918 ) | ( ~x30 & n7729 ) | ( n2918 & n7729 ) ;
  assign n18079 = ( n1001 & n2644 ) | ( n1001 & n5803 ) | ( n2644 & n5803 ) ;
  assign n18082 = n10874 ^ n2886 ^ n993 ;
  assign n18080 = ( n2247 & n2579 ) | ( n2247 & n4760 ) | ( n2579 & n4760 ) ;
  assign n18081 = ( n2876 & n4716 ) | ( n2876 & n18080 ) | ( n4716 & n18080 ) ;
  assign n18083 = n18082 ^ n18081 ^ n11426 ;
  assign n18084 = n12146 ^ n3295 ^ n3050 ;
  assign n18085 = ( n1359 & n2964 ) | ( n1359 & n18084 ) | ( n2964 & n18084 ) ;
  assign n18086 = ( ~n3968 & n18083 ) | ( ~n3968 & n18085 ) | ( n18083 & n18085 ) ;
  assign n18087 = n18086 ^ n14244 ^ n11681 ;
  assign n18088 = ( n2793 & n18079 ) | ( n2793 & n18087 ) | ( n18079 & n18087 ) ;
  assign n18089 = n15188 ^ n14094 ^ n1491 ;
  assign n18090 = ( ~n2313 & n3258 ) | ( ~n2313 & n4123 ) | ( n3258 & n4123 ) ;
  assign n18091 = ( n12420 & n13722 ) | ( n12420 & ~n18090 ) | ( n13722 & ~n18090 ) ;
  assign n18092 = ( n3488 & n9754 ) | ( n3488 & ~n17452 ) | ( n9754 & ~n17452 ) ;
  assign n18093 = ( n3801 & ~n7704 ) | ( n3801 & n15521 ) | ( ~n7704 & n15521 ) ;
  assign n18094 = ( ~n8060 & n9610 ) | ( ~n8060 & n9683 ) | ( n9610 & n9683 ) ;
  assign n18095 = n12889 ^ n4010 ^ n1396 ;
  assign n18096 = n18095 ^ n5504 ^ n1947 ;
  assign n18097 = ( n11186 & ~n11273 ) | ( n11186 & n18096 ) | ( ~n11273 & n18096 ) ;
  assign n18098 = ( n16606 & n18094 ) | ( n16606 & ~n18097 ) | ( n18094 & ~n18097 ) ;
  assign n18101 = n11648 ^ n5407 ^ n3514 ;
  assign n18099 = n16473 ^ n12904 ^ n7756 ;
  assign n18100 = ( n11974 & ~n14507 ) | ( n11974 & n18099 ) | ( ~n14507 & n18099 ) ;
  assign n18102 = n18101 ^ n18100 ^ n16041 ;
  assign n18103 = ( n1677 & n5600 ) | ( n1677 & ~n14595 ) | ( n5600 & ~n14595 ) ;
  assign n18104 = n18103 ^ n9885 ^ n7951 ;
  assign n18105 = ( n6443 & n6672 ) | ( n6443 & ~n10043 ) | ( n6672 & ~n10043 ) ;
  assign n18106 = n17633 ^ n15095 ^ n9408 ;
  assign n18107 = ( n12136 & n18105 ) | ( n12136 & ~n18106 ) | ( n18105 & ~n18106 ) ;
  assign n18112 = ( n3938 & ~n13706 ) | ( n3938 & n17256 ) | ( ~n13706 & n17256 ) ;
  assign n18113 = n18112 ^ n10171 ^ n8877 ;
  assign n18110 = n17368 ^ n12899 ^ n8170 ;
  assign n18111 = ( n12752 & ~n16149 ) | ( n12752 & n18110 ) | ( ~n16149 & n18110 ) ;
  assign n18114 = n18113 ^ n18111 ^ n9851 ;
  assign n18108 = ( n1661 & n4423 ) | ( n1661 & ~n17401 ) | ( n4423 & ~n17401 ) ;
  assign n18109 = n18108 ^ n13681 ^ n2820 ;
  assign n18115 = n18114 ^ n18109 ^ n15575 ;
  assign n18116 = ( n2022 & n6482 ) | ( n2022 & n10031 ) | ( n6482 & n10031 ) ;
  assign n18117 = n18116 ^ n5039 ^ n1798 ;
  assign n18118 = ( n4334 & n12019 ) | ( n4334 & ~n18117 ) | ( n12019 & ~n18117 ) ;
  assign n18119 = n18118 ^ n15147 ^ n13288 ;
  assign n18121 = ( n4845 & n10351 ) | ( n4845 & n11346 ) | ( n10351 & n11346 ) ;
  assign n18122 = ( n2772 & n10418 ) | ( n2772 & ~n18121 ) | ( n10418 & ~n18121 ) ;
  assign n18120 = ( n597 & n2619 ) | ( n597 & ~n12492 ) | ( n2619 & ~n12492 ) ;
  assign n18123 = n18122 ^ n18120 ^ n17494 ;
  assign n18124 = ( n14475 & ~n15293 ) | ( n14475 & n18123 ) | ( ~n15293 & n18123 ) ;
  assign n18125 = n17585 ^ n8585 ^ n7338 ;
  assign n18126 = ( ~n2244 & n16886 ) | ( ~n2244 & n18125 ) | ( n16886 & n18125 ) ;
  assign n18127 = n10557 ^ n4542 ^ n3981 ;
  assign n18128 = n18127 ^ n5084 ^ x0 ;
  assign n18129 = ( ~n683 & n1270 ) | ( ~n683 & n18128 ) | ( n1270 & n18128 ) ;
  assign n18130 = n17022 ^ n3509 ^ x46 ;
  assign n18136 = ( n3081 & n4097 ) | ( n3081 & n5205 ) | ( n4097 & n5205 ) ;
  assign n18131 = ( n277 & ~n12790 ) | ( n277 & n16064 ) | ( ~n12790 & n16064 ) ;
  assign n18132 = n5342 ^ n2870 ^ n1573 ;
  assign n18133 = n18132 ^ n6850 ^ n2759 ;
  assign n18134 = n16194 ^ n11945 ^ n11094 ;
  assign n18135 = ( n18131 & n18133 ) | ( n18131 & ~n18134 ) | ( n18133 & ~n18134 ) ;
  assign n18137 = n18136 ^ n18135 ^ n7455 ;
  assign n18138 = ( n4571 & n5064 ) | ( n4571 & ~n9790 ) | ( n5064 & ~n9790 ) ;
  assign n18139 = n18138 ^ n10417 ^ n4672 ;
  assign n18140 = ( ~n6386 & n11240 ) | ( ~n6386 & n17335 ) | ( n11240 & n17335 ) ;
  assign n18141 = n18140 ^ n9336 ^ n2581 ;
  assign n18142 = ( n7383 & n18139 ) | ( n7383 & ~n18141 ) | ( n18139 & ~n18141 ) ;
  assign n18143 = n18142 ^ n8162 ^ n5305 ;
  assign n18144 = n6313 ^ n3383 ^ n2419 ;
  assign n18145 = ( n7312 & n14941 ) | ( n7312 & n18144 ) | ( n14941 & n18144 ) ;
  assign n18146 = n18145 ^ n16085 ^ n2368 ;
  assign n18147 = ( n1809 & ~n6620 ) | ( n1809 & n18146 ) | ( ~n6620 & n18146 ) ;
  assign n18148 = ( n866 & n4092 ) | ( n866 & n4443 ) | ( n4092 & n4443 ) ;
  assign n18149 = n12293 ^ n11475 ^ n2794 ;
  assign n18152 = n9343 ^ n5451 ^ n2319 ;
  assign n18153 = ( n4692 & n7923 ) | ( n4692 & n18152 ) | ( n7923 & n18152 ) ;
  assign n18150 = n13292 ^ n8559 ^ n5978 ;
  assign n18151 = n18150 ^ n1359 ^ n810 ;
  assign n18154 = n18153 ^ n18151 ^ n779 ;
  assign n18155 = ( ~n18148 & n18149 ) | ( ~n18148 & n18154 ) | ( n18149 & n18154 ) ;
  assign n18156 = ( n675 & n9567 ) | ( n675 & ~n10298 ) | ( n9567 & ~n10298 ) ;
  assign n18157 = ( n1632 & ~n3225 ) | ( n1632 & n8849 ) | ( ~n3225 & n8849 ) ;
  assign n18158 = n18157 ^ n11819 ^ n11338 ;
  assign n18159 = n14343 ^ n8166 ^ n3190 ;
  assign n18160 = n18159 ^ n2596 ^ n2410 ;
  assign n18161 = n4800 ^ n3644 ^ n3078 ;
  assign n18162 = ( n5166 & n8753 ) | ( n5166 & ~n18161 ) | ( n8753 & ~n18161 ) ;
  assign n18163 = ( n13419 & n18160 ) | ( n13419 & n18162 ) | ( n18160 & n18162 ) ;
  assign n18164 = n18163 ^ n11168 ^ n986 ;
  assign n18167 = n8262 ^ n3223 ^ n1848 ;
  assign n18165 = n18090 ^ n17462 ^ n5709 ;
  assign n18166 = ( ~n2364 & n17056 ) | ( ~n2364 & n18165 ) | ( n17056 & n18165 ) ;
  assign n18168 = n18167 ^ n18166 ^ n9153 ;
  assign n18169 = n18168 ^ n13975 ^ n13387 ;
  assign n18170 = n2722 ^ n1428 ^ n477 ;
  assign n18171 = n18170 ^ n16187 ^ n11520 ;
  assign n18172 = ( n1740 & ~n15260 ) | ( n1740 & n18171 ) | ( ~n15260 & n18171 ) ;
  assign n18173 = ( ~x116 & n3661 ) | ( ~x116 & n7463 ) | ( n3661 & n7463 ) ;
  assign n18174 = ( n2242 & ~n11017 ) | ( n2242 & n18173 ) | ( ~n11017 & n18173 ) ;
  assign n18175 = n15459 ^ n13758 ^ n8260 ;
  assign n18176 = ( ~n871 & n5196 ) | ( ~n871 & n8759 ) | ( n5196 & n8759 ) ;
  assign n18178 = n13720 ^ n6515 ^ n988 ;
  assign n18177 = ( n1631 & n4994 ) | ( n1631 & n14356 ) | ( n4994 & n14356 ) ;
  assign n18179 = n18178 ^ n18177 ^ n16459 ;
  assign n18180 = ( n13864 & ~n16205 ) | ( n13864 & n16303 ) | ( ~n16205 & n16303 ) ;
  assign n18181 = ( n1489 & n1517 ) | ( n1489 & ~n18180 ) | ( n1517 & ~n18180 ) ;
  assign n18182 = n18181 ^ n13900 ^ n2718 ;
  assign n18183 = ( n3873 & n4259 ) | ( n3873 & ~n12829 ) | ( n4259 & ~n12829 ) ;
  assign n18184 = ( n2670 & ~n3785 ) | ( n2670 & n18183 ) | ( ~n3785 & n18183 ) ;
  assign n18185 = ( n528 & ~n10072 ) | ( n528 & n17244 ) | ( ~n10072 & n17244 ) ;
  assign n18186 = ( n3320 & ~n10370 ) | ( n3320 & n18185 ) | ( ~n10370 & n18185 ) ;
  assign n18187 = n11000 ^ n2384 ^ n1094 ;
  assign n18188 = ( n1209 & ~n1288 ) | ( n1209 & n18187 ) | ( ~n1288 & n18187 ) ;
  assign n18189 = n17374 ^ n14852 ^ n5110 ;
  assign n18190 = n18189 ^ n17536 ^ n12610 ;
  assign n18191 = n15751 ^ n4071 ^ n418 ;
  assign n18192 = ( n2529 & n5918 ) | ( n2529 & ~n18191 ) | ( n5918 & ~n18191 ) ;
  assign n18193 = ( n4184 & n4778 ) | ( n4184 & ~n18192 ) | ( n4778 & ~n18192 ) ;
  assign n18194 = n18193 ^ n14306 ^ n5153 ;
  assign n18198 = n14656 ^ n6277 ^ n465 ;
  assign n18196 = ( n4914 & n7215 ) | ( n4914 & ~n13338 ) | ( n7215 & ~n13338 ) ;
  assign n18195 = ( ~n316 & n8493 ) | ( ~n316 & n17882 ) | ( n8493 & n17882 ) ;
  assign n18197 = n18196 ^ n18195 ^ n8773 ;
  assign n18199 = n18198 ^ n18197 ^ n13479 ;
  assign n18200 = ( n5221 & ~n8569 ) | ( n5221 & n9134 ) | ( ~n8569 & n9134 ) ;
  assign n18201 = n16175 ^ n9562 ^ n7638 ;
  assign n18202 = n17361 ^ n16977 ^ n3747 ;
  assign n18203 = ( ~n8200 & n18201 ) | ( ~n8200 & n18202 ) | ( n18201 & n18202 ) ;
  assign n18204 = ( ~n2687 & n5818 ) | ( ~n2687 & n9701 ) | ( n5818 & n9701 ) ;
  assign n18205 = ( n6319 & n12394 ) | ( n6319 & ~n18058 ) | ( n12394 & ~n18058 ) ;
  assign n18206 = n18205 ^ n18100 ^ n13893 ;
  assign n18207 = ( n3076 & n11964 ) | ( n3076 & ~n16002 ) | ( n11964 & ~n16002 ) ;
  assign n18208 = ( n1955 & n2914 ) | ( n1955 & ~n3306 ) | ( n2914 & ~n3306 ) ;
  assign n18209 = ( n5387 & ~n9501 ) | ( n5387 & n18208 ) | ( ~n9501 & n18208 ) ;
  assign n18210 = ( n9256 & n9530 ) | ( n9256 & n18209 ) | ( n9530 & n18209 ) ;
  assign n18211 = ( n3047 & ~n7818 ) | ( n3047 & n10969 ) | ( ~n7818 & n10969 ) ;
  assign n18212 = ( n15156 & n18210 ) | ( n15156 & n18211 ) | ( n18210 & n18211 ) ;
  assign n18213 = ( n786 & n9628 ) | ( n786 & ~n18212 ) | ( n9628 & ~n18212 ) ;
  assign n18214 = ( n15441 & n17683 ) | ( n15441 & ~n18157 ) | ( n17683 & ~n18157 ) ;
  assign n18215 = n17839 ^ n9462 ^ n7689 ;
  assign n18216 = n18215 ^ n12284 ^ n7573 ;
  assign n18217 = ( ~n7835 & n10276 ) | ( ~n7835 & n13501 ) | ( n10276 & n13501 ) ;
  assign n18218 = ( n7072 & ~n7522 ) | ( n7072 & n18217 ) | ( ~n7522 & n18217 ) ;
  assign n18222 = n14570 ^ n9649 ^ n1024 ;
  assign n18221 = ( n2057 & ~n3790 ) | ( n2057 & n10283 ) | ( ~n3790 & n10283 ) ;
  assign n18219 = ( ~n1285 & n4312 ) | ( ~n1285 & n7310 ) | ( n4312 & n7310 ) ;
  assign n18220 = n18219 ^ n10559 ^ n918 ;
  assign n18223 = n18222 ^ n18221 ^ n18220 ;
  assign n18224 = n15742 ^ n15141 ^ n1792 ;
  assign n18225 = n18224 ^ n15609 ^ n3881 ;
  assign n18226 = ( n4024 & n6855 ) | ( n4024 & n8934 ) | ( n6855 & n8934 ) ;
  assign n18227 = n10956 ^ n783 ^ n588 ;
  assign n18228 = ( n1062 & ~n1571 ) | ( n1062 & n18227 ) | ( ~n1571 & n18227 ) ;
  assign n18229 = ( ~n8115 & n18226 ) | ( ~n8115 & n18228 ) | ( n18226 & n18228 ) ;
  assign n18235 = n8146 ^ n7840 ^ n4614 ;
  assign n18234 = ( n2230 & n5399 ) | ( n2230 & ~n6937 ) | ( n5399 & ~n6937 ) ;
  assign n18236 = n18235 ^ n18234 ^ n10466 ;
  assign n18232 = ( n6268 & ~n16323 ) | ( n6268 & n18219 ) | ( ~n16323 & n18219 ) ;
  assign n18233 = ( n10528 & n17146 ) | ( n10528 & ~n18232 ) | ( n17146 & ~n18232 ) ;
  assign n18230 = n6057 ^ n745 ^ n266 ;
  assign n18231 = n18230 ^ n13284 ^ n6448 ;
  assign n18237 = n18236 ^ n18233 ^ n18231 ;
  assign n18238 = ( n17525 & n18229 ) | ( n17525 & ~n18237 ) | ( n18229 & ~n18237 ) ;
  assign n18239 = n13048 ^ n9656 ^ n6299 ;
  assign n18240 = ( ~n296 & n2061 ) | ( ~n296 & n18239 ) | ( n2061 & n18239 ) ;
  assign n18241 = n10545 ^ n3071 ^ x93 ;
  assign n18242 = ( ~n694 & n9418 ) | ( ~n694 & n11281 ) | ( n9418 & n11281 ) ;
  assign n18243 = n18242 ^ n10474 ^ n5915 ;
  assign n18244 = n16358 ^ n8839 ^ n413 ;
  assign n18245 = n18244 ^ n8781 ^ n5053 ;
  assign n18246 = n16814 ^ n2409 ^ n1062 ;
  assign n18247 = n6344 ^ n3971 ^ n2797 ;
  assign n18248 = ( n1598 & n1613 ) | ( n1598 & ~n18247 ) | ( n1613 & ~n18247 ) ;
  assign n18249 = ( n7499 & ~n11763 ) | ( n7499 & n11778 ) | ( ~n11763 & n11778 ) ;
  assign n18250 = ( n6260 & n9073 ) | ( n6260 & n18249 ) | ( n9073 & n18249 ) ;
  assign n18251 = ( n7295 & n13710 ) | ( n7295 & ~n16721 ) | ( n13710 & ~n16721 ) ;
  assign n18252 = ( n6213 & n6769 ) | ( n6213 & n11679 ) | ( n6769 & n11679 ) ;
  assign n18253 = ( n9637 & n13483 ) | ( n9637 & ~n18252 ) | ( n13483 & ~n18252 ) ;
  assign n18254 = ( n18250 & n18251 ) | ( n18250 & n18253 ) | ( n18251 & n18253 ) ;
  assign n18255 = ( n3089 & n15655 ) | ( n3089 & ~n16481 ) | ( n15655 & ~n16481 ) ;
  assign n18256 = n15020 ^ n9892 ^ n7980 ;
  assign n18257 = n18256 ^ n12195 ^ n5160 ;
  assign n18258 = ( n1170 & n5963 ) | ( n1170 & n13232 ) | ( n5963 & n13232 ) ;
  assign n18259 = n18258 ^ n1452 ^ n622 ;
  assign n18260 = ( n3778 & ~n4679 ) | ( n3778 & n6351 ) | ( ~n4679 & n6351 ) ;
  assign n18261 = n18260 ^ n17434 ^ n15754 ;
  assign n18265 = n9051 ^ n7124 ^ n1704 ;
  assign n18263 = ( n1238 & n3280 ) | ( n1238 & n5887 ) | ( n3280 & n5887 ) ;
  assign n18262 = ( ~n3851 & n9601 ) | ( ~n3851 & n11172 ) | ( n9601 & n11172 ) ;
  assign n18264 = n18263 ^ n18262 ^ n11380 ;
  assign n18266 = n18265 ^ n18264 ^ n7972 ;
  assign n18275 = ( ~n278 & n585 ) | ( ~n278 & n9354 ) | ( n585 & n9354 ) ;
  assign n18273 = ( n1611 & n2518 ) | ( n1611 & ~n10813 ) | ( n2518 & ~n10813 ) ;
  assign n18274 = ( n7159 & n16356 ) | ( n7159 & ~n18273 ) | ( n16356 & ~n18273 ) ;
  assign n18276 = n18275 ^ n18274 ^ n3683 ;
  assign n18267 = ( n1944 & ~n5077 ) | ( n1944 & n10539 ) | ( ~n5077 & n10539 ) ;
  assign n18268 = n17621 ^ n12065 ^ n10927 ;
  assign n18269 = ( n8886 & n18267 ) | ( n8886 & n18268 ) | ( n18267 & n18268 ) ;
  assign n18270 = ( n701 & n8044 ) | ( n701 & ~n18269 ) | ( n8044 & ~n18269 ) ;
  assign n18271 = n18270 ^ n12962 ^ n7480 ;
  assign n18272 = ( ~n7137 & n9924 ) | ( ~n7137 & n18271 ) | ( n9924 & n18271 ) ;
  assign n18277 = n18276 ^ n18272 ^ n8675 ;
  assign n18278 = ( ~n1453 & n3878 ) | ( ~n1453 & n9162 ) | ( n3878 & n9162 ) ;
  assign n18279 = ( n1698 & n6448 ) | ( n1698 & ~n11029 ) | ( n6448 & ~n11029 ) ;
  assign n18280 = n17352 ^ n5182 ^ n908 ;
  assign n18281 = n9581 ^ n7329 ^ n1400 ;
  assign n18282 = ( ~n1524 & n3290 ) | ( ~n1524 & n18281 ) | ( n3290 & n18281 ) ;
  assign n18283 = n14276 ^ n9066 ^ n7175 ;
  assign n18284 = ( ~n9811 & n14094 ) | ( ~n9811 & n18283 ) | ( n14094 & n18283 ) ;
  assign n18285 = ( ~n3381 & n5001 ) | ( ~n3381 & n6250 ) | ( n5001 & n6250 ) ;
  assign n18286 = ( n2435 & n2932 ) | ( n2435 & n6891 ) | ( n2932 & n6891 ) ;
  assign n18287 = ( n1673 & n18285 ) | ( n1673 & ~n18286 ) | ( n18285 & ~n18286 ) ;
  assign n18293 = n13212 ^ n8065 ^ n3202 ;
  assign n18292 = n13087 ^ n11714 ^ n8027 ;
  assign n18288 = n12958 ^ n4718 ^ n2813 ;
  assign n18289 = ( x103 & n17494 ) | ( x103 & n18288 ) | ( n17494 & n18288 ) ;
  assign n18290 = ( ~n662 & n11903 ) | ( ~n662 & n18289 ) | ( n11903 & n18289 ) ;
  assign n18291 = n18290 ^ n5647 ^ n4328 ;
  assign n18294 = n18293 ^ n18292 ^ n18291 ;
  assign n18295 = n17717 ^ n16323 ^ n11567 ;
  assign n18296 = n18295 ^ n4326 ^ n1473 ;
  assign n18297 = ( n6130 & n8293 ) | ( n6130 & ~n15619 ) | ( n8293 & ~n15619 ) ;
  assign n18302 = n11513 ^ n10304 ^ n914 ;
  assign n18303 = n18302 ^ n2606 ^ n2541 ;
  assign n18298 = n14825 ^ n7334 ^ n2717 ;
  assign n18299 = ( ~n4640 & n9548 ) | ( ~n4640 & n10489 ) | ( n9548 & n10489 ) ;
  assign n18300 = ( n9690 & n18298 ) | ( n9690 & n18299 ) | ( n18298 & n18299 ) ;
  assign n18301 = n18300 ^ n16409 ^ n2873 ;
  assign n18304 = n18303 ^ n18301 ^ n16346 ;
  assign n18305 = ( ~n3406 & n17294 ) | ( ~n3406 & n17434 ) | ( n17294 & n17434 ) ;
  assign n18308 = n16711 ^ n11990 ^ n8617 ;
  assign n18306 = n17818 ^ n4589 ^ n2958 ;
  assign n18307 = n18306 ^ n13476 ^ n11021 ;
  assign n18309 = n18308 ^ n18307 ^ n14792 ;
  assign n18310 = n18309 ^ n16572 ^ n11262 ;
  assign n18311 = n8842 ^ n2316 ^ n1582 ;
  assign n18312 = n18311 ^ n4004 ^ n1759 ;
  assign n18313 = n14881 ^ n13868 ^ n497 ;
  assign n18314 = ( n789 & ~n9963 ) | ( n789 & n18313 ) | ( ~n9963 & n18313 ) ;
  assign n18315 = ( n4034 & n11454 ) | ( n4034 & n18314 ) | ( n11454 & n18314 ) ;
  assign n18319 = n8509 ^ n6405 ^ n2406 ;
  assign n18320 = ( n1714 & ~n5940 ) | ( n1714 & n13378 ) | ( ~n5940 & n13378 ) ;
  assign n18321 = ( n4538 & n15664 ) | ( n4538 & n18320 ) | ( n15664 & n18320 ) ;
  assign n18322 = ( n5440 & n18319 ) | ( n5440 & n18321 ) | ( n18319 & n18321 ) ;
  assign n18316 = n7246 ^ n1453 ^ n434 ;
  assign n18317 = ( n642 & n6299 ) | ( n642 & ~n8591 ) | ( n6299 & ~n8591 ) ;
  assign n18318 = ( n13189 & n18316 ) | ( n13189 & ~n18317 ) | ( n18316 & ~n18317 ) ;
  assign n18323 = n18322 ^ n18318 ^ n2857 ;
  assign n18324 = n6865 ^ n1934 ^ n150 ;
  assign n18332 = n14672 ^ n12156 ^ n1995 ;
  assign n18325 = n11928 ^ n8133 ^ n1941 ;
  assign n18326 = n11994 ^ n5183 ^ n2236 ;
  assign n18327 = ( ~n766 & n3233 ) | ( ~n766 & n6396 ) | ( n3233 & n6396 ) ;
  assign n18328 = ( n1491 & n6048 ) | ( n1491 & n18327 ) | ( n6048 & n18327 ) ;
  assign n18329 = ( ~n13548 & n18326 ) | ( ~n13548 & n18328 ) | ( n18326 & n18328 ) ;
  assign n18330 = ( n6269 & ~n10153 ) | ( n6269 & n18329 ) | ( ~n10153 & n18329 ) ;
  assign n18331 = ( n4167 & ~n18325 ) | ( n4167 & n18330 ) | ( ~n18325 & n18330 ) ;
  assign n18333 = n18332 ^ n18331 ^ n9070 ;
  assign n18342 = ( ~n746 & n2347 ) | ( ~n746 & n9847 ) | ( n2347 & n9847 ) ;
  assign n18343 = ( n2902 & n5683 ) | ( n2902 & n9667 ) | ( n5683 & n9667 ) ;
  assign n18344 = ( n2734 & n16280 ) | ( n2734 & n18343 ) | ( n16280 & n18343 ) ;
  assign n18345 = n18344 ^ n10874 ^ n5638 ;
  assign n18346 = ( n9545 & ~n18342 ) | ( n9545 & n18345 ) | ( ~n18342 & n18345 ) ;
  assign n18340 = ( n3342 & ~n3470 ) | ( n3342 & n8429 ) | ( ~n3470 & n8429 ) ;
  assign n18338 = n12170 ^ n4596 ^ n2648 ;
  assign n18337 = n16816 ^ n14552 ^ n5337 ;
  assign n18339 = n18338 ^ n18337 ^ n6227 ;
  assign n18334 = ( ~n4101 & n4403 ) | ( ~n4101 & n5967 ) | ( n4403 & n5967 ) ;
  assign n18335 = ( ~n7215 & n8959 ) | ( ~n7215 & n18334 ) | ( n8959 & n18334 ) ;
  assign n18336 = ( ~n2964 & n5473 ) | ( ~n2964 & n18335 ) | ( n5473 & n18335 ) ;
  assign n18341 = n18340 ^ n18339 ^ n18336 ;
  assign n18347 = n18346 ^ n18341 ^ n14062 ;
  assign n18351 = n9776 ^ n2475 ^ n2152 ;
  assign n18348 = n10418 ^ n973 ^ n363 ;
  assign n18349 = n10199 ^ n7471 ^ n3494 ;
  assign n18350 = ( ~n2023 & n18348 ) | ( ~n2023 & n18349 ) | ( n18348 & n18349 ) ;
  assign n18352 = n18351 ^ n18350 ^ n5799 ;
  assign n18353 = n12733 ^ n6160 ^ n651 ;
  assign n18354 = ( n1353 & ~n1922 ) | ( n1353 & n6999 ) | ( ~n1922 & n6999 ) ;
  assign n18355 = ( n3485 & ~n11447 ) | ( n3485 & n18354 ) | ( ~n11447 & n18354 ) ;
  assign n18356 = n14323 ^ n4564 ^ n3264 ;
  assign n18357 = n18356 ^ n11085 ^ n8434 ;
  assign n18358 = ( ~n353 & n18355 ) | ( ~n353 & n18357 ) | ( n18355 & n18357 ) ;
  assign n18359 = ( x125 & n10653 ) | ( x125 & n18358 ) | ( n10653 & n18358 ) ;
  assign n18362 = n11571 ^ n7990 ^ n1280 ;
  assign n18360 = ( x18 & n8441 ) | ( x18 & n9238 ) | ( n8441 & n9238 ) ;
  assign n18361 = ( n3758 & n8928 ) | ( n3758 & ~n18360 ) | ( n8928 & ~n18360 ) ;
  assign n18363 = n18362 ^ n18361 ^ n7023 ;
  assign n18364 = ( n10416 & n13931 ) | ( n10416 & ~n14888 ) | ( n13931 & ~n14888 ) ;
  assign n18365 = n18364 ^ n13990 ^ n7667 ;
  assign n18366 = n5468 ^ n4864 ^ n243 ;
  assign n18367 = ( n1470 & ~n1528 ) | ( n1470 & n13049 ) | ( ~n1528 & n13049 ) ;
  assign n18368 = ( n11583 & ~n18366 ) | ( n11583 & n18367 ) | ( ~n18366 & n18367 ) ;
  assign n18369 = ( ~n15683 & n18365 ) | ( ~n15683 & n18368 ) | ( n18365 & n18368 ) ;
  assign n18370 = n18369 ^ n16401 ^ n11640 ;
  assign n18371 = ( n903 & ~n3950 ) | ( n903 & n8688 ) | ( ~n3950 & n8688 ) ;
  assign n18372 = ( n11443 & n14554 ) | ( n11443 & ~n18371 ) | ( n14554 & ~n18371 ) ;
  assign n18373 = n5984 ^ n3838 ^ n1395 ;
  assign n18374 = ( n3212 & n10257 ) | ( n3212 & n18373 ) | ( n10257 & n18373 ) ;
  assign n18375 = ( n4514 & ~n8401 ) | ( n4514 & n14561 ) | ( ~n8401 & n14561 ) ;
  assign n18377 = n6751 ^ n4873 ^ n4452 ;
  assign n18376 = n12241 ^ n5934 ^ n5266 ;
  assign n18378 = n18377 ^ n18376 ^ n6140 ;
  assign n18379 = n18378 ^ n17021 ^ n4429 ;
  assign n18380 = n9460 ^ n1377 ^ n924 ;
  assign n18381 = ( n3479 & ~n3799 ) | ( n3479 & n7517 ) | ( ~n3799 & n7517 ) ;
  assign n18382 = ( ~n3716 & n3801 ) | ( ~n3716 & n4795 ) | ( n3801 & n4795 ) ;
  assign n18383 = ( n625 & ~n5725 ) | ( n625 & n18382 ) | ( ~n5725 & n18382 ) ;
  assign n18388 = n16874 ^ n10910 ^ n2306 ;
  assign n18386 = n16177 ^ n6583 ^ n1307 ;
  assign n18387 = n18386 ^ n14378 ^ n5863 ;
  assign n18389 = n18388 ^ n18387 ^ n12553 ;
  assign n18384 = ( n8618 & n11250 ) | ( n8618 & n14165 ) | ( n11250 & n14165 ) ;
  assign n18385 = n18384 ^ n10078 ^ n3732 ;
  assign n18390 = n18389 ^ n18385 ^ n10909 ;
  assign n18391 = ( ~n301 & n12904 ) | ( ~n301 & n14274 ) | ( n12904 & n14274 ) ;
  assign n18392 = ( n502 & ~n1318 ) | ( n502 & n4892 ) | ( ~n1318 & n4892 ) ;
  assign n18393 = n18392 ^ n5350 ^ n333 ;
  assign n18394 = ( n10224 & ~n16085 ) | ( n10224 & n18393 ) | ( ~n16085 & n18393 ) ;
  assign n18395 = ( ~n2203 & n8724 ) | ( ~n2203 & n18394 ) | ( n8724 & n18394 ) ;
  assign n18396 = n18395 ^ n8370 ^ n4132 ;
  assign n18397 = ( n17897 & ~n18391 ) | ( n17897 & n18396 ) | ( ~n18391 & n18396 ) ;
  assign n18403 = n12943 ^ n5322 ^ n3529 ;
  assign n18402 = ( n733 & n2210 ) | ( n733 & ~n6881 ) | ( n2210 & ~n6881 ) ;
  assign n18404 = n18403 ^ n18402 ^ n6093 ;
  assign n18405 = n18404 ^ n10260 ^ n2446 ;
  assign n18399 = n5091 ^ n4283 ^ n300 ;
  assign n18400 = n13982 ^ n1118 ^ n749 ;
  assign n18401 = ( n1467 & n18399 ) | ( n1467 & n18400 ) | ( n18399 & n18400 ) ;
  assign n18406 = n18405 ^ n18401 ^ n5067 ;
  assign n18398 = n10139 ^ n1699 ^ n356 ;
  assign n18407 = n18406 ^ n18398 ^ n15192 ;
  assign n18408 = ( ~n1674 & n5954 ) | ( ~n1674 & n11638 ) | ( n5954 & n11638 ) ;
  assign n18409 = ( n382 & n3052 ) | ( n382 & ~n18408 ) | ( n3052 & ~n18408 ) ;
  assign n18410 = ( n11079 & n13127 ) | ( n11079 & ~n18409 ) | ( n13127 & ~n18409 ) ;
  assign n18411 = ( ~n11320 & n15707 ) | ( ~n11320 & n18410 ) | ( n15707 & n18410 ) ;
  assign n18412 = ( n317 & n10441 ) | ( n317 & ~n15585 ) | ( n10441 & ~n15585 ) ;
  assign n18413 = ( n3248 & n18411 ) | ( n3248 & ~n18412 ) | ( n18411 & ~n18412 ) ;
  assign n18414 = n14518 ^ n3328 ^ n630 ;
  assign n18415 = ( n10926 & ~n12401 ) | ( n10926 & n18414 ) | ( ~n12401 & n18414 ) ;
  assign n18416 = ( n1413 & n4387 ) | ( n1413 & n13474 ) | ( n4387 & n13474 ) ;
  assign n18417 = ( n12817 & ~n13145 ) | ( n12817 & n18416 ) | ( ~n13145 & n18416 ) ;
  assign n18418 = n18417 ^ n14734 ^ n6632 ;
  assign n18423 = ( x120 & ~n9242 ) | ( x120 & n12097 ) | ( ~n9242 & n12097 ) ;
  assign n18424 = n18423 ^ n13269 ^ n3476 ;
  assign n18425 = ( n977 & ~n7943 ) | ( n977 & n18424 ) | ( ~n7943 & n18424 ) ;
  assign n18422 = ( n3475 & n7253 ) | ( n3475 & ~n14591 ) | ( n7253 & ~n14591 ) ;
  assign n18420 = ( n2460 & n2602 ) | ( n2460 & n7184 ) | ( n2602 & n7184 ) ;
  assign n18419 = ( ~n7015 & n9082 ) | ( ~n7015 & n13221 ) | ( n9082 & n13221 ) ;
  assign n18421 = n18420 ^ n18419 ^ n14954 ;
  assign n18426 = n18425 ^ n18422 ^ n18421 ;
  assign n18427 = ( n2243 & n6022 ) | ( n2243 & ~n9776 ) | ( n6022 & ~n9776 ) ;
  assign n18429 = n5460 ^ n4798 ^ n3323 ;
  assign n18428 = n12118 ^ n10607 ^ n3730 ;
  assign n18430 = n18429 ^ n18428 ^ n12422 ;
  assign n18431 = n4467 ^ n2628 ^ n574 ;
  assign n18432 = ( x110 & n525 ) | ( x110 & n8236 ) | ( n525 & n8236 ) ;
  assign n18433 = n18432 ^ n9851 ^ n2097 ;
  assign n18434 = ( n1907 & n1913 ) | ( n1907 & ~n2809 ) | ( n1913 & ~n2809 ) ;
  assign n18435 = ( n8266 & ~n8830 ) | ( n8266 & n9652 ) | ( ~n8830 & n9652 ) ;
  assign n18436 = ( n4291 & ~n5102 ) | ( n4291 & n10240 ) | ( ~n5102 & n10240 ) ;
  assign n18437 = ( ~n11084 & n17443 ) | ( ~n11084 & n18436 ) | ( n17443 & n18436 ) ;
  assign n18438 = n18437 ^ n12587 ^ n954 ;
  assign n18439 = ( n18434 & n18435 ) | ( n18434 & n18438 ) | ( n18435 & n18438 ) ;
  assign n18440 = ( n467 & n5763 ) | ( n467 & ~n18439 ) | ( n5763 & ~n18439 ) ;
  assign n18446 = n10153 ^ n4467 ^ n387 ;
  assign n18447 = n18446 ^ n16913 ^ n9880 ;
  assign n18441 = n6832 ^ n5422 ^ n5027 ;
  assign n18442 = ( n2832 & n15201 ) | ( n2832 & ~n18441 ) | ( n15201 & ~n18441 ) ;
  assign n18443 = n18442 ^ n16768 ^ n3248 ;
  assign n18444 = ( ~n3303 & n6028 ) | ( ~n3303 & n18443 ) | ( n6028 & n18443 ) ;
  assign n18445 = ( n10471 & ~n15628 ) | ( n10471 & n18444 ) | ( ~n15628 & n18444 ) ;
  assign n18448 = n18447 ^ n18445 ^ n13799 ;
  assign n18449 = ( n3018 & ~n3834 ) | ( n3018 & n15670 ) | ( ~n3834 & n15670 ) ;
  assign n18450 = ( n11568 & n16227 ) | ( n11568 & n17023 ) | ( n16227 & n17023 ) ;
  assign n18451 = n12240 ^ n8461 ^ n987 ;
  assign n18452 = ( n849 & ~n7427 ) | ( n849 & n12038 ) | ( ~n7427 & n12038 ) ;
  assign n18453 = n18452 ^ n14857 ^ n7495 ;
  assign n18454 = n18453 ^ n16404 ^ n10045 ;
  assign n18455 = ( n2362 & ~n18451 ) | ( n2362 & n18454 ) | ( ~n18451 & n18454 ) ;
  assign n18457 = ( n4780 & n5236 ) | ( n4780 & ~n6440 ) | ( n5236 & ~n6440 ) ;
  assign n18458 = ( n4568 & n10071 ) | ( n4568 & ~n18457 ) | ( n10071 & ~n18457 ) ;
  assign n18456 = ( n1105 & n6555 ) | ( n1105 & ~n14553 ) | ( n6555 & ~n14553 ) ;
  assign n18459 = n18458 ^ n18456 ^ n6500 ;
  assign n18460 = n18377 ^ n10954 ^ n1549 ;
  assign n18461 = n18460 ^ n7803 ^ n1156 ;
  assign n18462 = n18461 ^ n16553 ^ n400 ;
  assign n18463 = ( n4840 & n9205 ) | ( n4840 & ~n13041 ) | ( n9205 & ~n13041 ) ;
  assign n18464 = n7934 ^ n5426 ^ n4606 ;
  assign n18465 = ( ~n12802 & n18463 ) | ( ~n12802 & n18464 ) | ( n18463 & n18464 ) ;
  assign n18466 = n13686 ^ n5112 ^ x30 ;
  assign n18467 = n18466 ^ n18049 ^ n8941 ;
  assign n18468 = ( n3854 & n7037 ) | ( n3854 & n11228 ) | ( n7037 & n11228 ) ;
  assign n18469 = ( n3633 & ~n6856 ) | ( n3633 & n11297 ) | ( ~n6856 & n11297 ) ;
  assign n18470 = ( n15321 & ~n17700 ) | ( n15321 & n18469 ) | ( ~n17700 & n18469 ) ;
  assign n18471 = n15714 ^ n15189 ^ n521 ;
  assign n18472 = ( ~n909 & n2499 ) | ( ~n909 & n16445 ) | ( n2499 & n16445 ) ;
  assign n18473 = ( x122 & ~n8244 ) | ( x122 & n16834 ) | ( ~n8244 & n16834 ) ;
  assign n18474 = ( n901 & n2160 ) | ( n901 & ~n18473 ) | ( n2160 & ~n18473 ) ;
  assign n18475 = ( n9345 & n13563 ) | ( n9345 & ~n18474 ) | ( n13563 & ~n18474 ) ;
  assign n18476 = ( ~n18046 & n18472 ) | ( ~n18046 & n18475 ) | ( n18472 & n18475 ) ;
  assign n18477 = ( n12216 & n16714 ) | ( n12216 & ~n18476 ) | ( n16714 & ~n18476 ) ;
  assign n18478 = n15417 ^ n1943 ^ n1155 ;
  assign n18479 = n9321 ^ n6502 ^ n1690 ;
  assign n18480 = n18479 ^ n14627 ^ n768 ;
  assign n18481 = ( n14173 & n18478 ) | ( n14173 & ~n18480 ) | ( n18478 & ~n18480 ) ;
  assign n18482 = n6566 ^ n3824 ^ n536 ;
  assign n18483 = n13533 ^ n10415 ^ n584 ;
  assign n18484 = ( n10670 & n15727 ) | ( n10670 & ~n18483 ) | ( n15727 & ~n18483 ) ;
  assign n18485 = n18484 ^ n9974 ^ n1224 ;
  assign n18489 = n17789 ^ n11418 ^ n8538 ;
  assign n18490 = ( n3206 & ~n16127 ) | ( n3206 & n18489 ) | ( ~n16127 & n18489 ) ;
  assign n18486 = n6582 ^ n5991 ^ n4614 ;
  assign n18487 = ( n545 & ~n4327 ) | ( n545 & n8082 ) | ( ~n4327 & n8082 ) ;
  assign n18488 = ( n13685 & n18486 ) | ( n13685 & n18487 ) | ( n18486 & n18487 ) ;
  assign n18491 = n18490 ^ n18488 ^ n6843 ;
  assign n18492 = ( n379 & n2724 ) | ( n379 & ~n8001 ) | ( n2724 & ~n8001 ) ;
  assign n18493 = ( n965 & n7655 ) | ( n965 & ~n18492 ) | ( n7655 & ~n18492 ) ;
  assign n18494 = n18493 ^ n14140 ^ n3276 ;
  assign n18499 = n7615 ^ n2379 ^ x49 ;
  assign n18495 = n14118 ^ n11545 ^ n2557 ;
  assign n18496 = n18495 ^ n7966 ^ n4435 ;
  assign n18497 = ( n4003 & ~n7119 ) | ( n4003 & n18496 ) | ( ~n7119 & n18496 ) ;
  assign n18498 = ( n2164 & n7004 ) | ( n2164 & n18497 ) | ( n7004 & n18497 ) ;
  assign n18500 = n18499 ^ n18498 ^ n14495 ;
  assign n18501 = n17014 ^ n8848 ^ n6098 ;
  assign n18509 = ( n1163 & n2199 ) | ( n1163 & ~n12676 ) | ( n2199 & ~n12676 ) ;
  assign n18507 = n17991 ^ n6259 ^ n2094 ;
  assign n18508 = ( ~n11957 & n13920 ) | ( ~n11957 & n18507 ) | ( n13920 & n18507 ) ;
  assign n18504 = n16598 ^ n5370 ^ n2469 ;
  assign n18505 = n18504 ^ n3826 ^ x10 ;
  assign n18502 = ( n1288 & ~n12837 ) | ( n1288 & n14766 ) | ( ~n12837 & n14766 ) ;
  assign n18503 = n18502 ^ n5904 ^ n1385 ;
  assign n18506 = n18505 ^ n18503 ^ n9418 ;
  assign n18510 = n18509 ^ n18508 ^ n18506 ;
  assign n18511 = ( n7450 & n11327 ) | ( n7450 & ~n15625 ) | ( n11327 & ~n15625 ) ;
  assign n18512 = n18511 ^ n13265 ^ n11414 ;
  assign n18513 = n18512 ^ n4237 ^ n3186 ;
  assign n18514 = n12463 ^ n8647 ^ n5724 ;
  assign n18515 = ( n6673 & n10909 ) | ( n6673 & ~n18457 ) | ( n10909 & ~n18457 ) ;
  assign n18516 = ( n8725 & ~n9893 ) | ( n8725 & n18515 ) | ( ~n9893 & n18515 ) ;
  assign n18517 = n17536 ^ n16383 ^ n10190 ;
  assign n18518 = n11066 ^ n9144 ^ n2020 ;
  assign n18519 = ( ~n6572 & n7339 ) | ( ~n6572 & n18518 ) | ( n7339 & n18518 ) ;
  assign n18520 = ( ~n18516 & n18517 ) | ( ~n18516 & n18519 ) | ( n18517 & n18519 ) ;
  assign n18521 = ( n9217 & n10042 ) | ( n9217 & n11355 ) | ( n10042 & n11355 ) ;
  assign n18530 = n8529 ^ n2457 ^ n1899 ;
  assign n18531 = ( ~n6932 & n10310 ) | ( ~n6932 & n18530 ) | ( n10310 & n18530 ) ;
  assign n18528 = n13261 ^ n6542 ^ n3863 ;
  assign n18527 = ( n3309 & n4076 ) | ( n3309 & n10247 ) | ( n4076 & n10247 ) ;
  assign n18523 = ( n201 & ~n3913 ) | ( n201 & n4834 ) | ( ~n3913 & n4834 ) ;
  assign n18524 = n18523 ^ n14932 ^ n4677 ;
  assign n18525 = n18524 ^ n14590 ^ n12631 ;
  assign n18526 = n18525 ^ n13598 ^ n12591 ;
  assign n18529 = n18528 ^ n18527 ^ n18526 ;
  assign n18522 = ( ~n5989 & n12716 ) | ( ~n5989 & n13756 ) | ( n12716 & n13756 ) ;
  assign n18532 = n18531 ^ n18529 ^ n18522 ;
  assign n18536 = ( ~n155 & n712 ) | ( ~n155 & n3094 ) | ( n712 & n3094 ) ;
  assign n18537 = ( ~n11418 & n13080 ) | ( ~n11418 & n18536 ) | ( n13080 & n18536 ) ;
  assign n18533 = ( n11344 & n11578 ) | ( n11344 & n15521 ) | ( n11578 & n15521 ) ;
  assign n18534 = ( n11958 & n14190 ) | ( n11958 & ~n16090 ) | ( n14190 & ~n16090 ) ;
  assign n18535 = ( ~n6184 & n18533 ) | ( ~n6184 & n18534 ) | ( n18533 & n18534 ) ;
  assign n18538 = n18537 ^ n18535 ^ n4276 ;
  assign n18539 = ( n4192 & n14009 ) | ( n4192 & n15305 ) | ( n14009 & n15305 ) ;
  assign n18540 = n18539 ^ n5841 ^ n323 ;
  assign n18542 = n7943 ^ n6171 ^ n1628 ;
  assign n18543 = n18542 ^ n10997 ^ n7359 ;
  assign n18541 = ( n4113 & ~n8460 ) | ( n4113 & n9444 ) | ( ~n8460 & n9444 ) ;
  assign n18544 = n18543 ^ n18541 ^ n13707 ;
  assign n18545 = n18544 ^ n3892 ^ n3096 ;
  assign n18546 = ( n5655 & ~n15590 ) | ( n5655 & n16574 ) | ( ~n15590 & n16574 ) ;
  assign n18547 = n18546 ^ n8378 ^ n2464 ;
  assign n18548 = n16205 ^ n6108 ^ n5969 ;
  assign n18549 = n8770 ^ n1975 ^ x39 ;
  assign n18550 = n18549 ^ n11939 ^ n5522 ;
  assign n18551 = n16211 ^ n8212 ^ n2304 ;
  assign n18552 = ( n18548 & ~n18550 ) | ( n18548 & n18551 ) | ( ~n18550 & n18551 ) ;
  assign n18553 = ( n1490 & n2228 ) | ( n1490 & ~n15499 ) | ( n2228 & ~n15499 ) ;
  assign n18554 = n18553 ^ n8766 ^ n5763 ;
  assign n18555 = n14522 ^ n6056 ^ n240 ;
  assign n18556 = n10148 ^ n5520 ^ n3901 ;
  assign n18557 = n9892 ^ n4761 ^ n3141 ;
  assign n18558 = ( n6642 & n18556 ) | ( n6642 & n18557 ) | ( n18556 & n18557 ) ;
  assign n18559 = n4914 ^ n2156 ^ n1953 ;
  assign n18560 = n18559 ^ n11248 ^ n7159 ;
  assign n18561 = ( n7736 & ~n10521 ) | ( n7736 & n15256 ) | ( ~n10521 & n15256 ) ;
  assign n18562 = n18561 ^ n8160 ^ n2914 ;
  assign n18563 = ( ~x74 & n1201 ) | ( ~x74 & n4283 ) | ( n1201 & n4283 ) ;
  assign n18564 = ( x66 & n2896 ) | ( x66 & ~n4338 ) | ( n2896 & ~n4338 ) ;
  assign n18565 = n18564 ^ n5923 ^ n2359 ;
  assign n18566 = ( ~n6183 & n14939 ) | ( ~n6183 & n18565 ) | ( n14939 & n18565 ) ;
  assign n18567 = ( n1294 & n18563 ) | ( n1294 & n18566 ) | ( n18563 & n18566 ) ;
  assign n18568 = n13922 ^ n12352 ^ n11207 ;
  assign n18569 = ( n1470 & ~n7070 ) | ( n1470 & n18568 ) | ( ~n7070 & n18568 ) ;
  assign n18570 = ( n305 & n3296 ) | ( n305 & ~n3781 ) | ( n3296 & ~n3781 ) ;
  assign n18571 = ( n4425 & ~n9774 ) | ( n4425 & n18570 ) | ( ~n9774 & n18570 ) ;
  assign n18572 = ( n798 & n4191 ) | ( n798 & n10096 ) | ( n4191 & n10096 ) ;
  assign n18573 = ( n2269 & n6748 ) | ( n2269 & n18572 ) | ( n6748 & n18572 ) ;
  assign n18574 = ( n315 & n8777 ) | ( n315 & n10075 ) | ( n8777 & n10075 ) ;
  assign n18575 = n7861 ^ n4186 ^ n323 ;
  assign n18576 = n18575 ^ n8813 ^ n4136 ;
  assign n18577 = ( n3716 & ~n7908 ) | ( n3716 & n17248 ) | ( ~n7908 & n17248 ) ;
  assign n18578 = ( ~n3671 & n9203 ) | ( ~n3671 & n12705 ) | ( n9203 & n12705 ) ;
  assign n18579 = ( n3035 & ~n13255 ) | ( n3035 & n18578 ) | ( ~n13255 & n18578 ) ;
  assign n18580 = ( n2744 & n6845 ) | ( n2744 & n18579 ) | ( n6845 & n18579 ) ;
  assign n18586 = n8807 ^ n3365 ^ n2139 ;
  assign n18587 = ( n577 & n12042 ) | ( n577 & n18586 ) | ( n12042 & n18586 ) ;
  assign n18582 = n11742 ^ n6123 ^ n1068 ;
  assign n18583 = ( n1700 & n3119 ) | ( n1700 & ~n7116 ) | ( n3119 & ~n7116 ) ;
  assign n18584 = n18583 ^ n12054 ^ n10305 ;
  assign n18585 = ( ~n9239 & n18582 ) | ( ~n9239 & n18584 ) | ( n18582 & n18584 ) ;
  assign n18581 = n9255 ^ n1763 ^ n570 ;
  assign n18588 = n18587 ^ n18585 ^ n18581 ;
  assign n18589 = ( n2614 & ~n13619 ) | ( n2614 & n18588 ) | ( ~n13619 & n18588 ) ;
  assign n18591 = n12915 ^ n6068 ^ n667 ;
  assign n18592 = ( ~n825 & n952 ) | ( ~n825 & n18591 ) | ( n952 & n18591 ) ;
  assign n18590 = n16373 ^ n14396 ^ n10937 ;
  assign n18593 = n18592 ^ n18590 ^ n4110 ;
  assign n18594 = n18593 ^ n6595 ^ n1987 ;
  assign n18595 = ( n2497 & n6030 ) | ( n2497 & ~n16690 ) | ( n6030 & ~n16690 ) ;
  assign n18596 = n18595 ^ n3123 ^ n295 ;
  assign n18597 = n18596 ^ n15710 ^ n12811 ;
  assign n18598 = ( n1528 & ~n3877 ) | ( n1528 & n7499 ) | ( ~n3877 & n7499 ) ;
  assign n18599 = ( n204 & n379 ) | ( n204 & n9264 ) | ( n379 & n9264 ) ;
  assign n18600 = n18599 ^ n2358 ^ x75 ;
  assign n18601 = n18600 ^ n8898 ^ n3701 ;
  assign n18603 = n8843 ^ n7773 ^ n7253 ;
  assign n18604 = n18603 ^ n5069 ^ n476 ;
  assign n18602 = ( n824 & n7746 ) | ( n824 & n11764 ) | ( n7746 & n11764 ) ;
  assign n18605 = n18604 ^ n18602 ^ n2707 ;
  assign n18606 = n15161 ^ n11815 ^ n2274 ;
  assign n18607 = ( ~n13934 & n18605 ) | ( ~n13934 & n18606 ) | ( n18605 & n18606 ) ;
  assign n18608 = n7289 ^ n3255 ^ n796 ;
  assign n18609 = n14094 ^ n10735 ^ n1496 ;
  assign n18610 = n18609 ^ n17530 ^ n590 ;
  assign n18611 = ( n566 & ~n3125 ) | ( n566 & n18610 ) | ( ~n3125 & n18610 ) ;
  assign n18612 = ( ~n3211 & n12798 ) | ( ~n3211 & n16310 ) | ( n12798 & n16310 ) ;
  assign n18613 = ( n10665 & n13870 ) | ( n10665 & n18612 ) | ( n13870 & n18612 ) ;
  assign n18614 = ( ~n6067 & n8461 ) | ( ~n6067 & n8573 ) | ( n8461 & n8573 ) ;
  assign n18615 = ( ~n8974 & n12194 ) | ( ~n8974 & n17561 ) | ( n12194 & n17561 ) ;
  assign n18616 = n7421 ^ n4185 ^ n1029 ;
  assign n18617 = ( n4240 & n5806 ) | ( n4240 & ~n18616 ) | ( n5806 & ~n18616 ) ;
  assign n18618 = ( n7971 & n16870 ) | ( n7971 & n18617 ) | ( n16870 & n18617 ) ;
  assign n18619 = ( n5868 & n13834 ) | ( n5868 & n18618 ) | ( n13834 & n18618 ) ;
  assign n18620 = ( ~n8917 & n18615 ) | ( ~n8917 & n18619 ) | ( n18615 & n18619 ) ;
  assign n18621 = n13770 ^ n13454 ^ n10807 ;
  assign n18622 = n18621 ^ n13042 ^ n2686 ;
  assign n18623 = n9562 ^ n7525 ^ n4756 ;
  assign n18624 = ( n866 & n3962 ) | ( n866 & n7381 ) | ( n3962 & n7381 ) ;
  assign n18625 = ( n14812 & n18623 ) | ( n14812 & n18624 ) | ( n18623 & n18624 ) ;
  assign n18626 = ( n4835 & n8880 ) | ( n4835 & n18625 ) | ( n8880 & n18625 ) ;
  assign n18627 = n11475 ^ n10017 ^ n3305 ;
  assign n18628 = n11886 ^ n3486 ^ n2908 ;
  assign n18629 = n18628 ^ n11768 ^ n7961 ;
  assign n18635 = n4930 ^ n4120 ^ n3214 ;
  assign n18633 = n10771 ^ n6524 ^ n293 ;
  assign n18630 = n15028 ^ n837 ^ n425 ;
  assign n18631 = ( n2981 & n9399 ) | ( n2981 & ~n18630 ) | ( n9399 & ~n18630 ) ;
  assign n18632 = ( n4043 & n18178 ) | ( n4043 & ~n18631 ) | ( n18178 & ~n18631 ) ;
  assign n18634 = n18633 ^ n18632 ^ n8027 ;
  assign n18636 = n18635 ^ n18634 ^ n15925 ;
  assign n18639 = ( n458 & n12050 ) | ( n458 & ~n12693 ) | ( n12050 & ~n12693 ) ;
  assign n18640 = ( n1934 & n7096 ) | ( n1934 & ~n12856 ) | ( n7096 & ~n12856 ) ;
  assign n18641 = ( n5939 & n18074 ) | ( n5939 & ~n18640 ) | ( n18074 & ~n18640 ) ;
  assign n18642 = ( n17348 & n18639 ) | ( n17348 & ~n18641 ) | ( n18639 & ~n18641 ) ;
  assign n18637 = ( n1571 & n9756 ) | ( n1571 & n11173 ) | ( n9756 & n11173 ) ;
  assign n18638 = n18637 ^ n7655 ^ n7196 ;
  assign n18643 = n18642 ^ n18638 ^ n713 ;
  assign n18644 = ( n3007 & ~n9865 ) | ( n3007 & n15874 ) | ( ~n9865 & n15874 ) ;
  assign n18645 = ( n2600 & ~n10900 ) | ( n2600 & n18644 ) | ( ~n10900 & n18644 ) ;
  assign n18646 = n10895 ^ n7095 ^ n5484 ;
  assign n18647 = ( n9573 & ~n13436 ) | ( n9573 & n18646 ) | ( ~n13436 & n18646 ) ;
  assign n18648 = n7294 ^ n2987 ^ n360 ;
  assign n18649 = n18648 ^ n16183 ^ n4127 ;
  assign n18651 = ( x82 & ~n9956 ) | ( x82 & n12752 ) | ( ~n9956 & n12752 ) ;
  assign n18650 = ( ~n4546 & n9947 ) | ( ~n4546 & n14067 ) | ( n9947 & n14067 ) ;
  assign n18652 = n18651 ^ n18650 ^ n12216 ;
  assign n18655 = ( n1783 & n5131 ) | ( n1783 & n7901 ) | ( n5131 & n7901 ) ;
  assign n18653 = n7281 ^ n4916 ^ n1373 ;
  assign n18654 = n18653 ^ n13092 ^ n1952 ;
  assign n18656 = n18655 ^ n18654 ^ n12765 ;
  assign n18657 = ( n1292 & n13975 ) | ( n1292 & n14036 ) | ( n13975 & n14036 ) ;
  assign n18658 = ( ~n150 & n1046 ) | ( ~n150 & n1732 ) | ( n1046 & n1732 ) ;
  assign n18659 = ( ~n9789 & n14561 ) | ( ~n9789 & n18658 ) | ( n14561 & n18658 ) ;
  assign n18660 = n16870 ^ n13143 ^ n10232 ;
  assign n18661 = ( n18657 & n18659 ) | ( n18657 & ~n18660 ) | ( n18659 & ~n18660 ) ;
  assign n18662 = n11396 ^ n11178 ^ n1164 ;
  assign n18663 = ( n544 & n18316 ) | ( n544 & n18662 ) | ( n18316 & n18662 ) ;
  assign n18664 = n18663 ^ n14025 ^ n9896 ;
  assign n18665 = n18159 ^ n9884 ^ n3504 ;
  assign n18666 = ( n2974 & ~n9335 ) | ( n2974 & n11467 ) | ( ~n9335 & n11467 ) ;
  assign n18667 = ( n3262 & n18665 ) | ( n3262 & n18666 ) | ( n18665 & n18666 ) ;
  assign n18668 = ( x114 & n9662 ) | ( x114 & ~n18667 ) | ( n9662 & ~n18667 ) ;
  assign n18669 = ( ~n4963 & n9446 ) | ( ~n4963 & n10594 ) | ( n9446 & n10594 ) ;
  assign n18670 = ( n1065 & ~n12024 ) | ( n1065 & n14144 ) | ( ~n12024 & n14144 ) ;
  assign n18671 = n8858 ^ n7607 ^ n6639 ;
  assign n18672 = n18671 ^ n16635 ^ n9325 ;
  assign n18673 = n10434 ^ n1630 ^ x124 ;
  assign n18675 = n10439 ^ n3107 ^ n2749 ;
  assign n18674 = n2103 ^ n1309 ^ n587 ;
  assign n18676 = n18675 ^ n18674 ^ n1128 ;
  assign n18677 = n18676 ^ n12921 ^ n8189 ;
  assign n18678 = ( x11 & n11171 ) | ( x11 & ~n18677 ) | ( n11171 & ~n18677 ) ;
  assign n18679 = n8138 ^ n7650 ^ n6421 ;
  assign n18680 = n18679 ^ n6435 ^ n6384 ;
  assign n18681 = ( ~n331 & n4554 ) | ( ~n331 & n17080 ) | ( n4554 & n17080 ) ;
  assign n18682 = ( n4485 & n4901 ) | ( n4485 & ~n12643 ) | ( n4901 & ~n12643 ) ;
  assign n18683 = n18682 ^ n11311 ^ n4873 ;
  assign n18685 = n10056 ^ n5073 ^ n4673 ;
  assign n18684 = ( n9854 & n14062 ) | ( n9854 & n14492 ) | ( n14062 & n14492 ) ;
  assign n18686 = n18685 ^ n18684 ^ n8808 ;
  assign n18688 = ( n1983 & ~n10505 ) | ( n1983 & n17031 ) | ( ~n10505 & n17031 ) ;
  assign n18689 = ( n4515 & ~n14504 ) | ( n4515 & n18688 ) | ( ~n14504 & n18688 ) ;
  assign n18687 = n5372 ^ n5054 ^ n1032 ;
  assign n18690 = n18689 ^ n18687 ^ n8059 ;
  assign n18697 = n14724 ^ n7254 ^ n7165 ;
  assign n18691 = ( ~n2469 & n5077 ) | ( ~n2469 & n8341 ) | ( n5077 & n8341 ) ;
  assign n18692 = n18691 ^ n10244 ^ n3441 ;
  assign n18693 = n18692 ^ n10237 ^ n439 ;
  assign n18694 = n13185 ^ n9919 ^ n9000 ;
  assign n18695 = ( n4099 & ~n13904 ) | ( n4099 & n14248 ) | ( ~n13904 & n14248 ) ;
  assign n18696 = ( n18693 & ~n18694 ) | ( n18693 & n18695 ) | ( ~n18694 & n18695 ) ;
  assign n18698 = n18697 ^ n18696 ^ n6158 ;
  assign n18699 = ( ~n157 & n5435 ) | ( ~n157 & n8480 ) | ( n5435 & n8480 ) ;
  assign n18700 = n18699 ^ n15969 ^ n3017 ;
  assign n18701 = ( n9183 & n11910 ) | ( n9183 & n14777 ) | ( n11910 & n14777 ) ;
  assign n18702 = ( n13371 & n14965 ) | ( n13371 & ~n18701 ) | ( n14965 & ~n18701 ) ;
  assign n18704 = ( n2184 & n2564 ) | ( n2184 & ~n8084 ) | ( n2564 & ~n8084 ) ;
  assign n18703 = ( n1739 & n2003 ) | ( n1739 & ~n13360 ) | ( n2003 & ~n13360 ) ;
  assign n18705 = n18704 ^ n18703 ^ n14658 ;
  assign n18706 = ( n13324 & ~n18702 ) | ( n13324 & n18705 ) | ( ~n18702 & n18705 ) ;
  assign n18707 = n14009 ^ n3485 ^ n380 ;
  assign n18708 = n16003 ^ n8734 ^ n2910 ;
  assign n18709 = ( n4544 & n5286 ) | ( n4544 & ~n18708 ) | ( n5286 & ~n18708 ) ;
  assign n18710 = n8558 ^ n7576 ^ n221 ;
  assign n18711 = n18710 ^ n1092 ^ n461 ;
  assign n18712 = ( n2910 & ~n3470 ) | ( n2910 & n18711 ) | ( ~n3470 & n18711 ) ;
  assign n18713 = ( ~n5049 & n15351 ) | ( ~n5049 & n18712 ) | ( n15351 & n18712 ) ;
  assign n18714 = ( n325 & n4216 ) | ( n325 & n8276 ) | ( n4216 & n8276 ) ;
  assign n18715 = ( n4035 & ~n14334 ) | ( n4035 & n18714 ) | ( ~n14334 & n18714 ) ;
  assign n18716 = n13634 ^ n5415 ^ n2268 ;
  assign n18717 = ( ~n510 & n2397 ) | ( ~n510 & n6133 ) | ( n2397 & n6133 ) ;
  assign n18718 = ( n4621 & n5965 ) | ( n4621 & n18717 ) | ( n5965 & n18717 ) ;
  assign n18719 = n8938 ^ n7927 ^ n2589 ;
  assign n18720 = n18023 ^ n13776 ^ n1539 ;
  assign n18721 = n10590 ^ n4525 ^ n1022 ;
  assign n18722 = n18721 ^ n11235 ^ n10662 ;
  assign n18723 = ( n13966 & ~n18720 ) | ( n13966 & n18722 ) | ( ~n18720 & n18722 ) ;
  assign n18724 = n13711 ^ n11907 ^ n2351 ;
  assign n18725 = n13310 ^ n4012 ^ n585 ;
  assign n18726 = ( n1637 & n3164 ) | ( n1637 & ~n18725 ) | ( n3164 & ~n18725 ) ;
  assign n18727 = ( n4949 & n5505 ) | ( n4949 & ~n17787 ) | ( n5505 & ~n17787 ) ;
  assign n18732 = ( ~n2718 & n3107 ) | ( ~n2718 & n4671 ) | ( n3107 & n4671 ) ;
  assign n18730 = n12974 ^ n11932 ^ n4167 ;
  assign n18731 = ( n9676 & n15692 ) | ( n9676 & ~n18730 ) | ( n15692 & ~n18730 ) ;
  assign n18728 = ( ~n6981 & n13287 ) | ( ~n6981 & n16626 ) | ( n13287 & n16626 ) ;
  assign n18729 = n18728 ^ n15297 ^ n525 ;
  assign n18733 = n18732 ^ n18731 ^ n18729 ;
  assign n18734 = ( ~n1204 & n5329 ) | ( ~n1204 & n7778 ) | ( n5329 & n7778 ) ;
  assign n18735 = n5216 ^ n4451 ^ n3984 ;
  assign n18736 = n18735 ^ n14168 ^ n4597 ;
  assign n18737 = n18736 ^ n8032 ^ n5175 ;
  assign n18738 = ( n1671 & n11191 ) | ( n1671 & ~n18737 ) | ( n11191 & ~n18737 ) ;
  assign n18739 = n12841 ^ n10021 ^ n5521 ;
  assign n18740 = n18739 ^ n11997 ^ n1248 ;
  assign n18741 = ( n9619 & n18738 ) | ( n9619 & ~n18740 ) | ( n18738 & ~n18740 ) ;
  assign n18744 = ( n456 & n3940 ) | ( n456 & n4410 ) | ( n3940 & n4410 ) ;
  assign n18745 = n15063 ^ n9066 ^ n3209 ;
  assign n18746 = ( n5214 & ~n18744 ) | ( n5214 & n18745 ) | ( ~n18744 & n18745 ) ;
  assign n18742 = n15253 ^ n1878 ^ n248 ;
  assign n18743 = ( n6743 & n8925 ) | ( n6743 & n18742 ) | ( n8925 & n18742 ) ;
  assign n18747 = n18746 ^ n18743 ^ n10967 ;
  assign n18748 = n14283 ^ n12243 ^ n4881 ;
  assign n18749 = ( n3274 & n11171 ) | ( n3274 & n15083 ) | ( n11171 & n15083 ) ;
  assign n18751 = ( ~x58 & n11551 ) | ( ~x58 & n15843 ) | ( n11551 & n15843 ) ;
  assign n18752 = ( n5615 & ~n6818 ) | ( n5615 & n18751 ) | ( ~n6818 & n18751 ) ;
  assign n18753 = ( n4133 & ~n9855 ) | ( n4133 & n18752 ) | ( ~n9855 & n18752 ) ;
  assign n18754 = n18753 ^ n15875 ^ n6832 ;
  assign n18755 = n18754 ^ n7704 ^ n1099 ;
  assign n18750 = ( n2722 & ~n12229 ) | ( n2722 & n15028 ) | ( ~n12229 & n15028 ) ;
  assign n18756 = n18755 ^ n18750 ^ n1649 ;
  assign n18757 = n18756 ^ n17323 ^ n15519 ;
  assign n18758 = n18757 ^ n5593 ^ n5479 ;
  assign n18759 = n4640 ^ n4219 ^ n1941 ;
  assign n18760 = ( n2143 & ~n15291 ) | ( n2143 & n18759 ) | ( ~n15291 & n18759 ) ;
  assign n18761 = n17643 ^ n17146 ^ n4761 ;
  assign n18762 = ( n1640 & n9033 ) | ( n1640 & n18761 ) | ( n9033 & n18761 ) ;
  assign n18763 = ( n7148 & ~n12982 ) | ( n7148 & n18762 ) | ( ~n12982 & n18762 ) ;
  assign n18764 = n18498 ^ n11273 ^ n3133 ;
  assign n18765 = ( n4985 & n7032 ) | ( n4985 & n7057 ) | ( n7032 & n7057 ) ;
  assign n18766 = n18765 ^ n13216 ^ n5841 ;
  assign n18767 = n18766 ^ n12587 ^ n4248 ;
  assign n18768 = n13269 ^ n12555 ^ n5134 ;
  assign n18769 = ( n2231 & n6069 ) | ( n2231 & ~n14992 ) | ( n6069 & ~n14992 ) ;
  assign n18770 = n18769 ^ n9470 ^ n7979 ;
  assign n18771 = n18770 ^ n18529 ^ n7398 ;
  assign n18772 = ( n679 & ~n4468 ) | ( n679 & n16059 ) | ( ~n4468 & n16059 ) ;
  assign n18774 = ( n1968 & ~n3159 ) | ( n1968 & n8772 ) | ( ~n3159 & n8772 ) ;
  assign n18773 = n8368 ^ n2672 ^ n1272 ;
  assign n18775 = n18774 ^ n18773 ^ n11541 ;
  assign n18777 = ( n369 & ~n8970 ) | ( n369 & n10466 ) | ( ~n8970 & n10466 ) ;
  assign n18778 = ( n4898 & n5304 ) | ( n4898 & ~n18777 ) | ( n5304 & ~n18777 ) ;
  assign n18776 = ( n567 & n3295 ) | ( n567 & n8670 ) | ( n3295 & n8670 ) ;
  assign n18779 = n18778 ^ n18776 ^ n13482 ;
  assign n18780 = ( ~n4589 & n15102 ) | ( ~n4589 & n18779 ) | ( n15102 & n18779 ) ;
  assign n18781 = n5081 ^ n4492 ^ n1204 ;
  assign n18782 = ( ~n3987 & n7238 ) | ( ~n3987 & n7557 ) | ( n7238 & n7557 ) ;
  assign n18783 = ( ~n2081 & n4361 ) | ( ~n2081 & n18782 ) | ( n4361 & n18782 ) ;
  assign n18784 = ( n10602 & n18781 ) | ( n10602 & ~n18783 ) | ( n18781 & ~n18783 ) ;
  assign n18785 = n10087 ^ n2965 ^ n725 ;
  assign n18786 = n7041 ^ n4795 ^ x16 ;
  assign n18787 = ( n7455 & n9011 ) | ( n7455 & ~n18786 ) | ( n9011 & ~n18786 ) ;
  assign n18788 = ( n378 & n4412 ) | ( n378 & ~n18787 ) | ( n4412 & ~n18787 ) ;
  assign n18789 = ( n1615 & n12906 ) | ( n1615 & ~n16252 ) | ( n12906 & ~n16252 ) ;
  assign n18790 = n18789 ^ n17231 ^ n7960 ;
  assign n18791 = n11357 ^ n10821 ^ n7212 ;
  assign n18794 = n10282 ^ n6129 ^ n2890 ;
  assign n18792 = ( ~n7870 & n16314 ) | ( ~n7870 & n17626 ) | ( n16314 & n17626 ) ;
  assign n18793 = ( ~n6505 & n18666 ) | ( ~n6505 & n18792 ) | ( n18666 & n18792 ) ;
  assign n18795 = n18794 ^ n18793 ^ n8708 ;
  assign n18796 = n18069 ^ n10621 ^ n363 ;
  assign n18797 = ( n1136 & n1171 ) | ( n1136 & ~n6400 ) | ( n1171 & ~n6400 ) ;
  assign n18798 = n18797 ^ n7124 ^ n3010 ;
  assign n18799 = ( n8358 & ~n12576 ) | ( n8358 & n18798 ) | ( ~n12576 & n18798 ) ;
  assign n18800 = ( n5742 & n8397 ) | ( n5742 & n18799 ) | ( n8397 & n18799 ) ;
  assign n18801 = n8191 ^ n2070 ^ n1952 ;
  assign n18802 = ( n7360 & n14755 ) | ( n7360 & n18801 ) | ( n14755 & n18801 ) ;
  assign n18803 = n12734 ^ n6333 ^ n719 ;
  assign n18804 = ( n5715 & ~n18802 ) | ( n5715 & n18803 ) | ( ~n18802 & n18803 ) ;
  assign n18806 = ( n3231 & ~n10909 ) | ( n3231 & n16610 ) | ( ~n10909 & n16610 ) ;
  assign n18805 = ( ~n4067 & n4473 ) | ( ~n4067 & n11743 ) | ( n4473 & n11743 ) ;
  assign n18807 = n18806 ^ n18805 ^ n4867 ;
  assign n18808 = ( ~n4100 & n6614 ) | ( ~n4100 & n6633 ) | ( n6614 & n6633 ) ;
  assign n18809 = ( n3943 & n5867 ) | ( n3943 & ~n17717 ) | ( n5867 & ~n17717 ) ;
  assign n18810 = ( n10221 & n18808 ) | ( n10221 & ~n18809 ) | ( n18808 & ~n18809 ) ;
  assign n18811 = n18810 ^ n1937 ^ n697 ;
  assign n18812 = ( n3523 & n13722 ) | ( n3523 & n18811 ) | ( n13722 & n18811 ) ;
  assign n18813 = n12242 ^ n7884 ^ n4160 ;
  assign n18814 = ( n4470 & ~n11374 ) | ( n4470 & n13152 ) | ( ~n11374 & n13152 ) ;
  assign n18815 = ( x38 & n3422 ) | ( x38 & ~n18814 ) | ( n3422 & ~n18814 ) ;
  assign n18816 = n8734 ^ n7614 ^ n2259 ;
  assign n18817 = n18816 ^ n9791 ^ n6113 ;
  assign n18818 = n18817 ^ n7969 ^ n5779 ;
  assign n18819 = ( n1886 & n1988 ) | ( n1886 & n2733 ) | ( n1988 & n2733 ) ;
  assign n18820 = ( ~n4387 & n6281 ) | ( ~n4387 & n8334 ) | ( n6281 & n8334 ) ;
  assign n18821 = n18820 ^ n8981 ^ n5311 ;
  assign n18822 = ( n7374 & n18819 ) | ( n7374 & n18821 ) | ( n18819 & n18821 ) ;
  assign n18823 = ( n1162 & n2450 ) | ( n1162 & n6895 ) | ( n2450 & n6895 ) ;
  assign n18824 = ( n2766 & n7466 ) | ( n2766 & n11187 ) | ( n7466 & n11187 ) ;
  assign n18825 = ( n4999 & n6846 ) | ( n4999 & n18824 ) | ( n6846 & n18824 ) ;
  assign n18826 = ( n11506 & ~n18823 ) | ( n11506 & n18825 ) | ( ~n18823 & n18825 ) ;
  assign n18827 = ( n2861 & n17920 ) | ( n2861 & n18826 ) | ( n17920 & n18826 ) ;
  assign n18828 = ( n7435 & n9775 ) | ( n7435 & n11504 ) | ( n9775 & n11504 ) ;
  assign n18830 = n8616 ^ n4588 ^ n4232 ;
  assign n18831 = ( ~n2492 & n15773 ) | ( ~n2492 & n18830 ) | ( n15773 & n18830 ) ;
  assign n18829 = ( n3223 & n15888 ) | ( n3223 & n16930 ) | ( n15888 & n16930 ) ;
  assign n18832 = n18831 ^ n18829 ^ n16805 ;
  assign n18833 = ( n2494 & n5342 ) | ( n2494 & n10605 ) | ( n5342 & n10605 ) ;
  assign n18834 = ( n12916 & ~n15172 ) | ( n12916 & n18833 ) | ( ~n15172 & n18833 ) ;
  assign n18835 = n18834 ^ n8981 ^ n3100 ;
  assign n18836 = ( n2499 & n2506 ) | ( n2499 & n5556 ) | ( n2506 & n5556 ) ;
  assign n18837 = ( n3984 & ~n4396 ) | ( n3984 & n7770 ) | ( ~n4396 & n7770 ) ;
  assign n18838 = ( n1573 & ~n11654 ) | ( n1573 & n12265 ) | ( ~n11654 & n12265 ) ;
  assign n18839 = ( n18836 & n18837 ) | ( n18836 & n18838 ) | ( n18837 & n18838 ) ;
  assign n18846 = n6884 ^ n2384 ^ n587 ;
  assign n18843 = n8030 ^ n5823 ^ n1072 ;
  assign n18844 = ( n4544 & n8661 ) | ( n4544 & ~n18843 ) | ( n8661 & ~n18843 ) ;
  assign n18845 = ( n9651 & n15135 ) | ( n9651 & ~n18844 ) | ( n15135 & ~n18844 ) ;
  assign n18841 = n12541 ^ n4027 ^ n323 ;
  assign n18840 = n15271 ^ n6654 ^ n4963 ;
  assign n18842 = n18841 ^ n18840 ^ n15277 ;
  assign n18847 = n18846 ^ n18845 ^ n18842 ;
  assign n18848 = n18847 ^ n8189 ^ n2358 ;
  assign n18849 = n6362 ^ n5311 ^ n2760 ;
  assign n18853 = ( x116 & n5123 ) | ( x116 & ~n7343 ) | ( n5123 & ~n7343 ) ;
  assign n18850 = n7990 ^ n6966 ^ n645 ;
  assign n18851 = n18850 ^ n10072 ^ n1894 ;
  assign n18852 = n18851 ^ n17466 ^ n5719 ;
  assign n18854 = n18853 ^ n18852 ^ n18281 ;
  assign n18855 = n18854 ^ n6046 ^ n730 ;
  assign n18856 = ( ~n8072 & n18275 ) | ( ~n8072 & n18855 ) | ( n18275 & n18855 ) ;
  assign n18858 = n10350 ^ n4182 ^ n2299 ;
  assign n18859 = n18858 ^ n10088 ^ n4169 ;
  assign n18857 = n16364 ^ n15685 ^ n9698 ;
  assign n18860 = n18859 ^ n18857 ^ n1733 ;
  assign n18861 = ( x34 & n6789 ) | ( x34 & n18860 ) | ( n6789 & n18860 ) ;
  assign n18862 = ( n4586 & n10006 ) | ( n4586 & n11400 ) | ( n10006 & n11400 ) ;
  assign n18863 = n18862 ^ n14698 ^ n9008 ;
  assign n18864 = ( ~n3737 & n18861 ) | ( ~n3737 & n18863 ) | ( n18861 & n18863 ) ;
  assign n18869 = n8417 ^ n4280 ^ n1041 ;
  assign n18870 = ( n1514 & n9945 ) | ( n1514 & n18869 ) | ( n9945 & n18869 ) ;
  assign n18866 = n10446 ^ n7264 ^ n4782 ;
  assign n18867 = ( ~n718 & n3322 ) | ( ~n718 & n18866 ) | ( n3322 & n18866 ) ;
  assign n18865 = ( n1308 & n5236 ) | ( n1308 & ~n14111 ) | ( n5236 & ~n14111 ) ;
  assign n18868 = n18867 ^ n18865 ^ n3756 ;
  assign n18871 = n18870 ^ n18868 ^ n11320 ;
  assign n18872 = ( ~n4184 & n6295 ) | ( ~n4184 & n10476 ) | ( n6295 & n10476 ) ;
  assign n18873 = n18872 ^ n11702 ^ n292 ;
  assign n18874 = ( n636 & n18871 ) | ( n636 & n18873 ) | ( n18871 & n18873 ) ;
  assign n18875 = ( ~n685 & n2737 ) | ( ~n685 & n11485 ) | ( n2737 & n11485 ) ;
  assign n18876 = ( ~n1275 & n12373 ) | ( ~n1275 & n18875 ) | ( n12373 & n18875 ) ;
  assign n18877 = ( ~n3655 & n16950 ) | ( ~n3655 & n18876 ) | ( n16950 & n18876 ) ;
  assign n18879 = ( n1925 & ~n3064 ) | ( n1925 & n5307 ) | ( ~n3064 & n5307 ) ;
  assign n18878 = ( n1131 & n8698 ) | ( n1131 & n12247 ) | ( n8698 & n12247 ) ;
  assign n18880 = n18879 ^ n18878 ^ n15811 ;
  assign n18881 = ( n1143 & n2200 ) | ( n1143 & n7428 ) | ( n2200 & n7428 ) ;
  assign n18885 = n3490 ^ n2247 ^ n730 ;
  assign n18882 = n13761 ^ n6517 ^ n3342 ;
  assign n18883 = n18882 ^ n4117 ^ n1036 ;
  assign n18884 = n18883 ^ n7331 ^ n256 ;
  assign n18886 = n18885 ^ n18884 ^ n14823 ;
  assign n18887 = ( n9600 & n12177 ) | ( n9600 & n12545 ) | ( n12177 & n12545 ) ;
  assign n18888 = n16361 ^ n9380 ^ n3518 ;
  assign n18889 = n18888 ^ n18559 ^ n11645 ;
  assign n18890 = n10423 ^ n8667 ^ n3669 ;
  assign n18891 = ( n3157 & n18875 ) | ( n3157 & ~n18890 ) | ( n18875 & ~n18890 ) ;
  assign n18892 = ( n4026 & ~n17786 ) | ( n4026 & n18891 ) | ( ~n17786 & n18891 ) ;
  assign n18894 = n6021 ^ n5106 ^ n4242 ;
  assign n18895 = ( n3885 & n8230 ) | ( n3885 & n18894 ) | ( n8230 & n18894 ) ;
  assign n18893 = n5471 ^ n3295 ^ n935 ;
  assign n18896 = n18895 ^ n18893 ^ n4095 ;
  assign n18897 = ( ~n2384 & n5082 ) | ( ~n2384 & n18896 ) | ( n5082 & n18896 ) ;
  assign n18898 = n15367 ^ n11702 ^ n1716 ;
  assign n18899 = n13417 ^ n10724 ^ n8770 ;
  assign n18900 = ( n13329 & n17931 ) | ( n13329 & n18899 ) | ( n17931 & n18899 ) ;
  assign n18901 = n12651 ^ n8863 ^ n423 ;
  assign n18902 = n17822 ^ n17621 ^ n392 ;
  assign n18903 = ( n13466 & ~n16287 ) | ( n13466 & n18902 ) | ( ~n16287 & n18902 ) ;
  assign n18904 = n6302 ^ n3103 ^ n1101 ;
  assign n18905 = n18904 ^ n16337 ^ n13272 ;
  assign n18909 = n15519 ^ n14173 ^ n11654 ;
  assign n18910 = ( ~n6513 & n9294 ) | ( ~n6513 & n18909 ) | ( n9294 & n18909 ) ;
  assign n18908 = n18836 ^ n10471 ^ n2549 ;
  assign n18906 = n12738 ^ n6848 ^ n4387 ;
  assign n18907 = ( ~n571 & n2923 ) | ( ~n571 & n18906 ) | ( n2923 & n18906 ) ;
  assign n18911 = n18910 ^ n18908 ^ n18907 ;
  assign n18912 = ( n2363 & n4778 ) | ( n2363 & ~n8690 ) | ( n4778 & ~n8690 ) ;
  assign n18913 = ( n1060 & n9423 ) | ( n1060 & ~n11044 ) | ( n9423 & ~n11044 ) ;
  assign n18914 = ( n7716 & n12704 ) | ( n7716 & ~n18913 ) | ( n12704 & ~n18913 ) ;
  assign n18915 = ( n2676 & ~n3318 ) | ( n2676 & n17660 ) | ( ~n3318 & n17660 ) ;
  assign n18917 = n4484 ^ n3867 ^ n2920 ;
  assign n18916 = ( ~n2565 & n13814 ) | ( ~n2565 & n16620 ) | ( n13814 & n16620 ) ;
  assign n18918 = n18917 ^ n18916 ^ n8621 ;
  assign n18919 = n18918 ^ n10596 ^ n1247 ;
  assign n18920 = ( n5483 & n10066 ) | ( n5483 & n16044 ) | ( n10066 & n16044 ) ;
  assign n18921 = n18667 ^ n16290 ^ n5623 ;
  assign n18922 = ( n9127 & ~n18920 ) | ( n9127 & n18921 ) | ( ~n18920 & n18921 ) ;
  assign n18923 = ( ~n4280 & n8571 ) | ( ~n4280 & n17603 ) | ( n8571 & n17603 ) ;
  assign n18924 = n11343 ^ n9106 ^ n3331 ;
  assign n18925 = ( ~n10084 & n18572 ) | ( ~n10084 & n18924 ) | ( n18572 & n18924 ) ;
  assign n18926 = ( n3399 & n13914 ) | ( n3399 & ~n14198 ) | ( n13914 & ~n14198 ) ;
  assign n18927 = ( n347 & n4744 ) | ( n347 & ~n17799 ) | ( n4744 & ~n17799 ) ;
  assign n18928 = n18927 ^ n9992 ^ n1203 ;
  assign n18931 = n13194 ^ n7964 ^ n5853 ;
  assign n18932 = n18931 ^ n8905 ^ n3637 ;
  assign n18929 = n6652 ^ n3849 ^ n836 ;
  assign n18930 = n18929 ^ n7078 ^ n655 ;
  assign n18933 = n18932 ^ n18930 ^ n4130 ;
  assign n18934 = n16312 ^ n5035 ^ n3305 ;
  assign n18935 = n18934 ^ n17503 ^ n8622 ;
  assign n18940 = n5457 ^ n2741 ^ n509 ;
  assign n18936 = ( n5608 & ~n11692 ) | ( n5608 & n13951 ) | ( ~n11692 & n13951 ) ;
  assign n18937 = ( n2264 & ~n12638 ) | ( n2264 & n18936 ) | ( ~n12638 & n18936 ) ;
  assign n18938 = n18937 ^ n15936 ^ n8067 ;
  assign n18939 = n18938 ^ n16693 ^ n15353 ;
  assign n18941 = n18940 ^ n18939 ^ n3774 ;
  assign n18946 = ( ~n2210 & n7197 ) | ( ~n2210 & n16711 ) | ( n7197 & n16711 ) ;
  assign n18944 = ( n3879 & ~n6293 ) | ( n3879 & n16204 ) | ( ~n6293 & n16204 ) ;
  assign n18942 = ( n2029 & n2973 ) | ( n2029 & n6616 ) | ( n2973 & n6616 ) ;
  assign n18943 = ( ~n2207 & n11737 ) | ( ~n2207 & n18942 ) | ( n11737 & n18942 ) ;
  assign n18945 = n18944 ^ n18943 ^ n3450 ;
  assign n18947 = n18946 ^ n18945 ^ n13836 ;
  assign n18949 = n10976 ^ n9491 ^ n1557 ;
  assign n18948 = n13515 ^ n5817 ^ n4283 ;
  assign n18950 = n18949 ^ n18948 ^ n8574 ;
  assign n18951 = n8310 ^ n7076 ^ n515 ;
  assign n18952 = n18951 ^ n17846 ^ n12671 ;
  assign n18964 = n14768 ^ n11847 ^ n5538 ;
  assign n18955 = n11635 ^ n4099 ^ n3246 ;
  assign n18956 = n18955 ^ n5480 ^ x27 ;
  assign n18957 = ( ~n449 & n555 ) | ( ~n449 & n17473 ) | ( n555 & n17473 ) ;
  assign n18958 = ( n2039 & ~n3647 ) | ( n2039 & n5426 ) | ( ~n3647 & n5426 ) ;
  assign n18959 = n18958 ^ n18036 ^ n11704 ;
  assign n18960 = ( n3720 & n18957 ) | ( n3720 & n18959 ) | ( n18957 & n18959 ) ;
  assign n18961 = ( n1865 & n18956 ) | ( n1865 & n18960 ) | ( n18956 & n18960 ) ;
  assign n18953 = n15440 ^ n4665 ^ n1035 ;
  assign n18954 = ( ~n4375 & n14755 ) | ( ~n4375 & n18953 ) | ( n14755 & n18953 ) ;
  assign n18962 = n18961 ^ n18954 ^ n4284 ;
  assign n18963 = ( n2230 & ~n13745 ) | ( n2230 & n18962 ) | ( ~n13745 & n18962 ) ;
  assign n18965 = n18964 ^ n18963 ^ n16306 ;
  assign n18967 = n15000 ^ n9999 ^ n8234 ;
  assign n18966 = ( ~n6214 & n7336 ) | ( ~n6214 & n8824 ) | ( n7336 & n8824 ) ;
  assign n18968 = n18967 ^ n18966 ^ n1678 ;
  assign n18969 = ( n3498 & n6884 ) | ( n3498 & n7022 ) | ( n6884 & n7022 ) ;
  assign n18970 = n18969 ^ n13803 ^ n3942 ;
  assign n18971 = n18970 ^ n9928 ^ n6650 ;
  assign n18972 = n12338 ^ n6532 ^ n5956 ;
  assign n18973 = ( n160 & ~n6831 ) | ( n160 & n12708 ) | ( ~n6831 & n12708 ) ;
  assign n18974 = n16075 ^ n13404 ^ n8936 ;
  assign n18975 = ( n4954 & n18973 ) | ( n4954 & ~n18974 ) | ( n18973 & ~n18974 ) ;
  assign n18976 = n13338 ^ n9032 ^ n2948 ;
  assign n18981 = ( n6257 & ~n12059 ) | ( n6257 & n12228 ) | ( ~n12059 & n12228 ) ;
  assign n18979 = n2666 ^ n1221 ^ x94 ;
  assign n18980 = n18979 ^ n3840 ^ n3068 ;
  assign n18977 = ( n464 & n487 ) | ( n464 & ~n2218 ) | ( n487 & ~n2218 ) ;
  assign n18978 = n18977 ^ n8306 ^ n8166 ;
  assign n18982 = n18981 ^ n18980 ^ n18978 ;
  assign n18983 = ( n6611 & n9819 ) | ( n6611 & ~n11506 ) | ( n9819 & ~n11506 ) ;
  assign n18984 = ( n6320 & n13304 ) | ( n6320 & ~n18983 ) | ( n13304 & ~n18983 ) ;
  assign n18986 = n11642 ^ n10580 ^ n1048 ;
  assign n18985 = ( n1702 & ~n14909 ) | ( n1702 & n15068 ) | ( ~n14909 & n15068 ) ;
  assign n18987 = n18986 ^ n18985 ^ n8704 ;
  assign n18988 = ( n1322 & ~n1987 ) | ( n1322 & n4490 ) | ( ~n1987 & n4490 ) ;
  assign n18989 = ( n15746 & n15800 ) | ( n15746 & ~n18988 ) | ( n15800 & ~n18988 ) ;
  assign n18990 = ( n2201 & ~n3876 ) | ( n2201 & n12981 ) | ( ~n3876 & n12981 ) ;
  assign n18991 = ( n15433 & n18989 ) | ( n15433 & n18990 ) | ( n18989 & n18990 ) ;
  assign n18992 = n17114 ^ n8383 ^ n1401 ;
  assign n18993 = ( n1484 & n9581 ) | ( n1484 & n14011 ) | ( n9581 & n14011 ) ;
  assign n18994 = ( n5436 & n8718 ) | ( n5436 & n11834 ) | ( n8718 & n11834 ) ;
  assign n18995 = n11544 ^ n11238 ^ n921 ;
  assign n18996 = ( n4638 & ~n14931 ) | ( n4638 & n18995 ) | ( ~n14931 & n18995 ) ;
  assign n18997 = ( n7502 & ~n18994 ) | ( n7502 & n18996 ) | ( ~n18994 & n18996 ) ;
  assign n18998 = n18997 ^ n10816 ^ n9779 ;
  assign n18999 = ( n9264 & n11637 ) | ( n9264 & n15265 ) | ( n11637 & n15265 ) ;
  assign n19000 = n18999 ^ n11187 ^ n7331 ;
  assign n19001 = n19000 ^ n15153 ^ n13787 ;
  assign n19002 = n3655 ^ n1586 ^ n1081 ;
  assign n19003 = n19002 ^ n5089 ^ n3247 ;
  assign n19004 = n19003 ^ n12922 ^ n9788 ;
  assign n19005 = n13887 ^ n3204 ^ n1360 ;
  assign n19006 = n15605 ^ n6005 ^ n891 ;
  assign n19007 = ( n362 & n3756 ) | ( n362 & n12137 ) | ( n3756 & n12137 ) ;
  assign n19008 = ( n222 & ~n8234 ) | ( n222 & n19007 ) | ( ~n8234 & n19007 ) ;
  assign n19009 = ( n1528 & n3592 ) | ( n1528 & n18197 ) | ( n3592 & n18197 ) ;
  assign n19010 = ( n5634 & ~n8697 ) | ( n5634 & n14674 ) | ( ~n8697 & n14674 ) ;
  assign n19011 = ( ~n11042 & n12294 ) | ( ~n11042 & n19010 ) | ( n12294 & n19010 ) ;
  assign n19012 = n4188 ^ n2258 ^ n258 ;
  assign n19013 = ( ~n5954 & n6789 ) | ( ~n5954 & n19012 ) | ( n6789 & n19012 ) ;
  assign n19014 = ( n3278 & n3394 ) | ( n3278 & n19013 ) | ( n3394 & n19013 ) ;
  assign n19015 = ( n1127 & n17281 ) | ( n1127 & n19014 ) | ( n17281 & n19014 ) ;
  assign n19016 = ( ~n1246 & n8436 ) | ( ~n1246 & n14911 ) | ( n8436 & n14911 ) ;
  assign n19017 = n19016 ^ n12390 ^ n11849 ;
  assign n19018 = ( ~x112 & n330 ) | ( ~x112 & n8754 ) | ( n330 & n8754 ) ;
  assign n19019 = ( n202 & n745 ) | ( n202 & n19018 ) | ( n745 & n19018 ) ;
  assign n19020 = n11284 ^ n6562 ^ n3504 ;
  assign n19021 = n19020 ^ n10266 ^ n881 ;
  assign n19022 = ( ~n4717 & n7269 ) | ( ~n4717 & n7342 ) | ( n7269 & n7342 ) ;
  assign n19023 = n19022 ^ n3007 ^ x100 ;
  assign n19024 = n19023 ^ n16008 ^ n8649 ;
  assign n19025 = ( ~n6634 & n10417 ) | ( ~n6634 & n16055 ) | ( n10417 & n16055 ) ;
  assign n19026 = n19025 ^ n16224 ^ n3137 ;
  assign n19027 = n19026 ^ n18999 ^ n1203 ;
  assign n19028 = n16829 ^ n7185 ^ n1041 ;
  assign n19029 = ( n1352 & ~n18983 ) | ( n1352 & n19028 ) | ( ~n18983 & n19028 ) ;
  assign n19030 = ( n11005 & n11574 ) | ( n11005 & ~n19029 ) | ( n11574 & ~n19029 ) ;
  assign n19031 = n18358 ^ n10594 ^ n3636 ;
  assign n19032 = n13563 ^ n10274 ^ n4921 ;
  assign n19033 = n7920 ^ n5057 ^ n4062 ;
  assign n19034 = n19033 ^ n6466 ^ n1798 ;
  assign n19035 = ( n8930 & n16362 ) | ( n8930 & n19034 ) | ( n16362 & n19034 ) ;
  assign n19041 = ( n1821 & n6440 ) | ( n1821 & ~n7329 ) | ( n6440 & ~n7329 ) ;
  assign n19040 = ( n6761 & n12910 ) | ( n6761 & ~n17633 ) | ( n12910 & ~n17633 ) ;
  assign n19038 = ( n185 & n588 ) | ( n185 & ~n5177 ) | ( n588 & ~n5177 ) ;
  assign n19036 = n12342 ^ n162 ^ x78 ;
  assign n19037 = ( ~n9268 & n13843 ) | ( ~n9268 & n19036 ) | ( n13843 & n19036 ) ;
  assign n19039 = n19038 ^ n19037 ^ n5648 ;
  assign n19042 = n19041 ^ n19040 ^ n19039 ;
  assign n19043 = ( n9628 & n16352 ) | ( n9628 & ~n17627 ) | ( n16352 & ~n17627 ) ;
  assign n19044 = ( n6692 & ~n10161 ) | ( n6692 & n19043 ) | ( ~n10161 & n19043 ) ;
  assign n19049 = ( n12229 & n14534 ) | ( n12229 & n14986 ) | ( n14534 & n14986 ) ;
  assign n19050 = n19049 ^ n13062 ^ n9499 ;
  assign n19047 = ( n3479 & n4721 ) | ( n3479 & ~n6381 ) | ( n4721 & ~n6381 ) ;
  assign n19048 = ( n4475 & n14960 ) | ( n4475 & ~n19047 ) | ( n14960 & ~n19047 ) ;
  assign n19045 = n10571 ^ n5674 ^ n4885 ;
  assign n19046 = n19045 ^ n18489 ^ n9811 ;
  assign n19051 = n19050 ^ n19048 ^ n19046 ;
  assign n19052 = ( ~n2142 & n5218 ) | ( ~n2142 & n14075 ) | ( n5218 & n14075 ) ;
  assign n19053 = ( n989 & n2717 ) | ( n989 & ~n8571 ) | ( n2717 & ~n8571 ) ;
  assign n19054 = ( n3235 & n4089 ) | ( n3235 & n19053 ) | ( n4089 & n19053 ) ;
  assign n19055 = ( n14306 & n19052 ) | ( n14306 & n19054 ) | ( n19052 & n19054 ) ;
  assign n19057 = ( ~n1158 & n7381 ) | ( ~n1158 & n11168 ) | ( n7381 & n11168 ) ;
  assign n19056 = ( n2074 & n2506 ) | ( n2074 & ~n3795 ) | ( n2506 & ~n3795 ) ;
  assign n19058 = n19057 ^ n19056 ^ n5976 ;
  assign n19059 = ( n14378 & ~n19055 ) | ( n14378 & n19058 ) | ( ~n19055 & n19058 ) ;
  assign n19060 = n17815 ^ n6501 ^ n6236 ;
  assign n19061 = ( ~n7003 & n11769 ) | ( ~n7003 & n19060 ) | ( n11769 & n19060 ) ;
  assign n19062 = n17606 ^ n8844 ^ n5152 ;
  assign n19066 = n2937 ^ n1065 ^ n865 ;
  assign n19064 = n12609 ^ n2627 ^ n597 ;
  assign n19065 = n19064 ^ n14432 ^ n2462 ;
  assign n19063 = ( ~n8029 & n9553 ) | ( ~n8029 & n17494 ) | ( n9553 & n17494 ) ;
  assign n19067 = n19066 ^ n19065 ^ n19063 ;
  assign n19068 = ( n842 & ~n13798 ) | ( n842 & n15154 ) | ( ~n13798 & n15154 ) ;
  assign n19069 = ( n566 & n3316 ) | ( n566 & n15868 ) | ( n3316 & n15868 ) ;
  assign n19070 = ( n826 & ~n6011 ) | ( n826 & n19069 ) | ( ~n6011 & n19069 ) ;
  assign n19071 = ( n5175 & ~n6079 ) | ( n5175 & n18434 ) | ( ~n6079 & n18434 ) ;
  assign n19072 = ( n5082 & ~n6092 ) | ( n5082 & n18596 ) | ( ~n6092 & n18596 ) ;
  assign n19073 = ( n9437 & n19071 ) | ( n9437 & n19072 ) | ( n19071 & n19072 ) ;
  assign n19074 = ( n1512 & n4439 ) | ( n1512 & n5604 ) | ( n4439 & n5604 ) ;
  assign n19075 = ( n799 & ~n1483 ) | ( n799 & n1804 ) | ( ~n1483 & n1804 ) ;
  assign n19076 = n19075 ^ n17133 ^ n6615 ;
  assign n19077 = ( ~n14899 & n17727 ) | ( ~n14899 & n19076 ) | ( n17727 & n19076 ) ;
  assign n19081 = n16608 ^ n12973 ^ n12240 ;
  assign n19082 = ( n2481 & n3018 ) | ( n2481 & n19081 ) | ( n3018 & n19081 ) ;
  assign n19083 = ( ~n8303 & n14190 ) | ( ~n8303 & n19082 ) | ( n14190 & n19082 ) ;
  assign n19078 = ( n4181 & n11509 ) | ( n4181 & ~n12024 ) | ( n11509 & ~n12024 ) ;
  assign n19079 = ( n6752 & ~n12172 ) | ( n6752 & n19078 ) | ( ~n12172 & n19078 ) ;
  assign n19080 = ( ~n261 & n11513 ) | ( ~n261 & n19079 ) | ( n11513 & n19079 ) ;
  assign n19084 = n19083 ^ n19080 ^ n6111 ;
  assign n19085 = ( ~n3473 & n6445 ) | ( ~n3473 & n12213 ) | ( n6445 & n12213 ) ;
  assign n19086 = n12549 ^ n8694 ^ n412 ;
  assign n19087 = ( n10071 & n11429 ) | ( n10071 & ~n15865 ) | ( n11429 & ~n15865 ) ;
  assign n19088 = ( n12424 & n19086 ) | ( n12424 & n19087 ) | ( n19086 & n19087 ) ;
  assign n19089 = ( n15567 & ~n19085 ) | ( n15567 & n19088 ) | ( ~n19085 & n19088 ) ;
  assign n19090 = ( n355 & n2483 ) | ( n355 & ~n17161 ) | ( n2483 & ~n17161 ) ;
  assign n19091 = n10517 ^ n5803 ^ n4733 ;
  assign n19092 = n19091 ^ n14350 ^ n2269 ;
  assign n19093 = ( n754 & n5384 ) | ( n754 & n10713 ) | ( n5384 & n10713 ) ;
  assign n19094 = n15606 ^ n5136 ^ n2179 ;
  assign n19095 = ( n13178 & n13219 ) | ( n13178 & n19094 ) | ( n13219 & n19094 ) ;
  assign n19096 = ( n1045 & ~n3029 ) | ( n1045 & n18219 ) | ( ~n3029 & n18219 ) ;
  assign n19097 = n13583 ^ n12098 ^ n5489 ;
  assign n19098 = ( n3763 & n19096 ) | ( n3763 & ~n19097 ) | ( n19096 & ~n19097 ) ;
  assign n19099 = ( ~n1630 & n4226 ) | ( ~n1630 & n7814 ) | ( n4226 & n7814 ) ;
  assign n19100 = ( ~n4350 & n6062 ) | ( ~n4350 & n19099 ) | ( n6062 & n19099 ) ;
  assign n19101 = ( ~n8951 & n18476 ) | ( ~n8951 & n19100 ) | ( n18476 & n19100 ) ;
  assign n19102 = ( n11005 & n14026 ) | ( n11005 & ~n15781 ) | ( n14026 & ~n15781 ) ;
  assign n19103 = n8544 ^ n8167 ^ n7036 ;
  assign n19104 = ( n2512 & n4202 ) | ( n2512 & n19103 ) | ( n4202 & n19103 ) ;
  assign n19105 = ( n3927 & n5122 ) | ( n3927 & n19104 ) | ( n5122 & n19104 ) ;
  assign n19112 = n16151 ^ n5801 ^ n5644 ;
  assign n19109 = ( n488 & ~n1295 ) | ( n488 & n2110 ) | ( ~n1295 & n2110 ) ;
  assign n19110 = ( n5425 & ~n7598 ) | ( n5425 & n12028 ) | ( ~n7598 & n12028 ) ;
  assign n19111 = ( n5644 & n19109 ) | ( n5644 & ~n19110 ) | ( n19109 & ~n19110 ) ;
  assign n19113 = n19112 ^ n19111 ^ n6624 ;
  assign n19106 = ( n2092 & ~n2764 ) | ( n2092 & n8586 ) | ( ~n2764 & n8586 ) ;
  assign n19107 = ( n8162 & ~n9496 ) | ( n8162 & n19106 ) | ( ~n9496 & n19106 ) ;
  assign n19108 = n19107 ^ n13430 ^ n4786 ;
  assign n19114 = n19113 ^ n19108 ^ n12682 ;
  assign n19118 = ( n2002 & n4388 ) | ( n2002 & ~n8537 ) | ( n4388 & ~n8537 ) ;
  assign n19115 = ( n2141 & n4478 ) | ( n2141 & ~n10057 ) | ( n4478 & ~n10057 ) ;
  assign n19116 = ( n6388 & ~n9091 ) | ( n6388 & n19115 ) | ( ~n9091 & n19115 ) ;
  assign n19117 = n19116 ^ n15692 ^ n2305 ;
  assign n19119 = n19118 ^ n19117 ^ n12890 ;
  assign n19120 = n17315 ^ n9640 ^ n1180 ;
  assign n19121 = ( ~n11010 & n13170 ) | ( ~n11010 & n19120 ) | ( n13170 & n19120 ) ;
  assign n19139 = ( n668 & ~n10334 ) | ( n668 & n11130 ) | ( ~n10334 & n11130 ) ;
  assign n19140 = n19139 ^ n12347 ^ n7650 ;
  assign n19137 = ( n5016 & n7565 ) | ( n5016 & n8772 ) | ( n7565 & n8772 ) ;
  assign n19135 = n13051 ^ n11645 ^ n1464 ;
  assign n19136 = ( n8795 & ~n15905 ) | ( n8795 & n19135 ) | ( ~n15905 & n19135 ) ;
  assign n19138 = n19137 ^ n19136 ^ n4298 ;
  assign n19122 = n17793 ^ n12625 ^ n1869 ;
  assign n19123 = ( n4805 & n12544 ) | ( n4805 & n15245 ) | ( n12544 & n15245 ) ;
  assign n19124 = n10690 ^ n9773 ^ n2042 ;
  assign n19125 = ( ~n4840 & n6545 ) | ( ~n4840 & n9026 ) | ( n6545 & n9026 ) ;
  assign n19126 = ( n19123 & ~n19124 ) | ( n19123 & n19125 ) | ( ~n19124 & n19125 ) ;
  assign n19127 = n19126 ^ n18029 ^ n11126 ;
  assign n19128 = n8095 ^ n6898 ^ n4665 ;
  assign n19129 = n19128 ^ n5665 ^ n380 ;
  assign n19130 = n19129 ^ n10736 ^ n9306 ;
  assign n19131 = ( n6548 & ~n11875 ) | ( n6548 & n19130 ) | ( ~n11875 & n19130 ) ;
  assign n19132 = n19131 ^ n6521 ^ n6518 ;
  assign n19133 = n19132 ^ n10353 ^ n484 ;
  assign n19134 = ( n19122 & n19127 ) | ( n19122 & n19133 ) | ( n19127 & n19133 ) ;
  assign n19141 = n19140 ^ n19138 ^ n19134 ;
  assign n19144 = ( n1815 & n5159 ) | ( n1815 & n9503 ) | ( n5159 & n9503 ) ;
  assign n19142 = ( ~n673 & n2705 ) | ( ~n673 & n6618 ) | ( n2705 & n6618 ) ;
  assign n19143 = n19142 ^ n3992 ^ n900 ;
  assign n19145 = n19144 ^ n19143 ^ n7884 ;
  assign n19147 = n8621 ^ n2163 ^ n1663 ;
  assign n19148 = ( x79 & ~n677 ) | ( x79 & n15691 ) | ( ~n677 & n15691 ) ;
  assign n19149 = ( ~n1652 & n19147 ) | ( ~n1652 & n19148 ) | ( n19147 & n19148 ) ;
  assign n19146 = n15698 ^ n4816 ^ n1430 ;
  assign n19150 = n19149 ^ n19146 ^ n13959 ;
  assign n19157 = n12908 ^ n7363 ^ n5387 ;
  assign n19151 = n17484 ^ n8298 ^ n2751 ;
  assign n19152 = n12795 ^ n11306 ^ n1295 ;
  assign n19153 = ( ~n3984 & n11835 ) | ( ~n3984 & n19152 ) | ( n11835 & n19152 ) ;
  assign n19154 = n19153 ^ n12148 ^ n5073 ;
  assign n19155 = n19154 ^ n15279 ^ n12419 ;
  assign n19156 = ( n12135 & ~n19151 ) | ( n12135 & n19155 ) | ( ~n19151 & n19155 ) ;
  assign n19158 = n19157 ^ n19156 ^ n1863 ;
  assign n19159 = n18041 ^ n9833 ^ n3312 ;
  assign n19162 = n3627 ^ n1657 ^ n924 ;
  assign n19163 = n19162 ^ n8283 ^ n1260 ;
  assign n19164 = ( n6891 & n7460 ) | ( n6891 & ~n19163 ) | ( n7460 & ~n19163 ) ;
  assign n19161 = n3424 ^ n2722 ^ n2034 ;
  assign n19165 = n19164 ^ n19161 ^ n10308 ;
  assign n19160 = ( n2280 & n6399 ) | ( n2280 & ~n16440 ) | ( n6399 & ~n16440 ) ;
  assign n19166 = n19165 ^ n19160 ^ n17620 ;
  assign n19167 = n19166 ^ n7893 ^ n7325 ;
  assign n19168 = n18222 ^ n15405 ^ n5243 ;
  assign n19169 = ( n5164 & n8247 ) | ( n5164 & ~n19168 ) | ( n8247 & ~n19168 ) ;
  assign n19170 = n19169 ^ n15867 ^ n13129 ;
  assign n19171 = n19170 ^ n17226 ^ n2450 ;
  assign n19172 = ( ~n3590 & n10077 ) | ( ~n3590 & n11581 ) | ( n10077 & n11581 ) ;
  assign n19173 = n19172 ^ n12294 ^ n3042 ;
  assign n19174 = n6974 ^ n2706 ^ n1860 ;
  assign n19175 = ( n6230 & ~n9299 ) | ( n6230 & n19174 ) | ( ~n9299 & n19174 ) ;
  assign n19176 = n19175 ^ n17656 ^ n5942 ;
  assign n19177 = ( n1659 & n4369 ) | ( n1659 & n15540 ) | ( n4369 & n15540 ) ;
  assign n19179 = ( ~n3290 & n5647 ) | ( ~n3290 & n7725 ) | ( n5647 & n7725 ) ;
  assign n19180 = ( n2415 & n13301 ) | ( n2415 & ~n19179 ) | ( n13301 & ~n19179 ) ;
  assign n19178 = ( n6585 & n7214 ) | ( n6585 & n12040 ) | ( n7214 & n12040 ) ;
  assign n19181 = n19180 ^ n19178 ^ n5264 ;
  assign n19182 = n17166 ^ n3641 ^ n1471 ;
  assign n19183 = n16526 ^ n14860 ^ n8138 ;
  assign n19184 = ( n12135 & n19085 ) | ( n12135 & ~n19183 ) | ( n19085 & ~n19183 ) ;
  assign n19185 = ( n6878 & n19182 ) | ( n6878 & ~n19184 ) | ( n19182 & ~n19184 ) ;
  assign n19186 = n15326 ^ n8712 ^ n424 ;
  assign n19187 = ( n5811 & ~n15695 ) | ( n5811 & n18819 ) | ( ~n15695 & n18819 ) ;
  assign n19188 = ( ~n15872 & n19186 ) | ( ~n15872 & n19187 ) | ( n19186 & n19187 ) ;
  assign n19189 = ( n2229 & n11716 ) | ( n2229 & ~n13558 ) | ( n11716 & ~n13558 ) ;
  assign n19194 = ( n1514 & n3291 ) | ( n1514 & n13862 ) | ( n3291 & n13862 ) ;
  assign n19190 = n7407 ^ n3826 ^ n2366 ;
  assign n19191 = n19190 ^ n4671 ^ n1458 ;
  assign n19192 = ( ~n3492 & n9148 ) | ( ~n3492 & n19191 ) | ( n9148 & n19191 ) ;
  assign n19193 = n19192 ^ n6206 ^ n5170 ;
  assign n19195 = n19194 ^ n19193 ^ n14009 ;
  assign n19196 = n10589 ^ n6256 ^ n3765 ;
  assign n19198 = ( n3947 & ~n5224 ) | ( n3947 & n15435 ) | ( ~n5224 & n15435 ) ;
  assign n19197 = n13168 ^ n6959 ^ n4029 ;
  assign n19199 = n19198 ^ n19197 ^ n5024 ;
  assign n19200 = n19199 ^ n7156 ^ n7028 ;
  assign n19201 = ( x2 & n852 ) | ( x2 & n9249 ) | ( n852 & n9249 ) ;
  assign n19202 = ( n12347 & ~n19200 ) | ( n12347 & n19201 ) | ( ~n19200 & n19201 ) ;
  assign n19203 = ( ~n9623 & n19196 ) | ( ~n9623 & n19202 ) | ( n19196 & n19202 ) ;
  assign n19204 = n10734 ^ n9852 ^ n6107 ;
  assign n19205 = ( ~n8532 & n11393 ) | ( ~n8532 & n19204 ) | ( n11393 & n19204 ) ;
  assign n19206 = ( ~n6696 & n15261 ) | ( ~n6696 & n18615 ) | ( n15261 & n18615 ) ;
  assign n19208 = ( ~n3186 & n12556 ) | ( ~n3186 & n15470 ) | ( n12556 & n15470 ) ;
  assign n19207 = ( ~n2338 & n4076 ) | ( ~n2338 & n10969 ) | ( n4076 & n10969 ) ;
  assign n19209 = n19208 ^ n19207 ^ n16393 ;
  assign n19210 = n19209 ^ n2167 ^ n1347 ;
  assign n19211 = ( n4195 & ~n10704 ) | ( n4195 & n12146 ) | ( ~n10704 & n12146 ) ;
  assign n19212 = n19211 ^ n7264 ^ n2138 ;
  assign n19213 = n18509 ^ n6502 ^ n1491 ;
  assign n19214 = ( n12167 & ~n12921 ) | ( n12167 & n19213 ) | ( ~n12921 & n19213 ) ;
  assign n19215 = ( ~n4368 & n10397 ) | ( ~n4368 & n14328 ) | ( n10397 & n14328 ) ;
  assign n19216 = n4406 ^ n3704 ^ n2410 ;
  assign n19217 = n19216 ^ n12064 ^ n5726 ;
  assign n19218 = ( n8005 & n8112 ) | ( n8005 & n12824 ) | ( n8112 & n12824 ) ;
  assign n19219 = ( n8565 & n9392 ) | ( n8565 & ~n19218 ) | ( n9392 & ~n19218 ) ;
  assign n19220 = n12821 ^ n10795 ^ n3802 ;
  assign n19221 = n13251 ^ n11964 ^ n6838 ;
  assign n19222 = ( ~n10878 & n16243 ) | ( ~n10878 & n19221 ) | ( n16243 & n19221 ) ;
  assign n19223 = ( n8558 & n10575 ) | ( n8558 & ~n19222 ) | ( n10575 & ~n19222 ) ;
  assign n19226 = n3747 ^ n2780 ^ n2722 ;
  assign n19227 = n19226 ^ n16444 ^ n15063 ;
  assign n19225 = n9139 ^ n2198 ^ n929 ;
  assign n19224 = ( ~n305 & n3314 ) | ( ~n305 & n13479 ) | ( n3314 & n13479 ) ;
  assign n19228 = n19227 ^ n19225 ^ n19224 ;
  assign n19229 = ( n13055 & ~n19223 ) | ( n13055 & n19228 ) | ( ~n19223 & n19228 ) ;
  assign n19230 = ( n2213 & n4944 ) | ( n2213 & ~n11546 ) | ( n4944 & ~n11546 ) ;
  assign n19231 = ( n4530 & n6024 ) | ( n4530 & n19230 ) | ( n6024 & n19230 ) ;
  assign n19232 = ( n2990 & n4765 ) | ( n2990 & ~n15998 ) | ( n4765 & ~n15998 ) ;
  assign n19233 = ( n18270 & n18519 ) | ( n18270 & n19232 ) | ( n18519 & n19232 ) ;
  assign n19235 = n18679 ^ n13233 ^ n3434 ;
  assign n19236 = ( n7255 & ~n11707 ) | ( n7255 & n19235 ) | ( ~n11707 & n19235 ) ;
  assign n19234 = n11320 ^ n7418 ^ n7273 ;
  assign n19237 = n19236 ^ n19234 ^ n3973 ;
  assign n19238 = n19237 ^ n4994 ^ n1747 ;
  assign n19239 = n14607 ^ n8801 ^ n6666 ;
  assign n19240 = ( n766 & n11079 ) | ( n766 & n19085 ) | ( n11079 & n19085 ) ;
  assign n19241 = n19240 ^ n10962 ^ n7507 ;
  assign n19242 = n16617 ^ n13289 ^ n3635 ;
  assign n19243 = ( n783 & n17264 ) | ( n783 & ~n18212 ) | ( n17264 & ~n18212 ) ;
  assign n19244 = ( ~n6708 & n19242 ) | ( ~n6708 & n19243 ) | ( n19242 & n19243 ) ;
  assign n19245 = n2888 ^ n634 ^ n451 ;
  assign n19246 = n19245 ^ n12824 ^ n6999 ;
  assign n19247 = ( n6692 & n9360 ) | ( n6692 & ~n19246 ) | ( n9360 & ~n19246 ) ;
  assign n19248 = n7226 ^ n2394 ^ n1793 ;
  assign n19249 = n19248 ^ n8054 ^ n1302 ;
  assign n19250 = ( n12233 & n19247 ) | ( n12233 & n19249 ) | ( n19247 & n19249 ) ;
  assign n19251 = n12808 ^ n8327 ^ n7877 ;
  assign n19252 = ( n1441 & n10623 ) | ( n1441 & ~n17807 ) | ( n10623 & ~n17807 ) ;
  assign n19253 = ( n3205 & n17582 ) | ( n3205 & ~n18152 ) | ( n17582 & ~n18152 ) ;
  assign n19254 = ( n11456 & n13734 ) | ( n11456 & n19253 ) | ( n13734 & n19253 ) ;
  assign n19255 = n19254 ^ n11695 ^ n2437 ;
  assign n19256 = ( n4344 & n17208 ) | ( n4344 & n19255 ) | ( n17208 & n19255 ) ;
  assign n19257 = n15295 ^ n12557 ^ n10469 ;
  assign n19258 = ( n1369 & n3772 ) | ( n1369 & ~n5219 ) | ( n3772 & ~n5219 ) ;
  assign n19259 = n19258 ^ n11922 ^ n1699 ;
  assign n19260 = n19259 ^ n14167 ^ n13775 ;
  assign n19261 = ( n1315 & ~n19257 ) | ( n1315 & n19260 ) | ( ~n19257 & n19260 ) ;
  assign n19263 = n6466 ^ n4353 ^ n2215 ;
  assign n19262 = n17371 ^ n14311 ^ n12606 ;
  assign n19264 = n19263 ^ n19262 ^ n3572 ;
  assign n19265 = n6830 ^ n5721 ^ n282 ;
  assign n19266 = n19265 ^ n3374 ^ n2864 ;
  assign n19267 = n19266 ^ n4582 ^ n1204 ;
  assign n19268 = ( n4722 & n12804 ) | ( n4722 & ~n15274 ) | ( n12804 & ~n15274 ) ;
  assign n19269 = ( n15667 & n19267 ) | ( n15667 & ~n19268 ) | ( n19267 & ~n19268 ) ;
  assign n19270 = ( n495 & n9876 ) | ( n495 & ~n19269 ) | ( n9876 & ~n19269 ) ;
  assign n19271 = n13467 ^ n5196 ^ n4360 ;
  assign n19272 = n8634 ^ n3804 ^ n1431 ;
  assign n19273 = ( n15134 & ~n15544 ) | ( n15134 & n19272 ) | ( ~n15544 & n19272 ) ;
  assign n19274 = n19273 ^ n17626 ^ n14938 ;
  assign n19275 = n19107 ^ n13063 ^ n7991 ;
  assign n19276 = ( n350 & ~n852 ) | ( n350 & n19275 ) | ( ~n852 & n19275 ) ;
  assign n19278 = n3187 ^ n2128 ^ x105 ;
  assign n19277 = ( n2552 & n4372 ) | ( n2552 & n5962 ) | ( n4372 & n5962 ) ;
  assign n19279 = n19278 ^ n19277 ^ n1945 ;
  assign n19280 = n19279 ^ n15019 ^ n3499 ;
  assign n19281 = ( ~n7312 & n19276 ) | ( ~n7312 & n19280 ) | ( n19276 & n19280 ) ;
  assign n19282 = ( x7 & n2363 ) | ( x7 & n4376 ) | ( n2363 & n4376 ) ;
  assign n19283 = ( n11612 & n15898 ) | ( n11612 & n19282 ) | ( n15898 & n19282 ) ;
  assign n19284 = ( n6746 & n7897 ) | ( n6746 & ~n19283 ) | ( n7897 & ~n19283 ) ;
  assign n19285 = ( ~n3424 & n8889 ) | ( ~n3424 & n9985 ) | ( n8889 & n9985 ) ;
  assign n19286 = ( n13023 & n19242 ) | ( n13023 & ~n19285 ) | ( n19242 & ~n19285 ) ;
  assign n19287 = n11856 ^ n8447 ^ n1532 ;
  assign n19288 = n19287 ^ n7616 ^ n1442 ;
  assign n19289 = n19288 ^ n8719 ^ n4095 ;
  assign n19290 = ( ~n4280 & n9556 ) | ( ~n4280 & n18402 ) | ( n9556 & n18402 ) ;
  assign n19291 = ( n7979 & n13786 ) | ( n7979 & n19290 ) | ( n13786 & n19290 ) ;
  assign n19292 = n19291 ^ n13223 ^ n1018 ;
  assign n19293 = n2571 ^ n1590 ^ n1234 ;
  assign n19294 = n19293 ^ n18944 ^ n3281 ;
  assign n19295 = n9963 ^ n5087 ^ n1205 ;
  assign n19296 = n9658 ^ n3515 ^ n1335 ;
  assign n19297 = n19296 ^ n10525 ^ n3150 ;
  assign n19298 = ( n2676 & n9724 ) | ( n2676 & n19297 ) | ( n9724 & n19297 ) ;
  assign n19299 = ( n6773 & ~n9301 ) | ( n6773 & n19298 ) | ( ~n9301 & n19298 ) ;
  assign n19300 = ( n9520 & n19295 ) | ( n9520 & ~n19299 ) | ( n19295 & ~n19299 ) ;
  assign n19301 = ( ~n867 & n4476 ) | ( ~n867 & n18439 ) | ( n4476 & n18439 ) ;
  assign n19302 = n16468 ^ n13757 ^ n145 ;
  assign n19303 = ( n1159 & n4151 ) | ( n1159 & ~n15501 ) | ( n4151 & ~n15501 ) ;
  assign n19304 = ( n13932 & n19302 ) | ( n13932 & n19303 ) | ( n19302 & n19303 ) ;
  assign n19309 = n10435 ^ n6822 ^ n6692 ;
  assign n19305 = ( n2778 & ~n6745 ) | ( n2778 & n8036 ) | ( ~n6745 & n8036 ) ;
  assign n19306 = ( ~n2664 & n2818 ) | ( ~n2664 & n5908 ) | ( n2818 & n5908 ) ;
  assign n19307 = ( n4143 & ~n9010 ) | ( n4143 & n18556 ) | ( ~n9010 & n18556 ) ;
  assign n19308 = ( n19305 & n19306 ) | ( n19305 & ~n19307 ) | ( n19306 & ~n19307 ) ;
  assign n19310 = n19309 ^ n19308 ^ n6066 ;
  assign n19311 = ( n9312 & n19304 ) | ( n9312 & n19310 ) | ( n19304 & n19310 ) ;
  assign n19312 = ( ~n536 & n1622 ) | ( ~n536 & n7287 ) | ( n1622 & n7287 ) ;
  assign n19313 = n19312 ^ n8331 ^ n2617 ;
  assign n19314 = ( n5884 & ~n10708 ) | ( n5884 & n19313 ) | ( ~n10708 & n19313 ) ;
  assign n19316 = ( ~n3348 & n3729 ) | ( ~n3348 & n19248 ) | ( n3729 & n19248 ) ;
  assign n19315 = n14118 ^ n4377 ^ n715 ;
  assign n19317 = n19316 ^ n19315 ^ n2821 ;
  assign n19318 = n19317 ^ n17278 ^ n5492 ;
  assign n19319 = ( n3857 & n19314 ) | ( n3857 & ~n19318 ) | ( n19314 & ~n19318 ) ;
  assign n19320 = n12906 ^ n4264 ^ n3325 ;
  assign n19321 = n19320 ^ n5659 ^ n2965 ;
  assign n19322 = ( n6792 & n14331 ) | ( n6792 & n19321 ) | ( n14331 & n19321 ) ;
  assign n19323 = n19322 ^ n12215 ^ n11439 ;
  assign n19324 = ( n441 & ~n5388 ) | ( n441 & n6952 ) | ( ~n5388 & n6952 ) ;
  assign n19325 = n19324 ^ n9978 ^ n8600 ;
  assign n19326 = ( ~n6031 & n8242 ) | ( ~n6031 & n19325 ) | ( n8242 & n19325 ) ;
  assign n19327 = n19326 ^ n2721 ^ n181 ;
  assign n19328 = ( ~n4299 & n5544 ) | ( ~n4299 & n13127 ) | ( n5544 & n13127 ) ;
  assign n19329 = n19328 ^ n5372 ^ n4866 ;
  assign n19330 = n17489 ^ n11737 ^ n9235 ;
  assign n19331 = n19330 ^ n17548 ^ n15495 ;
  assign n19332 = ( n9156 & ~n12840 ) | ( n9156 & n13909 ) | ( ~n12840 & n13909 ) ;
  assign n19333 = n16967 ^ n16077 ^ n4297 ;
  assign n19335 = ( n1095 & n7116 ) | ( n1095 & ~n7320 ) | ( n7116 & ~n7320 ) ;
  assign n19334 = ( n7143 & n17708 ) | ( n7143 & n17956 ) | ( n17708 & n17956 ) ;
  assign n19336 = n19335 ^ n19334 ^ n8857 ;
  assign n19337 = n18878 ^ n9674 ^ n4127 ;
  assign n19338 = n10693 ^ n5459 ^ n3511 ;
  assign n19339 = ( n7321 & n14089 ) | ( n7321 & ~n19338 ) | ( n14089 & ~n19338 ) ;
  assign n19340 = n19339 ^ n13030 ^ n1670 ;
  assign n19341 = ( n2023 & n12235 ) | ( n2023 & ~n14552 ) | ( n12235 & ~n14552 ) ;
  assign n19342 = n17720 ^ n5881 ^ n3697 ;
  assign n19343 = ( n1511 & n6830 ) | ( n1511 & ~n19342 ) | ( n6830 & ~n19342 ) ;
  assign n19344 = n19343 ^ n9841 ^ n5540 ;
  assign n19345 = ( n8248 & n11549 ) | ( n8248 & n19344 ) | ( n11549 & n19344 ) ;
  assign n19346 = ( n158 & ~n6045 ) | ( n158 & n17775 ) | ( ~n6045 & n17775 ) ;
  assign n19347 = n15722 ^ n14293 ^ n6011 ;
  assign n19348 = n19347 ^ n5857 ^ n672 ;
  assign n19349 = ( n739 & ~n5782 ) | ( n739 & n12790 ) | ( ~n5782 & n12790 ) ;
  assign n19350 = ( n3007 & n6833 ) | ( n3007 & ~n12018 ) | ( n6833 & ~n12018 ) ;
  assign n19351 = n19350 ^ n11635 ^ n4413 ;
  assign n19352 = ( n3315 & ~n5702 ) | ( n3315 & n18152 ) | ( ~n5702 & n18152 ) ;
  assign n19353 = n19352 ^ n7007 ^ n1352 ;
  assign n19354 = ( n19349 & ~n19351 ) | ( n19349 & n19353 ) | ( ~n19351 & n19353 ) ;
  assign n19355 = n6872 ^ n1619 ^ n1095 ;
  assign n19356 = ( n5351 & n7054 ) | ( n5351 & n19355 ) | ( n7054 & n19355 ) ;
  assign n19363 = ( ~n601 & n3013 ) | ( ~n601 & n13819 ) | ( n3013 & n13819 ) ;
  assign n19364 = n8598 ^ n6522 ^ n4392 ;
  assign n19365 = ( n7821 & n19363 ) | ( n7821 & ~n19364 ) | ( n19363 & ~n19364 ) ;
  assign n19357 = ( n4233 & ~n4616 ) | ( n4233 & n6120 ) | ( ~n4616 & n6120 ) ;
  assign n19358 = n8333 ^ n3837 ^ n588 ;
  assign n19359 = ( n7711 & n19357 ) | ( n7711 & ~n19358 ) | ( n19357 & ~n19358 ) ;
  assign n19360 = ( n6430 & n11673 ) | ( n6430 & ~n19359 ) | ( n11673 & ~n19359 ) ;
  assign n19361 = ( n8479 & ~n15609 ) | ( n8479 & n19360 ) | ( ~n15609 & n19360 ) ;
  assign n19362 = n19361 ^ n8180 ^ n6896 ;
  assign n19366 = n19365 ^ n19362 ^ n707 ;
  assign n19367 = n11338 ^ n10151 ^ n1098 ;
  assign n19368 = ( n1858 & n10782 ) | ( n1858 & ~n14865 ) | ( n10782 & ~n14865 ) ;
  assign n19369 = n19368 ^ n9257 ^ n564 ;
  assign n19370 = ( n5533 & n12548 ) | ( n5533 & n19369 ) | ( n12548 & n19369 ) ;
  assign n19372 = ( n3577 & n7944 ) | ( n3577 & ~n8851 ) | ( n7944 & ~n8851 ) ;
  assign n19373 = ( n7214 & n9200 ) | ( n7214 & ~n19372 ) | ( n9200 & ~n19372 ) ;
  assign n19371 = ( ~n6311 & n9768 ) | ( ~n6311 & n17279 ) | ( n9768 & n17279 ) ;
  assign n19374 = n19373 ^ n19371 ^ n8286 ;
  assign n19375 = ( n6650 & n9877 ) | ( n6650 & n19374 ) | ( n9877 & n19374 ) ;
  assign n19376 = ( n5467 & ~n11723 ) | ( n5467 & n12734 ) | ( ~n11723 & n12734 ) ;
  assign n19377 = ( n8154 & ~n12277 ) | ( n8154 & n19376 ) | ( ~n12277 & n19376 ) ;
  assign n19378 = n19377 ^ n14883 ^ n3147 ;
  assign n19379 = n9208 ^ n7449 ^ n2295 ;
  assign n19380 = n17756 ^ n10995 ^ n5668 ;
  assign n19381 = ( ~n3353 & n7215 ) | ( ~n3353 & n15084 ) | ( n7215 & n15084 ) ;
  assign n19382 = n19381 ^ n18967 ^ n5937 ;
  assign n19383 = ( ~n19379 & n19380 ) | ( ~n19379 & n19382 ) | ( n19380 & n19382 ) ;
  assign n19384 = n19383 ^ n16796 ^ n3825 ;
  assign n19391 = ( ~n12481 & n12836 ) | ( ~n12481 & n14646 ) | ( n12836 & n14646 ) ;
  assign n19386 = n12192 ^ n7319 ^ n7222 ;
  assign n19387 = n19386 ^ n18316 ^ n16188 ;
  assign n19385 = ( ~n1823 & n3056 ) | ( ~n1823 & n3656 ) | ( n3056 & n3656 ) ;
  assign n19388 = n19387 ^ n19385 ^ n2128 ;
  assign n19389 = ( x46 & ~n11204 ) | ( x46 & n19388 ) | ( ~n11204 & n19388 ) ;
  assign n19390 = n19389 ^ n17107 ^ n13119 ;
  assign n19392 = n19391 ^ n19390 ^ n1082 ;
  assign n19393 = n19013 ^ n15661 ^ n3841 ;
  assign n19394 = n11240 ^ n6519 ^ n132 ;
  assign n19395 = n19394 ^ n13946 ^ n8653 ;
  assign n19396 = ( n8423 & n13667 ) | ( n8423 & ~n15726 ) | ( n13667 & ~n15726 ) ;
  assign n19397 = n10827 ^ n9883 ^ n5800 ;
  assign n19398 = n19397 ^ n15230 ^ n8594 ;
  assign n19399 = n15650 ^ n6241 ^ n1959 ;
  assign n19405 = n7798 ^ n2045 ^ n1641 ;
  assign n19406 = n19405 ^ n9489 ^ n9169 ;
  assign n19400 = n7850 ^ n4114 ^ n3597 ;
  assign n19401 = ( ~n8239 & n14250 ) | ( ~n8239 & n19400 ) | ( n14250 & n19400 ) ;
  assign n19402 = ( n5394 & n8150 ) | ( n5394 & n19401 ) | ( n8150 & n19401 ) ;
  assign n19403 = ( n2516 & n10095 ) | ( n2516 & n19402 ) | ( n10095 & n19402 ) ;
  assign n19404 = ( n10560 & n14485 ) | ( n10560 & n19403 ) | ( n14485 & n19403 ) ;
  assign n19407 = n19406 ^ n19404 ^ n4702 ;
  assign n19408 = n19369 ^ n18466 ^ n3901 ;
  assign n19412 = n9089 ^ n7560 ^ n639 ;
  assign n19410 = ( n1265 & n1465 ) | ( n1265 & ~n3990 ) | ( n1465 & ~n3990 ) ;
  assign n19409 = ( n1032 & n9236 ) | ( n1032 & n12479 ) | ( n9236 & n12479 ) ;
  assign n19411 = n19410 ^ n19409 ^ n8292 ;
  assign n19413 = n19412 ^ n19411 ^ n10574 ;
  assign n19414 = n15405 ^ n8559 ^ n6954 ;
  assign n19415 = ( n393 & n9200 ) | ( n393 & ~n13742 ) | ( n9200 & ~n13742 ) ;
  assign n19416 = ( n5729 & n19414 ) | ( n5729 & ~n19415 ) | ( n19414 & ~n19415 ) ;
  assign n19417 = ( n866 & n4861 ) | ( n866 & n12971 ) | ( n4861 & n12971 ) ;
  assign n19418 = ( n13887 & ~n17267 ) | ( n13887 & n19417 ) | ( ~n17267 & n19417 ) ;
  assign n19419 = ( n2229 & n3853 ) | ( n2229 & n5252 ) | ( n3853 & n5252 ) ;
  assign n19420 = n19419 ^ n8315 ^ n531 ;
  assign n19421 = ( n822 & ~n8351 ) | ( n822 & n19420 ) | ( ~n8351 & n19420 ) ;
  assign n19423 = ( x17 & n2674 ) | ( x17 & ~n13928 ) | ( n2674 & ~n13928 ) ;
  assign n19422 = ( ~n3147 & n3394 ) | ( ~n3147 & n13184 ) | ( n3394 & n13184 ) ;
  assign n19424 = n19423 ^ n19422 ^ n674 ;
  assign n19426 = ( ~n5089 & n6244 ) | ( ~n5089 & n9028 ) | ( n6244 & n9028 ) ;
  assign n19425 = n8392 ^ n5205 ^ n3909 ;
  assign n19427 = n19426 ^ n19425 ^ n14879 ;
  assign n19430 = ( n3325 & ~n5172 ) | ( n3325 & n8106 ) | ( ~n5172 & n8106 ) ;
  assign n19431 = n19430 ^ n13236 ^ n12134 ;
  assign n19428 = ( n3252 & n5183 ) | ( n3252 & n15946 ) | ( n5183 & n15946 ) ;
  assign n19429 = ( n5935 & n6419 ) | ( n5935 & n19428 ) | ( n6419 & n19428 ) ;
  assign n19432 = n19431 ^ n19429 ^ n9579 ;
  assign n19433 = ( n16135 & ~n19427 ) | ( n16135 & n19432 ) | ( ~n19427 & n19432 ) ;
  assign n19434 = n14454 ^ n3814 ^ n3444 ;
  assign n19435 = ( x123 & n4123 ) | ( x123 & ~n19023 ) | ( n4123 & ~n19023 ) ;
  assign n19436 = ( n798 & n8393 ) | ( n798 & ~n19435 ) | ( n8393 & ~n19435 ) ;
  assign n19437 = ( n2683 & n9633 ) | ( n2683 & n19436 ) | ( n9633 & n19436 ) ;
  assign n19438 = ( n2873 & n5954 ) | ( n2873 & ~n17293 ) | ( n5954 & ~n17293 ) ;
  assign n19439 = n9370 ^ n8838 ^ n5766 ;
  assign n19440 = n11035 ^ n5895 ^ n1811 ;
  assign n19441 = ( n19438 & n19439 ) | ( n19438 & ~n19440 ) | ( n19439 & ~n19440 ) ;
  assign n19442 = n19441 ^ n18679 ^ n2720 ;
  assign n19443 = n5410 ^ n1773 ^ n721 ;
  assign n19444 = n13338 ^ n2244 ^ n761 ;
  assign n19445 = ( n4136 & n6767 ) | ( n4136 & ~n19444 ) | ( n6767 & ~n19444 ) ;
  assign n19446 = ( n15300 & n19443 ) | ( n15300 & n19445 ) | ( n19443 & n19445 ) ;
  assign n19447 = ( n1979 & n3067 ) | ( n1979 & n6460 ) | ( n3067 & n6460 ) ;
  assign n19448 = n11204 ^ n6917 ^ n4586 ;
  assign n19449 = ( ~n4990 & n5899 ) | ( ~n4990 & n7414 ) | ( n5899 & n7414 ) ;
  assign n19450 = ( n994 & n3805 ) | ( n994 & ~n19449 ) | ( n3805 & ~n19449 ) ;
  assign n19451 = ( n19447 & n19448 ) | ( n19447 & ~n19450 ) | ( n19448 & ~n19450 ) ;
  assign n19452 = ( n586 & n766 ) | ( n586 & n10882 ) | ( n766 & n10882 ) ;
  assign n19456 = ( ~n6745 & n12814 ) | ( ~n6745 & n15700 ) | ( n12814 & n15700 ) ;
  assign n19454 = ( ~n741 & n2495 ) | ( ~n741 & n9125 ) | ( n2495 & n9125 ) ;
  assign n19453 = ( n4214 & n13993 ) | ( n4214 & n15797 ) | ( n13993 & n15797 ) ;
  assign n19455 = n19454 ^ n19453 ^ n9077 ;
  assign n19457 = n19456 ^ n19455 ^ n8039 ;
  assign n19458 = ( n18114 & n19452 ) | ( n18114 & n19457 ) | ( n19452 & n19457 ) ;
  assign n19459 = ( n1579 & ~n11338 ) | ( n1579 & n16487 ) | ( ~n11338 & n16487 ) ;
  assign n19460 = n10765 ^ n8542 ^ n6271 ;
  assign n19461 = ( n8427 & ~n12148 ) | ( n8427 & n13653 ) | ( ~n12148 & n13653 ) ;
  assign n19462 = n18752 ^ n2029 ^ n1550 ;
  assign n19463 = ( n1133 & n3620 ) | ( n1133 & ~n8230 ) | ( n3620 & ~n8230 ) ;
  assign n19464 = ( n8988 & n13398 ) | ( n8988 & n18946 ) | ( n13398 & n18946 ) ;
  assign n19465 = n944 ^ n682 ^ x53 ;
  assign n19466 = ( n4627 & ~n6685 ) | ( n4627 & n19465 ) | ( ~n6685 & n19465 ) ;
  assign n19467 = n2726 ^ n1504 ^ n718 ;
  assign n19468 = ( n4457 & ~n6441 ) | ( n4457 & n13232 ) | ( ~n6441 & n13232 ) ;
  assign n19469 = n16659 ^ n11638 ^ n3852 ;
  assign n19470 = ( ~n19467 & n19468 ) | ( ~n19467 & n19469 ) | ( n19468 & n19469 ) ;
  assign n19471 = ( n1780 & n11283 ) | ( n1780 & n19400 ) | ( n11283 & n19400 ) ;
  assign n19472 = n19471 ^ n11213 ^ n10111 ;
  assign n19473 = n19472 ^ n11578 ^ n1327 ;
  assign n19474 = n8145 ^ n5564 ^ n4937 ;
  assign n19475 = ( n252 & n15680 ) | ( n252 & n17408 ) | ( n15680 & n17408 ) ;
  assign n19478 = n10444 ^ n6240 ^ n3147 ;
  assign n19476 = ( n1953 & n6653 ) | ( n1953 & n9745 ) | ( n6653 & n9745 ) ;
  assign n19477 = ( n5032 & ~n5958 ) | ( n5032 & n19476 ) | ( ~n5958 & n19476 ) ;
  assign n19479 = n19478 ^ n19477 ^ n17553 ;
  assign n19480 = ( ~n3561 & n7826 ) | ( ~n3561 & n10631 ) | ( n7826 & n10631 ) ;
  assign n19481 = n14390 ^ n12690 ^ n427 ;
  assign n19482 = ( ~n1345 & n18334 ) | ( ~n1345 & n19481 ) | ( n18334 & n19481 ) ;
  assign n19483 = ( n10800 & n12297 ) | ( n10800 & ~n19482 ) | ( n12297 & ~n19482 ) ;
  assign n19484 = n18011 ^ n9091 ^ n3874 ;
  assign n19485 = n19484 ^ n18096 ^ n15869 ;
  assign n19486 = ( n3234 & n8026 ) | ( n3234 & n15898 ) | ( n8026 & n15898 ) ;
  assign n19487 = ( n2342 & n19454 ) | ( n2342 & n19486 ) | ( n19454 & n19486 ) ;
  assign n19488 = ( n287 & n980 ) | ( n287 & ~n12053 ) | ( n980 & ~n12053 ) ;
  assign n19489 = n19488 ^ n13178 ^ n6614 ;
  assign n19490 = n19489 ^ n12469 ^ n2417 ;
  assign n19491 = n6740 ^ n5933 ^ n4654 ;
  assign n19492 = ( n2062 & ~n9349 ) | ( n2062 & n19491 ) | ( ~n9349 & n19491 ) ;
  assign n19493 = n10157 ^ n9745 ^ n8302 ;
  assign n19494 = ( n4330 & ~n5967 ) | ( n4330 & n19493 ) | ( ~n5967 & n19493 ) ;
  assign n19495 = ( n13916 & ~n19492 ) | ( n13916 & n19494 ) | ( ~n19492 & n19494 ) ;
  assign n19496 = ( ~n6689 & n7879 ) | ( ~n6689 & n19495 ) | ( n7879 & n19495 ) ;
  assign n19498 = n11099 ^ n6835 ^ n3316 ;
  assign n19497 = ( n4543 & n10634 ) | ( n4543 & ~n13421 ) | ( n10634 & ~n13421 ) ;
  assign n19499 = n19498 ^ n19497 ^ n2075 ;
  assign n19501 = n14870 ^ n10931 ^ n6530 ;
  assign n19502 = ( n7169 & ~n19161 ) | ( n7169 & n19501 ) | ( ~n19161 & n19501 ) ;
  assign n19500 = ( n1011 & ~n3502 ) | ( n1011 & n10075 ) | ( ~n3502 & n10075 ) ;
  assign n19503 = n19502 ^ n19500 ^ n977 ;
  assign n19504 = ( n4572 & n18443 ) | ( n4572 & ~n19503 ) | ( n18443 & ~n19503 ) ;
  assign n19505 = n8980 ^ n5018 ^ n4381 ;
  assign n19511 = ( ~n900 & n1596 ) | ( ~n900 & n13745 ) | ( n1596 & n13745 ) ;
  assign n19512 = n9741 ^ n6967 ^ n1257 ;
  assign n19513 = n19512 ^ n18536 ^ n1357 ;
  assign n19514 = ( n14201 & n19511 ) | ( n14201 & ~n19513 ) | ( n19511 & ~n19513 ) ;
  assign n19509 = ( n1346 & n9087 ) | ( n1346 & ~n13195 ) | ( n9087 & ~n13195 ) ;
  assign n19510 = n19509 ^ n14835 ^ n2532 ;
  assign n19507 = n15388 ^ n13127 ^ n3627 ;
  assign n19506 = n12945 ^ n8325 ^ n6104 ;
  assign n19508 = n19507 ^ n19506 ^ n15574 ;
  assign n19515 = n19514 ^ n19510 ^ n19508 ;
  assign n19516 = n14167 ^ n12396 ^ n6887 ;
  assign n19517 = n13619 ^ n5871 ^ n4129 ;
  assign n19518 = n14248 ^ n7704 ^ n2348 ;
  assign n19519 = ( ~n12158 & n19517 ) | ( ~n12158 & n19518 ) | ( n19517 & n19518 ) ;
  assign n19520 = ( n9584 & ~n19516 ) | ( n9584 & n19519 ) | ( ~n19516 & n19519 ) ;
  assign n19521 = n14090 ^ n13403 ^ n1211 ;
  assign n19522 = n13456 ^ n9195 ^ n287 ;
  assign n19523 = n17093 ^ n8886 ^ n3356 ;
  assign n19524 = n16642 ^ n11895 ^ n9511 ;
  assign n19525 = n19524 ^ n13008 ^ n2887 ;
  assign n19526 = ( n1745 & n7571 ) | ( n1745 & ~n14865 ) | ( n7571 & ~n14865 ) ;
  assign n19527 = n5380 ^ n5295 ^ n3480 ;
  assign n19528 = ( ~n3427 & n8308 ) | ( ~n3427 & n19527 ) | ( n8308 & n19527 ) ;
  assign n19529 = ( ~n847 & n6336 ) | ( ~n847 & n19528 ) | ( n6336 & n19528 ) ;
  assign n19531 = ( ~n7796 & n10502 ) | ( ~n7796 & n12242 ) | ( n10502 & n12242 ) ;
  assign n19530 = n2946 ^ n1262 ^ n933 ;
  assign n19532 = n19531 ^ n19530 ^ n2631 ;
  assign n19533 = ( n1930 & n11166 ) | ( n1930 & n14139 ) | ( n11166 & n14139 ) ;
  assign n19534 = ( n6986 & ~n14734 ) | ( n6986 & n19533 ) | ( ~n14734 & n19533 ) ;
  assign n19535 = ( n6273 & n6357 ) | ( n6273 & ~n19534 ) | ( n6357 & ~n19534 ) ;
  assign n19536 = n14541 ^ n6240 ^ n3890 ;
  assign n19537 = n19536 ^ n13352 ^ n3179 ;
  assign n19538 = ( n8775 & ~n14037 ) | ( n8775 & n19494 ) | ( ~n14037 & n19494 ) ;
  assign n19539 = ( ~n3245 & n4944 ) | ( ~n3245 & n7356 ) | ( n4944 & n7356 ) ;
  assign n19540 = ( n15742 & n16381 ) | ( n15742 & n19539 ) | ( n16381 & n19539 ) ;
  assign n19541 = ( n6037 & n8438 ) | ( n6037 & n19540 ) | ( n8438 & n19540 ) ;
  assign n19542 = n13353 ^ n4808 ^ n3177 ;
  assign n19543 = n19542 ^ n12740 ^ n12538 ;
  assign n19544 = ( ~n642 & n16383 ) | ( ~n642 & n19055 ) | ( n16383 & n19055 ) ;
  assign n19545 = n5426 ^ n4944 ^ n353 ;
  assign n19546 = ( n11661 & n16239 ) | ( n11661 & ~n19545 ) | ( n16239 & ~n19545 ) ;
  assign n19547 = ( x92 & n910 ) | ( x92 & ~n19546 ) | ( n910 & ~n19546 ) ;
  assign n19548 = n8375 ^ n7760 ^ n4808 ;
  assign n19549 = ( ~n1809 & n4110 ) | ( ~n1809 & n19548 ) | ( n4110 & n19548 ) ;
  assign n19550 = ( ~n10802 & n15232 ) | ( ~n10802 & n19549 ) | ( n15232 & n19549 ) ;
  assign n19551 = n19550 ^ n18872 ^ n1011 ;
  assign n19552 = n14422 ^ n8063 ^ n4080 ;
  assign n19553 = ( n4764 & n18752 ) | ( n4764 & ~n19552 ) | ( n18752 & ~n19552 ) ;
  assign n19554 = ( n6502 & n7271 ) | ( n6502 & n8779 ) | ( n7271 & n8779 ) ;
  assign n19555 = ( n4855 & n14334 ) | ( n4855 & n19554 ) | ( n14334 & n19554 ) ;
  assign n19556 = n17260 ^ n14358 ^ n12005 ;
  assign n19557 = n6698 ^ n5476 ^ n1591 ;
  assign n19558 = n19557 ^ n13368 ^ n8314 ;
  assign n19559 = n13296 ^ n2900 ^ n2386 ;
  assign n19560 = ( n3847 & n3868 ) | ( n3847 & n10169 ) | ( n3868 & n10169 ) ;
  assign n19561 = ( n4045 & ~n19559 ) | ( n4045 & n19560 ) | ( ~n19559 & n19560 ) ;
  assign n19562 = ( n2232 & ~n7314 ) | ( n2232 & n7755 ) | ( ~n7314 & n7755 ) ;
  assign n19563 = ( n4479 & n12101 ) | ( n4479 & n19562 ) | ( n12101 & n19562 ) ;
  assign n19564 = ( ~n11809 & n18644 ) | ( ~n11809 & n19563 ) | ( n18644 & n19563 ) ;
  assign n19565 = n4612 ^ n1020 ^ n788 ;
  assign n19566 = ( ~n5161 & n8814 ) | ( ~n5161 & n19565 ) | ( n8814 & n19565 ) ;
  assign n19567 = ( n3175 & n12183 ) | ( n3175 & n12821 ) | ( n12183 & n12821 ) ;
  assign n19568 = n19567 ^ n15739 ^ n12925 ;
  assign n19569 = ( n154 & n19566 ) | ( n154 & ~n19568 ) | ( n19566 & ~n19568 ) ;
  assign n19573 = n7611 ^ n7198 ^ n5120 ;
  assign n19574 = n19573 ^ n7276 ^ n2073 ;
  assign n19572 = ( n5913 & n15418 ) | ( n5913 & ~n16919 ) | ( n15418 & ~n16919 ) ;
  assign n19575 = n19574 ^ n19572 ^ n16979 ;
  assign n19570 = ( n1752 & n7767 ) | ( n1752 & ~n9947 ) | ( n7767 & ~n9947 ) ;
  assign n19571 = n19570 ^ n10679 ^ x83 ;
  assign n19576 = n19575 ^ n19571 ^ n10913 ;
  assign n19578 = n11821 ^ n9119 ^ n7207 ;
  assign n19579 = ( ~n3295 & n4775 ) | ( ~n3295 & n19578 ) | ( n4775 & n19578 ) ;
  assign n19580 = n19579 ^ n19452 ^ n3058 ;
  assign n19577 = ( ~n4129 & n15802 ) | ( ~n4129 & n16773 ) | ( n15802 & n16773 ) ;
  assign n19581 = n19580 ^ n19577 ^ n13631 ;
  assign n19582 = ( n1184 & ~n5218 ) | ( n1184 & n5600 ) | ( ~n5218 & n5600 ) ;
  assign n19583 = n8595 ^ n5555 ^ n1990 ;
  assign n19584 = ( n13005 & n13991 ) | ( n13005 & ~n19583 ) | ( n13991 & ~n19583 ) ;
  assign n19585 = n17131 ^ n11829 ^ n6688 ;
  assign n19586 = ( ~n5566 & n6005 ) | ( ~n5566 & n8749 ) | ( n6005 & n8749 ) ;
  assign n19587 = n19586 ^ n14744 ^ n531 ;
  assign n19588 = ( ~n7513 & n9432 ) | ( ~n7513 & n15884 ) | ( n9432 & n15884 ) ;
  assign n19589 = ( n5071 & n15238 ) | ( n5071 & ~n19588 ) | ( n15238 & ~n19588 ) ;
  assign n19590 = ( n14285 & n19587 ) | ( n14285 & n19589 ) | ( n19587 & n19589 ) ;
  assign n19591 = ( ~n508 & n4360 ) | ( ~n508 & n6838 ) | ( n4360 & n6838 ) ;
  assign n19592 = ( ~n868 & n19590 ) | ( ~n868 & n19591 ) | ( n19590 & n19591 ) ;
  assign n19593 = n9211 ^ n8564 ^ n3914 ;
  assign n19594 = n19593 ^ n9626 ^ n8627 ;
  assign n19595 = ( n275 & n306 ) | ( n275 & n1047 ) | ( n306 & n1047 ) ;
  assign n19596 = n8254 ^ n7356 ^ n1115 ;
  assign n19597 = ( ~n8454 & n11311 ) | ( ~n8454 & n14644 ) | ( n11311 & n14644 ) ;
  assign n19598 = ( n10153 & n19596 ) | ( n10153 & n19597 ) | ( n19596 & n19597 ) ;
  assign n19599 = n6515 ^ n3800 ^ n203 ;
  assign n19600 = ( n1920 & ~n13714 ) | ( n1920 & n16275 ) | ( ~n13714 & n16275 ) ;
  assign n19601 = ( ~n2198 & n11450 ) | ( ~n2198 & n19600 ) | ( n11450 & n19600 ) ;
  assign n19602 = n7755 ^ n4950 ^ n4116 ;
  assign n19603 = ( n19599 & n19601 ) | ( n19599 & ~n19602 ) | ( n19601 & ~n19602 ) ;
  assign n19604 = n16587 ^ n14456 ^ n9453 ;
  assign n19605 = n6437 ^ n5219 ^ n3656 ;
  assign n19606 = ( n634 & ~n19604 ) | ( n634 & n19605 ) | ( ~n19604 & n19605 ) ;
  assign n19607 = n18133 ^ n9359 ^ n741 ;
  assign n19616 = n12013 ^ n10436 ^ n6282 ;
  assign n19614 = n17708 ^ n1354 ^ n1348 ;
  assign n19612 = n14994 ^ n14173 ^ n3170 ;
  assign n19613 = n19612 ^ n10251 ^ n3519 ;
  assign n19609 = ( n2518 & n6277 ) | ( n2518 & ~n13013 ) | ( n6277 & ~n13013 ) ;
  assign n19608 = n10447 ^ n1899 ^ n891 ;
  assign n19610 = n19609 ^ n19608 ^ n13064 ;
  assign n19611 = ( n13479 & n16247 ) | ( n13479 & ~n19610 ) | ( n16247 & ~n19610 ) ;
  assign n19615 = n19614 ^ n19613 ^ n19611 ;
  assign n19617 = n19616 ^ n19615 ^ n6204 ;
  assign n19618 = ( n5751 & ~n17115 ) | ( n5751 & n17686 ) | ( ~n17115 & n17686 ) ;
  assign n19619 = ( n6826 & ~n8077 ) | ( n6826 & n9954 ) | ( ~n8077 & n9954 ) ;
  assign n19620 = ( ~n172 & n499 ) | ( ~n172 & n1530 ) | ( n499 & n1530 ) ;
  assign n19621 = ( n6334 & ~n19619 ) | ( n6334 & n19620 ) | ( ~n19619 & n19620 ) ;
  assign n19622 = ( ~n13814 & n17775 ) | ( ~n13814 & n17855 ) | ( n17775 & n17855 ) ;
  assign n19623 = ( n697 & n2119 ) | ( n697 & n8697 ) | ( n2119 & n8697 ) ;
  assign n19624 = ( ~n5390 & n8204 ) | ( ~n5390 & n13894 ) | ( n8204 & n13894 ) ;
  assign n19625 = n14781 ^ n14285 ^ n7054 ;
  assign n19626 = ( ~n1824 & n14320 ) | ( ~n1824 & n19625 ) | ( n14320 & n19625 ) ;
  assign n19627 = ( n15265 & n19624 ) | ( n15265 & ~n19626 ) | ( n19624 & ~n19626 ) ;
  assign n19628 = ( ~n8773 & n19623 ) | ( ~n8773 & n19627 ) | ( n19623 & n19627 ) ;
  assign n19629 = ( n7481 & ~n19622 ) | ( n7481 & n19628 ) | ( ~n19622 & n19628 ) ;
  assign n19630 = n16480 ^ n13658 ^ n4250 ;
  assign n19631 = ( x2 & ~n6137 ) | ( x2 & n17165 ) | ( ~n6137 & n17165 ) ;
  assign n19632 = n14335 ^ n7715 ^ n3168 ;
  assign n19633 = ( n15653 & n19631 ) | ( n15653 & n19632 ) | ( n19631 & n19632 ) ;
  assign n19634 = n6281 ^ n3897 ^ n1193 ;
  assign n19635 = n19634 ^ n5042 ^ n1037 ;
  assign n19636 = ( n10720 & ~n13708 ) | ( n10720 & n16991 ) | ( ~n13708 & n16991 ) ;
  assign n19641 = n18132 ^ n6967 ^ n3262 ;
  assign n19638 = ( n3661 & n6215 ) | ( n3661 & n12365 ) | ( n6215 & n12365 ) ;
  assign n19639 = ( n295 & n931 ) | ( n295 & ~n7282 ) | ( n931 & ~n7282 ) ;
  assign n19640 = ( n15190 & n19638 ) | ( n15190 & ~n19639 ) | ( n19638 & ~n19639 ) ;
  assign n19642 = n19641 ^ n19640 ^ n10753 ;
  assign n19643 = ( ~n9456 & n10913 ) | ( ~n9456 & n19642 ) | ( n10913 & n19642 ) ;
  assign n19637 = ( n11796 & n12010 ) | ( n11796 & ~n16661 ) | ( n12010 & ~n16661 ) ;
  assign n19644 = n19643 ^ n19637 ^ n2216 ;
  assign n19645 = n19644 ^ n10991 ^ n3148 ;
  assign n19646 = n1496 ^ n809 ^ x43 ;
  assign n19647 = n19646 ^ n10063 ^ n3598 ;
  assign n19648 = n17930 ^ n17425 ^ n17069 ;
  assign n19651 = n15721 ^ n10416 ^ n836 ;
  assign n19652 = n19651 ^ n7720 ^ n3257 ;
  assign n19649 = n15193 ^ n6432 ^ n2247 ;
  assign n19650 = ( ~n3636 & n14865 ) | ( ~n3636 & n19649 ) | ( n14865 & n19649 ) ;
  assign n19653 = n19652 ^ n19650 ^ n11982 ;
  assign n19654 = n8427 ^ n6811 ^ n6518 ;
  assign n19655 = n19654 ^ n18402 ^ n5429 ;
  assign n19656 = n16132 ^ n10128 ^ n255 ;
  assign n19657 = ( n4957 & n7433 ) | ( n4957 & n19656 ) | ( n7433 & n19656 ) ;
  assign n19658 = ( n2482 & n4266 ) | ( n2482 & n4695 ) | ( n4266 & n4695 ) ;
  assign n19659 = ( n530 & n6299 ) | ( n530 & ~n17069 ) | ( n6299 & ~n17069 ) ;
  assign n19660 = n19659 ^ n17911 ^ n744 ;
  assign n19661 = n19660 ^ n18125 ^ n5467 ;
  assign n19662 = ( n2381 & n19658 ) | ( n2381 & ~n19661 ) | ( n19658 & ~n19661 ) ;
  assign n19663 = ( ~n6297 & n8352 ) | ( ~n6297 & n10278 ) | ( n8352 & n10278 ) ;
  assign n19664 = ( n12913 & n16231 ) | ( n12913 & n19046 ) | ( n16231 & n19046 ) ;
  assign n19665 = ( n13726 & n19663 ) | ( n13726 & n19664 ) | ( n19663 & n19664 ) ;
  assign n19668 = ( ~n6622 & n9652 ) | ( ~n6622 & n11096 ) | ( n9652 & n11096 ) ;
  assign n19666 = n12916 ^ n10477 ^ n2737 ;
  assign n19667 = ( ~n6128 & n14034 ) | ( ~n6128 & n19666 ) | ( n14034 & n19666 ) ;
  assign n19669 = n19668 ^ n19667 ^ n4385 ;
  assign n19670 = n19669 ^ n19574 ^ n4839 ;
  assign n19671 = ( n977 & ~n13372 ) | ( n977 & n13770 ) | ( ~n13372 & n13770 ) ;
  assign n19672 = n19671 ^ n5842 ^ n5058 ;
  assign n19673 = ( n4762 & ~n9795 ) | ( n4762 & n13811 ) | ( ~n9795 & n13811 ) ;
  assign n19674 = n19673 ^ n12399 ^ n1236 ;
  assign n19675 = ( ~n16370 & n19672 ) | ( ~n16370 & n19674 ) | ( n19672 & n19674 ) ;
  assign n19676 = ( ~n2048 & n12902 ) | ( ~n2048 & n19550 ) | ( n12902 & n19550 ) ;
  assign n19677 = n19355 ^ n17796 ^ n3360 ;
  assign n19680 = ( n390 & n3554 ) | ( n390 & ~n9100 ) | ( n3554 & ~n9100 ) ;
  assign n19681 = n19680 ^ n19162 ^ n4678 ;
  assign n19682 = n19681 ^ n12995 ^ n996 ;
  assign n19678 = ( n2678 & n7263 ) | ( n2678 & ~n12560 ) | ( n7263 & ~n12560 ) ;
  assign n19679 = ( n5741 & n17356 ) | ( n5741 & n19678 ) | ( n17356 & n19678 ) ;
  assign n19683 = n19682 ^ n19679 ^ n15592 ;
  assign n19684 = n10961 ^ n6885 ^ n205 ;
  assign n19685 = n17464 ^ n14809 ^ n6653 ;
  assign n19686 = ( n6711 & n19684 ) | ( n6711 & ~n19685 ) | ( n19684 & ~n19685 ) ;
  assign n19687 = n7137 ^ n4366 ^ n1777 ;
  assign n19688 = n19687 ^ n17323 ^ n4436 ;
  assign n19689 = ( n1495 & ~n3853 ) | ( n1495 & n6254 ) | ( ~n3853 & n6254 ) ;
  assign n19690 = n14181 ^ n3954 ^ n3636 ;
  assign n19691 = ( n8598 & ~n11196 ) | ( n8598 & n11796 ) | ( ~n11196 & n11796 ) ;
  assign n19692 = n19691 ^ n9804 ^ n7960 ;
  assign n19697 = n1473 ^ n841 ^ n635 ;
  assign n19698 = ( ~n7857 & n14438 ) | ( ~n7857 & n19697 ) | ( n14438 & n19697 ) ;
  assign n19693 = ( ~n2804 & n3290 ) | ( ~n2804 & n11538 ) | ( n3290 & n11538 ) ;
  assign n19694 = ( n2001 & n4300 ) | ( n2001 & ~n4612 ) | ( n4300 & ~n4612 ) ;
  assign n19695 = n19694 ^ n4298 ^ n3839 ;
  assign n19696 = ( n8051 & n19693 ) | ( n8051 & n19695 ) | ( n19693 & n19695 ) ;
  assign n19699 = n19698 ^ n19696 ^ n19448 ;
  assign n19700 = ( n1854 & ~n9748 ) | ( n1854 & n18404 ) | ( ~n9748 & n18404 ) ;
  assign n19702 = ( n1438 & ~n4221 ) | ( n1438 & n7285 ) | ( ~n4221 & n7285 ) ;
  assign n19701 = ( n6828 & n13023 ) | ( n6828 & n14869 ) | ( n13023 & n14869 ) ;
  assign n19703 = n19702 ^ n19701 ^ n4843 ;
  assign n19706 = n6860 ^ n4130 ^ n3003 ;
  assign n19704 = ( n870 & ~n2576 ) | ( n870 & n7734 ) | ( ~n2576 & n7734 ) ;
  assign n19705 = ( n2450 & ~n4182 ) | ( n2450 & n19704 ) | ( ~n4182 & n19704 ) ;
  assign n19707 = n19706 ^ n19705 ^ n9847 ;
  assign n19709 = ( n3559 & n3704 ) | ( n3559 & ~n7589 ) | ( n3704 & ~n7589 ) ;
  assign n19708 = ( n7171 & n17939 ) | ( n7171 & n19247 ) | ( n17939 & n19247 ) ;
  assign n19710 = n19709 ^ n19708 ^ n4572 ;
  assign n19711 = ( n6762 & ~n8605 ) | ( n6762 & n19710 ) | ( ~n8605 & n19710 ) ;
  assign n19712 = n14047 ^ n3244 ^ n961 ;
  assign n19715 = ( n466 & n6164 ) | ( n466 & n7402 ) | ( n6164 & n7402 ) ;
  assign n19713 = ( n1063 & ~n4704 ) | ( n1063 & n8557 ) | ( ~n4704 & n8557 ) ;
  assign n19714 = ( n9469 & n12801 ) | ( n9469 & n19713 ) | ( n12801 & n19713 ) ;
  assign n19716 = n19715 ^ n19714 ^ n1562 ;
  assign n19717 = ( n2596 & n8553 ) | ( n2596 & ~n12497 ) | ( n8553 & ~n12497 ) ;
  assign n19718 = ( n1368 & ~n1516 ) | ( n1368 & n17626 ) | ( ~n1516 & n17626 ) ;
  assign n19719 = ( n5155 & ~n19717 ) | ( n5155 & n19718 ) | ( ~n19717 & n19718 ) ;
  assign n19720 = n16076 ^ n7796 ^ n1090 ;
  assign n19721 = ( n11667 & n17993 ) | ( n11667 & n19720 ) | ( n17993 & n19720 ) ;
  assign n19722 = n17485 ^ n13184 ^ n7604 ;
  assign n19723 = ( n5072 & n19721 ) | ( n5072 & n19722 ) | ( n19721 & n19722 ) ;
  assign n19724 = n13671 ^ n9959 ^ n8598 ;
  assign n19728 = ( n5958 & n6203 ) | ( n5958 & ~n13789 ) | ( n6203 & ~n13789 ) ;
  assign n19729 = n19728 ^ n7265 ^ n485 ;
  assign n19730 = n14027 ^ n6714 ^ n1756 ;
  assign n19731 = ( n5155 & ~n19729 ) | ( n5155 & n19730 ) | ( ~n19729 & n19730 ) ;
  assign n19725 = n17950 ^ n3543 ^ n1571 ;
  assign n19726 = ( n991 & n1689 ) | ( n991 & ~n19725 ) | ( n1689 & ~n19725 ) ;
  assign n19727 = n19726 ^ n6983 ^ n2092 ;
  assign n19732 = n19731 ^ n19727 ^ n9501 ;
  assign n19733 = n8395 ^ n6030 ^ n868 ;
  assign n19734 = n7649 ^ n6241 ^ n993 ;
  assign n19735 = n19734 ^ n1987 ^ x74 ;
  assign n19736 = n19735 ^ n12837 ^ n197 ;
  assign n19737 = n15853 ^ n7458 ^ n4025 ;
  assign n19738 = n12494 ^ n11667 ^ n1320 ;
  assign n19739 = n19738 ^ n13848 ^ n1044 ;
  assign n19740 = ( n5130 & n14905 ) | ( n5130 & ~n19739 ) | ( n14905 & ~n19739 ) ;
  assign n19741 = ( n963 & ~n19737 ) | ( n963 & n19740 ) | ( ~n19737 & n19740 ) ;
  assign n19742 = ( x78 & ~n801 ) | ( x78 & n1883 ) | ( ~n801 & n1883 ) ;
  assign n19743 = n18994 ^ n4319 ^ n1835 ;
  assign n19744 = ( ~n4628 & n6731 ) | ( ~n4628 & n19743 ) | ( n6731 & n19743 ) ;
  assign n19745 = ( n550 & ~n6248 ) | ( n550 & n13228 ) | ( ~n6248 & n13228 ) ;
  assign n19746 = ( n19742 & n19744 ) | ( n19742 & n19745 ) | ( n19744 & n19745 ) ;
  assign n19749 = n13928 ^ n8555 ^ n1467 ;
  assign n19747 = n3876 ^ n2462 ^ n2399 ;
  assign n19748 = ( n2405 & ~n13061 ) | ( n2405 & n19747 ) | ( ~n13061 & n19747 ) ;
  assign n19750 = n19749 ^ n19748 ^ n18648 ;
  assign n19751 = n12831 ^ n6887 ^ n3687 ;
  assign n19752 = n3625 ^ n3281 ^ n1886 ;
  assign n19753 = n19752 ^ n8392 ^ n3837 ;
  assign n19754 = ( ~n794 & n2217 ) | ( ~n794 & n19753 ) | ( n2217 & n19753 ) ;
  assign n19755 = n19297 ^ n2817 ^ n1776 ;
  assign n19756 = ( n3935 & n5459 ) | ( n3935 & n9800 ) | ( n5459 & n9800 ) ;
  assign n19757 = ( n1855 & ~n7078 ) | ( n1855 & n13558 ) | ( ~n7078 & n13558 ) ;
  assign n19758 = ( ~n10641 & n19756 ) | ( ~n10641 & n19757 ) | ( n19756 & n19757 ) ;
  assign n19759 = ( n8415 & ~n11387 ) | ( n8415 & n16413 ) | ( ~n11387 & n16413 ) ;
  assign n19760 = ( n2313 & n18328 ) | ( n2313 & ~n19759 ) | ( n18328 & ~n19759 ) ;
  assign n19761 = ( n4128 & n6798 ) | ( n4128 & ~n19694 ) | ( n6798 & ~n19694 ) ;
  assign n19762 = ( n6087 & ~n18906 ) | ( n6087 & n19199 ) | ( ~n18906 & n19199 ) ;
  assign n19763 = ( n4491 & ~n16356 ) | ( n4491 & n19762 ) | ( ~n16356 & n19762 ) ;
  assign n19764 = n17598 ^ n15768 ^ n5369 ;
  assign n19765 = ( n5840 & n12942 ) | ( n5840 & n19764 ) | ( n12942 & n19764 ) ;
  assign n19766 = ( ~n1500 & n5370 ) | ( ~n1500 & n7459 ) | ( n5370 & n7459 ) ;
  assign n19767 = ( ~n594 & n1917 ) | ( ~n594 & n17838 ) | ( n1917 & n17838 ) ;
  assign n19768 = ( n4552 & n19766 ) | ( n4552 & n19767 ) | ( n19766 & n19767 ) ;
  assign n19769 = ( n2252 & n3453 ) | ( n2252 & ~n6506 ) | ( n3453 & ~n6506 ) ;
  assign n19770 = n10504 ^ n595 ^ n448 ;
  assign n19771 = n15278 ^ n14027 ^ n6016 ;
  assign n19774 = ( n2111 & ~n3097 ) | ( n2111 & n5315 ) | ( ~n3097 & n5315 ) ;
  assign n19772 = n13853 ^ n4112 ^ n2325 ;
  assign n19773 = ( ~n1857 & n18328 ) | ( ~n1857 & n19772 ) | ( n18328 & n19772 ) ;
  assign n19775 = n19774 ^ n19773 ^ n15988 ;
  assign n19776 = ( n1736 & n5314 ) | ( n1736 & n17802 ) | ( n5314 & n17802 ) ;
  assign n19777 = n19776 ^ n9245 ^ n2227 ;
  assign n19778 = ( ~n4425 & n6425 ) | ( ~n4425 & n13976 ) | ( n6425 & n13976 ) ;
  assign n19779 = n19778 ^ n15481 ^ n529 ;
  assign n19780 = ( ~n2931 & n7559 ) | ( ~n2931 & n7990 ) | ( n7559 & n7990 ) ;
  assign n19781 = ( n591 & n8278 ) | ( n591 & ~n11556 ) | ( n8278 & ~n11556 ) ;
  assign n19782 = ( n11378 & ~n19780 ) | ( n11378 & n19781 ) | ( ~n19780 & n19781 ) ;
  assign n19783 = ( ~n14867 & n19779 ) | ( ~n14867 & n19782 ) | ( n19779 & n19782 ) ;
  assign n19784 = ( n3969 & ~n12617 ) | ( n3969 & n18417 ) | ( ~n12617 & n18417 ) ;
  assign n19785 = n8905 ^ n1699 ^ n360 ;
  assign n19786 = ( ~n14743 & n19778 ) | ( ~n14743 & n19785 ) | ( n19778 & n19785 ) ;
  assign n19787 = n19786 ^ n15514 ^ n12042 ;
  assign n19788 = ( n3814 & ~n3838 ) | ( n3814 & n6581 ) | ( ~n3838 & n6581 ) ;
  assign n19789 = ( n1980 & ~n5516 ) | ( n1980 & n19788 ) | ( ~n5516 & n19788 ) ;
  assign n19790 = ( n1313 & ~n4401 ) | ( n1313 & n6676 ) | ( ~n4401 & n6676 ) ;
  assign n19791 = n12309 ^ n2943 ^ n1445 ;
  assign n19792 = ( n4387 & ~n19790 ) | ( n4387 & n19791 ) | ( ~n19790 & n19791 ) ;
  assign n19793 = n19792 ^ n6268 ^ n4780 ;
  assign n19794 = ( ~n5056 & n8363 ) | ( ~n5056 & n18522 ) | ( n8363 & n18522 ) ;
  assign n19795 = n17532 ^ n9696 ^ n2162 ;
  assign n19796 = n16124 ^ n4212 ^ n785 ;
  assign n19797 = n19796 ^ n18894 ^ n6289 ;
  assign n19798 = n19797 ^ n2336 ^ n1368 ;
  assign n19799 = n15308 ^ n13026 ^ n1239 ;
  assign n19800 = ( ~n17932 & n18054 ) | ( ~n17932 & n19799 ) | ( n18054 & n19799 ) ;
  assign n19801 = ( n17268 & n19798 ) | ( n17268 & n19800 ) | ( n19798 & n19800 ) ;
  assign n19802 = n8773 ^ n5511 ^ n5142 ;
  assign n19803 = n14666 ^ n11279 ^ n4863 ;
  assign n19804 = ( n6134 & n19802 ) | ( n6134 & n19803 ) | ( n19802 & n19803 ) ;
  assign n19805 = ( n1705 & ~n3105 ) | ( n1705 & n15953 ) | ( ~n3105 & n15953 ) ;
  assign n19806 = n19805 ^ n19347 ^ n6513 ;
  assign n19807 = n3986 ^ n2839 ^ n706 ;
  assign n19808 = ( n10182 & ~n19622 ) | ( n10182 & n19807 ) | ( ~n19622 & n19807 ) ;
  assign n19809 = ( n4044 & n12368 ) | ( n4044 & n19808 ) | ( n12368 & n19808 ) ;
  assign n19810 = n15813 ^ n14754 ^ n5163 ;
  assign n19811 = ( ~n4216 & n7685 ) | ( ~n4216 & n19530 ) | ( n7685 & n19530 ) ;
  assign n19812 = ( n13287 & ~n14126 ) | ( n13287 & n19811 ) | ( ~n14126 & n19811 ) ;
  assign n19813 = n13251 ^ n5580 ^ x13 ;
  assign n19814 = ( n12374 & ~n19109 ) | ( n12374 & n19813 ) | ( ~n19109 & n19813 ) ;
  assign n19815 = n6285 ^ n1554 ^ n982 ;
  assign n19816 = n17882 ^ n4865 ^ n3374 ;
  assign n19817 = ( n6710 & n19815 ) | ( n6710 & ~n19816 ) | ( n19815 & ~n19816 ) ;
  assign n19820 = ( ~n248 & n1692 ) | ( ~n248 & n12241 ) | ( n1692 & n12241 ) ;
  assign n19821 = n18073 ^ n2967 ^ n299 ;
  assign n19822 = ( n5053 & n19820 ) | ( n5053 & n19821 ) | ( n19820 & n19821 ) ;
  assign n19818 = ( n3117 & n5476 ) | ( n3117 & ~n10474 ) | ( n5476 & ~n10474 ) ;
  assign n19819 = ( n2796 & n13396 ) | ( n2796 & ~n19818 ) | ( n13396 & ~n19818 ) ;
  assign n19823 = n19822 ^ n19819 ^ n11235 ;
  assign n19824 = ( n2377 & ~n3020 ) | ( n2377 & n8729 ) | ( ~n3020 & n8729 ) ;
  assign n19825 = n19824 ^ n13682 ^ n9778 ;
  assign n19826 = n19825 ^ n18083 ^ n7680 ;
  assign n19827 = n12242 ^ n11838 ^ n4191 ;
  assign n19828 = n19827 ^ n18691 ^ n2600 ;
  assign n19829 = n6790 ^ n6440 ^ n3160 ;
  assign n19830 = n19829 ^ n16586 ^ n7714 ;
  assign n19831 = ( n301 & n13429 ) | ( n301 & ~n19830 ) | ( n13429 & ~n19830 ) ;
  assign n19832 = ( n2965 & n11213 ) | ( n2965 & n11418 ) | ( n11213 & n11418 ) ;
  assign n19833 = ( ~n19828 & n19831 ) | ( ~n19828 & n19832 ) | ( n19831 & n19832 ) ;
  assign n19834 = n9114 ^ n5626 ^ n1732 ;
  assign n19835 = n19834 ^ n8769 ^ n700 ;
  assign n19836 = ( ~n9189 & n12810 ) | ( ~n9189 & n19835 ) | ( n12810 & n19835 ) ;
  assign n19837 = ( ~n1481 & n1820 ) | ( ~n1481 & n3673 ) | ( n1820 & n3673 ) ;
  assign n19838 = n19837 ^ n13882 ^ n5340 ;
  assign n19839 = ( n7797 & n19836 ) | ( n7797 & n19838 ) | ( n19836 & n19838 ) ;
  assign n19840 = n17463 ^ n15385 ^ n6442 ;
  assign n19841 = n5850 ^ n2088 ^ n1447 ;
  assign n19842 = ( n14339 & n19632 ) | ( n14339 & n19841 ) | ( n19632 & n19841 ) ;
  assign n19844 = n18150 ^ n15495 ^ n2354 ;
  assign n19843 = n9674 ^ n2083 ^ n181 ;
  assign n19845 = n19844 ^ n19843 ^ n4281 ;
  assign n19846 = ( ~n2553 & n8450 ) | ( ~n2553 & n19845 ) | ( n8450 & n19845 ) ;
  assign n19847 = ( n3368 & n10895 ) | ( n3368 & n17022 ) | ( n10895 & n17022 ) ;
  assign n19848 = n9341 ^ n7901 ^ n1265 ;
  assign n19849 = ( ~n1554 & n1676 ) | ( ~n1554 & n11247 ) | ( n1676 & n11247 ) ;
  assign n19850 = ( n14124 & n19848 ) | ( n14124 & ~n19849 ) | ( n19848 & ~n19849 ) ;
  assign n19851 = n5448 ^ n5001 ^ n591 ;
  assign n19852 = ( n10404 & n11686 ) | ( n10404 & n17466 ) | ( n11686 & n17466 ) ;
  assign n19853 = ( n2285 & n19851 ) | ( n2285 & ~n19852 ) | ( n19851 & ~n19852 ) ;
  assign n19854 = n8501 ^ n7449 ^ n2390 ;
  assign n19855 = n5519 ^ n3358 ^ n1363 ;
  assign n19856 = ( n17068 & n18210 ) | ( n17068 & n19855 ) | ( n18210 & n19855 ) ;
  assign n19857 = ( n1868 & n5787 ) | ( n1868 & ~n9029 ) | ( n5787 & ~n9029 ) ;
  assign n19858 = n19857 ^ n14782 ^ n5530 ;
  assign n19859 = ( n2291 & n2516 ) | ( n2291 & ~n4328 ) | ( n2516 & ~n4328 ) ;
  assign n19860 = n19859 ^ n18603 ^ n1256 ;
  assign n19861 = n19860 ^ n15879 ^ n10946 ;
  assign n19862 = ( n1870 & ~n3496 ) | ( n1870 & n5005 ) | ( ~n3496 & n5005 ) ;
  assign n19863 = n13966 ^ n8774 ^ n8167 ;
  assign n19864 = ( n8827 & n16340 ) | ( n8827 & ~n19863 ) | ( n16340 & ~n19863 ) ;
  assign n19865 = ( n11445 & n19862 ) | ( n11445 & ~n19864 ) | ( n19862 & ~n19864 ) ;
  assign n19869 = ( n349 & ~n3671 ) | ( n349 & n8274 ) | ( ~n3671 & n8274 ) ;
  assign n19867 = ( n2164 & n2637 ) | ( n2164 & n7420 ) | ( n2637 & n7420 ) ;
  assign n19866 = n12426 ^ n11220 ^ n4312 ;
  assign n19868 = n19867 ^ n19866 ^ n433 ;
  assign n19870 = n19869 ^ n19868 ^ n3863 ;
  assign n19872 = n8047 ^ n7832 ^ n1014 ;
  assign n19871 = ( ~n4195 & n5512 ) | ( ~n4195 & n11235 ) | ( n5512 & n11235 ) ;
  assign n19873 = n19872 ^ n19871 ^ n3891 ;
  assign n19874 = n17443 ^ n13472 ^ n9656 ;
  assign n19875 = n9965 ^ n6002 ^ n4831 ;
  assign n19876 = ( n5372 & ~n9004 ) | ( n5372 & n19875 ) | ( ~n9004 & n19875 ) ;
  assign n19877 = n11948 ^ n10032 ^ n1419 ;
  assign n19878 = ( n11004 & ~n19495 ) | ( n11004 & n19877 ) | ( ~n19495 & n19877 ) ;
  assign n19879 = n14529 ^ n9948 ^ n7240 ;
  assign n19880 = n19879 ^ n17111 ^ n8212 ;
  assign n19881 = n14110 ^ n8195 ^ n7589 ;
  assign n19888 = n16226 ^ n14436 ^ n5047 ;
  assign n19885 = ( n7517 & ~n8061 ) | ( n7517 & n14278 ) | ( ~n8061 & n14278 ) ;
  assign n19883 = ( n874 & n1033 ) | ( n874 & n7636 ) | ( n1033 & n7636 ) ;
  assign n19884 = ( n2367 & n10146 ) | ( n2367 & n19883 ) | ( n10146 & n19883 ) ;
  assign n19882 = ( n1823 & n7636 ) | ( n1823 & ~n16641 ) | ( n7636 & ~n16641 ) ;
  assign n19886 = n19885 ^ n19884 ^ n19882 ;
  assign n19887 = ( n11328 & ~n16478 ) | ( n11328 & n19886 ) | ( ~n16478 & n19886 ) ;
  assign n19889 = n19888 ^ n19887 ^ n708 ;
  assign n19890 = ( n17349 & ~n18326 ) | ( n17349 & n18783 ) | ( ~n18326 & n18783 ) ;
  assign n19891 = ( n1106 & ~n11926 ) | ( n1106 & n14714 ) | ( ~n11926 & n14714 ) ;
  assign n19892 = n12397 ^ n6308 ^ n5593 ;
  assign n19893 = ( ~n422 & n8327 ) | ( ~n422 & n19892 ) | ( n8327 & n19892 ) ;
  assign n19894 = ( n8998 & n17108 ) | ( n8998 & n19893 ) | ( n17108 & n19893 ) ;
  assign n19898 = n10969 ^ n8296 ^ n8043 ;
  assign n19899 = ( n1920 & n2252 ) | ( n1920 & n19898 ) | ( n2252 & n19898 ) ;
  assign n19896 = ( n7904 & n10699 ) | ( n7904 & ~n13516 ) | ( n10699 & ~n13516 ) ;
  assign n19895 = n10758 ^ n4928 ^ n3649 ;
  assign n19897 = n19896 ^ n19895 ^ n16620 ;
  assign n19900 = n19899 ^ n19897 ^ n15900 ;
  assign n19901 = n5859 ^ n4443 ^ n2128 ;
  assign n19902 = n19901 ^ n14591 ^ n2446 ;
  assign n19907 = ( n4335 & ~n10175 ) | ( n4335 & n19527 ) | ( ~n10175 & n19527 ) ;
  assign n19904 = ( n235 & n4958 ) | ( n235 & n8298 ) | ( n4958 & n8298 ) ;
  assign n19905 = n19904 ^ n3497 ^ n1604 ;
  assign n19906 = ( n8804 & ~n13098 ) | ( n8804 & n19905 ) | ( ~n13098 & n19905 ) ;
  assign n19908 = n19907 ^ n19906 ^ n6804 ;
  assign n19903 = ( n673 & n9910 ) | ( n673 & n11056 ) | ( n9910 & n11056 ) ;
  assign n19909 = n19908 ^ n19903 ^ n5584 ;
  assign n19910 = n13646 ^ n3928 ^ n2329 ;
  assign n19911 = ( n3889 & n7954 ) | ( n3889 & ~n12414 ) | ( n7954 & ~n12414 ) ;
  assign n19912 = n19911 ^ n6484 ^ n2327 ;
  assign n19913 = n19912 ^ n19125 ^ n9175 ;
  assign n19914 = n16633 ^ n12875 ^ n1044 ;
  assign n19915 = n17204 ^ n11145 ^ n9346 ;
  assign n19916 = n10057 ^ n3295 ^ n1290 ;
  assign n19917 = n19916 ^ n13276 ^ n1601 ;
  assign n19918 = n9950 ^ n2731 ^ n2481 ;
  assign n19919 = n19918 ^ n19634 ^ n18160 ;
  assign n19920 = ( ~n10945 & n19917 ) | ( ~n10945 & n19919 ) | ( n19917 & n19919 ) ;
  assign n19921 = ( n4675 & n14183 ) | ( n4675 & ~n19920 ) | ( n14183 & ~n19920 ) ;
  assign n19922 = ( n408 & n3497 ) | ( n408 & ~n19908 ) | ( n3497 & ~n19908 ) ;
  assign n19923 = ( n4962 & n19143 ) | ( n4962 & ~n19922 ) | ( n19143 & ~n19922 ) ;
  assign n19924 = n17213 ^ n12414 ^ n8648 ;
  assign n19925 = n6701 ^ n3521 ^ n238 ;
  assign n19926 = ( n11022 & ~n19924 ) | ( n11022 & n19925 ) | ( ~n19924 & n19925 ) ;
  assign n19927 = n19926 ^ n14186 ^ n4878 ;
  assign n19928 = ( ~n3571 & n5387 ) | ( ~n3571 & n13072 ) | ( n5387 & n13072 ) ;
  assign n19930 = ( n2496 & ~n2787 ) | ( n2496 & n14841 ) | ( ~n2787 & n14841 ) ;
  assign n19931 = ( n1057 & n4725 ) | ( n1057 & n6218 ) | ( n4725 & n6218 ) ;
  assign n19932 = ( ~x63 & n19930 ) | ( ~x63 & n19931 ) | ( n19930 & n19931 ) ;
  assign n19929 = n9931 ^ n7181 ^ n309 ;
  assign n19933 = n19932 ^ n19929 ^ n15226 ;
  assign n19934 = n8118 ^ n4116 ^ n2943 ;
  assign n19935 = ( ~x7 & n859 ) | ( ~x7 & n19934 ) | ( n859 & n19934 ) ;
  assign n19936 = n19935 ^ n10265 ^ n2125 ;
  assign n19937 = ( ~n10620 & n12586 ) | ( ~n10620 & n19936 ) | ( n12586 & n19936 ) ;
  assign n19942 = ( n4239 & n10661 ) | ( n4239 & ~n10997 ) | ( n10661 & ~n10997 ) ;
  assign n19938 = ( n2238 & ~n2346 ) | ( n2238 & n8216 ) | ( ~n2346 & n8216 ) ;
  assign n19939 = n19938 ^ n10498 ^ x30 ;
  assign n19940 = ( ~n6562 & n12449 ) | ( ~n6562 & n19939 ) | ( n12449 & n19939 ) ;
  assign n19941 = ( n13615 & n18096 ) | ( n13615 & ~n19940 ) | ( n18096 & ~n19940 ) ;
  assign n19943 = n19942 ^ n19941 ^ n348 ;
  assign n19944 = n19604 ^ n18123 ^ n12581 ;
  assign n19945 = ( n2339 & ~n6620 ) | ( n2339 & n13227 ) | ( ~n6620 & n13227 ) ;
  assign n19946 = ( n573 & n9549 ) | ( n573 & n19945 ) | ( n9549 & n19945 ) ;
  assign n19947 = n19946 ^ n19728 ^ n4491 ;
  assign n19948 = ( ~n8733 & n12624 ) | ( ~n8733 & n19947 ) | ( n12624 & n19947 ) ;
  assign n19949 = n19056 ^ n16407 ^ n12341 ;
  assign n19950 = n15724 ^ n8795 ^ n4873 ;
  assign n19951 = ( n3134 & ~n5639 ) | ( n3134 & n7917 ) | ( ~n5639 & n7917 ) ;
  assign n19952 = n19951 ^ n2900 ^ n1768 ;
  assign n19953 = n14495 ^ n8565 ^ n3101 ;
  assign n19954 = n19953 ^ n2749 ^ n194 ;
  assign n19955 = ( n10099 & n11516 ) | ( n10099 & ~n18434 ) | ( n11516 & ~n18434 ) ;
  assign n19956 = ( n15743 & ~n19954 ) | ( n15743 & n19955 ) | ( ~n19954 & n19955 ) ;
  assign n19957 = n19956 ^ n12667 ^ n6736 ;
  assign n19958 = ( ~n6034 & n19952 ) | ( ~n6034 & n19957 ) | ( n19952 & n19957 ) ;
  assign n19959 = ( n5377 & ~n8014 ) | ( n5377 & n9369 ) | ( ~n8014 & n9369 ) ;
  assign n19960 = ( ~n2808 & n2868 ) | ( ~n2808 & n11217 ) | ( n2868 & n11217 ) ;
  assign n19961 = n8339 ^ n710 ^ n501 ;
  assign n19962 = n9561 ^ n2864 ^ n925 ;
  assign n19963 = ( n873 & ~n19961 ) | ( n873 & n19962 ) | ( ~n19961 & n19962 ) ;
  assign n19964 = ( n523 & n3324 ) | ( n523 & n5136 ) | ( n3324 & n5136 ) ;
  assign n19965 = ( n424 & n8673 ) | ( n424 & n19964 ) | ( n8673 & n19964 ) ;
  assign n19966 = n19965 ^ n9245 ^ n6991 ;
  assign n19967 = ( n15155 & n19963 ) | ( n15155 & ~n19966 ) | ( n19963 & ~n19966 ) ;
  assign n19968 = n19967 ^ n4478 ^ n3475 ;
  assign n19969 = n17804 ^ n9476 ^ n446 ;
  assign n19970 = ( n4758 & ~n18945 ) | ( n4758 & n19969 ) | ( ~n18945 & n19969 ) ;
  assign n19971 = n19970 ^ n8755 ^ x72 ;
  assign n19972 = n3633 ^ n3624 ^ n798 ;
  assign n19973 = ( ~n10131 & n11886 ) | ( ~n10131 & n19972 ) | ( n11886 & n19972 ) ;
  assign n19974 = ( ~n5479 & n17973 ) | ( ~n5479 & n19973 ) | ( n17973 & n19973 ) ;
  assign n19975 = ( ~n3910 & n4536 ) | ( ~n3910 & n8922 ) | ( n4536 & n8922 ) ;
  assign n19976 = ( n2977 & ~n4689 ) | ( n2977 & n19975 ) | ( ~n4689 & n19975 ) ;
  assign n19977 = ( n344 & n1294 ) | ( n344 & ~n3840 ) | ( n1294 & ~n3840 ) ;
  assign n19979 = n3772 ^ n1916 ^ n1180 ;
  assign n19978 = n18949 ^ n9985 ^ n4336 ;
  assign n19980 = n19979 ^ n19978 ^ n14050 ;
  assign n19981 = ( ~n3602 & n7148 ) | ( ~n3602 & n15515 ) | ( n7148 & n15515 ) ;
  assign n19982 = n19981 ^ n15895 ^ n4584 ;
  assign n19983 = ( n19977 & ~n19980 ) | ( n19977 & n19982 ) | ( ~n19980 & n19982 ) ;
  assign n19984 = n19983 ^ n12698 ^ n9113 ;
  assign n19985 = n5070 ^ n1193 ^ n441 ;
  assign n19986 = ( n1624 & n3417 ) | ( n1624 & n9135 ) | ( n3417 & n9135 ) ;
  assign n19987 = ( n4447 & ~n19985 ) | ( n4447 & n19986 ) | ( ~n19985 & n19986 ) ;
  assign n19988 = n19987 ^ n13713 ^ n12734 ;
  assign n19990 = n11681 ^ n10709 ^ n2400 ;
  assign n19991 = ( n9469 & n11250 ) | ( n9469 & ~n19990 ) | ( n11250 & ~n19990 ) ;
  assign n19989 = n19502 ^ n17655 ^ n2340 ;
  assign n19992 = n19991 ^ n19989 ^ n1274 ;
  assign n19993 = n18808 ^ n7755 ^ n6865 ;
  assign n19994 = ( n1295 & n3193 ) | ( n1295 & n6462 ) | ( n3193 & n6462 ) ;
  assign n19995 = ( n4626 & ~n11828 ) | ( n4626 & n19994 ) | ( ~n11828 & n19994 ) ;
  assign n19996 = ( n889 & n4460 ) | ( n889 & n5039 ) | ( n4460 & n5039 ) ;
  assign n19997 = ( n6352 & n19995 ) | ( n6352 & ~n19996 ) | ( n19995 & ~n19996 ) ;
  assign n19998 = ( ~n1152 & n4456 ) | ( ~n1152 & n6376 ) | ( n4456 & n6376 ) ;
  assign n19999 = ( n2358 & n5286 ) | ( n2358 & ~n15765 ) | ( n5286 & ~n15765 ) ;
  assign n20000 = n19999 ^ n5825 ^ n4718 ;
  assign n20001 = ( n6658 & n8583 ) | ( n6658 & n20000 ) | ( n8583 & n20000 ) ;
  assign n20002 = n14874 ^ n4914 ^ n1480 ;
  assign n20003 = ( ~n5471 & n18539 ) | ( ~n5471 & n20002 ) | ( n18539 & n20002 ) ;
  assign n20005 = n6838 ^ n3138 ^ n1791 ;
  assign n20004 = n10628 ^ n3804 ^ n1380 ;
  assign n20006 = n20005 ^ n20004 ^ n16515 ;
  assign n20007 = n20006 ^ n12717 ^ n4835 ;
  assign n20008 = n20005 ^ n19862 ^ n4620 ;
  assign n20009 = ( n1677 & n20007 ) | ( n1677 & ~n20008 ) | ( n20007 & ~n20008 ) ;
  assign n20011 = n9562 ^ n5209 ^ n1433 ;
  assign n20010 = n10312 ^ n6247 ^ n2609 ;
  assign n20012 = n20011 ^ n20010 ^ n13330 ;
  assign n20013 = n8543 ^ n8262 ^ n3515 ;
  assign n20014 = n20013 ^ n19742 ^ n16870 ;
  assign n20015 = n11778 ^ n5132 ^ n3162 ;
  assign n20016 = n4152 ^ n1967 ^ x127 ;
  assign n20017 = ( ~n999 & n20015 ) | ( ~n999 & n20016 ) | ( n20015 & n20016 ) ;
  assign n20018 = n20017 ^ n8406 ^ n580 ;
  assign n20019 = n17341 ^ n7726 ^ n6024 ;
  assign n20020 = n20019 ^ n4789 ^ n1423 ;
  assign n20021 = ( n8590 & ~n18842 ) | ( n8590 & n20020 ) | ( ~n18842 & n20020 ) ;
  assign n20022 = ( n13723 & ~n17494 ) | ( n13723 & n20021 ) | ( ~n17494 & n20021 ) ;
  assign n20023 = n4628 ^ n4469 ^ n836 ;
  assign n20024 = ( n1448 & n8549 ) | ( n1448 & n9373 ) | ( n8549 & n9373 ) ;
  assign n20025 = ( n17199 & n20023 ) | ( n17199 & ~n20024 ) | ( n20023 & ~n20024 ) ;
  assign n20026 = n13891 ^ n12287 ^ n2722 ;
  assign n20027 = ( ~n1343 & n2263 ) | ( ~n1343 & n20026 ) | ( n2263 & n20026 ) ;
  assign n20028 = n20027 ^ n5843 ^ n3694 ;
  assign n20029 = n6259 ^ n2260 ^ n1292 ;
  assign n20030 = ( n1390 & ~n12759 ) | ( n1390 & n20029 ) | ( ~n12759 & n20029 ) ;
  assign n20031 = ( n1153 & n10200 ) | ( n1153 & ~n20030 ) | ( n10200 & ~n20030 ) ;
  assign n20032 = n20031 ^ n19454 ^ n13759 ;
  assign n20033 = ( n8557 & ~n20028 ) | ( n8557 & n20032 ) | ( ~n20028 & n20032 ) ;
  assign n20034 = ( x34 & n9583 ) | ( x34 & n20033 ) | ( n9583 & n20033 ) ;
  assign n20036 = n13745 ^ n4582 ^ n3837 ;
  assign n20037 = n20036 ^ n9215 ^ n7769 ;
  assign n20035 = ( n2149 & ~n4886 ) | ( n2149 & n9815 ) | ( ~n4886 & n9815 ) ;
  assign n20038 = n20037 ^ n20035 ^ n14507 ;
  assign n20039 = ( n9711 & ~n12349 ) | ( n9711 & n19041 ) | ( ~n12349 & n19041 ) ;
  assign n20040 = ( n4276 & n5108 ) | ( n4276 & n14953 ) | ( n5108 & n14953 ) ;
  assign n20041 = ( n6623 & n19973 ) | ( n6623 & ~n20040 ) | ( n19973 & ~n20040 ) ;
  assign n20045 = n14668 ^ n9544 ^ n1501 ;
  assign n20044 = n9669 ^ n7827 ^ n1528 ;
  assign n20042 = ( n1283 & n6712 ) | ( n1283 & ~n8719 ) | ( n6712 & ~n8719 ) ;
  assign n20043 = ( ~n3343 & n14362 ) | ( ~n3343 & n20042 ) | ( n14362 & n20042 ) ;
  assign n20046 = n20045 ^ n20044 ^ n20043 ;
  assign n20047 = ( n3798 & n3862 ) | ( n3798 & n13803 ) | ( n3862 & n13803 ) ;
  assign n20048 = ( ~n3885 & n5720 ) | ( ~n3885 & n20047 ) | ( n5720 & n20047 ) ;
  assign n20049 = ( n6871 & n14758 ) | ( n6871 & ~n16573 ) | ( n14758 & ~n16573 ) ;
  assign n20050 = ( n18885 & n19165 ) | ( n18885 & n20049 ) | ( n19165 & n20049 ) ;
  assign n20051 = n16803 ^ n15284 ^ n10247 ;
  assign n20052 = ( n1264 & n8772 ) | ( n1264 & ~n11371 ) | ( n8772 & ~n11371 ) ;
  assign n20053 = ( n7158 & n18590 ) | ( n7158 & ~n20052 ) | ( n18590 & ~n20052 ) ;
  assign n20054 = ( n6776 & n20051 ) | ( n6776 & ~n20053 ) | ( n20051 & ~n20053 ) ;
  assign n20055 = ( n3408 & n14614 ) | ( n3408 & n20054 ) | ( n14614 & n20054 ) ;
  assign n20056 = ( ~n956 & n3260 ) | ( ~n956 & n6269 ) | ( n3260 & n6269 ) ;
  assign n20057 = ( n6100 & n7422 ) | ( n6100 & ~n20056 ) | ( n7422 & ~n20056 ) ;
  assign n20058 = n20057 ^ n14935 ^ n12847 ;
  assign n20059 = n18476 ^ n18168 ^ n1425 ;
  assign n20060 = n5118 ^ n4639 ^ n2338 ;
  assign n20061 = n15816 ^ n2367 ^ n858 ;
  assign n20062 = ( n1998 & ~n10164 ) | ( n1998 & n20061 ) | ( ~n10164 & n20061 ) ;
  assign n20063 = ( n3512 & ~n20060 ) | ( n3512 & n20062 ) | ( ~n20060 & n20062 ) ;
  assign n20064 = ( n154 & ~n10243 ) | ( n154 & n20063 ) | ( ~n10243 & n20063 ) ;
  assign n20065 = ( ~n2939 & n17562 ) | ( ~n2939 & n20064 ) | ( n17562 & n20064 ) ;
  assign n20066 = ( n1286 & ~n16107 ) | ( n1286 & n20065 ) | ( ~n16107 & n20065 ) ;
  assign n20067 = ( n831 & ~n1334 ) | ( n831 & n2566 ) | ( ~n1334 & n2566 ) ;
  assign n20068 = n20067 ^ n9801 ^ n9127 ;
  assign n20071 = n13109 ^ n9262 ^ n3469 ;
  assign n20069 = ( n2526 & n8904 ) | ( n2526 & ~n19161 ) | ( n8904 & ~n19161 ) ;
  assign n20070 = n20069 ^ n18416 ^ n8853 ;
  assign n20072 = n20071 ^ n20070 ^ n1501 ;
  assign n20074 = ( ~n3743 & n8714 ) | ( ~n3743 & n9548 ) | ( n8714 & n9548 ) ;
  assign n20073 = ( n9194 & n9611 ) | ( n9194 & n13203 ) | ( n9611 & n13203 ) ;
  assign n20075 = n20074 ^ n20073 ^ n8662 ;
  assign n20076 = ( ~n9195 & n19539 ) | ( ~n9195 & n20075 ) | ( n19539 & n20075 ) ;
  assign n20077 = ( ~n2231 & n3732 ) | ( ~n2231 & n17401 ) | ( n3732 & n17401 ) ;
  assign n20078 = ( ~n4274 & n19263 ) | ( ~n4274 & n20077 ) | ( n19263 & n20077 ) ;
  assign n20079 = ( n2589 & n9807 ) | ( n2589 & ~n14884 ) | ( n9807 & ~n14884 ) ;
  assign n20081 = n11395 ^ n10294 ^ n3937 ;
  assign n20080 = n13961 ^ n11903 ^ n11696 ;
  assign n20082 = n20081 ^ n20080 ^ n1390 ;
  assign n20083 = ( ~n3237 & n11795 ) | ( ~n3237 & n12738 ) | ( n11795 & n12738 ) ;
  assign n20084 = n17288 ^ n5142 ^ n2673 ;
  assign n20085 = ( n7494 & n13989 ) | ( n7494 & ~n14668 ) | ( n13989 & ~n14668 ) ;
  assign n20086 = ( n334 & ~n9863 ) | ( n334 & n20085 ) | ( ~n9863 & n20085 ) ;
  assign n20087 = n20086 ^ n18997 ^ n8900 ;
  assign n20088 = n15033 ^ n4625 ^ n187 ;
  assign n20089 = n11697 ^ n4566 ^ n736 ;
  assign n20090 = n9966 ^ n8821 ^ n6346 ;
  assign n20091 = ( n894 & n899 ) | ( n894 & n6819 ) | ( n899 & n6819 ) ;
  assign n20092 = n20091 ^ n13720 ^ n3931 ;
  assign n20093 = ( n3829 & n4697 ) | ( n3829 & n12591 ) | ( n4697 & n12591 ) ;
  assign n20096 = n7250 ^ n3189 ^ n1750 ;
  assign n20095 = ( n133 & ~n15202 ) | ( n133 & n16836 ) | ( ~n15202 & n16836 ) ;
  assign n20094 = ( ~n2786 & n9278 ) | ( ~n2786 & n10108 ) | ( n9278 & n10108 ) ;
  assign n20097 = n20096 ^ n20095 ^ n20094 ;
  assign n20106 = ( n4087 & ~n5195 ) | ( n4087 & n13072 ) | ( ~n5195 & n13072 ) ;
  assign n20107 = n20106 ^ n3820 ^ n3159 ;
  assign n20103 = ( ~n4318 & n5633 ) | ( ~n4318 & n9164 ) | ( n5633 & n9164 ) ;
  assign n20104 = n20103 ^ n10318 ^ n4675 ;
  assign n20100 = ( ~n2069 & n3063 ) | ( ~n2069 & n5518 ) | ( n3063 & n5518 ) ;
  assign n20099 = n13938 ^ n7043 ^ n1073 ;
  assign n20101 = n20100 ^ n20099 ^ n4700 ;
  assign n20098 = ( n3610 & n5900 ) | ( n3610 & n15268 ) | ( n5900 & n15268 ) ;
  assign n20102 = n20101 ^ n20098 ^ n3442 ;
  assign n20105 = n20104 ^ n20102 ^ n6174 ;
  assign n20108 = n20107 ^ n20105 ^ n14252 ;
  assign n20109 = n17069 ^ n6147 ^ n559 ;
  assign n20110 = n19414 ^ n18365 ^ n7660 ;
  assign n20111 = ( n19193 & ~n20109 ) | ( n19193 & n20110 ) | ( ~n20109 & n20110 ) ;
  assign n20112 = ( n1853 & ~n8497 ) | ( n1853 & n8789 ) | ( ~n8497 & n8789 ) ;
  assign n20113 = n20112 ^ n8998 ^ n4350 ;
  assign n20114 = ( n5402 & ~n5542 ) | ( n5402 & n20113 ) | ( ~n5542 & n20113 ) ;
  assign n20115 = ( ~n1388 & n3638 ) | ( ~n1388 & n20114 ) | ( n3638 & n20114 ) ;
  assign n20116 = ( n1973 & ~n12239 ) | ( n1973 & n13114 ) | ( ~n12239 & n13114 ) ;
  assign n20117 = n14762 ^ n12083 ^ n2297 ;
  assign n20118 = n13184 ^ n5736 ^ n4377 ;
  assign n20119 = n13909 ^ n10476 ^ n2074 ;
  assign n20120 = ( n6074 & n12824 ) | ( n6074 & ~n20119 ) | ( n12824 & ~n20119 ) ;
  assign n20121 = n7985 ^ n4531 ^ n1231 ;
  assign n20122 = ( n2185 & ~n8195 ) | ( n2185 & n20121 ) | ( ~n8195 & n20121 ) ;
  assign n20123 = ( n2122 & n20120 ) | ( n2122 & n20122 ) | ( n20120 & n20122 ) ;
  assign n20125 = n4756 ^ n4442 ^ x10 ;
  assign n20124 = n18267 ^ n9781 ^ n1807 ;
  assign n20126 = n20125 ^ n20124 ^ n13373 ;
  assign n20127 = n17080 ^ n515 ^ x117 ;
  assign n20128 = n13655 ^ n7346 ^ n186 ;
  assign n20129 = ( ~n2447 & n20127 ) | ( ~n2447 & n20128 ) | ( n20127 & n20128 ) ;
  assign n20130 = n17279 ^ n9493 ^ n5687 ;
  assign n20131 = ( n4494 & n7880 ) | ( n4494 & n8517 ) | ( n7880 & n8517 ) ;
  assign n20132 = ( n450 & n1515 ) | ( n450 & ~n10945 ) | ( n1515 & ~n10945 ) ;
  assign n20133 = n20132 ^ n17895 ^ n13944 ;
  assign n20134 = n20133 ^ n14739 ^ n7109 ;
  assign n20135 = ( ~n668 & n11080 ) | ( ~n668 & n20134 ) | ( n11080 & n20134 ) ;
  assign n20136 = n12228 ^ n4602 ^ n2110 ;
  assign n20137 = n20136 ^ n15336 ^ n5309 ;
  assign n20138 = ( ~n8638 & n11815 ) | ( ~n8638 & n18302 ) | ( n11815 & n18302 ) ;
  assign n20139 = ( n1553 & n3285 ) | ( n1553 & n20138 ) | ( n3285 & n20138 ) ;
  assign n20140 = ( n250 & n3710 ) | ( n250 & n4451 ) | ( n3710 & n4451 ) ;
  assign n20141 = ( n3827 & n8702 ) | ( n3827 & ~n9479 ) | ( n8702 & ~n9479 ) ;
  assign n20142 = ( n14654 & ~n20140 ) | ( n14654 & n20141 ) | ( ~n20140 & n20141 ) ;
  assign n20143 = n10902 ^ n8384 ^ n6723 ;
  assign n20144 = n20143 ^ n5291 ^ n3284 ;
  assign n20145 = ( n6913 & n12713 ) | ( n6913 & n16104 ) | ( n12713 & n16104 ) ;
  assign n20153 = ( n1162 & ~n5031 ) | ( n1162 & n15602 ) | ( ~n5031 & n15602 ) ;
  assign n20154 = n20153 ^ n10091 ^ n4415 ;
  assign n20155 = ( ~n3923 & n4462 ) | ( ~n3923 & n20154 ) | ( n4462 & n20154 ) ;
  assign n20146 = ( n1092 & ~n2981 ) | ( n1092 & n5110 ) | ( ~n2981 & n5110 ) ;
  assign n20147 = ( n5721 & ~n10319 ) | ( n5721 & n20146 ) | ( ~n10319 & n20146 ) ;
  assign n20148 = n5086 ^ n2366 ^ n1760 ;
  assign n20149 = ( n3047 & n20147 ) | ( n3047 & ~n20148 ) | ( n20147 & ~n20148 ) ;
  assign n20150 = ( n2103 & n12879 ) | ( n2103 & ~n20149 ) | ( n12879 & ~n20149 ) ;
  assign n20151 = ( ~n1492 & n14636 ) | ( ~n1492 & n20150 ) | ( n14636 & n20150 ) ;
  assign n20152 = ( n4440 & n5702 ) | ( n4440 & n20151 ) | ( n5702 & n20151 ) ;
  assign n20156 = n20155 ^ n20152 ^ n10803 ;
  assign n20160 = ( n2524 & n6501 ) | ( n2524 & n10690 ) | ( n6501 & n10690 ) ;
  assign n20157 = n6204 ^ n5505 ^ n4225 ;
  assign n20158 = n8435 ^ n2160 ^ n2028 ;
  assign n20159 = ( ~n4843 & n20157 ) | ( ~n4843 & n20158 ) | ( n20157 & n20158 ) ;
  assign n20161 = n20160 ^ n20159 ^ n423 ;
  assign n20163 = ( ~x119 & n4440 ) | ( ~x119 & n7253 ) | ( n4440 & n7253 ) ;
  assign n20162 = n10890 ^ n6406 ^ n3296 ;
  assign n20164 = n20163 ^ n20162 ^ n15120 ;
  assign n20165 = n20060 ^ n3434 ^ n1446 ;
  assign n20166 = ( n7501 & n9538 ) | ( n7501 & ~n20165 ) | ( n9538 & ~n20165 ) ;
  assign n20167 = ( n5364 & n9897 ) | ( n5364 & ~n19528 ) | ( n9897 & ~n19528 ) ;
  assign n20168 = ( ~n3373 & n5072 ) | ( ~n3373 & n20167 ) | ( n5072 & n20167 ) ;
  assign n20169 = ( ~n4919 & n14631 ) | ( ~n4919 & n16705 ) | ( n14631 & n16705 ) ;
  assign n20170 = ( n10649 & n15887 ) | ( n10649 & n20169 ) | ( n15887 & n20169 ) ;
  assign n20171 = ( ~n11615 & n18346 ) | ( ~n11615 & n20170 ) | ( n18346 & n20170 ) ;
  assign n20172 = n8900 ^ n8615 ^ n5200 ;
  assign n20173 = ( ~n5371 & n17655 ) | ( ~n5371 & n20172 ) | ( n17655 & n20172 ) ;
  assign n20174 = ( n18658 & n19064 ) | ( n18658 & ~n20173 ) | ( n19064 & ~n20173 ) ;
  assign n20175 = n20174 ^ n8521 ^ n2068 ;
  assign n20176 = n10949 ^ n10903 ^ n8778 ;
  assign n20177 = n20176 ^ n9617 ^ n1104 ;
  assign n20178 = n20177 ^ n7295 ^ n3716 ;
  assign n20179 = ( n8298 & n11516 ) | ( n8298 & ~n16586 ) | ( n11516 & ~n16586 ) ;
  assign n20180 = n20179 ^ n8230 ^ n2829 ;
  assign n20181 = ( ~x103 & n7410 ) | ( ~x103 & n10673 ) | ( n7410 & n10673 ) ;
  assign n20186 = ( n6054 & ~n11556 ) | ( n6054 & n16516 ) | ( ~n11556 & n16516 ) ;
  assign n20182 = ( n304 & ~n2108 ) | ( n304 & n7802 ) | ( ~n2108 & n7802 ) ;
  assign n20183 = ( n1941 & ~n9472 ) | ( n1941 & n10174 ) | ( ~n9472 & n10174 ) ;
  assign n20184 = ( n4065 & n7767 ) | ( n4065 & n20183 ) | ( n7767 & n20183 ) ;
  assign n20185 = ( n5150 & ~n20182 ) | ( n5150 & n20184 ) | ( ~n20182 & n20184 ) ;
  assign n20187 = n20186 ^ n20185 ^ n5625 ;
  assign n20188 = ( n8911 & n20181 ) | ( n8911 & n20187 ) | ( n20181 & n20187 ) ;
  assign n20189 = n20188 ^ n13944 ^ n11123 ;
  assign n20190 = ( n20178 & n20180 ) | ( n20178 & ~n20189 ) | ( n20180 & ~n20189 ) ;
  assign n20191 = n15435 ^ n12885 ^ n10451 ;
  assign n20192 = ( n3441 & ~n4466 ) | ( n3441 & n10050 ) | ( ~n4466 & n10050 ) ;
  assign n20193 = n20192 ^ n7248 ^ n5891 ;
  assign n20194 = ( n2006 & n15358 ) | ( n2006 & n20193 ) | ( n15358 & n20193 ) ;
  assign n20195 = n20194 ^ n3256 ^ n2388 ;
  assign n20196 = n20195 ^ n17708 ^ n11731 ;
  assign n20197 = ( ~n9413 & n20191 ) | ( ~n9413 & n20196 ) | ( n20191 & n20196 ) ;
  assign n20198 = ( n1475 & n10331 ) | ( n1475 & ~n20197 ) | ( n10331 & ~n20197 ) ;
  assign n20199 = ( n8199 & n8835 ) | ( n8199 & n11737 ) | ( n8835 & n11737 ) ;
  assign n20200 = n20199 ^ n8553 ^ n1069 ;
  assign n20201 = n16254 ^ n12733 ^ n355 ;
  assign n20202 = ( n215 & ~n6630 ) | ( n215 & n6989 ) | ( ~n6630 & n6989 ) ;
  assign n20203 = n20202 ^ n16075 ^ n13817 ;
  assign n20204 = ( n4783 & ~n14578 ) | ( n4783 & n19668 ) | ( ~n14578 & n19668 ) ;
  assign n20205 = ( n197 & n6997 ) | ( n197 & n10727 ) | ( n6997 & n10727 ) ;
  assign n20211 = n12859 ^ n2827 ^ n293 ;
  assign n20210 = n12444 ^ n8300 ^ n3892 ;
  assign n20206 = ( n1524 & ~n7564 ) | ( n1524 & n18496 ) | ( ~n7564 & n18496 ) ;
  assign n20207 = n20206 ^ n5825 ^ n897 ;
  assign n20208 = n20207 ^ n7745 ^ n5451 ;
  assign n20209 = n20208 ^ n5786 ^ n2827 ;
  assign n20212 = n20211 ^ n20210 ^ n20209 ;
  assign n20213 = ( n518 & ~n7315 ) | ( n518 & n14867 ) | ( ~n7315 & n14867 ) ;
  assign n20214 = n20213 ^ n5084 ^ n4785 ;
  assign n20215 = ( n6206 & ~n11519 ) | ( n6206 & n12767 ) | ( ~n11519 & n12767 ) ;
  assign n20216 = n20215 ^ n16630 ^ n14320 ;
  assign n20218 = ( n551 & ~n2529 ) | ( n551 & n3412 ) | ( ~n2529 & n3412 ) ;
  assign n20217 = ( n9138 & n14568 ) | ( n9138 & ~n15271 ) | ( n14568 & ~n15271 ) ;
  assign n20219 = n20218 ^ n20217 ^ n732 ;
  assign n20220 = ( n4415 & n10040 ) | ( n4415 & ~n15506 ) | ( n10040 & ~n15506 ) ;
  assign n20221 = ( ~n1555 & n4622 ) | ( ~n1555 & n20220 ) | ( n4622 & n20220 ) ;
  assign n20222 = ( ~n15727 & n20219 ) | ( ~n15727 & n20221 ) | ( n20219 & n20221 ) ;
  assign n20223 = ( n2212 & n2998 ) | ( n2212 & ~n7215 ) | ( n2998 & ~n7215 ) ;
  assign n20224 = n19052 ^ n2774 ^ n1642 ;
  assign n20225 = ( n15714 & n20223 ) | ( n15714 & n20224 ) | ( n20223 & n20224 ) ;
  assign n20231 = n11820 ^ n1236 ^ n730 ;
  assign n20227 = ( n4312 & n8000 ) | ( n4312 & n17165 ) | ( n8000 & n17165 ) ;
  assign n20228 = ( ~n8217 & n8557 ) | ( ~n8217 & n20227 ) | ( n8557 & n20227 ) ;
  assign n20226 = ( n3962 & ~n12276 ) | ( n3962 & n19780 ) | ( ~n12276 & n19780 ) ;
  assign n20229 = n20228 ^ n20226 ^ n7474 ;
  assign n20230 = ( ~n10248 & n13045 ) | ( ~n10248 & n20229 ) | ( n13045 & n20229 ) ;
  assign n20232 = n20231 ^ n20230 ^ n6806 ;
  assign n20237 = n16586 ^ n7347 ^ n3844 ;
  assign n20236 = ( n903 & n6216 ) | ( n903 & n12922 ) | ( n6216 & n12922 ) ;
  assign n20233 = n7655 ^ n3750 ^ n1927 ;
  assign n20234 = n20233 ^ n6826 ^ n1480 ;
  assign n20235 = n20234 ^ n6266 ^ n3973 ;
  assign n20238 = n20237 ^ n20236 ^ n20235 ;
  assign n20242 = n15680 ^ n13000 ^ n7489 ;
  assign n20239 = ( n3247 & ~n5862 ) | ( n3247 & n7712 ) | ( ~n5862 & n7712 ) ;
  assign n20240 = n20239 ^ n11318 ^ n1056 ;
  assign n20241 = n20240 ^ n12638 ^ n1387 ;
  assign n20243 = n20242 ^ n20241 ^ n11342 ;
  assign n20244 = n20243 ^ n17408 ^ n16453 ;
  assign n20246 = n4323 ^ n4003 ^ n811 ;
  assign n20245 = n10580 ^ n4613 ^ n3946 ;
  assign n20247 = n20246 ^ n20245 ^ n8386 ;
  assign n20248 = ( ~n4478 & n6111 ) | ( ~n4478 & n9525 ) | ( n6111 & n9525 ) ;
  assign n20249 = n11731 ^ n3939 ^ n791 ;
  assign n20250 = ( ~n5043 & n9488 ) | ( ~n5043 & n20249 ) | ( n9488 & n20249 ) ;
  assign n20251 = ( n5712 & ~n14129 ) | ( n5712 & n20250 ) | ( ~n14129 & n20250 ) ;
  assign n20252 = n11744 ^ n5832 ^ n1460 ;
  assign n20253 = ( n1978 & ~n2188 ) | ( n1978 & n6302 ) | ( ~n2188 & n6302 ) ;
  assign n20254 = n20253 ^ n19776 ^ n7593 ;
  assign n20255 = n20254 ^ n11344 ^ n3277 ;
  assign n20256 = ( n8980 & ~n9223 ) | ( n8980 & n20255 ) | ( ~n9223 & n20255 ) ;
  assign n20257 = ( n631 & ~n20252 ) | ( n631 & n20256 ) | ( ~n20252 & n20256 ) ;
  assign n20258 = n14974 ^ n12837 ^ n4507 ;
  assign n20259 = ( ~n3427 & n6315 ) | ( ~n3427 & n18066 ) | ( n6315 & n18066 ) ;
  assign n20260 = n20259 ^ n13713 ^ n8474 ;
  assign n20261 = ( n6937 & n10253 ) | ( n6937 & ~n14639 ) | ( n10253 & ~n14639 ) ;
  assign n20262 = ( n15814 & n15864 ) | ( n15814 & n20261 ) | ( n15864 & n20261 ) ;
  assign n20265 = n7615 ^ n7202 ^ n2126 ;
  assign n20263 = n10956 ^ n2874 ^ n1357 ;
  assign n20264 = n20263 ^ n8267 ^ n454 ;
  assign n20266 = n20265 ^ n20264 ^ n19857 ;
  assign n20267 = ( n4661 & ~n18293 ) | ( n4661 & n19934 ) | ( ~n18293 & n19934 ) ;
  assign n20268 = n20267 ^ n16376 ^ n15443 ;
  assign n20269 = n15046 ^ n12595 ^ n5013 ;
  assign n20270 = ( ~n1237 & n3244 ) | ( ~n1237 & n17551 ) | ( n3244 & n17551 ) ;
  assign n20271 = n17622 ^ n15175 ^ n6184 ;
  assign n20272 = ( n4055 & n8012 ) | ( n4055 & n18523 ) | ( n8012 & n18523 ) ;
  assign n20273 = ( ~n16069 & n20271 ) | ( ~n16069 & n20272 ) | ( n20271 & n20272 ) ;
  assign n20274 = ( x83 & ~n2608 ) | ( x83 & n16921 ) | ( ~n2608 & n16921 ) ;
  assign n20275 = n20274 ^ n6340 ^ n5991 ;
  assign n20276 = ( n1466 & n3085 ) | ( n1466 & n3655 ) | ( n3085 & n3655 ) ;
  assign n20277 = n20276 ^ n17744 ^ n17541 ;
  assign n20278 = n7570 ^ n1880 ^ n909 ;
  assign n20279 = ( ~n1521 & n7907 ) | ( ~n1521 & n20278 ) | ( n7907 & n20278 ) ;
  assign n20280 = ( n1400 & n1781 ) | ( n1400 & n15508 ) | ( n1781 & n15508 ) ;
  assign n20281 = ( n7980 & n14604 ) | ( n7980 & ~n20280 ) | ( n14604 & ~n20280 ) ;
  assign n20282 = ( ~n16182 & n20279 ) | ( ~n16182 & n20281 ) | ( n20279 & n20281 ) ;
  assign n20283 = ( n406 & n451 ) | ( n406 & ~n1835 ) | ( n451 & ~n1835 ) ;
  assign n20284 = ( n3327 & n3550 ) | ( n3327 & n20283 ) | ( n3550 & n20283 ) ;
  assign n20285 = n20284 ^ n14831 ^ n7263 ;
  assign n20286 = n20285 ^ n17640 ^ n2669 ;
  assign n20287 = ( n3349 & ~n6636 ) | ( n3349 & n20286 ) | ( ~n6636 & n20286 ) ;
  assign n20289 = ( n3461 & n3632 ) | ( n3461 & ~n5706 ) | ( n3632 & ~n5706 ) ;
  assign n20288 = ( n557 & ~n2357 ) | ( n557 & n7855 ) | ( ~n2357 & n7855 ) ;
  assign n20290 = n20289 ^ n20288 ^ n8088 ;
  assign n20291 = ( ~n6672 & n11981 ) | ( ~n6672 & n18478 ) | ( n11981 & n18478 ) ;
  assign n20292 = ( n549 & n4898 ) | ( n549 & n8723 ) | ( n4898 & n8723 ) ;
  assign n20295 = n11952 ^ n10829 ^ n130 ;
  assign n20294 = ( n11551 & n11813 ) | ( n11551 & n16630 ) | ( n11813 & n16630 ) ;
  assign n20293 = n18648 ^ n14152 ^ n8665 ;
  assign n20296 = n20295 ^ n20294 ^ n20293 ;
  assign n20297 = n9778 ^ n9028 ^ n3789 ;
  assign n20298 = ( ~n2539 & n2868 ) | ( ~n2539 & n16149 ) | ( n2868 & n16149 ) ;
  assign n20299 = ( n2660 & n5438 ) | ( n2660 & n10794 ) | ( n5438 & n10794 ) ;
  assign n20300 = ( n4207 & n20298 ) | ( n4207 & n20299 ) | ( n20298 & n20299 ) ;
  assign n20301 = n12615 ^ n10915 ^ n5967 ;
  assign n20302 = n20301 ^ n11681 ^ n2355 ;
  assign n20305 = ( n6531 & n6571 ) | ( n6531 & n16218 ) | ( n6571 & n16218 ) ;
  assign n20306 = n20305 ^ n19113 ^ n691 ;
  assign n20304 = ( n3139 & n12665 ) | ( n3139 & ~n12788 ) | ( n12665 & ~n12788 ) ;
  assign n20303 = ( n3978 & n10334 ) | ( n3978 & n14916 ) | ( n10334 & n14916 ) ;
  assign n20307 = n20306 ^ n20304 ^ n20303 ;
  assign n20308 = n18487 ^ n5819 ^ n3748 ;
  assign n20309 = n6836 ^ n2703 ^ n637 ;
  assign n20310 = ( x36 & ~n20308 ) | ( x36 & n20309 ) | ( ~n20308 & n20309 ) ;
  assign n20311 = n20310 ^ n9492 ^ n376 ;
  assign n20312 = ( n2724 & ~n18958 ) | ( n2724 & n19412 ) | ( ~n18958 & n19412 ) ;
  assign n20313 = ( ~n14651 & n20311 ) | ( ~n14651 & n20312 ) | ( n20311 & n20312 ) ;
  assign n20314 = n18122 ^ n12343 ^ n11378 ;
  assign n20315 = n20314 ^ n7183 ^ n1082 ;
  assign n20316 = n17439 ^ n14949 ^ n7331 ;
  assign n20317 = n20316 ^ n19747 ^ n4720 ;
  assign n20318 = ( n1834 & n14630 ) | ( n1834 & ~n17411 ) | ( n14630 & ~n17411 ) ;
  assign n20319 = ( n237 & n6392 ) | ( n237 & n20318 ) | ( n6392 & n20318 ) ;
  assign n20320 = ( ~n942 & n1327 ) | ( ~n942 & n7780 ) | ( n1327 & n7780 ) ;
  assign n20321 = n20320 ^ n8404 ^ n1613 ;
  assign n20322 = ( n4156 & ~n10120 ) | ( n4156 & n20321 ) | ( ~n10120 & n20321 ) ;
  assign n20323 = n20322 ^ n16282 ^ n15424 ;
  assign n20324 = ( n14973 & n14982 ) | ( n14973 & ~n20323 ) | ( n14982 & ~n20323 ) ;
  assign n20325 = n9545 ^ n7427 ^ n483 ;
  assign n20326 = ( n5954 & n6444 ) | ( n5954 & ~n20325 ) | ( n6444 & ~n20325 ) ;
  assign n20327 = ( n2362 & n3730 ) | ( n2362 & n10426 ) | ( n3730 & n10426 ) ;
  assign n20328 = ( n6771 & n7426 ) | ( n6771 & ~n15423 ) | ( n7426 & ~n15423 ) ;
  assign n20329 = ( ~n16881 & n18211 ) | ( ~n16881 & n20328 ) | ( n18211 & n20328 ) ;
  assign n20330 = ( n20326 & ~n20327 ) | ( n20326 & n20329 ) | ( ~n20327 & n20329 ) ;
  assign n20331 = ( n403 & n2088 ) | ( n403 & ~n6165 ) | ( n2088 & ~n6165 ) ;
  assign n20332 = ( ~n2459 & n8516 ) | ( ~n2459 & n11569 ) | ( n8516 & n11569 ) ;
  assign n20333 = ( n719 & n20331 ) | ( n719 & n20332 ) | ( n20331 & n20332 ) ;
  assign n20335 = ( n3321 & n3673 ) | ( n3321 & ~n5357 ) | ( n3673 & ~n5357 ) ;
  assign n20334 = n19312 ^ n12779 ^ n2327 ;
  assign n20336 = n20335 ^ n20334 ^ n7076 ;
  assign n20337 = ( n16689 & n18516 ) | ( n16689 & ~n20336 ) | ( n18516 & ~n20336 ) ;
  assign n20338 = n6093 ^ n1185 ^ n962 ;
  assign n20339 = n20338 ^ n19612 ^ n12100 ;
  assign n20340 = n20339 ^ n12185 ^ n7090 ;
  assign n20341 = ( n11947 & n20337 ) | ( n11947 & ~n20340 ) | ( n20337 & ~n20340 ) ;
  assign n20342 = n11871 ^ n6358 ^ n5480 ;
  assign n20343 = n20342 ^ n13815 ^ n7389 ;
  assign n20344 = ( n4454 & n5180 ) | ( n4454 & n11342 ) | ( n5180 & n11342 ) ;
  assign n20345 = n20344 ^ n5347 ^ n1132 ;
  assign n20346 = n18308 ^ n4587 ^ n2069 ;
  assign n20347 = n13023 ^ n10278 ^ n4378 ;
  assign n20348 = ( n1418 & ~n10013 ) | ( n1418 & n20347 ) | ( ~n10013 & n20347 ) ;
  assign n20349 = ( n686 & ~n12170 ) | ( n686 & n14692 ) | ( ~n12170 & n14692 ) ;
  assign n20350 = ( ~n5857 & n14058 ) | ( ~n5857 & n20349 ) | ( n14058 & n20349 ) ;
  assign n20351 = n20350 ^ n6829 ^ x23 ;
  assign n20352 = n17780 ^ n16229 ^ n12833 ;
  assign n20353 = ( n4661 & n7321 ) | ( n4661 & ~n9961 ) | ( n7321 & ~n9961 ) ;
  assign n20354 = n20353 ^ n5252 ^ n4156 ;
  assign n20355 = ( ~n2152 & n8899 ) | ( ~n2152 & n10788 ) | ( n8899 & n10788 ) ;
  assign n20356 = ( n1704 & n4301 ) | ( n1704 & n9438 ) | ( n4301 & n9438 ) ;
  assign n20357 = n20356 ^ n15841 ^ n4617 ;
  assign n20358 = n20357 ^ n4180 ^ n1820 ;
  assign n20359 = ( n6391 & n20355 ) | ( n6391 & ~n20358 ) | ( n20355 & ~n20358 ) ;
  assign n20360 = ( ~n12323 & n17722 ) | ( ~n12323 & n19276 ) | ( n17722 & n19276 ) ;
  assign n20361 = ( n443 & n484 ) | ( n443 & ~n16498 ) | ( n484 & ~n16498 ) ;
  assign n20362 = ( n4450 & n18265 ) | ( n4450 & ~n20361 ) | ( n18265 & ~n20361 ) ;
  assign n20363 = ( n1286 & n4518 ) | ( n1286 & n13139 ) | ( n4518 & n13139 ) ;
  assign n20364 = ( n789 & n2817 ) | ( n789 & n20363 ) | ( n2817 & n20363 ) ;
  assign n20365 = ( ~n4676 & n8648 ) | ( ~n4676 & n12260 ) | ( n8648 & n12260 ) ;
  assign n20366 = ( ~n5618 & n6987 ) | ( ~n5618 & n11641 ) | ( n6987 & n11641 ) ;
  assign n20367 = ( n5922 & n16158 ) | ( n5922 & ~n20366 ) | ( n16158 & ~n20366 ) ;
  assign n20370 = n5851 ^ n4266 ^ n1811 ;
  assign n20368 = n8242 ^ n6534 ^ n1851 ;
  assign n20369 = n20368 ^ n17850 ^ n8878 ;
  assign n20371 = n20370 ^ n20369 ^ n16168 ;
  assign n20372 = ( ~n6956 & n18997 ) | ( ~n6956 & n19053 ) | ( n18997 & n19053 ) ;
  assign n20373 = ( n1773 & n12099 ) | ( n1773 & ~n12590 ) | ( n12099 & ~n12590 ) ;
  assign n20374 = ( n3919 & n8163 ) | ( n3919 & ~n17555 ) | ( n8163 & ~n17555 ) ;
  assign n20375 = ( n1170 & n2195 ) | ( n1170 & ~n6631 ) | ( n2195 & ~n6631 ) ;
  assign n20376 = ( n6070 & n11020 ) | ( n6070 & n12875 ) | ( n11020 & n12875 ) ;
  assign n20377 = n17812 ^ n8559 ^ n6366 ;
  assign n20378 = ( ~n20375 & n20376 ) | ( ~n20375 & n20377 ) | ( n20376 & n20377 ) ;
  assign n20381 = n14445 ^ n14246 ^ n1361 ;
  assign n20382 = n20381 ^ n13835 ^ n5955 ;
  assign n20379 = ( n1273 & n1597 ) | ( n1273 & ~n3893 ) | ( n1597 & ~n3893 ) ;
  assign n20380 = ( ~n6869 & n18112 ) | ( ~n6869 & n20379 ) | ( n18112 & n20379 ) ;
  assign n20383 = n20382 ^ n20380 ^ n6857 ;
  assign n20384 = n3591 ^ n3220 ^ n1032 ;
  assign n20385 = ( n7256 & ~n14054 ) | ( n7256 & n16844 ) | ( ~n14054 & n16844 ) ;
  assign n20386 = ( n12632 & ~n20384 ) | ( n12632 & n20385 ) | ( ~n20384 & n20385 ) ;
  assign n20387 = n8349 ^ n6926 ^ n3806 ;
  assign n20388 = n19371 ^ n8767 ^ n8549 ;
  assign n20390 = ( n2092 & ~n5159 ) | ( n2092 & n8786 ) | ( ~n5159 & n8786 ) ;
  assign n20391 = ( ~n535 & n10521 ) | ( ~n535 & n15946 ) | ( n10521 & n15946 ) ;
  assign n20392 = ( n19047 & n20390 ) | ( n19047 & ~n20391 ) | ( n20390 & ~n20391 ) ;
  assign n20389 = n15694 ^ n3870 ^ n1681 ;
  assign n20393 = n20392 ^ n20389 ^ n1216 ;
  assign n20394 = ( n7751 & n9418 ) | ( n7751 & ~n19137 ) | ( n9418 & ~n19137 ) ;
  assign n20395 = ( ~n4608 & n16689 ) | ( ~n4608 & n19803 ) | ( n16689 & n19803 ) ;
  assign n20396 = ( ~n3938 & n13521 ) | ( ~n3938 & n17287 ) | ( n13521 & n17287 ) ;
  assign n20397 = n20396 ^ n12181 ^ n980 ;
  assign n20398 = ( ~n5111 & n12933 ) | ( ~n5111 & n15723 ) | ( n12933 & n15723 ) ;
  assign n20399 = ( n3585 & ~n11158 ) | ( n3585 & n20398 ) | ( ~n11158 & n20398 ) ;
  assign n20403 = n14312 ^ n3743 ^ n439 ;
  assign n20402 = ( n2609 & ~n6361 ) | ( n2609 & n13301 ) | ( ~n6361 & n13301 ) ;
  assign n20400 = ( n5555 & ~n6317 ) | ( n5555 & n17175 ) | ( ~n6317 & n17175 ) ;
  assign n20401 = ( n4422 & n6076 ) | ( n4422 & n20400 ) | ( n6076 & n20400 ) ;
  assign n20404 = n20403 ^ n20402 ^ n20401 ;
  assign n20405 = ( n5469 & ~n6234 ) | ( n5469 & n11623 ) | ( ~n6234 & n11623 ) ;
  assign n20406 = ( ~n8463 & n14501 ) | ( ~n8463 & n17006 ) | ( n14501 & n17006 ) ;
  assign n20407 = ( n10926 & n13923 ) | ( n10926 & ~n20406 ) | ( n13923 & ~n20406 ) ;
  assign n20408 = ( n341 & n12444 ) | ( n341 & ~n14191 ) | ( n12444 & ~n14191 ) ;
  assign n20409 = n17190 ^ n11202 ^ n867 ;
  assign n20410 = ( n15790 & n20408 ) | ( n15790 & ~n20409 ) | ( n20408 & ~n20409 ) ;
  assign n20411 = ( n1159 & ~n8570 ) | ( n1159 & n20410 ) | ( ~n8570 & n20410 ) ;
  assign n20412 = ( ~n20405 & n20407 ) | ( ~n20405 & n20411 ) | ( n20407 & n20411 ) ;
  assign n20413 = ( n2087 & n8392 ) | ( n2087 & ~n10224 ) | ( n8392 & ~n10224 ) ;
  assign n20414 = n9834 ^ n6981 ^ n4447 ;
  assign n20415 = n20414 ^ n18327 ^ n6047 ;
  assign n20416 = n12156 ^ n9113 ^ n7975 ;
  assign n20417 = ( n459 & n6191 ) | ( n459 & ~n17668 ) | ( n6191 & ~n17668 ) ;
  assign n20418 = ( n5972 & ~n20416 ) | ( n5972 & n20417 ) | ( ~n20416 & n20417 ) ;
  assign n20419 = ( ~n803 & n12897 ) | ( ~n803 & n19774 ) | ( n12897 & n19774 ) ;
  assign n20420 = n20419 ^ n18226 ^ n17484 ;
  assign n20421 = ( ~n6138 & n16927 ) | ( ~n6138 & n20420 ) | ( n16927 & n20420 ) ;
  assign n20422 = n13437 ^ n7813 ^ n3327 ;
  assign n20423 = n20422 ^ n12493 ^ n8011 ;
  assign n20424 = ( n3493 & n8601 ) | ( n3493 & n14109 ) | ( n8601 & n14109 ) ;
  assign n20425 = ( ~n4083 & n4084 ) | ( ~n4083 & n11215 ) | ( n4084 & n11215 ) ;
  assign n20426 = n20425 ^ n8745 ^ n1931 ;
  assign n20427 = n20426 ^ n19265 ^ n7845 ;
  assign n20428 = ( n713 & ~n10522 ) | ( n713 & n18403 ) | ( ~n10522 & n18403 ) ;
  assign n20429 = n20428 ^ n2050 ^ n1493 ;
  assign n20430 = ( n4929 & ~n16519 ) | ( n4929 & n20429 ) | ( ~n16519 & n20429 ) ;
  assign n20431 = n13022 ^ n5366 ^ n739 ;
  assign n20432 = ( n7200 & n10336 ) | ( n7200 & n20431 ) | ( n10336 & n20431 ) ;
  assign n20433 = ( n8905 & ~n13647 ) | ( n8905 & n15250 ) | ( ~n13647 & n15250 ) ;
  assign n20434 = n20433 ^ n12587 ^ n6274 ;
  assign n20435 = ( ~n782 & n2951 ) | ( ~n782 & n3355 ) | ( n2951 & n3355 ) ;
  assign n20436 = n20435 ^ n12349 ^ n7804 ;
  assign n20437 = ( ~n3114 & n4624 ) | ( ~n3114 & n13197 ) | ( n4624 & n13197 ) ;
  assign n20438 = ( n147 & n8790 ) | ( n147 & ~n10258 ) | ( n8790 & ~n10258 ) ;
  assign n20439 = ( n11793 & ~n15417 ) | ( n11793 & n20438 ) | ( ~n15417 & n20438 ) ;
  assign n20440 = n20439 ^ n2910 ^ n758 ;
  assign n20441 = n19306 ^ n19168 ^ n12528 ;
  assign n20442 = n20441 ^ n8878 ^ n5126 ;
  assign n20443 = n14887 ^ n6826 ^ n6304 ;
  assign n20444 = n2087 ^ n1584 ^ n1222 ;
  assign n20445 = ( n3185 & n18191 ) | ( n3185 & n20444 ) | ( n18191 & n20444 ) ;
  assign n20446 = n20445 ^ n18020 ^ n15284 ;
  assign n20448 = n15787 ^ n10879 ^ n10039 ;
  assign n20447 = n17460 ^ n13232 ^ x56 ;
  assign n20449 = n20448 ^ n20447 ^ n746 ;
  assign n20451 = ( n2591 & n9267 ) | ( n2591 & ~n9849 ) | ( n9267 & ~n9849 ) ;
  assign n20450 = ( n7685 & n12850 ) | ( n7685 & n20028 ) | ( n12850 & n20028 ) ;
  assign n20452 = n20451 ^ n20450 ^ n18209 ;
  assign n20454 = n4848 ^ n898 ^ n286 ;
  assign n20453 = ( ~n841 & n11534 ) | ( ~n841 & n13000 ) | ( n11534 & n13000 ) ;
  assign n20455 = n20454 ^ n20453 ^ n8227 ;
  assign n20456 = ( n18161 & n20452 ) | ( n18161 & n20455 ) | ( n20452 & n20455 ) ;
  assign n20457 = ( n683 & ~n20075 ) | ( n683 & n20456 ) | ( ~n20075 & n20456 ) ;
  assign n20458 = ( n2390 & n6975 ) | ( n2390 & n10851 ) | ( n6975 & n10851 ) ;
  assign n20459 = ( ~n12108 & n19931 ) | ( ~n12108 & n20458 ) | ( n19931 & n20458 ) ;
  assign n20460 = ( n10976 & ~n12147 ) | ( n10976 & n12292 ) | ( ~n12147 & n12292 ) ;
  assign n20461 = n20460 ^ n17197 ^ n1412 ;
  assign n20462 = ( n9449 & n11432 ) | ( n9449 & n19003 ) | ( n11432 & n19003 ) ;
  assign n20463 = n20462 ^ n13915 ^ n7360 ;
  assign n20464 = n20463 ^ n8328 ^ n7375 ;
  assign n20465 = n14871 ^ n12919 ^ n11145 ;
  assign n20466 = ( x4 & x48 ) | ( x4 & ~n1302 ) | ( x48 & ~n1302 ) ;
  assign n20467 = ( n4412 & n6227 ) | ( n4412 & n20466 ) | ( n6227 & n20466 ) ;
  assign n20468 = n8170 ^ n2875 ^ n333 ;
  assign n20469 = n20468 ^ n10424 ^ n6878 ;
  assign n20470 = ( ~n14842 & n20467 ) | ( ~n14842 & n20469 ) | ( n20467 & n20469 ) ;
  assign n20471 = ( n9857 & ~n20465 ) | ( n9857 & n20470 ) | ( ~n20465 & n20470 ) ;
  assign n20472 = ( ~n2340 & n13045 ) | ( ~n2340 & n18615 ) | ( n13045 & n18615 ) ;
  assign n20473 = n20472 ^ n6659 ^ n2855 ;
  assign n20475 = ( n2329 & ~n5623 ) | ( n2329 & n8215 ) | ( ~n5623 & n8215 ) ;
  assign n20476 = n20475 ^ n9269 ^ n9043 ;
  assign n20474 = n18843 ^ n5013 ^ n1095 ;
  assign n20477 = n20476 ^ n20474 ^ n16753 ;
  assign n20478 = ( n4159 & n9824 ) | ( n4159 & ~n12270 ) | ( n9824 & ~n12270 ) ;
  assign n20479 = n20478 ^ n6226 ^ n4589 ;
  assign n20480 = ( ~n2228 & n16226 ) | ( ~n2228 & n20479 ) | ( n16226 & n20479 ) ;
  assign n20481 = ( n4613 & n5897 ) | ( n4613 & n20480 ) | ( n5897 & n20480 ) ;
  assign n20482 = ( n3810 & n4143 ) | ( n3810 & n18754 ) | ( n4143 & n18754 ) ;
  assign n20483 = ( n3676 & n18666 ) | ( n3676 & ~n20482 ) | ( n18666 & ~n20482 ) ;
  assign n20484 = n10118 ^ n8668 ^ n8177 ;
  assign n20485 = n2591 ^ n2541 ^ n1613 ;
  assign n20486 = ( ~n7730 & n8277 ) | ( ~n7730 & n12647 ) | ( n8277 & n12647 ) ;
  assign n20487 = ( n3491 & n15718 ) | ( n3491 & n20486 ) | ( n15718 & n20486 ) ;
  assign n20488 = n10260 ^ n8789 ^ n1324 ;
  assign n20489 = n20488 ^ n13057 ^ n12537 ;
  assign n20490 = ( n2881 & ~n5333 ) | ( n2881 & n20489 ) | ( ~n5333 & n20489 ) ;
  assign n20491 = ( ~n20485 & n20487 ) | ( ~n20485 & n20490 ) | ( n20487 & n20490 ) ;
  assign n20492 = n20192 ^ n14364 ^ n13609 ;
  assign n20493 = ( n2112 & n8890 ) | ( n2112 & ~n10632 ) | ( n8890 & ~n10632 ) ;
  assign n20494 = ( n5308 & ~n15128 ) | ( n5308 & n18314 ) | ( ~n15128 & n18314 ) ;
  assign n20495 = ( n1783 & n20493 ) | ( n1783 & n20494 ) | ( n20493 & n20494 ) ;
  assign n20496 = ( n12644 & ~n12874 ) | ( n12644 & n19694 ) | ( ~n12874 & n19694 ) ;
  assign n20497 = n19265 ^ n15478 ^ n1007 ;
  assign n20498 = ( n15820 & ~n20496 ) | ( n15820 & n20497 ) | ( ~n20496 & n20497 ) ;
  assign n20499 = ( n20234 & ~n20495 ) | ( n20234 & n20498 ) | ( ~n20495 & n20498 ) ;
  assign n20500 = ( ~n5100 & n13279 ) | ( ~n5100 & n20355 ) | ( n13279 & n20355 ) ;
  assign n20503 = n4076 ^ n3397 ^ n1498 ;
  assign n20501 = ( n6371 & n8750 ) | ( n6371 & n18167 ) | ( n8750 & n18167 ) ;
  assign n20502 = ( n4463 & ~n8285 ) | ( n4463 & n20501 ) | ( ~n8285 & n20501 ) ;
  assign n20504 = n20503 ^ n20502 ^ n9174 ;
  assign n20505 = n3859 ^ n814 ^ n758 ;
  assign n20506 = ( ~n1740 & n7077 ) | ( ~n1740 & n20505 ) | ( n7077 & n20505 ) ;
  assign n20507 = ( n4368 & ~n6814 ) | ( n4368 & n20506 ) | ( ~n6814 & n20506 ) ;
  assign n20508 = n15779 ^ n14117 ^ n5320 ;
  assign n20509 = n20508 ^ n17426 ^ n9806 ;
  assign n20511 = ( n1977 & n6467 ) | ( n1977 & n18316 ) | ( n6467 & n18316 ) ;
  assign n20510 = n13756 ^ n6262 ^ n3449 ;
  assign n20512 = n20511 ^ n20510 ^ n19298 ;
  assign n20513 = ( n5007 & n19602 ) | ( n5007 & ~n20512 ) | ( n19602 & ~n20512 ) ;
  assign n20514 = ( n5622 & n13785 ) | ( n5622 & ~n20278 ) | ( n13785 & ~n20278 ) ;
  assign n20515 = n20514 ^ n7217 ^ n1567 ;
  assign n20516 = ( n2722 & n2747 ) | ( n2722 & ~n9008 ) | ( n2747 & ~n9008 ) ;
  assign n20517 = n9044 ^ n7547 ^ n3193 ;
  assign n20518 = ( ~n20515 & n20516 ) | ( ~n20515 & n20517 ) | ( n20516 & n20517 ) ;
  assign n20519 = ( x96 & n1953 ) | ( x96 & ~n5203 ) | ( n1953 & ~n5203 ) ;
  assign n20520 = ( ~n1287 & n9412 ) | ( ~n1287 & n20519 ) | ( n9412 & n20519 ) ;
  assign n20521 = n20520 ^ n16449 ^ n11843 ;
  assign n20522 = n20521 ^ n17822 ^ n15180 ;
  assign n20523 = n11660 ^ n3299 ^ n1505 ;
  assign n20524 = n17228 ^ n16711 ^ n6327 ;
  assign n20525 = ( ~n5263 & n20523 ) | ( ~n5263 & n20524 ) | ( n20523 & n20524 ) ;
  assign n20526 = n19465 ^ n10550 ^ n6318 ;
  assign n20527 = ( ~n2406 & n7335 ) | ( ~n2406 & n20526 ) | ( n7335 & n20526 ) ;
  assign n20528 = n13514 ^ n5791 ^ n1128 ;
  assign n20529 = ( ~n3531 & n6440 ) | ( ~n3531 & n20528 ) | ( n6440 & n20528 ) ;
  assign n20530 = ( n13514 & n19083 ) | ( n13514 & ~n20529 ) | ( n19083 & ~n20529 ) ;
  assign n20531 = ( n3400 & ~n18617 ) | ( n3400 & n20530 ) | ( ~n18617 & n20530 ) ;
  assign n20532 = n16334 ^ n3511 ^ n3113 ;
  assign n20533 = ( n637 & n15392 ) | ( n637 & ~n20532 ) | ( n15392 & ~n20532 ) ;
  assign n20534 = ( n14554 & n20531 ) | ( n14554 & n20533 ) | ( n20531 & n20533 ) ;
  assign n20535 = n15103 ^ n707 ^ n654 ;
  assign n20536 = n20535 ^ n10993 ^ n6300 ;
  assign n20538 = n5449 ^ n5138 ^ n1869 ;
  assign n20539 = n20538 ^ n13855 ^ n8660 ;
  assign n20540 = ( n9291 & n10098 ) | ( n9291 & ~n20539 ) | ( n10098 & ~n20539 ) ;
  assign n20537 = ( n12817 & n16635 ) | ( n12817 & ~n18966 ) | ( n16635 & ~n18966 ) ;
  assign n20541 = n20540 ^ n20537 ^ n10732 ;
  assign n20542 = n20208 ^ n6193 ^ n2198 ;
  assign n20543 = ( ~n670 & n2526 ) | ( ~n670 & n20542 ) | ( n2526 & n20542 ) ;
  assign n20544 = ( ~n5850 & n5923 ) | ( ~n5850 & n18360 ) | ( n5923 & n18360 ) ;
  assign n20545 = ( n20541 & n20543 ) | ( n20541 & n20544 ) | ( n20543 & n20544 ) ;
  assign n20546 = ( n2279 & ~n3196 ) | ( n2279 & n4261 ) | ( ~n3196 & n4261 ) ;
  assign n20547 = n20546 ^ n9158 ^ n6581 ;
  assign n20548 = n20547 ^ n16744 ^ n1716 ;
  assign n20549 = n20125 ^ n3000 ^ n1336 ;
  assign n20550 = ( n4373 & ~n7083 ) | ( n4373 & n12160 ) | ( ~n7083 & n12160 ) ;
  assign n20551 = ( n3068 & n7647 ) | ( n3068 & n20550 ) | ( n7647 & n20550 ) ;
  assign n20552 = n20551 ^ n13273 ^ n11843 ;
  assign n20553 = ( ~n18484 & n20549 ) | ( ~n18484 & n20552 ) | ( n20549 & n20552 ) ;
  assign n20554 = ( ~n1833 & n6733 ) | ( ~n1833 & n14431 ) | ( n6733 & n14431 ) ;
  assign n20555 = ( n2357 & ~n11321 ) | ( n2357 & n20554 ) | ( ~n11321 & n20554 ) ;
  assign n20556 = ( n597 & ~n9988 ) | ( n597 & n10515 ) | ( ~n9988 & n10515 ) ;
  assign n20558 = ( n7285 & n14595 ) | ( n7285 & ~n15896 ) | ( n14595 & ~n15896 ) ;
  assign n20557 = n17213 ^ n1324 ^ n405 ;
  assign n20559 = n20558 ^ n20557 ^ n881 ;
  assign n20560 = ( n1575 & n13251 ) | ( n1575 & n20559 ) | ( n13251 & n20559 ) ;
  assign n20561 = ( ~n5880 & n20556 ) | ( ~n5880 & n20560 ) | ( n20556 & n20560 ) ;
  assign n20583 = ( ~n2513 & n9519 ) | ( ~n2513 & n18590 ) | ( n9519 & n18590 ) ;
  assign n20584 = ( ~n9377 & n12066 ) | ( ~n9377 & n20583 ) | ( n12066 & n20583 ) ;
  assign n20562 = ( n10027 & n10294 ) | ( n10027 & n12491 ) | ( n10294 & n12491 ) ;
  assign n20563 = n20562 ^ n18657 ^ n17269 ;
  assign n20564 = n20563 ^ n15460 ^ n14520 ;
  assign n20565 = n20564 ^ n13246 ^ n6638 ;
  assign n20566 = n8191 ^ n328 ^ x66 ;
  assign n20567 = ( n10880 & n13236 ) | ( n10880 & n20566 ) | ( n13236 & n20566 ) ;
  assign n20568 = n20567 ^ n9199 ^ n467 ;
  assign n20569 = ( n1678 & ~n6784 ) | ( n1678 & n12738 ) | ( ~n6784 & n12738 ) ;
  assign n20570 = ( n581 & ~n14137 ) | ( n581 & n16682 ) | ( ~n14137 & n16682 ) ;
  assign n20571 = ( ~n20568 & n20569 ) | ( ~n20568 & n20570 ) | ( n20569 & n20570 ) ;
  assign n20572 = n15739 ^ n10753 ^ n5086 ;
  assign n20573 = n13846 ^ n6030 ^ n4308 ;
  assign n20574 = ( n3925 & ~n20572 ) | ( n3925 & n20573 ) | ( ~n20572 & n20573 ) ;
  assign n20575 = ( n1536 & ~n9104 ) | ( n1536 & n16151 ) | ( ~n9104 & n16151 ) ;
  assign n20576 = n20575 ^ n12962 ^ n1654 ;
  assign n20577 = n20576 ^ n7493 ^ n4240 ;
  assign n20578 = ( n1296 & n3123 ) | ( n1296 & ~n15172 ) | ( n3123 & ~n15172 ) ;
  assign n20579 = n20578 ^ n19680 ^ n9681 ;
  assign n20580 = ( n2585 & n10409 ) | ( n2585 & ~n20579 ) | ( n10409 & ~n20579 ) ;
  assign n20581 = ( n20574 & n20577 ) | ( n20574 & n20580 ) | ( n20577 & n20580 ) ;
  assign n20582 = ( ~n20565 & n20571 ) | ( ~n20565 & n20581 ) | ( n20571 & n20581 ) ;
  assign n20585 = n20584 ^ n20582 ^ n8963 ;
  assign n20591 = ( n8664 & n9615 ) | ( n8664 & n11669 ) | ( n9615 & n11669 ) ;
  assign n20586 = ( ~n6271 & n14063 ) | ( ~n6271 & n14701 ) | ( n14063 & n14701 ) ;
  assign n20587 = n13041 ^ n5133 ^ n2473 ;
  assign n20588 = ( n4900 & ~n6014 ) | ( n4900 & n20587 ) | ( ~n6014 & n20587 ) ;
  assign n20589 = ( n3427 & ~n15964 ) | ( n3427 & n20588 ) | ( ~n15964 & n20588 ) ;
  assign n20590 = ( n4951 & n20586 ) | ( n4951 & ~n20589 ) | ( n20586 & ~n20589 ) ;
  assign n20592 = n20591 ^ n20590 ^ n4936 ;
  assign n20593 = n15906 ^ n12750 ^ n11020 ;
  assign n20598 = ( ~n1917 & n3324 ) | ( ~n1917 & n5032 ) | ( n3324 & n5032 ) ;
  assign n20599 = ( n300 & ~n5531 ) | ( n300 & n20598 ) | ( ~n5531 & n20598 ) ;
  assign n20596 = n19706 ^ n6589 ^ n4195 ;
  assign n20594 = ( ~n6203 & n8405 ) | ( ~n6203 & n19671 ) | ( n8405 & n19671 ) ;
  assign n20595 = n20594 ^ n17022 ^ n11109 ;
  assign n20597 = n20596 ^ n20595 ^ n2013 ;
  assign n20600 = n20599 ^ n20597 ^ n4283 ;
  assign n20601 = n12306 ^ n9384 ^ n3198 ;
  assign n20602 = n20601 ^ n19343 ^ n4060 ;
  assign n20603 = ( n993 & ~n8728 ) | ( n993 & n20596 ) | ( ~n8728 & n20596 ) ;
  assign n20604 = ( ~n309 & n1430 ) | ( ~n309 & n5321 ) | ( n1430 & n5321 ) ;
  assign n20605 = ( n5335 & n9611 ) | ( n5335 & ~n11240 ) | ( n9611 & ~n11240 ) ;
  assign n20606 = ( ~n10129 & n20604 ) | ( ~n10129 & n20605 ) | ( n20604 & n20605 ) ;
  assign n20607 = ( n8182 & n10853 ) | ( n8182 & n20606 ) | ( n10853 & n20606 ) ;
  assign n20608 = n14051 ^ n10366 ^ n4044 ;
  assign n20609 = ( n2512 & n14276 ) | ( n2512 & ~n14362 ) | ( n14276 & ~n14362 ) ;
  assign n20610 = ( n12739 & n13174 ) | ( n12739 & n20609 ) | ( n13174 & n20609 ) ;
  assign n20611 = n8059 ^ n3518 ^ n1727 ;
  assign n20612 = n13223 ^ n9525 ^ n7565 ;
  assign n20613 = ( ~n1001 & n6724 ) | ( ~n1001 & n20612 ) | ( n6724 & n20612 ) ;
  assign n20614 = n20613 ^ n14472 ^ n6996 ;
  assign n20615 = n20614 ^ n12496 ^ n4438 ;
  assign n20618 = ( n6904 & n7723 ) | ( n6904 & n12663 ) | ( n7723 & n12663 ) ;
  assign n20616 = ( n2303 & ~n3017 ) | ( n2303 & n3206 ) | ( ~n3017 & n3206 ) ;
  assign n20617 = n20616 ^ n15701 ^ n7254 ;
  assign n20619 = n20618 ^ n20617 ^ n12880 ;
  assign n20620 = ( ~n10288 & n16830 ) | ( ~n10288 & n17561 ) | ( n16830 & n17561 ) ;
  assign n20621 = n20620 ^ n5387 ^ n4835 ;
  assign n20622 = ( n685 & n6701 ) | ( n685 & ~n20621 ) | ( n6701 & ~n20621 ) ;
  assign n20623 = ( n2250 & n11135 ) | ( n2250 & n16509 ) | ( n11135 & n16509 ) ;
  assign n20624 = ( ~n1124 & n5295 ) | ( ~n1124 & n20623 ) | ( n5295 & n20623 ) ;
  assign n20625 = ( n6434 & n15957 ) | ( n6434 & n20019 ) | ( n15957 & n20019 ) ;
  assign n20626 = ( n1045 & ~n5577 ) | ( n1045 & n12372 ) | ( ~n5577 & n12372 ) ;
  assign n20627 = ( n9865 & n13533 ) | ( n9865 & n20626 ) | ( n13533 & n20626 ) ;
  assign n20628 = ( n20624 & ~n20625 ) | ( n20624 & n20627 ) | ( ~n20625 & n20627 ) ;
  assign n20629 = ( n1597 & n11016 ) | ( n1597 & ~n11232 ) | ( n11016 & ~n11232 ) ;
  assign n20630 = n20629 ^ n17750 ^ n16647 ;
  assign n20632 = ( ~n8308 & n8873 ) | ( ~n8308 & n10773 ) | ( n8873 & n10773 ) ;
  assign n20631 = n19559 ^ n14638 ^ n10129 ;
  assign n20633 = n20632 ^ n20631 ^ n6697 ;
  assign n20635 = n11741 ^ n6169 ^ n6100 ;
  assign n20634 = n7574 ^ n7067 ^ n1853 ;
  assign n20636 = n20635 ^ n20634 ^ n6173 ;
  assign n20637 = n20408 ^ n20074 ^ n16511 ;
  assign n20638 = n20637 ^ n19872 ^ n17031 ;
  assign n20639 = ( ~n8549 & n12635 ) | ( ~n8549 & n14730 ) | ( n12635 & n14730 ) ;
  assign n20640 = n6736 ^ n4676 ^ n3482 ;
  assign n20641 = ( n2124 & ~n4291 ) | ( n2124 & n7241 ) | ( ~n4291 & n7241 ) ;
  assign n20642 = ( n9273 & ~n20640 ) | ( n9273 & n20641 ) | ( ~n20640 & n20641 ) ;
  assign n20643 = ( n20264 & n20639 ) | ( n20264 & ~n20642 ) | ( n20639 & ~n20642 ) ;
  assign n20644 = ( n3196 & n8378 ) | ( n3196 & ~n20643 ) | ( n8378 & ~n20643 ) ;
  assign n20645 = n16314 ^ n9055 ^ n3671 ;
  assign n20646 = n17709 ^ n13516 ^ n5755 ;
  assign n20647 = n20646 ^ n5632 ^ n2473 ;
  assign n20648 = ( n15094 & n20645 ) | ( n15094 & n20647 ) | ( n20645 & n20647 ) ;
  assign n20649 = ( ~n3880 & n10484 ) | ( ~n3880 & n17486 ) | ( n10484 & n17486 ) ;
  assign n20650 = ( n3054 & ~n5354 ) | ( n3054 & n7173 ) | ( ~n5354 & n7173 ) ;
  assign n20654 = ( ~n9836 & n10608 ) | ( ~n9836 & n17306 ) | ( n10608 & n17306 ) ;
  assign n20651 = ( n2202 & n3164 ) | ( n2202 & n10022 ) | ( n3164 & n10022 ) ;
  assign n20652 = ( n3787 & n6266 ) | ( n3787 & n20651 ) | ( n6266 & n20651 ) ;
  assign n20653 = ( n409 & n15578 ) | ( n409 & n20652 ) | ( n15578 & n20652 ) ;
  assign n20655 = n20654 ^ n20653 ^ n4957 ;
  assign n20656 = n19955 ^ n12356 ^ n10650 ;
  assign n20657 = n6379 ^ n5876 ^ n517 ;
  assign n20658 = ( n7753 & n20656 ) | ( n7753 & n20657 ) | ( n20656 & n20657 ) ;
  assign n20659 = n6128 ^ n4105 ^ n2153 ;
  assign n20660 = ( n4664 & n10739 ) | ( n4664 & n13045 ) | ( n10739 & n13045 ) ;
  assign n20661 = ( n16414 & ~n20659 ) | ( n16414 & n20660 ) | ( ~n20659 & n20660 ) ;
  assign n20662 = ( n3079 & ~n9360 ) | ( n3079 & n20661 ) | ( ~n9360 & n20661 ) ;
  assign n20663 = ( n2968 & n12575 ) | ( n2968 & ~n14618 ) | ( n12575 & ~n14618 ) ;
  assign n20664 = n19908 ^ n13522 ^ n7452 ;
  assign n20665 = ( n2884 & ~n12736 ) | ( n2884 & n13485 ) | ( ~n12736 & n13485 ) ;
  assign n20666 = ( n4833 & ~n10909 ) | ( n4833 & n20665 ) | ( ~n10909 & n20665 ) ;
  assign n20667 = n20666 ^ n17361 ^ n7017 ;
  assign n20668 = n14952 ^ n9861 ^ n7334 ;
  assign n20669 = n5271 ^ n4398 ^ n3084 ;
  assign n20670 = n20669 ^ n13325 ^ n3230 ;
  assign n20671 = n15690 ^ n4874 ^ n2331 ;
  assign n20672 = ( n3516 & n6689 ) | ( n3516 & n20671 ) | ( n6689 & n20671 ) ;
  assign n20673 = ( n2099 & n2683 ) | ( n2099 & ~n11948 ) | ( n2683 & ~n11948 ) ;
  assign n20674 = ( n12750 & n20350 ) | ( n12750 & ~n20673 ) | ( n20350 & ~n20673 ) ;
  assign n20675 = ( n6325 & ~n9440 ) | ( n6325 & n20674 ) | ( ~n9440 & n20674 ) ;
  assign n20676 = ( ~n1750 & n11549 ) | ( ~n1750 & n13249 ) | ( n11549 & n13249 ) ;
  assign n20679 = n15045 ^ n7109 ^ n5072 ;
  assign n20677 = n19429 ^ n11481 ^ n8290 ;
  assign n20678 = n20677 ^ n11815 ^ n4956 ;
  assign n20680 = n20679 ^ n20678 ^ n12659 ;
  assign n20681 = ( n1080 & n16446 ) | ( n1080 & ~n18205 ) | ( n16446 & ~n18205 ) ;
  assign n20682 = n20681 ^ n13022 ^ n6603 ;
  assign n20683 = n19128 ^ n18400 ^ n9191 ;
  assign n20684 = ( n3232 & n17718 ) | ( n3232 & ~n20683 ) | ( n17718 & ~n20683 ) ;
  assign n20685 = ( n6532 & n14563 ) | ( n6532 & n14653 ) | ( n14563 & n14653 ) ;
  assign n20686 = ( ~n10763 & n14336 ) | ( ~n10763 & n15238 ) | ( n14336 & n15238 ) ;
  assign n20687 = n17534 ^ n15322 ^ n5479 ;
  assign n20688 = ( n15496 & n16700 ) | ( n15496 & ~n20687 ) | ( n16700 & ~n20687 ) ;
  assign n20689 = ( n3405 & n12868 ) | ( n3405 & n18349 ) | ( n12868 & n18349 ) ;
  assign n20690 = ( n673 & ~n13969 ) | ( n673 & n20689 ) | ( ~n13969 & n20689 ) ;
  assign n20691 = n5077 ^ n3524 ^ n177 ;
  assign n20692 = n20691 ^ n14917 ^ n6094 ;
  assign n20693 = ( ~n4552 & n8684 ) | ( ~n4552 & n9291 ) | ( n8684 & n9291 ) ;
  assign n20694 = n20693 ^ n20496 ^ n4485 ;
  assign n20695 = n20694 ^ n15491 ^ n7210 ;
  assign n20696 = n20695 ^ n13793 ^ n12503 ;
  assign n20697 = ( n535 & ~n8011 ) | ( n535 & n16573 ) | ( ~n8011 & n16573 ) ;
  assign n20698 = ( n4675 & ~n5009 ) | ( n4675 & n5183 ) | ( ~n5009 & n5183 ) ;
  assign n20699 = n19360 ^ n12357 ^ n7990 ;
  assign n20700 = ( n15384 & ~n20698 ) | ( n15384 & n20699 ) | ( ~n20698 & n20699 ) ;
  assign n20701 = ( ~n642 & n2661 ) | ( ~n642 & n16633 ) | ( n2661 & n16633 ) ;
  assign n20702 = n20701 ^ n13358 ^ n11371 ;
  assign n20703 = ( ~x32 & n4465 ) | ( ~x32 & n16023 ) | ( n4465 & n16023 ) ;
  assign n20704 = n7337 ^ n4616 ^ n3196 ;
  assign n20705 = n20704 ^ n5731 ^ n1029 ;
  assign n20706 = ( n17428 & n20293 ) | ( n17428 & ~n20705 ) | ( n20293 & ~n20705 ) ;
  assign n20707 = ( ~n243 & n2147 ) | ( ~n243 & n2249 ) | ( n2147 & n2249 ) ;
  assign n20708 = n20707 ^ n10054 ^ n9652 ;
  assign n20709 = ( ~x116 & n8075 ) | ( ~x116 & n20708 ) | ( n8075 & n20708 ) ;
  assign n20710 = ( n2197 & n6719 ) | ( n2197 & ~n14849 ) | ( n6719 & ~n14849 ) ;
  assign n20711 = ( n617 & ~n20709 ) | ( n617 & n20710 ) | ( ~n20709 & n20710 ) ;
  assign n20712 = ( n8739 & n15078 ) | ( n8739 & ~n15644 ) | ( n15078 & ~n15644 ) ;
  assign n20713 = ( n8867 & n11941 ) | ( n8867 & ~n20712 ) | ( n11941 & ~n20712 ) ;
  assign n20714 = ( n2080 & ~n12576 ) | ( n2080 & n19715 ) | ( ~n12576 & n19715 ) ;
  assign n20715 = ( n996 & n20713 ) | ( n996 & ~n20714 ) | ( n20713 & ~n20714 ) ;
  assign n20716 = ( n9968 & ~n18177 ) | ( n9968 & n20715 ) | ( ~n18177 & n20715 ) ;
  assign n20717 = ( n6124 & n13985 ) | ( n6124 & n19342 ) | ( n13985 & n19342 ) ;
  assign n20718 = ( n8082 & n9104 ) | ( n8082 & n12694 ) | ( n9104 & n12694 ) ;
  assign n20719 = n20718 ^ n9659 ^ n2252 ;
  assign n20720 = n14917 ^ n11560 ^ n7180 ;
  assign n20729 = n13036 ^ n9299 ^ n5345 ;
  assign n20732 = ( n5026 & n8876 ) | ( n5026 & n13369 ) | ( n8876 & n13369 ) ;
  assign n20730 = ( n5527 & ~n9302 ) | ( n5527 & n19985 ) | ( ~n9302 & n19985 ) ;
  assign n20731 = ( ~n1005 & n7738 ) | ( ~n1005 & n20730 ) | ( n7738 & n20730 ) ;
  assign n20733 = n20732 ^ n20731 ^ n8335 ;
  assign n20734 = ( ~n5931 & n20729 ) | ( ~n5931 & n20733 ) | ( n20729 & n20733 ) ;
  assign n20726 = ( n8883 & n9370 ) | ( n8883 & ~n9966 ) | ( n9370 & ~n9966 ) ;
  assign n20727 = ( ~n1174 & n5474 ) | ( ~n1174 & n20726 ) | ( n5474 & n20726 ) ;
  assign n20725 = n11754 ^ n1247 ^ n748 ;
  assign n20724 = ( ~n4473 & n8009 ) | ( ~n4473 & n14842 ) | ( n8009 & n14842 ) ;
  assign n20728 = n20727 ^ n20725 ^ n20724 ;
  assign n20735 = n20734 ^ n20728 ^ n3824 ;
  assign n20721 = n18942 ^ n4378 ^ n940 ;
  assign n20722 = n20721 ^ n11310 ^ n2484 ;
  assign n20723 = n20722 ^ n7094 ^ n1283 ;
  assign n20736 = n20735 ^ n20723 ^ n1335 ;
  assign n20737 = ( n5297 & n12263 ) | ( n5297 & ~n16270 ) | ( n12263 & ~n16270 ) ;
  assign n20738 = n13301 ^ n1730 ^ n1137 ;
  assign n20739 = ( n6567 & n20737 ) | ( n6567 & n20738 ) | ( n20737 & n20738 ) ;
  assign n20740 = n20739 ^ n14232 ^ n4255 ;
  assign n20741 = ( n2448 & ~n14243 ) | ( n2448 & n18808 ) | ( ~n14243 & n18808 ) ;
  assign n20742 = ( n8702 & n10459 ) | ( n8702 & ~n20741 ) | ( n10459 & ~n20741 ) ;
  assign n20743 = ( n3784 & n14419 ) | ( n3784 & n15754 ) | ( n14419 & n15754 ) ;
  assign n20744 = n20743 ^ n19879 ^ n3493 ;
  assign n20745 = ( n12749 & ~n18300 ) | ( n12749 & n20591 ) | ( ~n18300 & n20591 ) ;
  assign n20746 = n20745 ^ n8717 ^ n3084 ;
  assign n20747 = n20746 ^ n15058 ^ n2767 ;
  assign n20748 = ( n3228 & ~n10319 ) | ( n3228 & n13114 ) | ( ~n10319 & n13114 ) ;
  assign n20749 = n15420 ^ n11794 ^ n4963 ;
  assign n20750 = ( ~n3692 & n20748 ) | ( ~n3692 & n20749 ) | ( n20748 & n20749 ) ;
  assign n20751 = n16469 ^ n16090 ^ n14737 ;
  assign n20752 = ( ~n7760 & n13145 ) | ( ~n7760 & n20751 ) | ( n13145 & n20751 ) ;
  assign n20753 = n13314 ^ n5081 ^ n391 ;
  assign n20754 = n20753 ^ n9062 ^ n5171 ;
  assign n20757 = ( n3002 & n3207 ) | ( n3002 & n17756 ) | ( n3207 & n17756 ) ;
  assign n20755 = ( ~n2229 & n2926 ) | ( ~n2229 & n8932 ) | ( n2926 & n8932 ) ;
  assign n20756 = ( n4502 & n5578 ) | ( n4502 & n20755 ) | ( n5578 & n20755 ) ;
  assign n20758 = n20757 ^ n20756 ^ n18939 ;
  assign n20759 = n17860 ^ n9249 ^ x96 ;
  assign n20760 = n19749 ^ n17561 ^ n3292 ;
  assign n20761 = n20760 ^ n12648 ^ n651 ;
  assign n20762 = ( ~n934 & n3904 ) | ( ~n934 & n20761 ) | ( n3904 & n20761 ) ;
  assign n20763 = ( ~n7024 & n17860 ) | ( ~n7024 & n20762 ) | ( n17860 & n20762 ) ;
  assign n20764 = ( n1121 & n9460 ) | ( n1121 & n17957 ) | ( n9460 & n17957 ) ;
  assign n20765 = n13356 ^ n2231 ^ n574 ;
  assign n20766 = ( n939 & ~n4833 ) | ( n939 & n20765 ) | ( ~n4833 & n20765 ) ;
  assign n20767 = ( ~n13952 & n14154 ) | ( ~n13952 & n15743 ) | ( n14154 & n15743 ) ;
  assign n20768 = ( ~n5248 & n7432 ) | ( ~n5248 & n19465 ) | ( n7432 & n19465 ) ;
  assign n20769 = ( n3209 & n4193 ) | ( n3209 & n7358 ) | ( n4193 & n7358 ) ;
  assign n20770 = ( n9211 & ~n16967 ) | ( n9211 & n20769 ) | ( ~n16967 & n20769 ) ;
  assign n20772 = n19916 ^ n13421 ^ n8207 ;
  assign n20771 = ( ~n9889 & n12535 ) | ( ~n9889 & n20520 ) | ( n12535 & n20520 ) ;
  assign n20773 = n20772 ^ n20771 ^ n13262 ;
  assign n20774 = n11749 ^ n2354 ^ n664 ;
  assign n20775 = ( n3346 & n14335 ) | ( n3346 & n20774 ) | ( n14335 & n20774 ) ;
  assign n20776 = ( ~n782 & n3763 ) | ( ~n782 & n20775 ) | ( n3763 & n20775 ) ;
  assign n20777 = ( n4778 & n5144 ) | ( n4778 & n17275 ) | ( n5144 & n17275 ) ;
  assign n20778 = n18275 ^ n9900 ^ n6581 ;
  assign n20779 = n20778 ^ n14971 ^ n8387 ;
  assign n20780 = n14744 ^ n13983 ^ n12494 ;
  assign n20781 = n8977 ^ n8913 ^ n6143 ;
  assign n20782 = ( x67 & ~n6320 ) | ( x67 & n7807 ) | ( ~n6320 & n7807 ) ;
  assign n20783 = ( n3110 & ~n20781 ) | ( n3110 & n20782 ) | ( ~n20781 & n20782 ) ;
  assign n20784 = ( n466 & n3731 ) | ( n466 & ~n4847 ) | ( n3731 & ~n4847 ) ;
  assign n20785 = ( n18286 & ~n20506 ) | ( n18286 & n20784 ) | ( ~n20506 & n20784 ) ;
  assign n20786 = ( n7192 & n16509 ) | ( n7192 & ~n16731 ) | ( n16509 & ~n16731 ) ;
  assign n20787 = n20272 ^ n10589 ^ n5578 ;
  assign n20788 = n6358 ^ n5486 ^ n3362 ;
  assign n20789 = ( n6854 & ~n14220 ) | ( n6854 & n17458 ) | ( ~n14220 & n17458 ) ;
  assign n20797 = n12544 ^ n11910 ^ n9190 ;
  assign n20794 = ( x4 & n1294 ) | ( x4 & n3392 ) | ( n1294 & n3392 ) ;
  assign n20793 = n12665 ^ n8044 ^ n5823 ;
  assign n20795 = n20794 ^ n20793 ^ n18442 ;
  assign n20796 = n20795 ^ n16489 ^ n8225 ;
  assign n20791 = ( x31 & ~n1333 ) | ( x31 & n2343 ) | ( ~n1333 & n2343 ) ;
  assign n20790 = n13344 ^ n4782 ^ n3141 ;
  assign n20792 = n20791 ^ n20790 ^ n20176 ;
  assign n20798 = n20797 ^ n20796 ^ n20792 ;
  assign n20799 = ( n6807 & n9900 ) | ( n6807 & ~n19516 ) | ( n9900 & ~n19516 ) ;
  assign n20800 = n19232 ^ n4069 ^ n3153 ;
  assign n20801 = n7310 ^ n5175 ^ n2098 ;
  assign n20802 = n20801 ^ n1296 ^ n1030 ;
  assign n20803 = ( ~n1657 & n1827 ) | ( ~n1657 & n10852 ) | ( n1827 & n10852 ) ;
  assign n20804 = n20803 ^ n13994 ^ n2634 ;
  assign n20805 = n17598 ^ n7609 ^ n2896 ;
  assign n20806 = ( ~n20802 & n20804 ) | ( ~n20802 & n20805 ) | ( n20804 & n20805 ) ;
  assign n20808 = n17248 ^ n8943 ^ n2582 ;
  assign n20809 = ( ~n2933 & n12440 ) | ( ~n2933 & n16963 ) | ( n12440 & n16963 ) ;
  assign n20810 = ( n9110 & n20808 ) | ( n9110 & n20809 ) | ( n20808 & n20809 ) ;
  assign n20807 = ( ~n4890 & n8285 ) | ( ~n4890 & n12503 ) | ( n8285 & n12503 ) ;
  assign n20811 = n20810 ^ n20807 ^ n1962 ;
  assign n20812 = n12559 ^ n8523 ^ n2028 ;
  assign n20813 = ( ~n379 & n877 ) | ( ~n379 & n1169 ) | ( n877 & n1169 ) ;
  assign n20814 = ( n7687 & ~n18502 ) | ( n7687 & n20722 ) | ( ~n18502 & n20722 ) ;
  assign n20815 = n17262 ^ n14005 ^ n2043 ;
  assign n20816 = n20815 ^ n17160 ^ n10810 ;
  assign n20817 = n15886 ^ n14349 ^ n14004 ;
  assign n20818 = ( ~n3541 & n18671 ) | ( ~n3541 & n20817 ) | ( n18671 & n20817 ) ;
  assign n20819 = ( n7752 & n9862 ) | ( n7752 & n20818 ) | ( n9862 & n20818 ) ;
  assign n20820 = n5432 ^ n2174 ^ n850 ;
  assign n20821 = ( n4813 & ~n5410 ) | ( n4813 & n8423 ) | ( ~n5410 & n8423 ) ;
  assign n20822 = ( n3851 & n14660 ) | ( n3851 & n20821 ) | ( n14660 & n20821 ) ;
  assign n20823 = n17791 ^ n3757 ^ n2361 ;
  assign n20824 = ( n3670 & n9383 ) | ( n3670 & ~n20823 ) | ( n9383 & ~n20823 ) ;
  assign n20825 = n4739 ^ n4270 ^ n2332 ;
  assign n20826 = ( n8019 & ~n12749 ) | ( n8019 & n20825 ) | ( ~n12749 & n20825 ) ;
  assign n20828 = ( n5394 & n8007 ) | ( n5394 & ~n8220 ) | ( n8007 & ~n8220 ) ;
  assign n20827 = ( n7165 & n15472 ) | ( n7165 & ~n16366 ) | ( n15472 & ~n16366 ) ;
  assign n20829 = n20828 ^ n20827 ^ n12372 ;
  assign n20830 = n19290 ^ n15590 ^ n14113 ;
  assign n20831 = n12079 ^ n11927 ^ n10859 ;
  assign n20834 = n12962 ^ n11666 ^ n2451 ;
  assign n20832 = ( n3344 & n8882 ) | ( n3344 & ~n10905 ) | ( n8882 & ~n10905 ) ;
  assign n20833 = n20832 ^ n10078 ^ n8133 ;
  assign n20835 = n20834 ^ n20833 ^ n5518 ;
  assign n20836 = n17625 ^ n16630 ^ n4454 ;
  assign n20837 = n8203 ^ n3762 ^ n3710 ;
  assign n20838 = n20837 ^ n5029 ^ n1995 ;
  assign n20839 = ( n177 & n1373 ) | ( n177 & ~n9565 ) | ( n1373 & ~n9565 ) ;
  assign n20840 = ( n5139 & n5823 ) | ( n5139 & ~n6742 ) | ( n5823 & ~n6742 ) ;
  assign n20841 = n20840 ^ n2363 ^ n1753 ;
  assign n20842 = ( ~n5786 & n15744 ) | ( ~n5786 & n20841 ) | ( n15744 & n20841 ) ;
  assign n20843 = ( ~n16207 & n20839 ) | ( ~n16207 & n20842 ) | ( n20839 & n20842 ) ;
  assign n20844 = ( n7722 & n9369 ) | ( n7722 & ~n14875 ) | ( n9369 & ~n14875 ) ;
  assign n20845 = ( n11383 & ~n14526 ) | ( n11383 & n20844 ) | ( ~n14526 & n20844 ) ;
  assign n20846 = n20845 ^ n15142 ^ n5167 ;
  assign n20847 = n9645 ^ n7957 ^ n1299 ;
  assign n20848 = ( n2586 & n9160 ) | ( n2586 & n20847 ) | ( n9160 & n20847 ) ;
  assign n20849 = ( n2170 & ~n8377 ) | ( n2170 & n16838 ) | ( ~n8377 & n16838 ) ;
  assign n20850 = ( ~n8745 & n14058 ) | ( ~n8745 & n17811 ) | ( n14058 & n17811 ) ;
  assign n20851 = ( n14332 & n19050 ) | ( n14332 & n20850 ) | ( n19050 & n20850 ) ;
  assign n20852 = n13439 ^ n12604 ^ x28 ;
  assign n20853 = ( ~n8739 & n11605 ) | ( ~n8739 & n16142 ) | ( n11605 & n16142 ) ;
  assign n20854 = n9850 ^ n7197 ^ n429 ;
  assign n20855 = ( n1917 & n3786 ) | ( n1917 & ~n20854 ) | ( n3786 & ~n20854 ) ;
  assign n20856 = ( n9957 & ~n20853 ) | ( n9957 & n20855 ) | ( ~n20853 & n20855 ) ;
  assign n20857 = ( ~n7328 & n20852 ) | ( ~n7328 & n20856 ) | ( n20852 & n20856 ) ;
  assign n20858 = ( n10054 & n14449 ) | ( n10054 & ~n14722 ) | ( n14449 & ~n14722 ) ;
  assign n20859 = n13745 ^ n13280 ^ n2136 ;
  assign n20860 = n20859 ^ n18270 ^ n10599 ;
  assign n20861 = ( n7443 & ~n8058 ) | ( n7443 & n20860 ) | ( ~n8058 & n20860 ) ;
  assign n20862 = n19045 ^ n7076 ^ n6771 ;
  assign n20863 = n20862 ^ n10976 ^ n9516 ;
  assign n20864 = ( n3397 & ~n8360 ) | ( n3397 & n20863 ) | ( ~n8360 & n20863 ) ;
  assign n20865 = ( n297 & n8327 ) | ( n297 & ~n12918 ) | ( n8327 & ~n12918 ) ;
  assign n20866 = n15779 ^ n14923 ^ n6681 ;
  assign n20867 = ( n15953 & n20865 ) | ( n15953 & ~n20866 ) | ( n20865 & ~n20866 ) ;
  assign n20868 = ( ~n499 & n1156 ) | ( ~n499 & n5405 ) | ( n1156 & n5405 ) ;
  assign n20869 = ( ~n1178 & n6031 ) | ( ~n1178 & n20868 ) | ( n6031 & n20868 ) ;
  assign n20870 = n20869 ^ n7556 ^ n3478 ;
  assign n20871 = n17021 ^ n3886 ^ n3238 ;
  assign n20872 = ( n6071 & n14923 ) | ( n6071 & n20871 ) | ( n14923 & n20871 ) ;
  assign n20873 = ( n1460 & n20870 ) | ( n1460 & ~n20872 ) | ( n20870 & ~n20872 ) ;
  assign n20874 = ( n13225 & n14696 ) | ( n13225 & ~n17907 ) | ( n14696 & ~n17907 ) ;
  assign n20875 = n20874 ^ n9633 ^ n8558 ;
  assign n20876 = ( n2356 & n5570 ) | ( n2356 & n20875 ) | ( n5570 & n20875 ) ;
  assign n20877 = n19734 ^ n13904 ^ n3058 ;
  assign n20878 = n8658 ^ n5346 ^ n2302 ;
  assign n20879 = ( n9857 & n14566 ) | ( n9857 & ~n20878 ) | ( n14566 & ~n20878 ) ;
  assign n20880 = n12616 ^ n7756 ^ n3964 ;
  assign n20881 = n20880 ^ n9887 ^ n6183 ;
  assign n20882 = ( ~n20877 & n20879 ) | ( ~n20877 & n20881 ) | ( n20879 & n20881 ) ;
  assign n20883 = ( n3840 & n6803 ) | ( n3840 & ~n10715 ) | ( n6803 & ~n10715 ) ;
  assign n20884 = ( ~n1109 & n11767 ) | ( ~n1109 & n20704 ) | ( n11767 & n20704 ) ;
  assign n20885 = n20884 ^ n7508 ^ n6320 ;
  assign n20886 = ( ~n1738 & n1990 ) | ( ~n1738 & n2916 ) | ( n1990 & n2916 ) ;
  assign n20887 = ( n4641 & n20885 ) | ( n4641 & n20886 ) | ( n20885 & n20886 ) ;
  assign n20890 = n3735 ^ n3446 ^ n2846 ;
  assign n20891 = n20890 ^ n15073 ^ x80 ;
  assign n20888 = n11020 ^ n9203 ^ x65 ;
  assign n20889 = n20888 ^ n12732 ^ n10025 ;
  assign n20892 = n20891 ^ n20889 ^ n19979 ;
  assign n20893 = n16485 ^ n10180 ^ n2813 ;
  assign n20894 = ( n2121 & ~n3039 ) | ( n2121 & n20893 ) | ( ~n3039 & n20893 ) ;
  assign n20895 = ( n9764 & n11336 ) | ( n9764 & ~n20019 ) | ( n11336 & ~n20019 ) ;
  assign n20896 = n20895 ^ n1999 ^ n1875 ;
  assign n20897 = n16167 ^ n6859 ^ n3068 ;
  assign n20898 = ( n1597 & ~n12466 ) | ( n1597 & n14766 ) | ( ~n12466 & n14766 ) ;
  assign n20899 = ( n2535 & ~n10967 ) | ( n2535 & n20898 ) | ( ~n10967 & n20898 ) ;
  assign n20900 = ( ~n7339 & n18999 ) | ( ~n7339 & n20899 ) | ( n18999 & n20899 ) ;
  assign n20903 = n12074 ^ n7744 ^ n763 ;
  assign n20901 = n7257 ^ n6579 ^ n4621 ;
  assign n20902 = n20901 ^ n10715 ^ n372 ;
  assign n20904 = n20903 ^ n20902 ^ n14471 ;
  assign n20905 = n20904 ^ n13180 ^ n1734 ;
  assign n20906 = ( n992 & n6190 ) | ( n992 & n6714 ) | ( n6190 & n6714 ) ;
  assign n20907 = n15473 ^ n11059 ^ n1901 ;
  assign n20908 = n7317 ^ n4085 ^ n3091 ;
  assign n20909 = ( n6276 & ~n6717 ) | ( n6276 & n20908 ) | ( ~n6717 & n20908 ) ;
  assign n20910 = ( n20906 & n20907 ) | ( n20906 & n20909 ) | ( n20907 & n20909 ) ;
  assign n20911 = ( n697 & ~n4487 ) | ( n697 & n10359 ) | ( ~n4487 & n10359 ) ;
  assign n20912 = ( ~n15991 & n17092 ) | ( ~n15991 & n20911 ) | ( n17092 & n20911 ) ;
  assign n20913 = n20912 ^ n15316 ^ n14948 ;
  assign n20914 = n16411 ^ n15007 ^ n864 ;
  assign n20915 = n20914 ^ n10368 ^ n9891 ;
  assign n20916 = n7379 ^ n7038 ^ n1546 ;
  assign n20917 = ( n10666 & n20915 ) | ( n10666 & n20916 ) | ( n20915 & n20916 ) ;
  assign n20918 = n20917 ^ n7275 ^ n6967 ;
  assign n20919 = n14740 ^ n14264 ^ n11876 ;
  assign n20920 = n20919 ^ n17179 ^ n11387 ;
  assign n20921 = n16799 ^ n10312 ^ n6896 ;
  assign n20922 = n19118 ^ n12513 ^ n4040 ;
  assign n20923 = ( n6664 & n9460 ) | ( n6664 & n18020 ) | ( n9460 & n18020 ) ;
  assign n20924 = ( ~n8466 & n15393 ) | ( ~n8466 & n18055 ) | ( n15393 & n18055 ) ;
  assign n20925 = ( n10901 & n17376 ) | ( n10901 & ~n18644 ) | ( n17376 & ~n18644 ) ;
  assign n20926 = ( n20923 & ~n20924 ) | ( n20923 & n20925 ) | ( ~n20924 & n20925 ) ;
  assign n20927 = n17655 ^ n9424 ^ n1415 ;
  assign n20928 = n20794 ^ n7667 ^ n3649 ;
  assign n20929 = ( n13115 & ~n20927 ) | ( n13115 & n20928 ) | ( ~n20927 & n20928 ) ;
  assign n20930 = ( n4053 & n11661 ) | ( n4053 & ~n13663 ) | ( n11661 & ~n13663 ) ;
  assign n20931 = ( n504 & n5237 ) | ( n504 & ~n8123 ) | ( n5237 & ~n8123 ) ;
  assign n20932 = n20931 ^ n20677 ^ n15759 ;
  assign n20933 = ( n2327 & ~n4590 ) | ( n2327 & n10548 ) | ( ~n4590 & n10548 ) ;
  assign n20935 = n14952 ^ n13626 ^ n2957 ;
  assign n20934 = ( n6830 & n10638 ) | ( n6830 & ~n11370 ) | ( n10638 & ~n11370 ) ;
  assign n20936 = n20935 ^ n20934 ^ n9387 ;
  assign n20937 = n20936 ^ n11429 ^ n9389 ;
  assign n20938 = ( ~n1993 & n11843 ) | ( ~n1993 & n14384 ) | ( n11843 & n14384 ) ;
  assign n20939 = n15135 ^ n5477 ^ n4759 ;
  assign n20940 = n20774 ^ n13239 ^ n3550 ;
  assign n20941 = n15704 ^ n10562 ^ n611 ;
  assign n20942 = n20941 ^ n14026 ^ n2927 ;
  assign n20943 = n19112 ^ n15320 ^ n11923 ;
  assign n20944 = n15418 ^ n11982 ^ n6194 ;
  assign n20945 = n20944 ^ n20803 ^ n8765 ;
  assign n20946 = ( ~n8496 & n18691 ) | ( ~n8496 & n20945 ) | ( n18691 & n20945 ) ;
  assign n20947 = ( ~n18957 & n20943 ) | ( ~n18957 & n20946 ) | ( n20943 & n20946 ) ;
  assign n20948 = n4733 ^ n1986 ^ n1404 ;
  assign n20949 = n20948 ^ n17193 ^ n776 ;
  assign n20950 = ( n7810 & n13388 ) | ( n7810 & n18969 ) | ( n13388 & n18969 ) ;
  assign n20951 = n16270 ^ n14589 ^ n5860 ;
  assign n20952 = ( ~n6489 & n7320 ) | ( ~n6489 & n18544 ) | ( n7320 & n18544 ) ;
  assign n20953 = ( n2505 & ~n9402 ) | ( n2505 & n20952 ) | ( ~n9402 & n20952 ) ;
  assign n20954 = ( ~n18317 & n20951 ) | ( ~n18317 & n20953 ) | ( n20951 & n20953 ) ;
  assign n20955 = ( n462 & n6876 ) | ( n462 & ~n19995 ) | ( n6876 & ~n19995 ) ;
  assign n20956 = n11652 ^ n7930 ^ n2271 ;
  assign n20957 = n13540 ^ n12766 ^ n5865 ;
  assign n20958 = ( ~n1215 & n8688 ) | ( ~n1215 & n20957 ) | ( n8688 & n20957 ) ;
  assign n20959 = n19445 ^ n10920 ^ n10245 ;
  assign n20961 = n10067 ^ n6423 ^ n5238 ;
  assign n20962 = n20961 ^ n10699 ^ n6202 ;
  assign n20960 = n12433 ^ n11486 ^ n5980 ;
  assign n20963 = n20962 ^ n20960 ^ n5326 ;
  assign n20965 = n10433 ^ n3785 ^ n1757 ;
  assign n20964 = ( n154 & n4557 ) | ( n154 & ~n17841 ) | ( n4557 & ~n17841 ) ;
  assign n20966 = n20965 ^ n20964 ^ n9391 ;
  assign n20967 = n19002 ^ n5893 ^ n871 ;
  assign n20968 = ( n2205 & n13440 ) | ( n2205 & n20967 ) | ( n13440 & n20967 ) ;
  assign n20969 = n14684 ^ n10051 ^ n6987 ;
  assign n20970 = ( n3160 & n5101 ) | ( n3160 & n10489 ) | ( n5101 & n10489 ) ;
  assign n20971 = ( n4604 & n14733 ) | ( n4604 & n20970 ) | ( n14733 & n20970 ) ;
  assign n20972 = ( n9795 & n12386 ) | ( n9795 & ~n20755 ) | ( n12386 & ~n20755 ) ;
  assign n20973 = ( n9439 & ~n10972 ) | ( n9439 & n13870 ) | ( ~n10972 & n13870 ) ;
  assign n20974 = n20973 ^ n14397 ^ n2460 ;
  assign n20975 = n6598 ^ n5498 ^ n616 ;
  assign n20976 = ( ~n8684 & n17279 ) | ( ~n8684 & n18342 ) | ( n17279 & n18342 ) ;
  assign n20977 = ( n16897 & ~n20975 ) | ( n16897 & n20976 ) | ( ~n20975 & n20976 ) ;
  assign n20978 = ( n4451 & ~n12324 ) | ( n4451 & n20977 ) | ( ~n12324 & n20977 ) ;
  assign n20979 = ( ~n14184 & n14240 ) | ( ~n14184 & n20451 ) | ( n14240 & n20451 ) ;
  assign n20980 = n17618 ^ n7483 ^ n3491 ;
  assign n20981 = ( n13809 & ~n20338 ) | ( n13809 & n20980 ) | ( ~n20338 & n20980 ) ;
  assign n20982 = ( ~n3811 & n11541 ) | ( ~n3811 & n17190 ) | ( n11541 & n17190 ) ;
  assign n20983 = n8651 ^ n6480 ^ n5841 ;
  assign n20984 = n20983 ^ n19738 ^ n7057 ;
  assign n20985 = ( n9442 & ~n16255 ) | ( n9442 & n20984 ) | ( ~n16255 & n20984 ) ;
  assign n20986 = n18377 ^ n9092 ^ n4749 ;
  assign n20988 = ( ~n1230 & n3103 ) | ( ~n1230 & n4584 ) | ( n3103 & n4584 ) ;
  assign n20987 = ( n2538 & ~n5761 ) | ( n2538 & n19578 ) | ( ~n5761 & n19578 ) ;
  assign n20989 = n20988 ^ n20987 ^ n1375 ;
  assign n20990 = ( n470 & n1556 ) | ( n470 & n20989 ) | ( n1556 & n20989 ) ;
  assign n20991 = n20990 ^ n18852 ^ n6181 ;
  assign n20992 = n16963 ^ n7647 ^ n1035 ;
  assign n20993 = ( n3045 & ~n9128 ) | ( n3045 & n9592 ) | ( ~n9128 & n9592 ) ;
  assign n20994 = n20993 ^ n15112 ^ n13617 ;
  assign n20995 = n20994 ^ n9487 ^ n3309 ;
  assign n20996 = n19096 ^ n7763 ^ n4847 ;
  assign n20997 = n10771 ^ n10268 ^ n4673 ;
  assign n20998 = ( n1733 & n3218 ) | ( n1733 & ~n20997 ) | ( n3218 & ~n20997 ) ;
  assign n20999 = ( ~n6224 & n20996 ) | ( ~n6224 & n20998 ) | ( n20996 & n20998 ) ;
  assign n21000 = ( n4224 & n6498 ) | ( n4224 & n15054 ) | ( n6498 & n15054 ) ;
  assign n21001 = ( ~n8805 & n17846 ) | ( ~n8805 & n21000 ) | ( n17846 & n21000 ) ;
  assign n21002 = ( n2622 & ~n7033 ) | ( n2622 & n15413 ) | ( ~n7033 & n15413 ) ;
  assign n21003 = n15712 ^ n10153 ^ n1185 ;
  assign n21004 = ( n7863 & ~n21002 ) | ( n7863 & n21003 ) | ( ~n21002 & n21003 ) ;
  assign n21005 = ( n5090 & n8801 ) | ( n5090 & n20199 ) | ( n8801 & n20199 ) ;
  assign n21006 = ( ~n9936 & n10609 ) | ( ~n9936 & n16731 ) | ( n10609 & n16731 ) ;
  assign n21007 = n21006 ^ n8532 ^ n1931 ;
  assign n21008 = n21007 ^ n11984 ^ n7937 ;
  assign n21009 = n21008 ^ n20794 ^ n10332 ;
  assign n21010 = ( n12581 & n16319 ) | ( n12581 & n18762 ) | ( n16319 & n18762 ) ;
  assign n21011 = ( n2744 & ~n4974 ) | ( n2744 & n17771 ) | ( ~n4974 & n17771 ) ;
  assign n21012 = n10736 ^ n6502 ^ n2582 ;
  assign n21013 = n10545 ^ n6341 ^ n5204 ;
  assign n21014 = ( n6409 & ~n13429 ) | ( n6409 & n21013 ) | ( ~n13429 & n21013 ) ;
  assign n21015 = ( ~n473 & n13598 ) | ( ~n473 & n21014 ) | ( n13598 & n21014 ) ;
  assign n21016 = n15746 ^ n10615 ^ n8141 ;
  assign n21017 = n16888 ^ n8635 ^ n2505 ;
  assign n21018 = n16987 ^ n11222 ^ n6651 ;
  assign n21019 = n6165 ^ n5720 ^ n3053 ;
  assign n21020 = ( n3214 & ~n10867 ) | ( n3214 & n21019 ) | ( ~n10867 & n21019 ) ;
  assign n21021 = ( n3663 & ~n12836 ) | ( n3663 & n21020 ) | ( ~n12836 & n21020 ) ;
  assign n21022 = ( n16272 & n21018 ) | ( n16272 & n21021 ) | ( n21018 & n21021 ) ;
  assign n21023 = n17343 ^ n5775 ^ n5377 ;
  assign n21024 = ( n2122 & n7164 ) | ( n2122 & ~n21023 ) | ( n7164 & ~n21023 ) ;
  assign n21025 = n21024 ^ n4617 ^ n1386 ;
  assign n21026 = n3174 ^ n2877 ^ n2805 ;
  assign n21027 = ( n4189 & ~n6263 ) | ( n4189 & n21026 ) | ( ~n6263 & n21026 ) ;
  assign n21028 = ( n367 & n2077 ) | ( n367 & ~n8825 ) | ( n2077 & ~n8825 ) ;
  assign n21029 = n21028 ^ n14285 ^ n309 ;
  assign n21030 = n21029 ^ n16488 ^ n10025 ;
  assign n21031 = n21030 ^ n19111 ^ n16572 ;
  assign n21032 = n7722 ^ n934 ^ n711 ;
  assign n21033 = ( n15971 & n16090 ) | ( n15971 & ~n16119 ) | ( n16090 & ~n16119 ) ;
  assign n21034 = n21033 ^ n9855 ^ n7285 ;
  assign n21035 = n13519 ^ n12293 ^ n7680 ;
  assign n21036 = ( n1181 & ~n6069 ) | ( n1181 & n14869 ) | ( ~n6069 & n14869 ) ;
  assign n21037 = n21036 ^ n19752 ^ n3601 ;
  assign n21038 = ( n1356 & n11562 ) | ( n1356 & ~n21037 ) | ( n11562 & ~n21037 ) ;
  assign n21039 = ( ~n3306 & n3663 ) | ( ~n3306 & n21038 ) | ( n3663 & n21038 ) ;
  assign n21040 = ( n6133 & n10583 ) | ( n6133 & ~n21039 ) | ( n10583 & ~n21039 ) ;
  assign n21041 = n12407 ^ n6747 ^ n2171 ;
  assign n21042 = n21041 ^ n11936 ^ n11849 ;
  assign n21043 = n14006 ^ n11142 ^ n6019 ;
  assign n21044 = n5477 ^ n4210 ^ n1959 ;
  assign n21045 = n21044 ^ n13010 ^ n3659 ;
  assign n21046 = n9895 ^ n4537 ^ n1143 ;
  assign n21047 = n16606 ^ n9811 ^ n4945 ;
  assign n21048 = ( n6568 & n21046 ) | ( n6568 & n21047 ) | ( n21046 & n21047 ) ;
  assign n21049 = n9747 ^ n7357 ^ n892 ;
  assign n21050 = ( ~n4734 & n10979 ) | ( ~n4734 & n21049 ) | ( n10979 & n21049 ) ;
  assign n21051 = ( n819 & n8154 ) | ( n819 & n11760 ) | ( n8154 & n11760 ) ;
  assign n21052 = ( n20532 & n21050 ) | ( n20532 & ~n21051 ) | ( n21050 & ~n21051 ) ;
  assign n21053 = ( n6918 & n10161 ) | ( n6918 & n13459 ) | ( n10161 & n13459 ) ;
  assign n21054 = ( n2665 & n5588 ) | ( n2665 & n14220 ) | ( n5588 & n14220 ) ;
  assign n21055 = n7572 ^ n3102 ^ n1059 ;
  assign n21056 = ( ~n1868 & n3426 ) | ( ~n1868 & n12454 ) | ( n3426 & n12454 ) ;
  assign n21057 = ( n17352 & n21055 ) | ( n17352 & n21056 ) | ( n21055 & n21056 ) ;
  assign n21058 = ( n5515 & n21054 ) | ( n5515 & n21057 ) | ( n21054 & n21057 ) ;
  assign n21059 = ( n2234 & n3707 ) | ( n2234 & ~n11350 ) | ( n3707 & ~n11350 ) ;
  assign n21060 = ( n837 & n15883 ) | ( n837 & ~n21059 ) | ( n15883 & ~n21059 ) ;
  assign n21061 = n21060 ^ n10351 ^ n6241 ;
  assign n21063 = n4009 ^ n3437 ^ n2308 ;
  assign n21062 = ( n1056 & n4682 ) | ( n1056 & ~n7163 ) | ( n4682 & ~n7163 ) ;
  assign n21064 = n21063 ^ n21062 ^ n4823 ;
  assign n21065 = n21064 ^ n8122 ^ n6567 ;
  assign n21066 = n21065 ^ n20531 ^ n459 ;
  assign n21067 = n6704 ^ n4114 ^ n280 ;
  assign n21068 = n19072 ^ n18159 ^ n1619 ;
  assign n21069 = n21068 ^ n15998 ^ n5079 ;
  assign n21070 = ( n196 & n16757 ) | ( n196 & ~n21069 ) | ( n16757 & ~n21069 ) ;
  assign n21071 = n21070 ^ n15998 ^ n13189 ;
  assign n21072 = ( ~n672 & n9665 ) | ( ~n672 & n20186 ) | ( n9665 & n20186 ) ;
  assign n21073 = n21072 ^ n14801 ^ n5685 ;
  assign n21074 = ( n21067 & n21071 ) | ( n21067 & ~n21073 ) | ( n21071 & ~n21073 ) ;
  assign n21075 = ( ~n6541 & n8228 ) | ( ~n6541 & n9551 ) | ( n8228 & n9551 ) ;
  assign n21076 = ( n2748 & n3388 ) | ( n2748 & n6866 ) | ( n3388 & n6866 ) ;
  assign n21077 = n21076 ^ n2617 ^ n1162 ;
  assign n21078 = n11431 ^ n767 ^ n600 ;
  assign n21079 = ( n3749 & n4374 ) | ( n3749 & n17613 ) | ( n4374 & n17613 ) ;
  assign n21080 = n12344 ^ n9947 ^ n8236 ;
  assign n21081 = ( n3247 & n16219 ) | ( n3247 & ~n16438 ) | ( n16219 & ~n16438 ) ;
  assign n21082 = ( n12818 & n21080 ) | ( n12818 & n21081 ) | ( n21080 & n21081 ) ;
  assign n21083 = ( n3069 & ~n19194 ) | ( n3069 & n19897 ) | ( ~n19194 & n19897 ) ;
  assign n21084 = n11073 ^ n8502 ^ n3248 ;
  assign n21085 = ( n10636 & n11610 ) | ( n10636 & ~n21084 ) | ( n11610 & ~n21084 ) ;
  assign n21086 = ( ~n3851 & n11202 ) | ( ~n3851 & n21085 ) | ( n11202 & n21085 ) ;
  assign n21087 = n6471 ^ n2934 ^ n199 ;
  assign n21088 = ( ~n4838 & n6920 ) | ( ~n4838 & n21087 ) | ( n6920 & n21087 ) ;
  assign n21089 = n8951 ^ n2424 ^ n1419 ;
  assign n21090 = ( n3634 & n21088 ) | ( n3634 & n21089 ) | ( n21088 & n21089 ) ;
  assign n21091 = ( ~n3272 & n3422 ) | ( ~n3272 & n4756 ) | ( n3422 & n4756 ) ;
  assign n21092 = n21091 ^ n4995 ^ n1293 ;
  assign n21093 = n21092 ^ n9478 ^ n2744 ;
  assign n21094 = ( n15452 & ~n20565 ) | ( n15452 & n21093 ) | ( ~n20565 & n21093 ) ;
  assign n21097 = n17756 ^ n2630 ^ n1553 ;
  assign n21098 = ( n8215 & n10040 ) | ( n8215 & ~n21097 ) | ( n10040 & ~n21097 ) ;
  assign n21099 = n21098 ^ n15476 ^ n3431 ;
  assign n21095 = ( n2665 & ~n5898 ) | ( n2665 & n17343 ) | ( ~n5898 & n17343 ) ;
  assign n21096 = n21095 ^ n12947 ^ n1383 ;
  assign n21100 = n21099 ^ n21096 ^ n18298 ;
  assign n21101 = ( ~n3902 & n7551 ) | ( ~n3902 & n9222 ) | ( n7551 & n9222 ) ;
  assign n21102 = ( n9257 & ~n12263 ) | ( n9257 & n21101 ) | ( ~n12263 & n21101 ) ;
  assign n21103 = n21102 ^ n10319 ^ n7660 ;
  assign n21104 = ( n1075 & n6855 ) | ( n1075 & ~n8705 ) | ( n6855 & ~n8705 ) ;
  assign n21105 = ( ~n14847 & n16115 ) | ( ~n14847 & n21104 ) | ( n16115 & n21104 ) ;
  assign n21106 = ( n940 & n9795 ) | ( n940 & n11811 ) | ( n9795 & n11811 ) ;
  assign n21107 = ( ~n482 & n10108 ) | ( ~n482 & n17126 ) | ( n10108 & n17126 ) ;
  assign n21108 = n13789 ^ n12097 ^ n3954 ;
  assign n21109 = n21108 ^ n14762 ^ n7756 ;
  assign n21110 = ( n2134 & n21107 ) | ( n2134 & n21109 ) | ( n21107 & n21109 ) ;
  assign n21111 = n21110 ^ n15915 ^ n12905 ;
  assign n21112 = ( n10429 & ~n14514 ) | ( n10429 & n21111 ) | ( ~n14514 & n21111 ) ;
  assign n21116 = ( n6114 & n7781 ) | ( n6114 & n10264 ) | ( n7781 & n10264 ) ;
  assign n21117 = n21116 ^ n16381 ^ n10495 ;
  assign n21118 = n21117 ^ n12317 ^ n6592 ;
  assign n21113 = n17399 ^ n7102 ^ n2964 ;
  assign n21114 = ( ~n7375 & n8385 ) | ( ~n7375 & n13608 ) | ( n8385 & n13608 ) ;
  assign n21115 = ( n3440 & n21113 ) | ( n3440 & ~n21114 ) | ( n21113 & ~n21114 ) ;
  assign n21119 = n21118 ^ n21115 ^ n9593 ;
  assign n21120 = ( n17264 & n18276 ) | ( n17264 & n21119 ) | ( n18276 & n21119 ) ;
  assign n21121 = n9673 ^ n1971 ^ n1274 ;
  assign n21125 = n7187 ^ n6164 ^ n5839 ;
  assign n21124 = n7969 ^ n2604 ^ n2432 ;
  assign n21122 = ( n1998 & ~n3594 ) | ( n1998 & n6108 ) | ( ~n3594 & n6108 ) ;
  assign n21123 = n21122 ^ n11021 ^ n1028 ;
  assign n21126 = n21125 ^ n21124 ^ n21123 ;
  assign n21127 = ( n1328 & ~n4819 ) | ( n1328 & n5588 ) | ( ~n4819 & n5588 ) ;
  assign n21128 = n21127 ^ n10406 ^ n2754 ;
  assign n21129 = n21128 ^ n20810 ^ n14018 ;
  assign n21132 = n15666 ^ n8053 ^ n5363 ;
  assign n21133 = n21132 ^ n5736 ^ n4758 ;
  assign n21130 = n15840 ^ n1857 ^ n334 ;
  assign n21131 = n21130 ^ n20621 ^ n15392 ;
  assign n21134 = n21133 ^ n21131 ^ n12088 ;
  assign n21135 = n16815 ^ n5362 ^ n354 ;
  assign n21136 = n11673 ^ n7483 ^ n6074 ;
  assign n21137 = ( ~n5483 & n17979 ) | ( ~n5483 & n21136 ) | ( n17979 & n21136 ) ;
  assign n21138 = n21137 ^ n19148 ^ n10532 ;
  assign n21139 = ( n10173 & n16438 ) | ( n10173 & ~n21138 ) | ( n16438 & ~n21138 ) ;
  assign n21140 = ( n981 & n1884 ) | ( n981 & n6096 ) | ( n1884 & n6096 ) ;
  assign n21141 = n9471 ^ n5132 ^ n135 ;
  assign n21142 = ( n10844 & ~n15148 ) | ( n10844 & n21141 ) | ( ~n15148 & n21141 ) ;
  assign n21143 = ( n6854 & ~n10549 ) | ( n6854 & n21142 ) | ( ~n10549 & n21142 ) ;
  assign n21144 = ( n6086 & n19023 ) | ( n6086 & ~n21143 ) | ( n19023 & ~n21143 ) ;
  assign n21145 = n20841 ^ n16456 ^ n9266 ;
  assign n21148 = n4236 ^ n715 ^ n336 ;
  assign n21146 = n11395 ^ n1353 ^ n429 ;
  assign n21147 = n21146 ^ n3230 ^ n454 ;
  assign n21149 = n21148 ^ n21147 ^ n4753 ;
  assign n21150 = n18486 ^ n7190 ^ n5834 ;
  assign n21151 = n21150 ^ n10650 ^ n9434 ;
  assign n21152 = ( n3566 & n4157 ) | ( n3566 & ~n14911 ) | ( n4157 & ~n14911 ) ;
  assign n21153 = ( n1690 & n10889 ) | ( n1690 & n15066 ) | ( n10889 & n15066 ) ;
  assign n21154 = n21153 ^ n20908 ^ n20054 ;
  assign n21155 = n4397 ^ n219 ^ x29 ;
  assign n21156 = ( n5248 & n5682 ) | ( n5248 & ~n21155 ) | ( n5682 & ~n21155 ) ;
  assign n21157 = n21156 ^ n19351 ^ n13507 ;
  assign n21158 = ( n1034 & ~n12780 ) | ( n1034 & n21157 ) | ( ~n12780 & n21157 ) ;
  assign n21159 = ( ~n5577 & n18769 ) | ( ~n5577 & n21158 ) | ( n18769 & n21158 ) ;
  assign n21160 = n9968 ^ n6376 ^ n5524 ;
  assign n21161 = ( n1944 & ~n3187 ) | ( n1944 & n12744 ) | ( ~n3187 & n12744 ) ;
  assign n21162 = ( n6331 & ~n16779 ) | ( n6331 & n21161 ) | ( ~n16779 & n21161 ) ;
  assign n21163 = ( n13004 & ~n21160 ) | ( n13004 & n21162 ) | ( ~n21160 & n21162 ) ;
  assign n21164 = n18288 ^ n9751 ^ n5553 ;
  assign n21165 = ( n6948 & ~n10013 ) | ( n6948 & n13436 ) | ( ~n10013 & n13436 ) ;
  assign n21166 = ( ~n3574 & n3744 ) | ( ~n3574 & n4045 ) | ( n3744 & n4045 ) ;
  assign n21167 = n21166 ^ n2406 ^ n318 ;
  assign n21168 = ( n3212 & n21165 ) | ( n3212 & ~n21167 ) | ( n21165 & ~n21167 ) ;
  assign n21169 = ( ~n9263 & n12001 ) | ( ~n9263 & n21168 ) | ( n12001 & n21168 ) ;
  assign n21170 = ( ~n3478 & n12448 ) | ( ~n3478 & n12659 ) | ( n12448 & n12659 ) ;
  assign n21171 = n21170 ^ n7043 ^ n2862 ;
  assign n21175 = ( n2396 & n14102 ) | ( n2396 & n14644 ) | ( n14102 & n14644 ) ;
  assign n21172 = ( n2529 & ~n4639 ) | ( n2529 & n12763 ) | ( ~n4639 & n12763 ) ;
  assign n21173 = n21172 ^ n2612 ^ n1259 ;
  assign n21174 = n21173 ^ n5274 ^ n1378 ;
  assign n21176 = n21175 ^ n21174 ^ n18489 ;
  assign n21177 = n20904 ^ n5973 ^ n3450 ;
  assign n21178 = ( ~n6229 & n10687 ) | ( ~n6229 & n20230 ) | ( n10687 & n20230 ) ;
  assign n21179 = ( n1502 & n1955 ) | ( n1502 & n2769 ) | ( n1955 & n2769 ) ;
  assign n21180 = ( n10605 & ~n12975 ) | ( n10605 & n21179 ) | ( ~n12975 & n21179 ) ;
  assign n21181 = ( n1773 & n2279 ) | ( n1773 & ~n3453 ) | ( n2279 & ~n3453 ) ;
  assign n21182 = n15844 ^ n9410 ^ n3061 ;
  assign n21183 = ( n15040 & n21181 ) | ( n15040 & n21182 ) | ( n21181 & n21182 ) ;
  assign n21184 = n20727 ^ n14683 ^ n13700 ;
  assign n21185 = n21184 ^ n14371 ^ n7186 ;
  assign n21186 = ( ~n1386 & n13088 ) | ( ~n1386 & n14680 ) | ( n13088 & n14680 ) ;
  assign n21187 = n21186 ^ n12523 ^ n11031 ;
  assign n21188 = ( ~n7879 & n10664 ) | ( ~n7879 & n14197 ) | ( n10664 & n14197 ) ;
  assign n21189 = n19020 ^ n10403 ^ n327 ;
  assign n21190 = ( n3622 & n9090 ) | ( n3622 & ~n10539 ) | ( n9090 & ~n10539 ) ;
  assign n21191 = n21190 ^ n10547 ^ n1136 ;
  assign n21192 = ( n2601 & n5100 ) | ( n2601 & ~n21191 ) | ( n5100 & ~n21191 ) ;
  assign n21193 = ( n807 & n1245 ) | ( n807 & ~n5758 ) | ( n1245 & ~n5758 ) ;
  assign n21194 = n19897 ^ n11469 ^ n2290 ;
  assign n21195 = n21194 ^ n16722 ^ n8296 ;
  assign n21196 = n10412 ^ n7798 ^ n1149 ;
  assign n21197 = n21196 ^ n13828 ^ n12239 ;
  assign n21198 = n11878 ^ n10688 ^ n7186 ;
  assign n21199 = ( n7421 & ~n12078 ) | ( n7421 & n21198 ) | ( ~n12078 & n21198 ) ;
  assign n21200 = ( n686 & n12606 ) | ( n686 & n21199 ) | ( n12606 & n21199 ) ;
  assign n21205 = ( n1952 & n3476 ) | ( n1952 & n9778 ) | ( n3476 & n9778 ) ;
  assign n21206 = n21205 ^ n5701 ^ n1505 ;
  assign n21204 = ( n651 & ~n900 ) | ( n651 & n11334 ) | ( ~n900 & n11334 ) ;
  assign n21207 = n21206 ^ n21204 ^ n9582 ;
  assign n21203 = n11737 ^ n5573 ^ n1769 ;
  assign n21201 = ( n2860 & n5295 ) | ( n2860 & ~n12061 ) | ( n5295 & ~n12061 ) ;
  assign n21202 = n21201 ^ n20215 ^ n10875 ;
  assign n21208 = n21207 ^ n21203 ^ n21202 ;
  assign n21212 = n6616 ^ n5734 ^ n2543 ;
  assign n21209 = ( n3105 & ~n6639 ) | ( n3105 & n14127 ) | ( ~n6639 & n14127 ) ;
  assign n21210 = n21209 ^ n10571 ^ n6039 ;
  assign n21211 = ( n8288 & n13759 ) | ( n8288 & ~n21210 ) | ( n13759 & ~n21210 ) ;
  assign n21213 = n21212 ^ n21211 ^ n10485 ;
  assign n21214 = n21213 ^ n18041 ^ n3524 ;
  assign n21215 = n17466 ^ n3025 ^ x20 ;
  assign n21216 = ( ~n13329 & n15379 ) | ( ~n13329 & n20192 ) | ( n15379 & n20192 ) ;
  assign n21217 = n21216 ^ n11481 ^ n9755 ;
  assign n21218 = n21217 ^ n11038 ^ n8112 ;
  assign n21219 = n20475 ^ n16237 ^ n11285 ;
  assign n21220 = n21219 ^ n7185 ^ n7154 ;
  assign n21221 = ( n3216 & n4328 ) | ( n3216 & ~n21220 ) | ( n4328 & ~n21220 ) ;
  assign n21222 = ( n10557 & ~n15936 ) | ( n10557 & n16420 ) | ( ~n15936 & n16420 ) ;
  assign n21223 = n12961 ^ n11952 ^ n9541 ;
  assign n21224 = ( n8800 & n18810 ) | ( n8800 & ~n21223 ) | ( n18810 & ~n21223 ) ;
  assign n21225 = ( n2273 & n2409 ) | ( n2273 & n15130 ) | ( n2409 & n15130 ) ;
  assign n21226 = n21225 ^ n12967 ^ n2138 ;
  assign n21227 = n11749 ^ n10911 ^ n1914 ;
  assign n21228 = n21227 ^ n17232 ^ n5455 ;
  assign n21229 = n19565 ^ n15439 ^ n12321 ;
  assign n21230 = ( n6531 & ~n17989 ) | ( n6531 & n21229 ) | ( ~n17989 & n21229 ) ;
  assign n21231 = n21230 ^ n5721 ^ n3260 ;
  assign n21232 = n12544 ^ n5530 ^ n284 ;
  assign n21233 = n21232 ^ n3221 ^ n3149 ;
  assign n21236 = n18150 ^ n14710 ^ n12294 ;
  assign n21234 = ( n2662 & ~n9521 ) | ( n2662 & n12784 ) | ( ~n9521 & n12784 ) ;
  assign n21235 = n21234 ^ n18173 ^ n2481 ;
  assign n21237 = n21236 ^ n21235 ^ n16105 ;
  assign n21238 = ( ~n2414 & n4282 ) | ( ~n2414 & n10693 ) | ( n4282 & n10693 ) ;
  assign n21239 = ( n5827 & ~n10881 ) | ( n5827 & n15391 ) | ( ~n10881 & n15391 ) ;
  assign n21240 = ( n5231 & n14009 ) | ( n5231 & n20951 ) | ( n14009 & n20951 ) ;
  assign n21241 = ( n12112 & n17343 ) | ( n12112 & n19818 ) | ( n17343 & n19818 ) ;
  assign n21242 = ( n11491 & n13106 ) | ( n11491 & n21241 ) | ( n13106 & n21241 ) ;
  assign n21243 = n21242 ^ n17987 ^ n3303 ;
  assign n21244 = ( ~n6726 & n10962 ) | ( ~n6726 & n12804 ) | ( n10962 & n12804 ) ;
  assign n21245 = n17671 ^ n14018 ^ n10054 ;
  assign n21246 = ( ~n2386 & n9201 ) | ( ~n2386 & n9937 ) | ( n9201 & n9937 ) ;
  assign n21247 = n21246 ^ n18144 ^ n3200 ;
  assign n21248 = n6746 ^ n5406 ^ n2058 ;
  assign n21250 = n11047 ^ n6357 ^ n5829 ;
  assign n21249 = n15514 ^ n8404 ^ n1258 ;
  assign n21251 = n21250 ^ n21249 ^ n11623 ;
  assign n21252 = n20263 ^ n2946 ^ n2117 ;
  assign n21253 = ( n21248 & n21251 ) | ( n21248 & ~n21252 ) | ( n21251 & ~n21252 ) ;
  assign n21254 = ( n4151 & n10154 ) | ( n4151 & ~n21253 ) | ( n10154 & ~n21253 ) ;
  assign n21255 = ( ~n1425 & n10171 ) | ( ~n1425 & n20753 ) | ( n10171 & n20753 ) ;
  assign n21256 = n8087 ^ n3951 ^ n1156 ;
  assign n21257 = ( n1630 & ~n11835 ) | ( n1630 & n21256 ) | ( ~n11835 & n21256 ) ;
  assign n21261 = ( n1709 & n10828 ) | ( n1709 & n16834 ) | ( n10828 & n16834 ) ;
  assign n21259 = ( n7867 & n9141 ) | ( n7867 & ~n13686 ) | ( n9141 & ~n13686 ) ;
  assign n21258 = ( n513 & n5845 ) | ( n513 & n6070 ) | ( n5845 & n6070 ) ;
  assign n21260 = n21259 ^ n21258 ^ n18012 ;
  assign n21262 = n21261 ^ n21260 ^ n6583 ;
  assign n21263 = n21262 ^ n20451 ^ n6808 ;
  assign n21269 = ( n2896 & n8770 ) | ( n2896 & n9473 ) | ( n8770 & n9473 ) ;
  assign n21264 = ( n1080 & ~n2852 ) | ( n1080 & n3763 ) | ( ~n2852 & n3763 ) ;
  assign n21265 = n21264 ^ n5410 ^ n1174 ;
  assign n21266 = n21265 ^ n11418 ^ n10148 ;
  assign n21267 = n16667 ^ n6288 ^ n602 ;
  assign n21268 = ( n19277 & n21266 ) | ( n19277 & n21267 ) | ( n21266 & n21267 ) ;
  assign n21270 = n21269 ^ n21268 ^ n19230 ;
  assign n21271 = n16911 ^ n12642 ^ n11621 ;
  assign n21272 = ( n3210 & n21270 ) | ( n3210 & ~n21271 ) | ( n21270 & ~n21271 ) ;
  assign n21273 = ( ~n2692 & n6221 ) | ( ~n2692 & n8904 ) | ( n6221 & n8904 ) ;
  assign n21274 = ( ~n4693 & n6217 ) | ( ~n4693 & n20520 ) | ( n6217 & n20520 ) ;
  assign n21275 = ( n260 & n5952 ) | ( n260 & ~n21274 ) | ( n5952 & ~n21274 ) ;
  assign n21276 = ( n20850 & n21273 ) | ( n20850 & ~n21275 ) | ( n21273 & ~n21275 ) ;
  assign n21279 = ( n712 & ~n11292 ) | ( n712 & n13578 ) | ( ~n11292 & n13578 ) ;
  assign n21277 = n7734 ^ n7503 ^ n1503 ;
  assign n21278 = ( ~n1245 & n19299 ) | ( ~n1245 & n21277 ) | ( n19299 & n21277 ) ;
  assign n21280 = n21279 ^ n21278 ^ n2110 ;
  assign n21281 = ( n13216 & n20035 ) | ( n13216 & ~n21280 ) | ( n20035 & ~n21280 ) ;
  assign n21282 = n13376 ^ n1444 ^ n892 ;
  assign n21283 = ( n159 & ~n3539 ) | ( n159 & n18559 ) | ( ~n3539 & n18559 ) ;
  assign n21284 = n21283 ^ n8203 ^ n1774 ;
  assign n21285 = ( n15220 & n21282 ) | ( n15220 & ~n21284 ) | ( n21282 & ~n21284 ) ;
  assign n21286 = ( n5768 & n17379 ) | ( n5768 & n21285 ) | ( n17379 & n21285 ) ;
  assign n21287 = ( n2836 & n5945 ) | ( n2836 & n10071 ) | ( n5945 & n10071 ) ;
  assign n21288 = n21287 ^ n19550 ^ n5905 ;
  assign n21289 = ( n6063 & ~n7006 ) | ( n6063 & n13646 ) | ( ~n7006 & n13646 ) ;
  assign n21290 = ( n7715 & n15952 ) | ( n7715 & n21289 ) | ( n15952 & n21289 ) ;
  assign n21291 = ( n3446 & n10000 ) | ( n3446 & n14567 ) | ( n10000 & n14567 ) ;
  assign n21292 = n9373 ^ n4463 ^ n938 ;
  assign n21294 = ( n5046 & ~n9133 ) | ( n5046 & n18528 ) | ( ~n9133 & n18528 ) ;
  assign n21293 = n16628 ^ n9007 ^ n7419 ;
  assign n21295 = n21294 ^ n21293 ^ n15908 ;
  assign n21296 = ( n12964 & n21292 ) | ( n12964 & ~n21295 ) | ( n21292 & ~n21295 ) ;
  assign n21297 = ( n2014 & n21291 ) | ( n2014 & ~n21296 ) | ( n21291 & ~n21296 ) ;
  assign n21298 = n18823 ^ n5544 ^ n3275 ;
  assign n21299 = ( n3617 & n13626 ) | ( n3617 & n21298 ) | ( n13626 & n21298 ) ;
  assign n21300 = n1957 ^ n1132 ^ n993 ;
  assign n21301 = ( ~n3156 & n11560 ) | ( ~n3156 & n21300 ) | ( n11560 & n21300 ) ;
  assign n21302 = ( n4656 & n21299 ) | ( n4656 & ~n21301 ) | ( n21299 & ~n21301 ) ;
  assign n21303 = ( n5232 & n11475 ) | ( n5232 & n21302 ) | ( n11475 & n21302 ) ;
  assign n21304 = n18392 ^ n18250 ^ n4154 ;
  assign n21305 = n21304 ^ n15263 ^ n4679 ;
  assign n21306 = n15868 ^ n9076 ^ n7484 ;
  assign n21307 = n9801 ^ n9630 ^ n2560 ;
  assign n21308 = n21307 ^ n10040 ^ n7831 ;
  assign n21309 = ( ~n953 & n7868 ) | ( ~n953 & n12420 ) | ( n7868 & n12420 ) ;
  assign n21310 = ( n1905 & n4609 ) | ( n1905 & ~n13546 ) | ( n4609 & ~n13546 ) ;
  assign n21311 = n21310 ^ n21170 ^ n17525 ;
  assign n21314 = n8639 ^ n7635 ^ n583 ;
  assign n21315 = n21314 ^ n15159 ^ n2633 ;
  assign n21316 = n21315 ^ n6693 ^ n821 ;
  assign n21312 = n17958 ^ n14632 ^ n4278 ;
  assign n21313 = n21312 ^ n8202 ^ n5785 ;
  assign n21317 = n21316 ^ n21313 ^ n1133 ;
  assign n21319 = ( ~n2735 & n3462 ) | ( ~n2735 & n11906 ) | ( n3462 & n11906 ) ;
  assign n21318 = ( n7276 & n13873 ) | ( n7276 & n16987 ) | ( n13873 & n16987 ) ;
  assign n21320 = n21319 ^ n21318 ^ n595 ;
  assign n21321 = ( n4391 & n4626 ) | ( n4391 & n4983 ) | ( n4626 & n4983 ) ;
  assign n21322 = ( ~n4151 & n6981 ) | ( ~n4151 & n21321 ) | ( n6981 & n21321 ) ;
  assign n21323 = ( n2265 & n7454 ) | ( n2265 & ~n13852 ) | ( n7454 & ~n13852 ) ;
  assign n21324 = n7616 ^ n7192 ^ n2344 ;
  assign n21325 = ( n5376 & n5785 ) | ( n5376 & ~n7774 ) | ( n5785 & ~n7774 ) ;
  assign n21326 = n13601 ^ n7760 ^ n798 ;
  assign n21327 = ( n1863 & n4944 ) | ( n1863 & ~n21326 ) | ( n4944 & ~n21326 ) ;
  assign n21328 = ( n5683 & n8818 ) | ( n5683 & ~n21327 ) | ( n8818 & ~n21327 ) ;
  assign n21333 = n12100 ^ n3897 ^ n3476 ;
  assign n21329 = ( n3850 & n6512 ) | ( n3850 & n7396 ) | ( n6512 & n7396 ) ;
  assign n21330 = ( n2260 & n7917 ) | ( n2260 & ~n21329 ) | ( n7917 & ~n21329 ) ;
  assign n21331 = ( ~n6209 & n13136 ) | ( ~n6209 & n21330 ) | ( n13136 & n21330 ) ;
  assign n21332 = n21331 ^ n15202 ^ n352 ;
  assign n21334 = n21333 ^ n21332 ^ n6267 ;
  assign n21337 = n12833 ^ n6214 ^ n4644 ;
  assign n21335 = ( ~n2548 & n3181 ) | ( ~n2548 & n7923 ) | ( n3181 & n7923 ) ;
  assign n21336 = n21335 ^ n5470 ^ n2944 ;
  assign n21338 = n21337 ^ n21336 ^ n8155 ;
  assign n21339 = n21338 ^ n12942 ^ n12769 ;
  assign n21340 = n15838 ^ n8322 ^ n2157 ;
  assign n21341 = ( ~n10715 & n21182 ) | ( ~n10715 & n21340 ) | ( n21182 & n21340 ) ;
  assign n21342 = n11330 ^ n10360 ^ n10223 ;
  assign n21343 = n21342 ^ n14141 ^ n9554 ;
  assign n21344 = ( ~n6623 & n13571 ) | ( ~n6623 & n20390 ) | ( n13571 & n20390 ) ;
  assign n21345 = ( ~n886 & n2923 ) | ( ~n886 & n14296 ) | ( n2923 & n14296 ) ;
  assign n21346 = ( n9952 & n11784 ) | ( n9952 & n13044 ) | ( n11784 & n13044 ) ;
  assign n21347 = ( n791 & ~n2972 ) | ( n791 & n8216 ) | ( ~n2972 & n8216 ) ;
  assign n21348 = ( n19208 & n21346 ) | ( n19208 & n21347 ) | ( n21346 & n21347 ) ;
  assign n21349 = ( x121 & n3037 ) | ( x121 & n7613 ) | ( n3037 & n7613 ) ;
  assign n21350 = ( n4353 & n8546 ) | ( n4353 & ~n21349 ) | ( n8546 & ~n21349 ) ;
  assign n21351 = n18632 ^ n11242 ^ n9778 ;
  assign n21352 = ( n6125 & n8406 ) | ( n6125 & n21351 ) | ( n8406 & n21351 ) ;
  assign n21353 = n21076 ^ n7299 ^ n3187 ;
  assign n21354 = n21353 ^ n17013 ^ n16984 ;
  assign n21355 = n21354 ^ n21207 ^ n4222 ;
  assign n21356 = n17315 ^ n5555 ^ n752 ;
  assign n21357 = n20605 ^ n16253 ^ n10409 ;
  assign n21358 = ( n3221 & ~n5401 ) | ( n3221 & n21357 ) | ( ~n5401 & n21357 ) ;
  assign n21359 = n7919 ^ n1911 ^ n721 ;
  assign n21360 = ( ~n1205 & n4617 ) | ( ~n1205 & n21359 ) | ( n4617 & n21359 ) ;
  assign n21361 = n20551 ^ n11118 ^ n135 ;
  assign n21362 = ( n2391 & ~n9015 ) | ( n2391 & n21361 ) | ( ~n9015 & n21361 ) ;
  assign n21365 = n3138 ^ n802 ^ n245 ;
  assign n21363 = ( n3072 & n5959 ) | ( n3072 & n12465 ) | ( n5959 & n12465 ) ;
  assign n21364 = n21363 ^ n3886 ^ n1951 ;
  assign n21366 = n21365 ^ n21364 ^ n18139 ;
  assign n21367 = ( n4353 & n7382 ) | ( n4353 & ~n21366 ) | ( n7382 & ~n21366 ) ;
  assign n21368 = n19930 ^ n2403 ^ n639 ;
  assign n21369 = ( n4504 & ~n13900 ) | ( n4504 & n15106 ) | ( ~n13900 & n15106 ) ;
  assign n21370 = ( n15890 & ~n21368 ) | ( n15890 & n21369 ) | ( ~n21368 & n21369 ) ;
  assign n21371 = ( n3018 & n18581 ) | ( n3018 & n21370 ) | ( n18581 & n21370 ) ;
  assign n21372 = ( ~n1122 & n1896 ) | ( ~n1122 & n3674 ) | ( n1896 & n3674 ) ;
  assign n21373 = n21372 ^ n12367 ^ n1291 ;
  assign n21374 = ( n5282 & n16749 ) | ( n5282 & n21373 ) | ( n16749 & n21373 ) ;
  assign n21375 = n10763 ^ n10283 ^ n6080 ;
  assign n21376 = ( n4420 & ~n17240 ) | ( n4420 & n21375 ) | ( ~n17240 & n21375 ) ;
  assign n21377 = n12532 ^ n8502 ^ n2933 ;
  assign n21378 = n21377 ^ n19798 ^ n16370 ;
  assign n21379 = n21378 ^ n4748 ^ n350 ;
  assign n21380 = n21056 ^ n7078 ^ n6254 ;
  assign n21381 = ( ~n14062 & n18951 ) | ( ~n14062 & n21380 ) | ( n18951 & n21380 ) ;
  assign n21382 = ( n7972 & ~n8524 ) | ( n7972 & n14313 ) | ( ~n8524 & n14313 ) ;
  assign n21383 = ( n1001 & n10320 ) | ( n1001 & n13238 ) | ( n10320 & n13238 ) ;
  assign n21384 = ( n944 & ~n1032 ) | ( n944 & n14655 ) | ( ~n1032 & n14655 ) ;
  assign n21385 = ( ~n10606 & n18866 ) | ( ~n10606 & n21384 ) | ( n18866 & n21384 ) ;
  assign n21386 = ( n2084 & ~n15758 ) | ( n2084 & n21385 ) | ( ~n15758 & n21385 ) ;
  assign n21387 = ( ~n450 & n8843 ) | ( ~n450 & n21386 ) | ( n8843 & n21386 ) ;
  assign n21388 = ( n21382 & ~n21383 ) | ( n21382 & n21387 ) | ( ~n21383 & n21387 ) ;
  assign n21389 = n15481 ^ n11613 ^ n4605 ;
  assign n21390 = n18299 ^ n14687 ^ n6747 ;
  assign n21391 = ( ~n15444 & n18002 ) | ( ~n15444 & n21390 ) | ( n18002 & n21390 ) ;
  assign n21392 = ( n1612 & n11406 ) | ( n1612 & ~n16379 ) | ( n11406 & ~n16379 ) ;
  assign n21393 = n21392 ^ n12558 ^ n2994 ;
  assign n21394 = ( ~n18125 & n20011 ) | ( ~n18125 & n21393 ) | ( n20011 & n21393 ) ;
  assign n21395 = ( n4703 & n13404 ) | ( n4703 & n19517 ) | ( n13404 & n19517 ) ;
  assign n21396 = n15496 ^ n8304 ^ n7734 ;
  assign n21397 = ( n7423 & n11119 ) | ( n7423 & n17240 ) | ( n11119 & n17240 ) ;
  assign n21398 = ( n19355 & ~n21396 ) | ( n19355 & n21397 ) | ( ~n21396 & n21397 ) ;
  assign n21399 = ( n10950 & n16339 ) | ( n10950 & ~n21398 ) | ( n16339 & ~n21398 ) ;
  assign n21400 = n20051 ^ n4306 ^ n3980 ;
  assign n21401 = ( ~n600 & n3617 ) | ( ~n600 & n5675 ) | ( n3617 & n5675 ) ;
  assign n21402 = n21401 ^ n12045 ^ n7651 ;
  assign n21403 = ( ~n4612 & n10057 ) | ( ~n4612 & n21402 ) | ( n10057 & n21402 ) ;
  assign n21404 = ( n7406 & n18401 ) | ( n7406 & ~n21403 ) | ( n18401 & ~n21403 ) ;
  assign n21405 = ( ~n667 & n5833 ) | ( ~n667 & n6306 ) | ( n5833 & n6306 ) ;
  assign n21406 = n21405 ^ n9565 ^ n2218 ;
  assign n21407 = ( n178 & n4800 ) | ( n178 & ~n21406 ) | ( n4800 & ~n21406 ) ;
  assign n21408 = n21407 ^ n9440 ^ n4104 ;
  assign n21409 = ( n936 & ~n9008 ) | ( n936 & n14650 ) | ( ~n9008 & n14650 ) ;
  assign n21410 = ( n5233 & ~n14327 ) | ( n5233 & n18090 ) | ( ~n14327 & n18090 ) ;
  assign n21411 = ( n19339 & n21409 ) | ( n19339 & n21410 ) | ( n21409 & n21410 ) ;
  assign n21412 = ( n10189 & n10360 ) | ( n10189 & ~n21411 ) | ( n10360 & ~n21411 ) ;
  assign n21413 = ( n882 & n6868 ) | ( n882 & n7922 ) | ( n6868 & n7922 ) ;
  assign n21414 = n21413 ^ n20406 ^ n15849 ;
  assign n21415 = n21414 ^ n18086 ^ n3838 ;
  assign n21416 = n9658 ^ n8799 ^ n678 ;
  assign n21417 = n11908 ^ n1109 ^ x69 ;
  assign n21418 = n21417 ^ n13053 ^ n6714 ;
  assign n21419 = n21418 ^ n17894 ^ n2944 ;
  assign n21420 = ( n5249 & ~n21416 ) | ( n5249 & n21419 ) | ( ~n21416 & n21419 ) ;
  assign n21421 = n11069 ^ n2532 ^ n955 ;
  assign n21422 = ( n1312 & ~n2430 ) | ( n1312 & n5273 ) | ( ~n2430 & n5273 ) ;
  assign n21423 = ( n6845 & ~n15499 ) | ( n6845 & n21422 ) | ( ~n15499 & n21422 ) ;
  assign n21424 = n12882 ^ n4097 ^ n3860 ;
  assign n21425 = ( ~n7493 & n13360 ) | ( ~n7493 & n21424 ) | ( n13360 & n21424 ) ;
  assign n21426 = ( n1556 & n20748 ) | ( n1556 & n21160 ) | ( n20748 & n21160 ) ;
  assign n21427 = ( n1111 & n5172 ) | ( n1111 & n14455 ) | ( n5172 & n14455 ) ;
  assign n21428 = n21427 ^ n15683 ^ n4000 ;
  assign n21429 = n4006 ^ n2381 ^ n638 ;
  assign n21430 = ( n1082 & n20289 ) | ( n1082 & n21429 ) | ( n20289 & n21429 ) ;
  assign n21431 = n21430 ^ n18469 ^ n15121 ;
  assign n21433 = n8865 ^ n6463 ^ n723 ;
  assign n21432 = ( ~n6666 & n10380 ) | ( ~n6666 & n14549 ) | ( n10380 & n14549 ) ;
  assign n21434 = n21433 ^ n21432 ^ n12576 ;
  assign n21435 = ( ~n2177 & n2603 ) | ( ~n2177 & n5262 ) | ( n2603 & n5262 ) ;
  assign n21436 = ( n2928 & ~n3297 ) | ( n2928 & n10207 ) | ( ~n3297 & n10207 ) ;
  assign n21437 = ( ~n15180 & n21435 ) | ( ~n15180 & n21436 ) | ( n21435 & n21436 ) ;
  assign n21438 = n21437 ^ n11364 ^ n3399 ;
  assign n21439 = n7132 ^ n5050 ^ n2178 ;
  assign n21440 = n11623 ^ n9199 ^ n1155 ;
  assign n21441 = ( ~n9717 & n10095 ) | ( ~n9717 & n13091 ) | ( n10095 & n13091 ) ;
  assign n21442 = ( n8655 & ~n21440 ) | ( n8655 & n21441 ) | ( ~n21440 & n21441 ) ;
  assign n21443 = n21442 ^ n15827 ^ n7202 ;
  assign n21444 = ( n1869 & n12787 ) | ( n1869 & ~n14806 ) | ( n12787 & ~n14806 ) ;
  assign n21445 = n21444 ^ n11449 ^ n1352 ;
  assign n21446 = n21445 ^ n17973 ^ n729 ;
  assign n21447 = ( n7456 & n17426 ) | ( n7456 & n21446 ) | ( n17426 & n21446 ) ;
  assign n21448 = n21256 ^ n10139 ^ n2748 ;
  assign n21449 = ( ~n268 & n3734 ) | ( ~n268 & n5280 ) | ( n3734 & n5280 ) ;
  assign n21450 = ( n3175 & n11181 ) | ( n3175 & n21449 ) | ( n11181 & n21449 ) ;
  assign n21451 = n21450 ^ n9252 ^ n9026 ;
  assign n21452 = ( ~n1034 & n7741 ) | ( ~n1034 & n10657 ) | ( n7741 & n10657 ) ;
  assign n21453 = n21452 ^ n11455 ^ n7988 ;
  assign n21454 = n17121 ^ n3865 ^ n474 ;
  assign n21455 = ( n10864 & n19631 ) | ( n10864 & ~n21454 ) | ( n19631 & ~n21454 ) ;
  assign n21456 = n21455 ^ n20029 ^ n9285 ;
  assign n21457 = ( ~n2305 & n10115 ) | ( ~n2305 & n20011 ) | ( n10115 & n20011 ) ;
  assign n21458 = n8660 ^ n7803 ^ n5808 ;
  assign n21459 = n21458 ^ n13323 ^ n12852 ;
  assign n21461 = n16124 ^ n14579 ^ n460 ;
  assign n21460 = ( n6285 & n17832 ) | ( n6285 & n18766 ) | ( n17832 & n18766 ) ;
  assign n21462 = n21461 ^ n21460 ^ n3089 ;
  assign n21463 = n21462 ^ n9731 ^ n9289 ;
  assign n21464 = ( n3275 & ~n9445 ) | ( n3275 & n13548 ) | ( ~n9445 & n13548 ) ;
  assign n21465 = n15034 ^ n13734 ^ n6050 ;
  assign n21466 = ( n2040 & n12506 ) | ( n2040 & n21465 ) | ( n12506 & n21465 ) ;
  assign n21467 = ( n1392 & ~n21464 ) | ( n1392 & n21466 ) | ( ~n21464 & n21466 ) ;
  assign n21468 = ( n7609 & n21463 ) | ( n7609 & ~n21467 ) | ( n21463 & ~n21467 ) ;
  assign n21469 = ( n11980 & ~n13123 ) | ( n11980 & n18653 ) | ( ~n13123 & n18653 ) ;
  assign n21470 = ( n557 & n8960 ) | ( n557 & n13593 ) | ( n8960 & n13593 ) ;
  assign n21471 = ( n9145 & n14494 ) | ( n9145 & n21470 ) | ( n14494 & n21470 ) ;
  assign n21472 = n21471 ^ n8886 ^ n5706 ;
  assign n21473 = ( n3672 & n4478 ) | ( n3672 & n12294 ) | ( n4478 & n12294 ) ;
  assign n21474 = n21473 ^ n15872 ^ n3014 ;
  assign n21476 = n20237 ^ n13352 ^ n12234 ;
  assign n21475 = n8231 ^ n6147 ^ n2877 ;
  assign n21477 = n21476 ^ n21475 ^ n13773 ;
  assign n21479 = ( ~n5761 & n13265 ) | ( ~n5761 & n17872 ) | ( n13265 & n17872 ) ;
  assign n21478 = ( n475 & ~n2374 ) | ( n475 & n7090 ) | ( ~n2374 & n7090 ) ;
  assign n21480 = n21479 ^ n21478 ^ n11769 ;
  assign n21481 = n7801 ^ n6726 ^ n466 ;
  assign n21482 = n21481 ^ n16793 ^ n7016 ;
  assign n21483 = n17177 ^ n13457 ^ n389 ;
  assign n21484 = ( n11209 & n21067 ) | ( n11209 & n21483 ) | ( n21067 & n21483 ) ;
  assign n21485 = ( ~n2353 & n10464 ) | ( ~n2353 & n13561 ) | ( n10464 & n13561 ) ;
  assign n21486 = n11029 ^ n10589 ^ n8749 ;
  assign n21487 = ( n4071 & n9364 ) | ( n4071 & n21486 ) | ( n9364 & n21486 ) ;
  assign n21488 = ( n6498 & n13411 ) | ( n6498 & n21487 ) | ( n13411 & n21487 ) ;
  assign n21489 = n21488 ^ n10948 ^ n7869 ;
  assign n21490 = ( n4550 & ~n16409 ) | ( n4550 & n21489 ) | ( ~n16409 & n21489 ) ;
  assign n21491 = n18262 ^ n17523 ^ n3284 ;
  assign n21492 = ( n948 & ~n8058 ) | ( n948 & n12185 ) | ( ~n8058 & n12185 ) ;
  assign n21493 = n21492 ^ n2454 ^ n1096 ;
  assign n21494 = ( n4279 & ~n6864 ) | ( n4279 & n10098 ) | ( ~n6864 & n10098 ) ;
  assign n21495 = n21494 ^ n15909 ^ n12828 ;
  assign n21496 = n13942 ^ n5827 ^ n952 ;
  assign n21497 = ( ~n7830 & n14019 ) | ( ~n7830 & n21496 ) | ( n14019 & n21496 ) ;
  assign n21503 = ( n8790 & n9270 ) | ( n8790 & ~n20868 ) | ( n9270 & ~n20868 ) ;
  assign n21501 = ( n6686 & n8066 ) | ( n6686 & ~n13552 ) | ( n8066 & ~n13552 ) ;
  assign n21502 = ( n6866 & n13912 ) | ( n6866 & n21501 ) | ( n13912 & n21501 ) ;
  assign n21504 = n21503 ^ n21502 ^ n3691 ;
  assign n21498 = ( ~n3409 & n4689 ) | ( ~n3409 & n9196 ) | ( n4689 & n9196 ) ;
  assign n21499 = n21498 ^ n18730 ^ n6142 ;
  assign n21500 = n21499 ^ n15422 ^ n7503 ;
  assign n21505 = n21504 ^ n21500 ^ n13590 ;
  assign n21508 = n20505 ^ n6906 ^ x98 ;
  assign n21506 = ( ~n3973 & n6177 ) | ( ~n3973 & n13872 ) | ( n6177 & n13872 ) ;
  assign n21507 = ( n5314 & n8889 ) | ( n5314 & ~n21506 ) | ( n8889 & ~n21506 ) ;
  assign n21509 = n21508 ^ n21507 ^ n15336 ;
  assign n21510 = ( n5665 & n12751 ) | ( n5665 & n21509 ) | ( n12751 & n21509 ) ;
  assign n21511 = n7985 ^ n7347 ^ n4592 ;
  assign n21512 = ( n9070 & n20519 ) | ( n9070 & ~n21511 ) | ( n20519 & ~n21511 ) ;
  assign n21513 = ( n12970 & n14838 ) | ( n12970 & n15343 ) | ( n14838 & n15343 ) ;
  assign n21514 = ( n1274 & n2092 ) | ( n1274 & n7506 ) | ( n2092 & n7506 ) ;
  assign n21515 = n21514 ^ n3855 ^ n3233 ;
  assign n21516 = ( n4584 & ~n4673 ) | ( n4584 & n15393 ) | ( ~n4673 & n15393 ) ;
  assign n21517 = ( n3203 & n18408 ) | ( n3203 & ~n21516 ) | ( n18408 & ~n21516 ) ;
  assign n21518 = ( n987 & ~n2225 ) | ( n987 & n5213 ) | ( ~n2225 & n5213 ) ;
  assign n21519 = ( ~n6553 & n11082 ) | ( ~n6553 & n21518 ) | ( n11082 & n21518 ) ;
  assign n21520 = ( n4171 & n9074 ) | ( n4171 & ~n21519 ) | ( n9074 & ~n21519 ) ;
  assign n21521 = n21354 ^ n12750 ^ n901 ;
  assign n21522 = ( n15972 & n16098 ) | ( n15972 & ~n21521 ) | ( n16098 & ~n21521 ) ;
  assign n21523 = ( n14437 & n20575 ) | ( n14437 & n21216 ) | ( n20575 & n21216 ) ;
  assign n21524 = ( n4716 & n7847 ) | ( n4716 & ~n21523 ) | ( n7847 & ~n21523 ) ;
  assign n21525 = n21524 ^ n17326 ^ n10811 ;
  assign n21526 = ( n3451 & ~n5465 ) | ( n3451 & n21525 ) | ( ~n5465 & n21525 ) ;
  assign n21527 = n20320 ^ n12385 ^ n4130 ;
  assign n21528 = ( n8743 & ~n14363 ) | ( n8743 & n18604 ) | ( ~n14363 & n18604 ) ;
  assign n21529 = ( ~n2305 & n17053 ) | ( ~n2305 & n21528 ) | ( n17053 & n21528 ) ;
  assign n21532 = n2910 ^ n1547 ^ n1224 ;
  assign n21530 = ( ~n4935 & n5478 ) | ( ~n4935 & n18563 ) | ( n5478 & n18563 ) ;
  assign n21531 = ( n2404 & n10749 ) | ( n2404 & n21530 ) | ( n10749 & n21530 ) ;
  assign n21533 = n21532 ^ n21531 ^ n6140 ;
  assign n21534 = ( n3717 & n6555 ) | ( n3717 & n9425 ) | ( n6555 & n9425 ) ;
  assign n21535 = ( n1457 & ~n3303 ) | ( n1457 & n21534 ) | ( ~n3303 & n21534 ) ;
  assign n21536 = n21535 ^ n8084 ^ n4087 ;
  assign n21537 = n7426 ^ n1791 ^ n1195 ;
  assign n21538 = ( ~n3723 & n21036 ) | ( ~n3723 & n21537 ) | ( n21036 & n21537 ) ;
  assign n21539 = n8267 ^ n2464 ^ n2234 ;
  assign n21540 = n16871 ^ n12568 ^ n5134 ;
  assign n21541 = ( ~n4768 & n19866 ) | ( ~n4768 & n21540 ) | ( n19866 & n21540 ) ;
  assign n21542 = ( n4989 & ~n7308 ) | ( n4989 & n15886 ) | ( ~n7308 & n15886 ) ;
  assign n21543 = ( ~n3625 & n7108 ) | ( ~n3625 & n8163 ) | ( n7108 & n8163 ) ;
  assign n21544 = n21543 ^ n12292 ^ n3172 ;
  assign n21545 = ( n1184 & ~n5887 ) | ( n1184 & n14896 ) | ( ~n5887 & n14896 ) ;
  assign n21546 = n21545 ^ n4060 ^ n3579 ;
  assign n21547 = n11871 ^ n8846 ^ n4171 ;
  assign n21551 = ( n312 & n14969 ) | ( n312 & n21264 ) | ( n14969 & n21264 ) ;
  assign n21549 = n14021 ^ n7333 ^ n6322 ;
  assign n21548 = ( ~n680 & n6025 ) | ( ~n680 & n14268 ) | ( n6025 & n14268 ) ;
  assign n21550 = n21549 ^ n21548 ^ n5022 ;
  assign n21552 = n21551 ^ n21550 ^ n382 ;
  assign n21553 = ( ~n2602 & n7560 ) | ( ~n2602 & n7852 ) | ( n7560 & n7852 ) ;
  assign n21554 = n21553 ^ n1893 ^ n886 ;
  assign n21555 = ( n21547 & n21552 ) | ( n21547 & ~n21554 ) | ( n21552 & ~n21554 ) ;
  assign n21556 = ( ~n21544 & n21546 ) | ( ~n21544 & n21555 ) | ( n21546 & n21555 ) ;
  assign n21557 = ( n1052 & n12848 ) | ( n1052 & ~n16700 ) | ( n12848 & ~n16700 ) ;
  assign n21558 = ( n2027 & n7466 ) | ( n2027 & ~n10780 ) | ( n7466 & ~n10780 ) ;
  assign n21559 = n21558 ^ n12974 ^ n1437 ;
  assign n21562 = ( n537 & n1056 ) | ( n537 & ~n8527 ) | ( n1056 & ~n8527 ) ;
  assign n21560 = ( n1316 & n3910 ) | ( n1316 & ~n4235 ) | ( n3910 & ~n4235 ) ;
  assign n21561 = ( n7240 & n20091 ) | ( n7240 & n21560 ) | ( n20091 & n21560 ) ;
  assign n21563 = n21562 ^ n21561 ^ n7849 ;
  assign n21568 = n12806 ^ n9127 ^ n5344 ;
  assign n21566 = ( n525 & n8285 ) | ( n525 & ~n17349 ) | ( n8285 & ~n17349 ) ;
  assign n21567 = ( n7181 & n16983 ) | ( n7181 & ~n21566 ) | ( n16983 & ~n21566 ) ;
  assign n21564 = ( n2062 & n4982 ) | ( n2062 & ~n5078 ) | ( n4982 & ~n5078 ) ;
  assign n21565 = n21564 ^ n16304 ^ n9666 ;
  assign n21569 = n21568 ^ n21567 ^ n21565 ;
  assign n21572 = n14860 ^ n4793 ^ n1866 ;
  assign n21570 = n15304 ^ n5399 ^ n4441 ;
  assign n21571 = ( n1453 & n3288 ) | ( n1453 & n21570 ) | ( n3288 & n21570 ) ;
  assign n21573 = n21572 ^ n21571 ^ n20635 ;
  assign n21574 = n21573 ^ n19778 ^ n14405 ;
  assign n21576 = ( n394 & n2395 ) | ( n394 & ~n2424 ) | ( n2395 & ~n2424 ) ;
  assign n21577 = n21576 ^ n16378 ^ n8828 ;
  assign n21575 = n20134 ^ n7648 ^ n2376 ;
  assign n21578 = n21577 ^ n21575 ^ n20327 ;
  assign n21579 = ( n2087 & ~n3896 ) | ( n2087 & n5161 ) | ( ~n3896 & n5161 ) ;
  assign n21580 = n21579 ^ n12841 ^ n5816 ;
  assign n21581 = ( ~n955 & n6875 ) | ( ~n955 & n8583 ) | ( n6875 & n8583 ) ;
  assign n21582 = ( ~n8733 & n20402 ) | ( ~n8733 & n21581 ) | ( n20402 & n21581 ) ;
  assign n21583 = ( n2053 & n18356 ) | ( n2053 & n21582 ) | ( n18356 & n21582 ) ;
  assign n21584 = ( n3987 & ~n15473 ) | ( n3987 & n21437 ) | ( ~n15473 & n21437 ) ;
  assign n21585 = n6403 ^ n1843 ^ n1040 ;
  assign n21586 = n16171 ^ n13360 ^ n5814 ;
  assign n21587 = ( n6063 & n21585 ) | ( n6063 & n21586 ) | ( n21585 & n21586 ) ;
  assign n21588 = ( n3981 & n12535 ) | ( n3981 & ~n20143 ) | ( n12535 & ~n20143 ) ;
  assign n21589 = ( n2146 & n5797 ) | ( n2146 & n21588 ) | ( n5797 & n21588 ) ;
  assign n21590 = n10121 ^ n2737 ^ n2333 ;
  assign n21591 = n21590 ^ n15118 ^ n2549 ;
  assign n21592 = ( ~n15308 & n21589 ) | ( ~n15308 & n21591 ) | ( n21589 & n21591 ) ;
  assign n21594 = ( n1046 & n4077 ) | ( n1046 & n8037 ) | ( n4077 & n8037 ) ;
  assign n21595 = n21594 ^ n17278 ^ n6849 ;
  assign n21593 = n11648 ^ n10738 ^ n4266 ;
  assign n21596 = n21595 ^ n21593 ^ n10435 ;
  assign n21597 = ( n13073 & ~n19679 ) | ( n13073 & n21373 ) | ( ~n19679 & n21373 ) ;
  assign n21598 = n17131 ^ n12755 ^ n2943 ;
  assign n21611 = ( ~n6362 & n7646 ) | ( ~n6362 & n11773 ) | ( n7646 & n11773 ) ;
  assign n21610 = ( n12831 & ~n14218 ) | ( n12831 & n14941 ) | ( ~n14218 & n14941 ) ;
  assign n21612 = n21611 ^ n21610 ^ n10222 ;
  assign n21607 = n12834 ^ n3181 ^ n2638 ;
  assign n21608 = ( n3800 & n9508 ) | ( n3800 & n21607 ) | ( n9508 & n21607 ) ;
  assign n21604 = ( ~n300 & n10049 ) | ( ~n300 & n12478 ) | ( n10049 & n12478 ) ;
  assign n21605 = n21604 ^ n8390 ^ n3937 ;
  assign n21606 = ( n12386 & n21107 ) | ( n12386 & ~n21605 ) | ( n21107 & ~n21605 ) ;
  assign n21609 = n21608 ^ n21606 ^ n17357 ;
  assign n21613 = n21612 ^ n21609 ^ n9097 ;
  assign n21599 = n9883 ^ n2581 ^ n1450 ;
  assign n21600 = ( n3691 & n4652 ) | ( n3691 & n6869 ) | ( n4652 & n6869 ) ;
  assign n21601 = ( n3742 & n12764 ) | ( n3742 & n21600 ) | ( n12764 & n21600 ) ;
  assign n21602 = ( ~n13871 & n21599 ) | ( ~n13871 & n21601 ) | ( n21599 & n21601 ) ;
  assign n21603 = ( n2949 & ~n4950 ) | ( n2949 & n21602 ) | ( ~n4950 & n21602 ) ;
  assign n21614 = n21613 ^ n21603 ^ n15336 ;
  assign n21615 = ( n5550 & ~n7202 ) | ( n5550 & n16641 ) | ( ~n7202 & n16641 ) ;
  assign n21616 = n14807 ^ n14149 ^ n10643 ;
  assign n21617 = n21616 ^ n7367 ^ n3869 ;
  assign n21618 = ( ~n2329 & n12936 ) | ( ~n2329 & n18528 ) | ( n12936 & n18528 ) ;
  assign n21619 = n21618 ^ n18934 ^ n7632 ;
  assign n21620 = n21619 ^ n15667 ^ n7914 ;
  assign n21621 = ( n4466 & n21617 ) | ( n4466 & ~n21620 ) | ( n21617 & ~n21620 ) ;
  assign n21622 = n21621 ^ n18222 ^ n658 ;
  assign n21624 = n8334 ^ n4401 ^ n518 ;
  assign n21623 = ( ~n3497 & n7583 ) | ( ~n3497 & n17986 ) | ( n7583 & n17986 ) ;
  assign n21625 = n21624 ^ n21623 ^ n241 ;
  assign n21627 = ( ~n2322 & n4944 ) | ( ~n2322 & n11928 ) | ( n4944 & n11928 ) ;
  assign n21628 = ( n3086 & n7298 ) | ( n3086 & n21627 ) | ( n7298 & n21627 ) ;
  assign n21629 = ( ~n10093 & n20718 ) | ( ~n10093 & n21628 ) | ( n20718 & n21628 ) ;
  assign n21630 = n21629 ^ n6956 ^ n5779 ;
  assign n21626 = n21098 ^ n10567 ^ n9393 ;
  assign n21631 = n21630 ^ n21626 ^ n11104 ;
  assign n21632 = ( n1247 & n11908 ) | ( n1247 & ~n18360 ) | ( n11908 & ~n18360 ) ;
  assign n21633 = ( ~n1564 & n16235 ) | ( ~n1564 & n21632 ) | ( n16235 & n21632 ) ;
  assign n21634 = n21633 ^ n9798 ^ n8622 ;
  assign n21635 = n20769 ^ n13642 ^ n2548 ;
  assign n21636 = ( ~n2214 & n2767 ) | ( ~n2214 & n12688 ) | ( n2767 & n12688 ) ;
  assign n21637 = n21636 ^ n9444 ^ n3568 ;
  assign n21638 = n15856 ^ n3125 ^ n452 ;
  assign n21639 = ( n7086 & n21107 ) | ( n7086 & n21638 ) | ( n21107 & n21638 ) ;
  assign n21640 = n19164 ^ n13585 ^ n9781 ;
  assign n21641 = ( n14653 & n16160 ) | ( n14653 & ~n17479 ) | ( n16160 & ~n17479 ) ;
  assign n21642 = ( n1050 & n11252 ) | ( n1050 & ~n11343 ) | ( n11252 & ~n11343 ) ;
  assign n21643 = n1933 ^ n1619 ^ x36 ;
  assign n21644 = n21643 ^ n13372 ^ n4590 ;
  assign n21645 = ( n6065 & n17792 ) | ( n6065 & ~n21644 ) | ( n17792 & ~n21644 ) ;
  assign n21646 = ( n4732 & n8848 ) | ( n4732 & ~n14993 ) | ( n8848 & ~n14993 ) ;
  assign n21647 = ( n4981 & ~n11358 ) | ( n4981 & n21646 ) | ( ~n11358 & n21646 ) ;
  assign n21648 = n21647 ^ n19097 ^ n6552 ;
  assign n21649 = ( n836 & n21645 ) | ( n836 & n21648 ) | ( n21645 & n21648 ) ;
  assign n21650 = n21649 ^ n19439 ^ n7374 ;
  assign n21651 = ( n4869 & n5926 ) | ( n4869 & ~n6064 ) | ( n5926 & ~n6064 ) ;
  assign n21652 = n6215 ^ n5768 ^ n3434 ;
  assign n21653 = n21652 ^ n16811 ^ n5104 ;
  assign n21654 = ( n4765 & ~n21651 ) | ( n4765 & n21653 ) | ( ~n21651 & n21653 ) ;
  assign n21655 = ( n6069 & n9116 ) | ( n6069 & ~n17589 ) | ( n9116 & ~n17589 ) ;
  assign n21656 = ( n438 & n7603 ) | ( n438 & ~n8100 ) | ( n7603 & ~n8100 ) ;
  assign n21657 = ( n8272 & n10690 ) | ( n8272 & n21656 ) | ( n10690 & n21656 ) ;
  assign n21658 = ( n18321 & ~n21655 ) | ( n18321 & n21657 ) | ( ~n21655 & n21657 ) ;
  assign n21659 = n16757 ^ n7536 ^ n690 ;
  assign n21660 = ( n8845 & n18583 ) | ( n8845 & ~n21659 ) | ( n18583 & ~n21659 ) ;
  assign n21663 = ( n4121 & n5172 ) | ( n4121 & n9281 ) | ( n5172 & n9281 ) ;
  assign n21662 = n6988 ^ n1078 ^ n937 ;
  assign n21661 = ( n1778 & ~n12379 ) | ( n1778 & n15929 ) | ( ~n12379 & n15929 ) ;
  assign n21664 = n21663 ^ n21662 ^ n21661 ;
  assign n21665 = ( n1967 & n19405 ) | ( n1967 & ~n21664 ) | ( n19405 & ~n21664 ) ;
  assign n21666 = n21665 ^ n2639 ^ n702 ;
  assign n21671 = ( ~n2535 & n3618 ) | ( ~n2535 & n18820 ) | ( n3618 & n18820 ) ;
  assign n21672 = n21671 ^ n13846 ^ n2027 ;
  assign n21668 = n5262 ^ n3618 ^ n2601 ;
  assign n21667 = ( ~n1134 & n1977 ) | ( ~n1134 & n12613 ) | ( n1977 & n12613 ) ;
  assign n21669 = n21668 ^ n21667 ^ n19501 ;
  assign n21670 = n21669 ^ n11897 ^ x75 ;
  assign n21673 = n21672 ^ n21670 ^ n4928 ;
  assign n21674 = n16510 ^ n14495 ^ n1318 ;
  assign n21675 = n21674 ^ n20165 ^ n9794 ;
  assign n21676 = ( ~n1561 & n6646 ) | ( ~n1561 & n8080 ) | ( n6646 & n8080 ) ;
  assign n21677 = ( n1589 & n3353 ) | ( n1589 & n4030 ) | ( n3353 & n4030 ) ;
  assign n21678 = ( n13123 & n21676 ) | ( n13123 & ~n21677 ) | ( n21676 & ~n21677 ) ;
  assign n21679 = n19534 ^ n12866 ^ n10304 ;
  assign n21680 = ( n16462 & n16791 ) | ( n16462 & n20138 ) | ( n16791 & n20138 ) ;
  assign n21681 = n11237 ^ n3162 ^ n352 ;
  assign n21682 = ( n3495 & n12269 ) | ( n3495 & n21681 ) | ( n12269 & n21681 ) ;
  assign n21683 = n21682 ^ n12565 ^ n10777 ;
  assign n21684 = n7011 ^ n4855 ^ n1749 ;
  assign n21685 = n21684 ^ n14419 ^ n6957 ;
  assign n21686 = ( n1424 & n11127 ) | ( n1424 & ~n21685 ) | ( n11127 & ~n21685 ) ;
  assign n21687 = ( n4061 & n16829 ) | ( n4061 & n21686 ) | ( n16829 & n21686 ) ;
  assign n21688 = n15393 ^ n8711 ^ n6983 ;
  assign n21689 = ( n755 & ~n3253 ) | ( n755 & n4623 ) | ( ~n3253 & n4623 ) ;
  assign n21690 = ( n1537 & ~n12153 ) | ( n1537 & n21689 ) | ( ~n12153 & n21689 ) ;
  assign n21691 = ( n855 & ~n21688 ) | ( n855 & n21690 ) | ( ~n21688 & n21690 ) ;
  assign n21692 = ( x111 & ~n355 ) | ( x111 & n12694 ) | ( ~n355 & n12694 ) ;
  assign n21693 = ( n4531 & n19192 ) | ( n4531 & n21692 ) | ( n19192 & n21692 ) ;
  assign n21694 = n21693 ^ n8226 ^ n4019 ;
  assign n21695 = ( n1132 & ~n18217 ) | ( n1132 & n18677 ) | ( ~n18217 & n18677 ) ;
  assign n21696 = ( ~n771 & n2281 ) | ( ~n771 & n21695 ) | ( n2281 & n21695 ) ;
  assign n21707 = ( n4825 & n5076 ) | ( n4825 & ~n10556 ) | ( n5076 & ~n10556 ) ;
  assign n21705 = n14041 ^ n9530 ^ n625 ;
  assign n21706 = n21705 ^ n9891 ^ n418 ;
  assign n21708 = n21707 ^ n21706 ^ n3371 ;
  assign n21697 = n7940 ^ n6296 ^ n862 ;
  assign n21698 = ( ~n9789 & n16353 ) | ( ~n9789 & n21697 ) | ( n16353 & n21697 ) ;
  assign n21699 = n21698 ^ n11894 ^ n1087 ;
  assign n21702 = n7033 ^ n5440 ^ n5279 ;
  assign n21701 = ( n837 & n2699 ) | ( n837 & n14627 ) | ( n2699 & n14627 ) ;
  assign n21700 = n20734 ^ n2452 ^ n2120 ;
  assign n21703 = n21702 ^ n21701 ^ n21700 ;
  assign n21704 = ( ~n6919 & n21699 ) | ( ~n6919 & n21703 ) | ( n21699 & n21703 ) ;
  assign n21709 = n21708 ^ n21704 ^ n16382 ;
  assign n21710 = n21521 ^ n17170 ^ n10755 ;
  assign n21711 = n19994 ^ n14948 ^ n5209 ;
  assign n21712 = n9727 ^ n7615 ^ n1742 ;
  assign n21713 = n15397 ^ n9039 ^ n5372 ;
  assign n21714 = n18406 ^ n10035 ^ n1858 ;
  assign n21715 = n21714 ^ n7975 ^ n6176 ;
  assign n21716 = n13424 ^ n4222 ^ n1188 ;
  assign n21717 = ( ~n1614 & n16264 ) | ( ~n1614 & n21716 ) | ( n16264 & n21716 ) ;
  assign n21718 = ( n1439 & n6741 ) | ( n1439 & ~n15733 ) | ( n6741 & ~n15733 ) ;
  assign n21719 = ( n2506 & n16991 ) | ( n2506 & ~n21718 ) | ( n16991 & ~n21718 ) ;
  assign n21720 = ( n7585 & n21717 ) | ( n7585 & n21719 ) | ( n21717 & n21719 ) ;
  assign n21724 = n14670 ^ n11945 ^ n3551 ;
  assign n21725 = n21724 ^ n12062 ^ n2054 ;
  assign n21723 = n10534 ^ n4872 ^ n1707 ;
  assign n21721 = ( n3689 & ~n12163 ) | ( n3689 & n13855 ) | ( ~n12163 & n13855 ) ;
  assign n21722 = ( n4580 & n11913 ) | ( n4580 & ~n21721 ) | ( n11913 & ~n21721 ) ;
  assign n21726 = n21725 ^ n21723 ^ n21722 ;
  assign n21727 = ( n1026 & ~n3476 ) | ( n1026 & n4627 ) | ( ~n3476 & n4627 ) ;
  assign n21728 = n16041 ^ n13103 ^ n5797 ;
  assign n21729 = ( n13386 & ~n21727 ) | ( n13386 & n21728 ) | ( ~n21727 & n21728 ) ;
  assign n21730 = n12005 ^ n8583 ^ n3532 ;
  assign n21731 = n19174 ^ n2516 ^ n2329 ;
  assign n21732 = n21731 ^ n19469 ^ n16410 ;
  assign n21733 = ( n21249 & ~n21730 ) | ( n21249 & n21732 ) | ( ~n21730 & n21732 ) ;
  assign n21734 = n19828 ^ n10392 ^ n2297 ;
  assign n21735 = n10905 ^ n3334 ^ n2622 ;
  assign n21736 = n21735 ^ n13705 ^ n6495 ;
  assign n21737 = n14510 ^ n2569 ^ n628 ;
  assign n21738 = ( n3586 & n17449 ) | ( n3586 & n21737 ) | ( n17449 & n21737 ) ;
  assign n21739 = n17381 ^ n6218 ^ n2220 ;
  assign n21740 = ( ~n2999 & n20250 ) | ( ~n2999 & n21739 ) | ( n20250 & n21739 ) ;
  assign n21741 = n15112 ^ n3304 ^ n730 ;
  assign n21744 = ( ~n3539 & n14067 ) | ( ~n3539 & n20983 ) | ( n14067 & n20983 ) ;
  assign n21742 = n13223 ^ n12183 ^ n11676 ;
  assign n21743 = ( ~n6795 & n6809 ) | ( ~n6795 & n21742 ) | ( n6809 & n21742 ) ;
  assign n21745 = n21744 ^ n21743 ^ n5993 ;
  assign n21746 = n21745 ^ n9161 ^ n2942 ;
  assign n21747 = ( n3051 & n3142 ) | ( n3051 & ~n21746 ) | ( n3142 & ~n21746 ) ;
  assign n21748 = n21396 ^ n11563 ^ n995 ;
  assign n21749 = ( n14973 & n19668 ) | ( n14973 & n21748 ) | ( n19668 & n21748 ) ;
  assign n21750 = ( ~n2228 & n7221 ) | ( ~n2228 & n21749 ) | ( n7221 & n21749 ) ;
  assign n21751 = n12617 ^ n7190 ^ n6627 ;
  assign n21752 = n13627 ^ n5323 ^ n2591 ;
  assign n21753 = ( ~n2636 & n8055 ) | ( ~n2636 & n21752 ) | ( n8055 & n21752 ) ;
  assign n21754 = n14636 ^ n9782 ^ n9359 ;
  assign n21755 = ( n3777 & n11917 ) | ( n3777 & n14541 ) | ( n11917 & n14541 ) ;
  assign n21756 = ( ~n21753 & n21754 ) | ( ~n21753 & n21755 ) | ( n21754 & n21755 ) ;
  assign n21757 = ( n661 & n11732 ) | ( n661 & ~n17524 ) | ( n11732 & ~n17524 ) ;
  assign n21758 = ( ~n4019 & n16152 ) | ( ~n4019 & n21757 ) | ( n16152 & n21757 ) ;
  assign n21759 = ( ~n7434 & n10960 ) | ( ~n7434 & n21758 ) | ( n10960 & n21758 ) ;
  assign n21760 = ( n2865 & ~n3818 ) | ( n2865 & n7240 ) | ( ~n3818 & n7240 ) ;
  assign n21761 = n21760 ^ n6922 ^ n3542 ;
  assign n21762 = n6658 ^ n4083 ^ n3656 ;
  assign n21763 = n15157 ^ n13139 ^ n6176 ;
  assign n21764 = ( n7813 & n21142 ) | ( n7813 & ~n21763 ) | ( n21142 & ~n21763 ) ;
  assign n21765 = ( n15128 & n21762 ) | ( n15128 & n21764 ) | ( n21762 & n21764 ) ;
  assign n21772 = ( n1959 & ~n2536 ) | ( n1959 & n10874 ) | ( ~n2536 & n10874 ) ;
  assign n21768 = ( ~n750 & n1891 ) | ( ~n750 & n10058 ) | ( n1891 & n10058 ) ;
  assign n21769 = ( n8079 & ~n8930 ) | ( n8079 & n21768 ) | ( ~n8930 & n21768 ) ;
  assign n21770 = n21769 ^ n15027 ^ n6345 ;
  assign n21766 = n20384 ^ n12428 ^ n2185 ;
  assign n21767 = n21766 ^ n7322 ^ n2124 ;
  assign n21771 = n21770 ^ n21767 ^ n21670 ;
  assign n21773 = n21772 ^ n21771 ^ n4314 ;
  assign n21774 = n8189 ^ n6253 ^ n2870 ;
  assign n21775 = n21774 ^ n14142 ^ n3378 ;
  assign n21776 = ( ~n1866 & n2861 ) | ( ~n1866 & n6125 ) | ( n2861 & n6125 ) ;
  assign n21777 = ( n1632 & n2095 ) | ( n1632 & n21776 ) | ( n2095 & n21776 ) ;
  assign n21778 = n16659 ^ n13088 ^ n8750 ;
  assign n21780 = n8429 ^ n4475 ^ x104 ;
  assign n21779 = n13871 ^ n12406 ^ n10731 ;
  assign n21781 = n21780 ^ n21779 ^ n20862 ;
  assign n21782 = n21781 ^ n20823 ^ n4269 ;
  assign n21783 = n8486 ^ n4617 ^ n2349 ;
  assign n21784 = n21783 ^ n16851 ^ n1656 ;
  assign n21785 = ( n5460 & ~n10648 ) | ( n5460 & n21784 ) | ( ~n10648 & n21784 ) ;
  assign n21786 = ( n344 & ~n760 ) | ( n344 & n10823 ) | ( ~n760 & n10823 ) ;
  assign n21787 = n10529 ^ n5297 ^ n4448 ;
  assign n21788 = ( n5857 & n7501 ) | ( n5857 & ~n21787 ) | ( n7501 & ~n21787 ) ;
  assign n21789 = n21788 ^ n7023 ^ n4401 ;
  assign n21790 = n15090 ^ n9082 ^ n3320 ;
  assign n21791 = n21790 ^ n8042 ^ n2276 ;
  assign n21792 = n21791 ^ n21609 ^ n446 ;
  assign n21794 = ( n687 & n2715 ) | ( n687 & ~n13015 ) | ( n2715 & ~n13015 ) ;
  assign n21793 = n8858 ^ n8118 ^ n4372 ;
  assign n21795 = n21794 ^ n21793 ^ n20781 ;
  assign n21796 = ( n2514 & n7321 ) | ( n2514 & ~n12100 ) | ( n7321 & ~n12100 ) ;
  assign n21797 = n8827 ^ n4607 ^ n3618 ;
  assign n21798 = n21797 ^ n20408 ^ n4165 ;
  assign n21799 = n21798 ^ n11310 ^ n1808 ;
  assign n21800 = ( n362 & n10979 ) | ( n362 & n13187 ) | ( n10979 & n13187 ) ;
  assign n21801 = ( n2227 & n21799 ) | ( n2227 & ~n21800 ) | ( n21799 & ~n21800 ) ;
  assign n21802 = ( n1767 & n2491 ) | ( n1767 & n21801 ) | ( n2491 & n21801 ) ;
  assign n21803 = ( ~n10310 & n21796 ) | ( ~n10310 & n21802 ) | ( n21796 & n21802 ) ;
  assign n21804 = n21803 ^ n19076 ^ n17792 ;
  assign n21805 = n17770 ^ n13807 ^ n4542 ;
  assign n21806 = ( ~n2200 & n2213 ) | ( ~n2200 & n7822 ) | ( n2213 & n7822 ) ;
  assign n21807 = ( n3836 & ~n20908 ) | ( n3836 & n21806 ) | ( ~n20908 & n21806 ) ;
  assign n21808 = n16810 ^ n12171 ^ n1511 ;
  assign n21809 = ( n5741 & ~n18623 ) | ( n5741 & n21808 ) | ( ~n18623 & n21808 ) ;
  assign n21811 = n8074 ^ n2848 ^ n2599 ;
  assign n21812 = ( n2056 & n3739 ) | ( n2056 & n21811 ) | ( n3739 & n21811 ) ;
  assign n21810 = n19276 ^ n18602 ^ n4800 ;
  assign n21813 = n21812 ^ n21810 ^ n18389 ;
  assign n21814 = n9145 ^ n4399 ^ n2453 ;
  assign n21815 = ( n3327 & n14643 ) | ( n3327 & n18285 ) | ( n14643 & n18285 ) ;
  assign n21816 = ( n945 & ~n21814 ) | ( n945 & n21815 ) | ( ~n21814 & n21815 ) ;
  assign n21817 = n6886 ^ n3275 ^ n1071 ;
  assign n21818 = n18229 ^ n16810 ^ n16733 ;
  assign n21819 = ( n7153 & n21387 ) | ( n7153 & ~n21818 ) | ( n21387 & ~n21818 ) ;
  assign n21820 = ( n5725 & n7187 ) | ( n5725 & ~n10350 ) | ( n7187 & ~n10350 ) ;
  assign n21821 = ( n3937 & n10623 ) | ( n3937 & ~n13120 ) | ( n10623 & ~n13120 ) ;
  assign n21822 = ( n2662 & n4786 ) | ( n2662 & n5774 ) | ( n4786 & n5774 ) ;
  assign n21823 = n21822 ^ n18412 ^ n11711 ;
  assign n21826 = ( n7516 & ~n16064 ) | ( n7516 & n17631 ) | ( ~n16064 & n17631 ) ;
  assign n21827 = ( n1858 & ~n6731 ) | ( n1858 & n21826 ) | ( ~n6731 & n21826 ) ;
  assign n21828 = n21827 ^ n16485 ^ n5266 ;
  assign n21824 = n14504 ^ n1858 ^ n382 ;
  assign n21825 = n21824 ^ n9655 ^ n3374 ;
  assign n21829 = n21828 ^ n21825 ^ n13261 ;
  assign n21830 = n21829 ^ n17199 ^ n11770 ;
  assign n21831 = n5270 ^ n4488 ^ n137 ;
  assign n21832 = n21831 ^ n18732 ^ n3655 ;
  assign n21833 = n21832 ^ n14329 ^ n2621 ;
  assign n21834 = n21833 ^ n12397 ^ n9698 ;
  assign n21835 = n11541 ^ n7273 ^ n890 ;
  assign n21836 = ( x96 & ~n7614 ) | ( x96 & n8361 ) | ( ~n7614 & n8361 ) ;
  assign n21837 = n21754 ^ n7215 ^ n2862 ;
  assign n21838 = n21824 ^ n14600 ^ n2918 ;
  assign n21839 = ( n8951 & ~n21837 ) | ( n8951 & n21838 ) | ( ~n21837 & n21838 ) ;
  assign n21840 = n21839 ^ n9961 ^ n3078 ;
  assign n21841 = ( ~n8192 & n14263 ) | ( ~n8192 & n21170 ) | ( n14263 & n21170 ) ;
  assign n21842 = n7696 ^ n3885 ^ n2315 ;
  assign n21843 = ( ~n732 & n961 ) | ( ~n732 & n21842 ) | ( n961 & n21842 ) ;
  assign n21844 = ( ~n10653 & n17262 ) | ( ~n10653 & n21843 ) | ( n17262 & n21843 ) ;
  assign n21845 = ( n3667 & n11439 ) | ( n3667 & n12468 ) | ( n11439 & n12468 ) ;
  assign n21846 = ( n2386 & n3568 ) | ( n2386 & n21845 ) | ( n3568 & n21845 ) ;
  assign n21847 = n21846 ^ n21463 ^ n4789 ;
  assign n21848 = ( n443 & n5854 ) | ( n443 & n7896 ) | ( n5854 & n7896 ) ;
  assign n21849 = ( n198 & ~n12294 ) | ( n198 & n21848 ) | ( ~n12294 & n21848 ) ;
  assign n21850 = n10685 ^ n8532 ^ n705 ;
  assign n21851 = ( ~n2323 & n18489 ) | ( ~n2323 & n21850 ) | ( n18489 & n21850 ) ;
  assign n21852 = ( n4555 & ~n6090 ) | ( n4555 & n17884 ) | ( ~n6090 & n17884 ) ;
  assign n21853 = ( n17213 & ~n21851 ) | ( n17213 & n21852 ) | ( ~n21851 & n21852 ) ;
  assign n21854 = ( n3879 & ~n7479 ) | ( n3879 & n15164 ) | ( ~n7479 & n15164 ) ;
  assign n21855 = n21854 ^ n17585 ^ n6627 ;
  assign n21856 = n21855 ^ n17965 ^ n5849 ;
  assign n21857 = ( n2001 & ~n13250 ) | ( n2001 & n21856 ) | ( ~n13250 & n21856 ) ;
  assign n21858 = ( n1884 & n5615 ) | ( n1884 & n14096 ) | ( n5615 & n14096 ) ;
  assign n21859 = n21742 ^ n18841 ^ n7093 ;
  assign n21860 = n21859 ^ n3630 ^ n846 ;
  assign n21861 = ( n10126 & n15004 ) | ( n10126 & n19678 ) | ( n15004 & n19678 ) ;
  assign n21862 = ( n2654 & ~n10908 ) | ( n2654 & n21649 ) | ( ~n10908 & n21649 ) ;
  assign n21869 = n20308 ^ n1419 ^ n605 ;
  assign n21870 = n16259 ^ n10570 ^ x62 ;
  assign n21871 = ( ~n519 & n21869 ) | ( ~n519 & n21870 ) | ( n21869 & n21870 ) ;
  assign n21865 = n10308 ^ n5386 ^ n4927 ;
  assign n21866 = n21865 ^ n9816 ^ n8207 ;
  assign n21867 = ( n7531 & ~n8802 ) | ( n7531 & n21866 ) | ( ~n8802 & n21866 ) ;
  assign n21863 = ( n3717 & n12165 ) | ( n3717 & ~n13258 ) | ( n12165 & ~n13258 ) ;
  assign n21864 = n21863 ^ n20098 ^ n16047 ;
  assign n21868 = n21867 ^ n21864 ^ n2744 ;
  assign n21872 = n21871 ^ n21868 ^ n11664 ;
  assign n21873 = n11032 ^ n11002 ^ n4180 ;
  assign n21874 = ( ~n7569 & n11103 ) | ( ~n7569 & n21873 ) | ( n11103 & n21873 ) ;
  assign n21876 = ( n1579 & ~n5052 ) | ( n1579 & n10336 ) | ( ~n5052 & n10336 ) ;
  assign n21875 = ( n2328 & n8714 ) | ( n2328 & n10788 ) | ( n8714 & n10788 ) ;
  assign n21877 = n21876 ^ n21875 ^ n11866 ;
  assign n21879 = ( x15 & n1374 ) | ( x15 & ~n15261 ) | ( n1374 & ~n15261 ) ;
  assign n21878 = n12907 ^ n9435 ^ n3253 ;
  assign n21880 = n21879 ^ n21878 ^ n9513 ;
  assign n21881 = n21880 ^ n17411 ^ n12910 ;
  assign n21882 = ( n4151 & n4960 ) | ( n4151 & n11286 ) | ( n4960 & n11286 ) ;
  assign n21883 = ( n1020 & n2666 ) | ( n1020 & ~n21882 ) | ( n2666 & ~n21882 ) ;
  assign n21884 = ( n6422 & n12040 ) | ( n6422 & n19260 ) | ( n12040 & n19260 ) ;
  assign n21885 = ( n171 & n11248 ) | ( n171 & n12620 ) | ( n11248 & n12620 ) ;
  assign n21886 = ( n14793 & n21884 ) | ( n14793 & ~n21885 ) | ( n21884 & ~n21885 ) ;
  assign n21887 = ( n17504 & ~n21883 ) | ( n17504 & n21886 ) | ( ~n21883 & n21886 ) ;
  assign n21890 = ( ~n3652 & n4241 ) | ( ~n3652 & n6540 ) | ( n4241 & n6540 ) ;
  assign n21891 = ( n6943 & n9806 ) | ( n6943 & ~n21890 ) | ( n9806 & ~n21890 ) ;
  assign n21888 = n14086 ^ n3169 ^ n969 ;
  assign n21889 = ( ~n6113 & n14164 ) | ( ~n6113 & n21888 ) | ( n14164 & n21888 ) ;
  assign n21892 = n21891 ^ n21889 ^ n16626 ;
  assign n21893 = n21892 ^ n18268 ^ n11240 ;
  assign n21894 = ( n3493 & ~n8796 ) | ( n3493 & n16495 ) | ( ~n8796 & n16495 ) ;
  assign n21895 = ( n1479 & n10106 ) | ( n1479 & n12862 ) | ( n10106 & n12862 ) ;
  assign n21896 = n19297 ^ n8376 ^ n5603 ;
  assign n21897 = ( n761 & n8537 ) | ( n761 & ~n9251 ) | ( n8537 & ~n9251 ) ;
  assign n21898 = ( n21895 & ~n21896 ) | ( n21895 & n21897 ) | ( ~n21896 & n21897 ) ;
  assign n21899 = n18236 ^ n12553 ^ n7531 ;
  assign n21900 = ( n5117 & n7686 ) | ( n5117 & n21899 ) | ( n7686 & n21899 ) ;
  assign n21901 = n21879 ^ n6287 ^ n1784 ;
  assign n21902 = ( ~n15650 & n21818 ) | ( ~n15650 & n21901 ) | ( n21818 & n21901 ) ;
  assign n21903 = ( ~n9080 & n9519 ) | ( ~n9080 & n21902 ) | ( n9519 & n21902 ) ;
  assign n21904 = ( n2313 & ~n4326 ) | ( n2313 & n15174 ) | ( ~n4326 & n15174 ) ;
  assign n21905 = ( n2127 & n3037 ) | ( n2127 & ~n21904 ) | ( n3037 & ~n21904 ) ;
  assign n21906 = n6181 ^ n5078 ^ n979 ;
  assign n21907 = ( n2560 & n21905 ) | ( n2560 & n21906 ) | ( n21905 & n21906 ) ;
  assign n21908 = n8727 ^ n7551 ^ n611 ;
  assign n21909 = n20964 ^ n16700 ^ n14688 ;
  assign n21910 = ( x124 & n14081 ) | ( x124 & ~n16939 ) | ( n14081 & ~n16939 ) ;
  assign n21911 = n21910 ^ n17434 ^ n4312 ;
  assign n21912 = ( n3635 & n18609 ) | ( n3635 & ~n21911 ) | ( n18609 & ~n21911 ) ;
  assign n21913 = ( n1164 & ~n11449 ) | ( n1164 & n21912 ) | ( ~n11449 & n21912 ) ;
  assign n21914 = n20594 ^ n19123 ^ n14089 ;
  assign n21915 = ( n9458 & n14771 ) | ( n9458 & n21914 ) | ( n14771 & n21914 ) ;
  assign n21916 = ( n1427 & ~n6406 ) | ( n1427 & n16053 ) | ( ~n6406 & n16053 ) ;
  assign n21918 = ( n1614 & n2881 ) | ( n1614 & n7832 ) | ( n2881 & n7832 ) ;
  assign n21917 = ( ~n11034 & n12190 ) | ( ~n11034 & n14414 ) | ( n12190 & n14414 ) ;
  assign n21919 = n21918 ^ n21917 ^ n3648 ;
  assign n21920 = ( ~n1734 & n2330 ) | ( ~n1734 & n3181 ) | ( n2330 & n3181 ) ;
  assign n21921 = n19373 ^ n19353 ^ n3661 ;
  assign n21922 = ( n2509 & n4470 ) | ( n2509 & ~n5818 ) | ( n4470 & ~n5818 ) ;
  assign n21923 = n21922 ^ n8375 ^ n7220 ;
  assign n21924 = ( n18476 & ~n21921 ) | ( n18476 & n21923 ) | ( ~n21921 & n21923 ) ;
  assign n21925 = n12929 ^ n2634 ^ x124 ;
  assign n21926 = ( n7674 & n21924 ) | ( n7674 & ~n21925 ) | ( n21924 & ~n21925 ) ;
  assign n21927 = ( n835 & n9656 ) | ( n835 & n12821 ) | ( n9656 & n12821 ) ;
  assign n21929 = ( n12291 & ~n12738 ) | ( n12291 & n19296 ) | ( ~n12738 & n19296 ) ;
  assign n21930 = n21929 ^ n16787 ^ n12068 ;
  assign n21928 = n15890 ^ n7061 ^ n4858 ;
  assign n21931 = n21930 ^ n21928 ^ n4526 ;
  assign n21932 = n7183 ^ n4921 ^ n4298 ;
  assign n21933 = ( n2644 & ~n4410 ) | ( n2644 & n7801 ) | ( ~n4410 & n7801 ) ;
  assign n21934 = ( ~n6417 & n13871 ) | ( ~n6417 & n21933 ) | ( n13871 & n21933 ) ;
  assign n21935 = n16226 ^ n14671 ^ n9415 ;
  assign n21936 = ( n21932 & n21934 ) | ( n21932 & n21935 ) | ( n21934 & n21935 ) ;
  assign n21937 = n21936 ^ n11062 ^ n10781 ;
  assign n21938 = n19669 ^ n16780 ^ n1954 ;
  assign n21939 = n21938 ^ n20825 ^ n8919 ;
  assign n21940 = ( n11380 & n17586 ) | ( n11380 & n20469 ) | ( n17586 & n20469 ) ;
  assign n21941 = ( n1090 & n4515 ) | ( n1090 & n8419 ) | ( n4515 & n8419 ) ;
  assign n21942 = ( n11082 & n17838 ) | ( n11082 & ~n20708 ) | ( n17838 & ~n20708 ) ;
  assign n21943 = ( ~n1137 & n17228 ) | ( ~n1137 & n21942 ) | ( n17228 & n21942 ) ;
  assign n21944 = ( ~n18844 & n21941 ) | ( ~n18844 & n21943 ) | ( n21941 & n21943 ) ;
  assign n21945 = n21944 ^ n18391 ^ n7431 ;
  assign n21946 = n9198 ^ n4219 ^ n1832 ;
  assign n21947 = n20723 ^ n14905 ^ n811 ;
  assign n21948 = n11639 ^ n8900 ^ n3492 ;
  assign n21949 = n21948 ^ n21110 ^ n300 ;
  assign n21950 = ( n8538 & ~n15143 ) | ( n8538 & n21949 ) | ( ~n15143 & n21949 ) ;
  assign n21957 = n9636 ^ n4019 ^ n3850 ;
  assign n21958 = n5590 ^ n3314 ^ n1639 ;
  assign n21959 = ( n4171 & n21957 ) | ( n4171 & n21958 ) | ( n21957 & n21958 ) ;
  assign n21956 = ( n6263 & n15418 ) | ( n6263 & n15480 ) | ( n15418 & n15480 ) ;
  assign n21954 = ( n6584 & n10909 ) | ( n6584 & ~n17276 ) | ( n10909 & ~n17276 ) ;
  assign n21951 = ( n2060 & n5465 ) | ( n2060 & n8584 ) | ( n5465 & n8584 ) ;
  assign n21952 = ( n4596 & ~n6963 ) | ( n4596 & n21951 ) | ( ~n6963 & n21951 ) ;
  assign n21953 = n21952 ^ n20693 ^ n13155 ;
  assign n21955 = n21954 ^ n21953 ^ n8836 ;
  assign n21960 = n21959 ^ n21956 ^ n21955 ;
  assign n21961 = ( n1025 & n4351 ) | ( n1025 & n14566 ) | ( n4351 & n14566 ) ;
  assign n21962 = ( ~n1865 & n8775 ) | ( ~n1865 & n12214 ) | ( n8775 & n12214 ) ;
  assign n21963 = n20239 ^ n15548 ^ n10868 ;
  assign n21964 = n21963 ^ n14333 ^ n9017 ;
  assign n21965 = ( n10941 & n21697 ) | ( n10941 & ~n21964 ) | ( n21697 & ~n21964 ) ;
  assign n21966 = n21965 ^ n7278 ^ n2112 ;
  assign n21967 = ( n3663 & n8727 ) | ( n3663 & n20832 ) | ( n8727 & n20832 ) ;
  assign n21968 = ( n5783 & ~n21966 ) | ( n5783 & n21967 ) | ( ~n21966 & n21967 ) ;
  assign n21969 = ( ~n15579 & n16286 ) | ( ~n15579 & n18720 ) | ( n16286 & n18720 ) ;
  assign n21970 = ( n6231 & n9947 ) | ( n6231 & ~n21969 ) | ( n9947 & ~n21969 ) ;
  assign n21971 = ( ~n6953 & n8227 ) | ( ~n6953 & n11178 ) | ( n8227 & n11178 ) ;
  assign n21972 = n21971 ^ n9942 ^ n5692 ;
  assign n21974 = n14325 ^ n8185 ^ n3945 ;
  assign n21973 = ( n5056 & n5449 ) | ( n5056 & ~n5999 ) | ( n5449 & ~n5999 ) ;
  assign n21975 = n21974 ^ n21973 ^ n2436 ;
  assign n21976 = ( ~n9731 & n10223 ) | ( ~n9731 & n21175 ) | ( n10223 & n21175 ) ;
  assign n21977 = ( n8879 & n17194 ) | ( n8879 & ~n21976 ) | ( n17194 & ~n21976 ) ;
  assign n21978 = ( n8415 & n8473 ) | ( n8415 & n10396 ) | ( n8473 & n10396 ) ;
  assign n21979 = n21978 ^ n18264 ^ n7867 ;
  assign n21980 = n14707 ^ n8244 ^ n4842 ;
  assign n21981 = n6065 ^ n2413 ^ n986 ;
  assign n21982 = n21981 ^ n17987 ^ n7181 ;
  assign n21983 = ( n3668 & n5506 ) | ( n3668 & n21982 ) | ( n5506 & n21982 ) ;
  assign n21984 = ( ~n15028 & n21980 ) | ( ~n15028 & n21983 ) | ( n21980 & n21983 ) ;
  assign n21985 = ( n10438 & n10890 ) | ( n10438 & ~n20448 ) | ( n10890 & ~n20448 ) ;
  assign n21986 = ( n8635 & ~n15283 ) | ( n8635 & n21985 ) | ( ~n15283 & n21985 ) ;
  assign n21987 = ( n624 & n8717 ) | ( n624 & ~n14374 ) | ( n8717 & ~n14374 ) ;
  assign n21988 = ( n639 & ~n6210 ) | ( n639 & n21987 ) | ( ~n6210 & n21987 ) ;
  assign n21989 = n5633 ^ n2800 ^ x103 ;
  assign n21990 = ( n1418 & n13867 ) | ( n1418 & ~n20192 ) | ( n13867 & ~n20192 ) ;
  assign n21991 = n14648 ^ n9430 ^ n788 ;
  assign n21992 = n15717 ^ n8576 ^ n2617 ;
  assign n21993 = n12491 ^ n6919 ^ n2349 ;
  assign n21994 = ( n6100 & n7597 ) | ( n6100 & n21993 ) | ( n7597 & n21993 ) ;
  assign n21995 = n9316 ^ n9045 ^ n6881 ;
  assign n21996 = ( n2089 & ~n9795 ) | ( n2089 & n21995 ) | ( ~n9795 & n21995 ) ;
  assign n21997 = ( n2201 & n21994 ) | ( n2201 & n21996 ) | ( n21994 & n21996 ) ;
  assign n21998 = ( x48 & n3262 ) | ( x48 & ~n7131 ) | ( n3262 & ~n7131 ) ;
  assign n21999 = n17186 ^ n8004 ^ n3981 ;
  assign n22000 = ( n9144 & n11193 ) | ( n9144 & ~n15909 ) | ( n11193 & ~n15909 ) ;
  assign n22001 = ( n3117 & ~n3813 ) | ( n3117 & n9509 ) | ( ~n3813 & n9509 ) ;
  assign n22002 = ( n15142 & n16969 ) | ( n15142 & ~n22001 ) | ( n16969 & ~n22001 ) ;
  assign n22003 = ( ~n2651 & n13596 ) | ( ~n2651 & n22002 ) | ( n13596 & n22002 ) ;
  assign n22004 = n8008 ^ n3036 ^ n2719 ;
  assign n22005 = ( n699 & n8210 ) | ( n699 & n22004 ) | ( n8210 & n22004 ) ;
  assign n22006 = ( n575 & ~n7472 ) | ( n575 & n22005 ) | ( ~n7472 & n22005 ) ;
  assign n22007 = ( n186 & n18189 ) | ( n186 & n22006 ) | ( n18189 & n22006 ) ;
  assign n22008 = ( n4564 & n11006 ) | ( n4564 & n12241 ) | ( n11006 & n12241 ) ;
  assign n22009 = ( ~n5827 & n10787 ) | ( ~n5827 & n17627 ) | ( n10787 & n17627 ) ;
  assign n22010 = ( n7717 & n11988 ) | ( n7717 & ~n20996 ) | ( n11988 & ~n20996 ) ;
  assign n22011 = ( n8918 & n9198 ) | ( n8918 & ~n22010 ) | ( n9198 & ~n22010 ) ;
  assign n22012 = n21703 ^ n7814 ^ n5208 ;
  assign n22013 = n12929 ^ n10450 ^ n1997 ;
  assign n22014 = ( n2186 & n4747 ) | ( n2186 & ~n7172 ) | ( n4747 & ~n7172 ) ;
  assign n22015 = ( n4206 & ~n6830 ) | ( n4206 & n9558 ) | ( ~n6830 & n9558 ) ;
  assign n22016 = ( n22013 & ~n22014 ) | ( n22013 & n22015 ) | ( ~n22014 & n22015 ) ;
  assign n22018 = ( n1152 & n5233 ) | ( n1152 & ~n19867 ) | ( n5233 & ~n19867 ) ;
  assign n22019 = n22018 ^ n14849 ^ n5874 ;
  assign n22017 = n18958 ^ n7216 ^ n6519 ;
  assign n22020 = n22019 ^ n22017 ^ n15254 ;
  assign n22026 = n20727 ^ n10073 ^ n718 ;
  assign n22021 = n20575 ^ n12151 ^ n572 ;
  assign n22022 = n16502 ^ n6581 ^ n3704 ;
  assign n22023 = n22022 ^ n18754 ^ n13717 ;
  assign n22024 = ( n4488 & n22021 ) | ( n4488 & n22023 ) | ( n22021 & n22023 ) ;
  assign n22025 = ( n8870 & n17633 ) | ( n8870 & ~n22024 ) | ( n17633 & ~n22024 ) ;
  assign n22027 = n22026 ^ n22025 ^ n13511 ;
  assign n22031 = n7526 ^ n3970 ^ n2513 ;
  assign n22032 = n22031 ^ n12833 ^ n2224 ;
  assign n22033 = n8643 ^ n4060 ^ n1140 ;
  assign n22034 = n22033 ^ n18217 ^ n1774 ;
  assign n22035 = ( n312 & n14849 ) | ( n312 & n22034 ) | ( n14849 & n22034 ) ;
  assign n22036 = ( n14070 & ~n22032 ) | ( n14070 & n22035 ) | ( ~n22032 & n22035 ) ;
  assign n22029 = ( n947 & n1268 ) | ( n947 & ~n10282 ) | ( n1268 & ~n10282 ) ;
  assign n22030 = ( n3485 & n20104 ) | ( n3485 & n22029 ) | ( n20104 & n22029 ) ;
  assign n22028 = ( n1738 & ~n16772 ) | ( n1738 & n18977 ) | ( ~n16772 & n18977 ) ;
  assign n22037 = n22036 ^ n22030 ^ n22028 ;
  assign n22038 = ( n4323 & n4541 ) | ( n4323 & ~n5174 ) | ( n4541 & ~n5174 ) ;
  assign n22039 = n22038 ^ n17758 ^ n9599 ;
  assign n22040 = n22039 ^ n19128 ^ n511 ;
  assign n22041 = n22040 ^ n10391 ^ n10087 ;
  assign n22042 = n22041 ^ n18492 ^ n13026 ;
  assign n22043 = n14075 ^ n7862 ^ n6174 ;
  assign n22044 = n9115 ^ n1107 ^ n798 ;
  assign n22045 = ( n7022 & n8604 ) | ( n7022 & n22044 ) | ( n8604 & n22044 ) ;
  assign n22046 = ( n1915 & n22043 ) | ( n1915 & ~n22045 ) | ( n22043 & ~n22045 ) ;
  assign n22047 = n22046 ^ n9131 ^ n2920 ;
  assign n22052 = ( n8277 & n12289 ) | ( n8277 & n16916 ) | ( n12289 & n16916 ) ;
  assign n22048 = n7624 ^ n6737 ^ n3289 ;
  assign n22049 = ( ~n6339 & n15680 ) | ( ~n6339 & n22048 ) | ( n15680 & n22048 ) ;
  assign n22050 = n22049 ^ n8312 ^ n1082 ;
  assign n22051 = n22050 ^ n6034 ^ n6021 ;
  assign n22053 = n22052 ^ n22051 ^ n12810 ;
  assign n22054 = ( ~n11910 & n21980 ) | ( ~n11910 & n22053 ) | ( n21980 & n22053 ) ;
  assign n22056 = ( n6751 & n14659 ) | ( n6751 & n19226 ) | ( n14659 & n19226 ) ;
  assign n22057 = ( n4927 & n7516 ) | ( n4927 & n22056 ) | ( n7516 & n22056 ) ;
  assign n22055 = ( ~n1059 & n8039 ) | ( ~n1059 & n14423 ) | ( n8039 & n14423 ) ;
  assign n22058 = n22057 ^ n22055 ^ n18985 ;
  assign n22059 = ( n1942 & ~n14108 ) | ( n1942 & n21298 ) | ( ~n14108 & n21298 ) ;
  assign n22060 = ( n10608 & n15441 ) | ( n10608 & ~n15951 ) | ( n15441 & ~n15951 ) ;
  assign n22061 = ( n3936 & ~n8060 ) | ( n3936 & n22060 ) | ( ~n8060 & n22060 ) ;
  assign n22063 = ( ~n665 & n16361 ) | ( ~n665 & n19447 ) | ( n16361 & n19447 ) ;
  assign n22062 = ( n669 & n10959 ) | ( n669 & ~n18655 ) | ( n10959 & ~n18655 ) ;
  assign n22064 = n22063 ^ n22062 ^ n1126 ;
  assign n22065 = n22064 ^ n20478 ^ n9473 ;
  assign n22066 = ( n7995 & n12507 ) | ( n7995 & ~n16466 ) | ( n12507 & ~n16466 ) ;
  assign n22067 = ( ~n5218 & n7314 ) | ( ~n5218 & n22066 ) | ( n7314 & n22066 ) ;
  assign n22068 = n16999 ^ n11124 ^ n6501 ;
  assign n22069 = ( n13541 & n19922 ) | ( n13541 & ~n22068 ) | ( n19922 & ~n22068 ) ;
  assign n22070 = n13809 ^ n8286 ^ n6355 ;
  assign n22071 = ( n4303 & n22069 ) | ( n4303 & ~n22070 ) | ( n22069 & ~n22070 ) ;
  assign n22072 = ( n16814 & ~n19260 ) | ( n16814 & n22071 ) | ( ~n19260 & n22071 ) ;
  assign n22073 = n11040 ^ n2706 ^ n1331 ;
  assign n22074 = n22073 ^ n13194 ^ n5802 ;
  assign n22075 = ( n5287 & n10629 ) | ( n5287 & ~n13277 ) | ( n10629 & ~n13277 ) ;
  assign n22076 = n22075 ^ n6950 ^ n2906 ;
  assign n22077 = n22076 ^ n14282 ^ n2243 ;
  assign n22081 = n10618 ^ n7779 ^ n5107 ;
  assign n22080 = ( n1617 & n7499 ) | ( n1617 & ~n18011 ) | ( n7499 & ~n18011 ) ;
  assign n22078 = ( n353 & ~n3878 ) | ( n353 & n7264 ) | ( ~n3878 & n7264 ) ;
  assign n22079 = ( n3459 & n13376 ) | ( n3459 & ~n22078 ) | ( n13376 & ~n22078 ) ;
  assign n22082 = n22081 ^ n22080 ^ n22079 ;
  assign n22083 = n19258 ^ n12330 ^ n10377 ;
  assign n22084 = ( n137 & ~n3585 ) | ( n137 & n22083 ) | ( ~n3585 & n22083 ) ;
  assign n22085 = ( n707 & n6754 ) | ( n707 & n22084 ) | ( n6754 & n22084 ) ;
  assign n22086 = n10256 ^ n8177 ^ n4582 ;
  assign n22087 = n10893 ^ n9300 ^ n6341 ;
  assign n22088 = ( n1421 & ~n1824 ) | ( n1421 & n8649 ) | ( ~n1824 & n8649 ) ;
  assign n22089 = ( n2437 & ~n22087 ) | ( n2437 & n22088 ) | ( ~n22087 & n22088 ) ;
  assign n22090 = n22089 ^ n7232 ^ n3228 ;
  assign n22091 = ( n4292 & n22086 ) | ( n4292 & n22090 ) | ( n22086 & n22090 ) ;
  assign n22092 = n21294 ^ n13660 ^ n8997 ;
  assign n22093 = n22092 ^ n18595 ^ n12642 ;
  assign n22094 = ( n3850 & n10897 ) | ( n3850 & ~n22093 ) | ( n10897 & ~n22093 ) ;
  assign n22095 = ( n2284 & n4428 ) | ( n2284 & ~n22094 ) | ( n4428 & ~n22094 ) ;
  assign n22096 = n22095 ^ n14997 ^ n4886 ;
  assign n22097 = n6914 ^ n4172 ^ n4123 ;
  assign n22098 = ( n7913 & ~n21656 ) | ( n7913 & n22097 ) | ( ~n21656 & n22097 ) ;
  assign n22099 = n22098 ^ n10588 ^ n4596 ;
  assign n22100 = ( n10897 & n11906 ) | ( n10897 & n22099 ) | ( n11906 & n22099 ) ;
  assign n22101 = n3734 ^ n2420 ^ n522 ;
  assign n22102 = n22101 ^ n14534 ^ n4406 ;
  assign n22104 = n15431 ^ n1154 ^ n892 ;
  assign n22105 = n22104 ^ n4938 ^ n4102 ;
  assign n22106 = n9048 ^ n6098 ^ n1992 ;
  assign n22107 = ( n4589 & ~n9184 ) | ( n4589 & n22106 ) | ( ~n9184 & n22106 ) ;
  assign n22108 = n19293 ^ n12601 ^ n2289 ;
  assign n22109 = ( n2563 & n14729 ) | ( n2563 & ~n22108 ) | ( n14729 & ~n22108 ) ;
  assign n22110 = n22109 ^ n4387 ^ n3094 ;
  assign n22111 = ( ~n2508 & n17383 ) | ( ~n2508 & n22110 ) | ( n17383 & n22110 ) ;
  assign n22112 = n22111 ^ n10694 ^ n5102 ;
  assign n22113 = ( n9020 & ~n22107 ) | ( n9020 & n22112 ) | ( ~n22107 & n22112 ) ;
  assign n22114 = ( n1078 & n22105 ) | ( n1078 & ~n22113 ) | ( n22105 & ~n22113 ) ;
  assign n22103 = n13780 ^ n1206 ^ n824 ;
  assign n22115 = n22114 ^ n22103 ^ n14119 ;
  assign n22116 = ( ~n20242 & n22102 ) | ( ~n20242 & n22115 ) | ( n22102 & n22115 ) ;
  assign n22118 = ( n3492 & ~n7420 ) | ( n3492 & n13882 ) | ( ~n7420 & n13882 ) ;
  assign n22119 = n22118 ^ n14471 ^ n2826 ;
  assign n22117 = n11800 ^ n2189 ^ n656 ;
  assign n22120 = n22119 ^ n22117 ^ n16110 ;
  assign n22121 = ( ~n506 & n4129 ) | ( ~n506 & n7178 ) | ( n4129 & n7178 ) ;
  assign n22122 = ( n2512 & ~n7397 ) | ( n2512 & n11380 ) | ( ~n7397 & n11380 ) ;
  assign n22123 = n9174 ^ n7775 ^ n7059 ;
  assign n22124 = n5230 ^ n4166 ^ n1153 ;
  assign n22125 = ( n3235 & n8144 ) | ( n3235 & n22124 ) | ( n8144 & n22124 ) ;
  assign n22126 = ( n7114 & ~n22123 ) | ( n7114 & n22125 ) | ( ~n22123 & n22125 ) ;
  assign n22127 = ( n4888 & ~n9463 ) | ( n4888 & n22126 ) | ( ~n9463 & n22126 ) ;
  assign n22128 = n15424 ^ n13635 ^ n593 ;
  assign n22129 = n22128 ^ n14771 ^ n13383 ;
  assign n22130 = n16665 ^ n12356 ^ n347 ;
  assign n22131 = ( ~n4437 & n10596 ) | ( ~n4437 & n13422 ) | ( n10596 & n13422 ) ;
  assign n22132 = n10742 ^ n6971 ^ n1381 ;
  assign n22133 = n22132 ^ n6331 ^ n1831 ;
  assign n22134 = ( n7336 & n16885 ) | ( n7336 & n22133 ) | ( n16885 & n22133 ) ;
  assign n22135 = ( n1432 & n22131 ) | ( n1432 & ~n22134 ) | ( n22131 & ~n22134 ) ;
  assign n22136 = n16540 ^ n12094 ^ n7421 ;
  assign n22141 = ( n2601 & n7391 ) | ( n2601 & n16204 ) | ( n7391 & n16204 ) ;
  assign n22137 = ( ~n3522 & n11491 ) | ( ~n3522 & n15897 ) | ( n11491 & n15897 ) ;
  assign n22138 = ( n10698 & ~n11612 ) | ( n10698 & n22137 ) | ( ~n11612 & n22137 ) ;
  assign n22139 = n22138 ^ n8484 ^ n4711 ;
  assign n22140 = ( n1536 & n20419 ) | ( n1536 & ~n22139 ) | ( n20419 & ~n22139 ) ;
  assign n22142 = n22141 ^ n22140 ^ n7766 ;
  assign n22143 = n9054 ^ n3532 ^ n1289 ;
  assign n22144 = n21911 ^ n4490 ^ x81 ;
  assign n22145 = n14234 ^ n11356 ^ n887 ;
  assign n22146 = n14274 ^ n12767 ^ n10931 ;
  assign n22147 = n19213 ^ n18879 ^ n13867 ;
  assign n22148 = n12915 ^ n7189 ^ n1639 ;
  assign n22149 = ( n2632 & n4789 ) | ( n2632 & ~n22148 ) | ( n4789 & ~n22148 ) ;
  assign n22150 = ( ~n5421 & n6373 ) | ( ~n5421 & n14541 ) | ( n6373 & n14541 ) ;
  assign n22151 = n20032 ^ n12509 ^ n2614 ;
  assign n22152 = ( n946 & n15378 ) | ( n946 & ~n22151 ) | ( n15378 & ~n22151 ) ;
  assign n22153 = ( n3568 & n22150 ) | ( n3568 & n22152 ) | ( n22150 & n22152 ) ;
  assign n22154 = n18829 ^ n16044 ^ n6066 ;
  assign n22155 = ( n17522 & n17535 ) | ( n17522 & n22154 ) | ( n17535 & n22154 ) ;
  assign n22156 = ( n3483 & n5197 ) | ( n3483 & n7357 ) | ( n5197 & n7357 ) ;
  assign n22157 = ( ~n3025 & n10825 ) | ( ~n3025 & n18943 ) | ( n10825 & n18943 ) ;
  assign n22158 = n22157 ^ n4011 ^ n3726 ;
  assign n22159 = n13475 ^ n10713 ^ n6575 ;
  assign n22160 = ( n5206 & ~n12571 ) | ( n5206 & n22159 ) | ( ~n12571 & n22159 ) ;
  assign n22161 = n22160 ^ n11777 ^ n8798 ;
  assign n22162 = ( n5455 & n7407 ) | ( n5455 & ~n22161 ) | ( n7407 & ~n22161 ) ;
  assign n22163 = n20163 ^ n13606 ^ n2553 ;
  assign n22164 = n4136 ^ n3021 ^ n1223 ;
  assign n22165 = ( ~n21427 & n22163 ) | ( ~n21427 & n22164 ) | ( n22163 & n22164 ) ;
  assign n22166 = ( n15791 & n16606 ) | ( n15791 & ~n21483 ) | ( n16606 & ~n21483 ) ;
  assign n22167 = n16485 ^ n1883 ^ n1195 ;
  assign n22168 = ( n877 & n2951 ) | ( n877 & ~n22167 ) | ( n2951 & ~n22167 ) ;
  assign n22169 = n22168 ^ n3656 ^ n1387 ;
  assign n22170 = n22169 ^ n13634 ^ n3451 ;
  assign n22171 = n12248 ^ n3918 ^ n3844 ;
  assign n22172 = ( n11303 & n18264 ) | ( n11303 & n22171 ) | ( n18264 & n22171 ) ;
  assign n22173 = ( n1079 & n11845 ) | ( n1079 & n16816 ) | ( n11845 & n16816 ) ;
  assign n22174 = n22173 ^ n21494 ^ n21361 ;
  assign n22175 = ( n7362 & n8542 ) | ( n7362 & ~n11407 ) | ( n8542 & ~n11407 ) ;
  assign n22176 = ( n1778 & n14583 ) | ( n1778 & ~n22175 ) | ( n14583 & ~n22175 ) ;
  assign n22177 = ( n2093 & n9169 ) | ( n2093 & ~n22176 ) | ( n9169 & ~n22176 ) ;
  assign n22178 = ( n3074 & n13256 ) | ( n3074 & n22076 ) | ( n13256 & n22076 ) ;
  assign n22179 = ( n4454 & n4743 ) | ( n4454 & ~n7251 ) | ( n4743 & ~n7251 ) ;
  assign n22180 = ( n11130 & n12902 ) | ( n11130 & ~n22179 ) | ( n12902 & ~n22179 ) ;
  assign n22181 = ( ~n8829 & n9602 ) | ( ~n8829 & n16854 ) | ( n9602 & n16854 ) ;
  assign n22182 = n16433 ^ n4611 ^ n1615 ;
  assign n22183 = ( n1954 & n7048 ) | ( n1954 & n21380 ) | ( n7048 & n21380 ) ;
  assign n22184 = ( n627 & ~n6594 ) | ( n627 & n22183 ) | ( ~n6594 & n22183 ) ;
  assign n22185 = n16635 ^ n16206 ^ n5276 ;
  assign n22186 = ( n14288 & ~n16464 ) | ( n14288 & n22185 ) | ( ~n16464 & n22185 ) ;
  assign n22187 = ( n7816 & n14280 ) | ( n7816 & n22186 ) | ( n14280 & n22186 ) ;
  assign n22188 = ( n9780 & n13444 ) | ( n9780 & n22187 ) | ( n13444 & n22187 ) ;
  assign n22194 = n18557 ^ n15119 ^ n9420 ;
  assign n22195 = ( n3030 & ~n10801 ) | ( n3030 & n22194 ) | ( ~n10801 & n22194 ) ;
  assign n22191 = n10579 ^ n3401 ^ x24 ;
  assign n22192 = ( n484 & ~n7922 ) | ( n484 & n22191 ) | ( ~n7922 & n22191 ) ;
  assign n22190 = n20877 ^ n7283 ^ n1808 ;
  assign n22189 = n12507 ^ n5072 ^ n3286 ;
  assign n22193 = n22192 ^ n22190 ^ n22189 ;
  assign n22196 = n22195 ^ n22193 ^ n14735 ;
  assign n22205 = n15974 ^ n15326 ^ n6839 ;
  assign n22202 = ( n960 & n4481 ) | ( n960 & ~n16115 ) | ( n4481 & ~n16115 ) ;
  assign n22203 = ( n2278 & ~n8252 ) | ( n2278 & n22202 ) | ( ~n8252 & n22202 ) ;
  assign n22204 = n22203 ^ n19966 ^ n17955 ;
  assign n22206 = n22205 ^ n22204 ^ n11334 ;
  assign n22199 = n11129 ^ n1769 ^ n792 ;
  assign n22200 = ( n1827 & ~n16216 ) | ( n1827 & n22199 ) | ( ~n16216 & n22199 ) ;
  assign n22197 = n13051 ^ n8094 ^ n1469 ;
  assign n22198 = ( n2571 & n6426 ) | ( n2571 & n22197 ) | ( n6426 & n22197 ) ;
  assign n22201 = n22200 ^ n22198 ^ n15416 ;
  assign n22207 = n22206 ^ n22201 ^ n6826 ;
  assign n22208 = n9220 ^ n7897 ^ n6208 ;
  assign n22209 = n22208 ^ n12388 ^ n4966 ;
  assign n22210 = n22209 ^ n4895 ^ n2705 ;
  assign n22211 = ( ~n716 & n2509 ) | ( ~n716 & n19324 ) | ( n2509 & n19324 ) ;
  assign n22212 = ( n10190 & n18863 ) | ( n10190 & n22211 ) | ( n18863 & n22211 ) ;
  assign n22213 = ( n8032 & ~n10687 ) | ( n8032 & n12187 ) | ( ~n10687 & n12187 ) ;
  assign n22214 = n22213 ^ n4833 ^ n2371 ;
  assign n22217 = n19361 ^ n13352 ^ n12690 ;
  assign n22215 = n6406 ^ n3884 ^ n3161 ;
  assign n22216 = ( n1877 & ~n21604 ) | ( n1877 & n22215 ) | ( ~n21604 & n22215 ) ;
  assign n22218 = n22217 ^ n22216 ^ x66 ;
  assign n22219 = ( n8371 & n9262 ) | ( n8371 & n21212 ) | ( n9262 & n21212 ) ;
  assign n22220 = n22219 ^ n9508 ^ n7966 ;
  assign n22221 = n22220 ^ n13367 ^ n6971 ;
  assign n22222 = n9684 ^ n5587 ^ n5251 ;
  assign n22223 = ( n1956 & n6759 ) | ( n1956 & ~n8169 ) | ( n6759 & ~n8169 ) ;
  assign n22224 = ( ~n5059 & n5408 ) | ( ~n5059 & n12541 ) | ( n5408 & n12541 ) ;
  assign n22225 = ( n8225 & n9354 ) | ( n8225 & n22224 ) | ( n9354 & n22224 ) ;
  assign n22226 = ( n1343 & n22223 ) | ( n1343 & ~n22225 ) | ( n22223 & ~n22225 ) ;
  assign n22227 = ( n194 & n14408 ) | ( n194 & n22226 ) | ( n14408 & n22226 ) ;
  assign n22228 = n12406 ^ n5766 ^ n2616 ;
  assign n22229 = ( n16954 & n20060 ) | ( n16954 & n22228 ) | ( n20060 & n22228 ) ;
  assign n22234 = ( n4193 & n6651 ) | ( n4193 & ~n7255 ) | ( n6651 & ~n7255 ) ;
  assign n22230 = ( n5567 & ~n8745 ) | ( n5567 & n16687 ) | ( ~n8745 & n16687 ) ;
  assign n22231 = n22230 ^ n7389 ^ n7063 ;
  assign n22232 = n22231 ^ n8618 ^ n7159 ;
  assign n22233 = n22232 ^ n9103 ^ n3858 ;
  assign n22235 = n22234 ^ n22233 ^ n4036 ;
  assign n22239 = n18073 ^ n16665 ^ n6257 ;
  assign n22240 = ( ~n1299 & n7056 ) | ( ~n1299 & n22239 ) | ( n7056 & n22239 ) ;
  assign n22236 = ( n6922 & n7897 ) | ( n6922 & n18273 ) | ( n7897 & n18273 ) ;
  assign n22237 = ( n1647 & ~n20195 ) | ( n1647 & n22236 ) | ( ~n20195 & n22236 ) ;
  assign n22238 = n22237 ^ n21194 ^ x95 ;
  assign n22241 = n22240 ^ n22238 ^ n13055 ;
  assign n22242 = ( x33 & ~n4435 ) | ( x33 & n5630 ) | ( ~n4435 & n5630 ) ;
  assign n22243 = n11297 ^ n9095 ^ n6739 ;
  assign n22244 = n22243 ^ n5829 ^ n5178 ;
  assign n22245 = ( n11584 & n22231 ) | ( n11584 & ~n22244 ) | ( n22231 & ~n22244 ) ;
  assign n22250 = n18824 ^ n11438 ^ n8741 ;
  assign n22246 = ( n4722 & n9761 ) | ( n4722 & ~n19129 ) | ( n9761 & ~n19129 ) ;
  assign n22247 = ( n2416 & n8494 ) | ( n2416 & ~n9787 ) | ( n8494 & ~n9787 ) ;
  assign n22248 = ( n625 & n22246 ) | ( n625 & n22247 ) | ( n22246 & n22247 ) ;
  assign n22249 = n22248 ^ n3898 ^ n1510 ;
  assign n22251 = n22250 ^ n22249 ^ n2925 ;
  assign n22252 = ( ~n9132 & n22245 ) | ( ~n9132 & n22251 ) | ( n22245 & n22251 ) ;
  assign n22255 = ( n7720 & ~n10185 ) | ( n7720 & n13134 ) | ( ~n10185 & n13134 ) ;
  assign n22256 = n22255 ^ n10136 ^ n6461 ;
  assign n22253 = n7336 ^ n5770 ^ n1710 ;
  assign n22254 = n22253 ^ n10688 ^ n820 ;
  assign n22257 = n22256 ^ n22254 ^ n16225 ;
  assign n22258 = ( n3170 & n5802 ) | ( n3170 & n16041 ) | ( n5802 & n16041 ) ;
  assign n22259 = ( ~n1474 & n2575 ) | ( ~n1474 & n7403 ) | ( n2575 & n7403 ) ;
  assign n22260 = n22259 ^ n11735 ^ n4352 ;
  assign n22261 = ( ~n1476 & n20325 ) | ( ~n1476 & n22260 ) | ( n20325 & n22260 ) ;
  assign n22263 = ( n3131 & n3529 ) | ( n3131 & ~n3842 ) | ( n3529 & ~n3842 ) ;
  assign n22262 = n21848 ^ n14353 ^ n4281 ;
  assign n22264 = n22263 ^ n22262 ^ n1278 ;
  assign n22265 = ( n6018 & ~n21833 ) | ( n6018 & n22264 ) | ( ~n21833 & n22264 ) ;
  assign n22268 = ( ~n5281 & n5859 ) | ( ~n5281 & n6043 ) | ( n5859 & n6043 ) ;
  assign n22269 = ( n217 & ~n7804 ) | ( n217 & n17659 ) | ( ~n7804 & n17659 ) ;
  assign n22270 = ( n8457 & n22268 ) | ( n8457 & n22269 ) | ( n22268 & n22269 ) ;
  assign n22266 = ( n190 & n3429 ) | ( n190 & n5823 ) | ( n3429 & n5823 ) ;
  assign n22267 = n22266 ^ n6314 ^ n4536 ;
  assign n22271 = n22270 ^ n22267 ^ n8761 ;
  assign n22272 = n17025 ^ n13825 ^ n3326 ;
  assign n22276 = ( n3638 & n11944 ) | ( n3638 & ~n12033 ) | ( n11944 & ~n12033 ) ;
  assign n22275 = n16012 ^ n12936 ^ n3590 ;
  assign n22273 = n19278 ^ n2635 ^ n2328 ;
  assign n22274 = ( ~n8480 & n14052 ) | ( ~n8480 & n22273 ) | ( n14052 & n22273 ) ;
  assign n22277 = n22276 ^ n22275 ^ n22274 ;
  assign n22278 = n22277 ^ n4548 ^ n3635 ;
  assign n22279 = n11173 ^ n10222 ^ n4615 ;
  assign n22280 = n12845 ^ n6877 ^ n1290 ;
  assign n22281 = n22280 ^ n20121 ^ n9952 ;
  assign n22282 = n19727 ^ n4307 ^ n1099 ;
  assign n22283 = ( n5031 & n22281 ) | ( n5031 & n22282 ) | ( n22281 & n22282 ) ;
  assign n22286 = ( n794 & ~n3080 ) | ( n794 & n10237 ) | ( ~n3080 & n10237 ) ;
  assign n22284 = n11071 ^ n4155 ^ n2289 ;
  assign n22285 = n22284 ^ n5864 ^ n5021 ;
  assign n22287 = n22286 ^ n22285 ^ n19625 ;
  assign n22288 = ( ~n3229 & n15979 ) | ( ~n3229 & n22287 ) | ( n15979 & n22287 ) ;
  assign n22289 = n22288 ^ n21636 ^ n16603 ;
  assign n22294 = ( n3418 & ~n5099 ) | ( n3418 & n7329 ) | ( ~n5099 & n7329 ) ;
  assign n22290 = ( n5721 & n6220 ) | ( n5721 & ~n21289 ) | ( n6220 & ~n21289 ) ;
  assign n22291 = n15701 ^ n14689 ^ n994 ;
  assign n22292 = ( n1265 & n11381 ) | ( n1265 & ~n22291 ) | ( n11381 & ~n22291 ) ;
  assign n22293 = ( n13238 & n22290 ) | ( n13238 & ~n22292 ) | ( n22290 & ~n22292 ) ;
  assign n22295 = n22294 ^ n22293 ^ n4237 ;
  assign n22296 = ( n6039 & n10140 ) | ( n6039 & n14819 ) | ( n10140 & n14819 ) ;
  assign n22298 = ( n1383 & n3341 ) | ( n1383 & n10496 ) | ( n3341 & n10496 ) ;
  assign n22299 = n22298 ^ n16492 ^ n6394 ;
  assign n22297 = n13102 ^ n10626 ^ n4146 ;
  assign n22300 = n22299 ^ n22297 ^ n21983 ;
  assign n22301 = n22300 ^ n1728 ^ n1359 ;
  assign n22302 = n3720 ^ n3285 ^ n1551 ;
  assign n22303 = n10050 ^ n7115 ^ n6211 ;
  assign n22306 = n12635 ^ n5822 ^ n2667 ;
  assign n22307 = n22306 ^ n9043 ^ n3326 ;
  assign n22304 = ( n556 & ~n1699 ) | ( n556 & n2222 ) | ( ~n1699 & n2222 ) ;
  assign n22305 = ( n14595 & n16033 ) | ( n14595 & n22304 ) | ( n16033 & n22304 ) ;
  assign n22308 = n22307 ^ n22305 ^ n13114 ;
  assign n22309 = ( n7145 & n21535 ) | ( n7145 & ~n22308 ) | ( n21535 & ~n22308 ) ;
  assign n22310 = n20546 ^ n12241 ^ n8408 ;
  assign n22311 = ( n8955 & n20625 ) | ( n8955 & ~n22310 ) | ( n20625 & ~n22310 ) ;
  assign n22312 = ( n2296 & n4774 ) | ( n2296 & n11945 ) | ( n4774 & n11945 ) ;
  assign n22313 = n3743 ^ n3695 ^ n3088 ;
  assign n22314 = ( n5232 & n22312 ) | ( n5232 & n22313 ) | ( n22312 & n22313 ) ;
  assign n22315 = n21667 ^ n15074 ^ n2531 ;
  assign n22316 = ( n13411 & ~n18743 ) | ( n13411 & n22315 ) | ( ~n18743 & n22315 ) ;
  assign n22317 = ( n7565 & ~n13522 ) | ( n7565 & n20008 ) | ( ~n13522 & n20008 ) ;
  assign n22318 = ( n5125 & n12149 ) | ( n5125 & ~n22087 ) | ( n12149 & ~n22087 ) ;
  assign n22319 = n22318 ^ n10329 ^ n2088 ;
  assign n22320 = n22319 ^ n4307 ^ n2452 ;
  assign n22321 = ( n3091 & n7226 ) | ( n3091 & ~n8945 ) | ( n7226 & ~n8945 ) ;
  assign n22322 = n22321 ^ n6231 ^ n3081 ;
  assign n22323 = ( n4605 & n8067 ) | ( n4605 & ~n17416 ) | ( n8067 & ~n17416 ) ;
  assign n22324 = n14790 ^ n10501 ^ n8253 ;
  assign n22325 = ( n301 & n17039 ) | ( n301 & ~n22324 ) | ( n17039 & ~n22324 ) ;
  assign n22326 = ( n181 & n4616 ) | ( n181 & n22325 ) | ( n4616 & n22325 ) ;
  assign n22327 = n22326 ^ n21342 ^ n19163 ;
  assign n22329 = n19258 ^ n16047 ^ n9072 ;
  assign n22328 = ( n13356 & n16150 ) | ( n13356 & ~n17459 ) | ( n16150 & ~n17459 ) ;
  assign n22330 = n22329 ^ n22328 ^ n13585 ;
  assign n22331 = ( ~n1353 & n2028 ) | ( ~n1353 & n9291 ) | ( n2028 & n9291 ) ;
  assign n22332 = n20815 ^ n18783 ^ n347 ;
  assign n22333 = ( n12135 & n22286 ) | ( n12135 & ~n22332 ) | ( n22286 & ~n22332 ) ;
  assign n22334 = ( n4070 & n12537 ) | ( n4070 & n13534 ) | ( n12537 & n13534 ) ;
  assign n22335 = n22334 ^ n14793 ^ n6803 ;
  assign n22336 = ( n2455 & n5813 ) | ( n2455 & ~n7778 ) | ( n5813 & ~n7778 ) ;
  assign n22337 = ( n11529 & n19694 ) | ( n11529 & n22336 ) | ( n19694 & n22336 ) ;
  assign n22338 = n22337 ^ n20392 ^ n1236 ;
  assign n22339 = ( n6490 & ~n11493 ) | ( n6490 & n12138 ) | ( ~n11493 & n12138 ) ;
  assign n22340 = ( ~n7140 & n9094 ) | ( ~n7140 & n22339 ) | ( n9094 & n22339 ) ;
  assign n22341 = ( n483 & ~n1700 ) | ( n483 & n6562 ) | ( ~n1700 & n6562 ) ;
  assign n22342 = n22341 ^ n19864 ^ n19596 ;
  assign n22343 = n15509 ^ n15175 ^ n6125 ;
  assign n22344 = n22343 ^ n11476 ^ n4572 ;
  assign n22345 = n18386 ^ n12540 ^ n11542 ;
  assign n22346 = ( ~n1488 & n7093 ) | ( ~n1488 & n17092 ) | ( n7093 & n17092 ) ;
  assign n22347 = n22346 ^ n21219 ^ n4421 ;
  assign n22348 = ( n484 & n12767 ) | ( n484 & n21295 ) | ( n12767 & n21295 ) ;
  assign n22350 = n17750 ^ n9855 ^ n8879 ;
  assign n22349 = ( n5919 & n7793 ) | ( n5919 & n17049 ) | ( n7793 & n17049 ) ;
  assign n22351 = n22350 ^ n22349 ^ n9208 ;
  assign n22352 = n17538 ^ n6575 ^ n711 ;
  assign n22353 = ( n5840 & n7743 ) | ( n5840 & ~n22352 ) | ( n7743 & ~n22352 ) ;
  assign n22354 = ( ~n8405 & n10940 ) | ( ~n8405 & n22353 ) | ( n10940 & n22353 ) ;
  assign n22355 = n16741 ^ n8712 ^ n368 ;
  assign n22356 = n22057 ^ n14862 ^ n4879 ;
  assign n22357 = ( n2127 & n6472 ) | ( n2127 & n18692 ) | ( n6472 & n18692 ) ;
  assign n22360 = n14273 ^ n9491 ^ n2333 ;
  assign n22358 = ( n7573 & ~n14800 ) | ( n7573 & n16099 ) | ( ~n14800 & n16099 ) ;
  assign n22359 = n22358 ^ n17158 ^ n17070 ;
  assign n22361 = n22360 ^ n22359 ^ n16889 ;
  assign n22362 = ( n1466 & n3761 ) | ( n1466 & ~n3929 ) | ( n3761 & ~n3929 ) ;
  assign n22363 = n22362 ^ n7394 ^ n424 ;
  assign n22364 = n22363 ^ n22336 ^ n16412 ;
  assign n22365 = ( n837 & ~n15638 ) | ( n837 & n22364 ) | ( ~n15638 & n22364 ) ;
  assign n22366 = ( n4171 & n5185 ) | ( n4171 & ~n18444 ) | ( n5185 & ~n18444 ) ;
  assign n22367 = n15265 ^ n13104 ^ n737 ;
  assign n22368 = ( n4372 & n8172 ) | ( n4372 & ~n13269 ) | ( n8172 & ~n13269 ) ;
  assign n22369 = n19697 ^ n13053 ^ n5734 ;
  assign n22370 = n19980 ^ n9025 ^ n3000 ;
  assign n22371 = n22370 ^ n12658 ^ n5604 ;
  assign n22372 = ( n7247 & n16564 ) | ( n7247 & ~n19573 ) | ( n16564 & ~n19573 ) ;
  assign n22373 = n17419 ^ n6423 ^ n3575 ;
  assign n22374 = n22373 ^ n9307 ^ n8583 ;
  assign n22375 = ( n10411 & n14099 ) | ( n10411 & ~n15244 ) | ( n14099 & ~n15244 ) ;
  assign n22376 = n22375 ^ n11404 ^ n6915 ;
  assign n22377 = n22376 ^ n5161 ^ n4620 ;
  assign n22378 = n10243 ^ n5315 ^ n661 ;
  assign n22379 = n17559 ^ n8198 ^ n1941 ;
  assign n22380 = n22379 ^ n20975 ^ n20177 ;
  assign n22381 = n6562 ^ n4795 ^ n943 ;
  assign n22382 = n20879 ^ n17249 ^ n14012 ;
  assign n22383 = ( n11515 & ~n21748 ) | ( n11515 & n22382 ) | ( ~n21748 & n22382 ) ;
  assign n22384 = ( n754 & ~n1466 ) | ( n754 & n6248 ) | ( ~n1466 & n6248 ) ;
  assign n22385 = ( n4902 & ~n7699 ) | ( n4902 & n11794 ) | ( ~n7699 & n11794 ) ;
  assign n22386 = ( ~n7778 & n11956 ) | ( ~n7778 & n22385 ) | ( n11956 & n22385 ) ;
  assign n22387 = ( n11886 & n17121 ) | ( n11886 & n22386 ) | ( n17121 & n22386 ) ;
  assign n22388 = n13654 ^ n11574 ^ n8668 ;
  assign n22389 = ( ~n4248 & n6088 ) | ( ~n4248 & n22388 ) | ( n6088 & n22388 ) ;
  assign n22390 = n17544 ^ n15852 ^ n979 ;
  assign n22391 = ( n5066 & n10856 ) | ( n5066 & ~n19565 ) | ( n10856 & ~n19565 ) ;
  assign n22392 = n13292 ^ n5854 ^ n5221 ;
  assign n22393 = ( ~n4602 & n5997 ) | ( ~n4602 & n6570 ) | ( n5997 & n6570 ) ;
  assign n22394 = ( n14605 & n22392 ) | ( n14605 & n22393 ) | ( n22392 & n22393 ) ;
  assign n22395 = ( ~n22390 & n22391 ) | ( ~n22390 & n22394 ) | ( n22391 & n22394 ) ;
  assign n22396 = n10513 ^ n6461 ^ n5079 ;
  assign n22397 = ( n17467 & n22385 ) | ( n17467 & n22396 ) | ( n22385 & n22396 ) ;
  assign n22398 = ( n2099 & n12435 ) | ( n2099 & n19118 ) | ( n12435 & n19118 ) ;
  assign n22399 = n10819 ^ n3591 ^ n2642 ;
  assign n22400 = ( n12077 & n22398 ) | ( n12077 & n22399 ) | ( n22398 & n22399 ) ;
  assign n22401 = ( n21697 & n22397 ) | ( n21697 & n22400 ) | ( n22397 & n22400 ) ;
  assign n22402 = ( n2134 & n6715 ) | ( n2134 & ~n12739 ) | ( n6715 & ~n12739 ) ;
  assign n22403 = ( n3368 & ~n9270 ) | ( n3368 & n22402 ) | ( ~n9270 & n22402 ) ;
  assign n22404 = ( ~n17623 & n20543 ) | ( ~n17623 & n22403 ) | ( n20543 & n22403 ) ;
  assign n22405 = ( n2453 & n6681 ) | ( n2453 & ~n13218 ) | ( n6681 & ~n13218 ) ;
  assign n22406 = n13641 ^ n7799 ^ n4489 ;
  assign n22407 = n22406 ^ n16599 ^ n14606 ;
  assign n22408 = ( n11363 & ~n14308 ) | ( n11363 & n20946 ) | ( ~n14308 & n20946 ) ;
  assign n22410 = ( n7420 & ~n8094 ) | ( n7420 & n9112 ) | ( ~n8094 & n9112 ) ;
  assign n22411 = ( n7296 & n15574 ) | ( n7296 & ~n22410 ) | ( n15574 & ~n22410 ) ;
  assign n22412 = ( ~n3593 & n8204 ) | ( ~n3593 & n22411 ) | ( n8204 & n22411 ) ;
  assign n22409 = ( n1050 & n13104 ) | ( n1050 & n14705 ) | ( n13104 & n14705 ) ;
  assign n22413 = n22412 ^ n22409 ^ n18152 ;
  assign n22414 = ( n7133 & n12399 ) | ( n7133 & n17339 ) | ( n12399 & n17339 ) ;
  assign n22415 = n9365 ^ n4131 ^ n1364 ;
  assign n22416 = n22230 ^ n20757 ^ n1008 ;
  assign n22417 = ( n9989 & n15668 ) | ( n9989 & n22416 ) | ( n15668 & n22416 ) ;
  assign n22418 = ( n22414 & n22415 ) | ( n22414 & ~n22417 ) | ( n22415 & ~n22417 ) ;
  assign n22419 = ( n1586 & n7428 ) | ( n1586 & n18075 ) | ( n7428 & n18075 ) ;
  assign n22420 = n14448 ^ n10607 ^ n4914 ;
  assign n22421 = ( ~n10931 & n22419 ) | ( ~n10931 & n22420 ) | ( n22419 & n22420 ) ;
  assign n22422 = ( n8410 & n11454 ) | ( n8410 & n22421 ) | ( n11454 & n22421 ) ;
  assign n22423 = n22422 ^ n19916 ^ n3811 ;
  assign n22426 = ( n4756 & n6275 ) | ( n4756 & n14754 ) | ( n6275 & n14754 ) ;
  assign n22424 = ( n1205 & n1476 ) | ( n1205 & n10089 ) | ( n1476 & n10089 ) ;
  assign n22425 = n22424 ^ n11418 ^ n10657 ;
  assign n22427 = n22426 ^ n22425 ^ n13991 ;
  assign n22428 = ( n1045 & ~n9249 ) | ( n1045 & n15825 ) | ( ~n9249 & n15825 ) ;
  assign n22429 = n18579 ^ n17105 ^ n523 ;
  assign n22434 = n11428 ^ n6094 ^ n197 ;
  assign n22433 = n6955 ^ n5685 ^ n2228 ;
  assign n22430 = ( n2590 & ~n7136 ) | ( n2590 & n11077 ) | ( ~n7136 & n11077 ) ;
  assign n22431 = ( n12849 & n21416 ) | ( n12849 & n22430 ) | ( n21416 & n22430 ) ;
  assign n22432 = ( n4556 & n5130 ) | ( n4556 & n22431 ) | ( n5130 & n22431 ) ;
  assign n22435 = n22434 ^ n22433 ^ n22432 ;
  assign n22436 = ( ~n2615 & n4783 ) | ( ~n2615 & n8770 ) | ( n4783 & n8770 ) ;
  assign n22437 = ( n8801 & n9377 ) | ( n8801 & n12150 ) | ( n9377 & n12150 ) ;
  assign n22438 = ( n3321 & ~n11604 ) | ( n3321 & n16240 ) | ( ~n11604 & n16240 ) ;
  assign n22439 = ( ~n514 & n22437 ) | ( ~n514 & n22438 ) | ( n22437 & n22438 ) ;
  assign n22442 = n20182 ^ n17779 ^ n2857 ;
  assign n22440 = n11847 ^ n7484 ^ n6500 ;
  assign n22441 = ( ~n12672 & n16702 ) | ( ~n12672 & n22440 ) | ( n16702 & n22440 ) ;
  assign n22443 = n22442 ^ n22441 ^ n16834 ;
  assign n22445 = n10117 ^ n9797 ^ n9349 ;
  assign n22444 = n9133 ^ n6015 ^ n5068 ;
  assign n22446 = n22445 ^ n22444 ^ n2436 ;
  assign n22447 = ( n2115 & n20566 ) | ( n2115 & ~n22446 ) | ( n20566 & ~n22446 ) ;
  assign n22448 = n22447 ^ n20599 ^ n15778 ;
  assign n22449 = n20957 ^ n10960 ^ n2298 ;
  assign n22450 = n6629 ^ n5061 ^ x55 ;
  assign n22451 = n18801 ^ n10432 ^ n1035 ;
  assign n22452 = ( n21912 & n22450 ) | ( n21912 & n22451 ) | ( n22450 & n22451 ) ;
  assign n22453 = ( ~n2427 & n7920 ) | ( ~n2427 & n22360 ) | ( n7920 & n22360 ) ;
  assign n22454 = ( ~n9421 & n18391 ) | ( ~n9421 & n22453 ) | ( n18391 & n22453 ) ;
  assign n22455 = n19596 ^ n10682 ^ n3242 ;
  assign n22456 = ( n14881 & n17298 ) | ( n14881 & ~n22455 ) | ( n17298 & ~n22455 ) ;
  assign n22459 = ( n2303 & n9024 ) | ( n2303 & ~n13698 ) | ( n9024 & ~n13698 ) ;
  assign n22460 = n22459 ^ n15893 ^ n8529 ;
  assign n22457 = ( n3198 & ~n3686 ) | ( n3198 & n10467 ) | ( ~n3686 & n10467 ) ;
  assign n22458 = n22457 ^ n5639 ^ n5471 ;
  assign n22461 = n22460 ^ n22458 ^ n13472 ;
  assign n22462 = ( n9472 & ~n22456 ) | ( n9472 & n22461 ) | ( ~n22456 & n22461 ) ;
  assign n22463 = n5469 ^ n2987 ^ n2009 ;
  assign n22464 = ( n4600 & n7459 ) | ( n4600 & ~n14169 ) | ( n7459 & ~n14169 ) ;
  assign n22465 = n18810 ^ n12071 ^ n406 ;
  assign n22466 = ( n22463 & n22464 ) | ( n22463 & n22465 ) | ( n22464 & n22465 ) ;
  assign n22467 = ( ~n768 & n2504 ) | ( ~n768 & n6688 ) | ( n2504 & n6688 ) ;
  assign n22468 = n22467 ^ n2493 ^ n500 ;
  assign n22469 = n15875 ^ n6397 ^ n727 ;
  assign n22470 = ( n17844 & n22468 ) | ( n17844 & n22469 ) | ( n22468 & n22469 ) ;
  assign n22471 = ( n7388 & ~n11879 ) | ( n7388 & n15669 ) | ( ~n11879 & n15669 ) ;
  assign n22472 = n22471 ^ n20474 ^ n15627 ;
  assign n22473 = ( n2807 & ~n5753 ) | ( n2807 & n20169 ) | ( ~n5753 & n20169 ) ;
  assign n22474 = ( n3079 & n7772 ) | ( n3079 & n10401 ) | ( n7772 & n10401 ) ;
  assign n22475 = n22474 ^ n19605 ^ n4568 ;
  assign n22476 = ( n2214 & ~n3260 ) | ( n2214 & n20462 ) | ( ~n3260 & n20462 ) ;
  assign n22477 = n22476 ^ n13756 ^ n7165 ;
  assign n22478 = n7452 ^ n4982 ^ n3407 ;
  assign n22479 = n22478 ^ n8166 ^ n4402 ;
  assign n22480 = n22262 ^ n13965 ^ n1539 ;
  assign n22481 = ( n2349 & n2533 ) | ( n2349 & n7057 ) | ( n2533 & n7057 ) ;
  assign n22482 = ( n5171 & n21039 ) | ( n5171 & n21217 ) | ( n21039 & n21217 ) ;
  assign n22483 = ( n5220 & ~n22481 ) | ( n5220 & n22482 ) | ( ~n22481 & n22482 ) ;
  assign n22484 = n9963 ^ n7464 ^ n1376 ;
  assign n22485 = n22484 ^ n4611 ^ n3470 ;
  assign n22486 = n22485 ^ n21062 ^ n7970 ;
  assign n22487 = ( n4594 & n4861 ) | ( n4594 & n13726 ) | ( n4861 & n13726 ) ;
  assign n22488 = n22487 ^ n18995 ^ n569 ;
  assign n22489 = ( n376 & n12360 ) | ( n376 & n22488 ) | ( n12360 & n22488 ) ;
  assign n22490 = ( ~n6199 & n19939 ) | ( ~n6199 & n22489 ) | ( n19939 & n22489 ) ;
  assign n22491 = ( n2207 & ~n3550 ) | ( n2207 & n4791 ) | ( ~n3550 & n4791 ) ;
  assign n22492 = n12796 ^ n9654 ^ n9224 ;
  assign n22493 = ( n5402 & n13541 ) | ( n5402 & ~n22492 ) | ( n13541 & ~n22492 ) ;
  assign n22494 = ( n13183 & n18787 ) | ( n13183 & ~n22493 ) | ( n18787 & ~n22493 ) ;
  assign n22495 = ( n840 & n17993 ) | ( n840 & n21230 ) | ( n17993 & n21230 ) ;
  assign n22496 = ( n6701 & ~n22013 ) | ( n6701 & n22495 ) | ( ~n22013 & n22495 ) ;
  assign n22497 = ( n2562 & n9187 ) | ( n2562 & n9443 ) | ( n9187 & n9443 ) ;
  assign n22498 = ( n6573 & n21509 ) | ( n6573 & n22497 ) | ( n21509 & n22497 ) ;
  assign n22499 = ( n6461 & n8244 ) | ( n6461 & n22498 ) | ( n8244 & n22498 ) ;
  assign n22500 = n22499 ^ n21186 ^ n1926 ;
  assign n22501 = ( n2747 & ~n6462 ) | ( n2747 & n9319 ) | ( ~n6462 & n9319 ) ;
  assign n22502 = ( n3563 & ~n15560 ) | ( n3563 & n22501 ) | ( ~n15560 & n22501 ) ;
  assign n22503 = ( n2723 & ~n8107 ) | ( n2723 & n15800 ) | ( ~n8107 & n15800 ) ;
  assign n22504 = ( n613 & ~n22502 ) | ( n613 & n22503 ) | ( ~n22502 & n22503 ) ;
  assign n22505 = ( ~n2477 & n4487 ) | ( ~n2477 & n20195 ) | ( n4487 & n20195 ) ;
  assign n22506 = n11321 ^ n9363 ^ n3076 ;
  assign n22507 = ( ~n13668 & n17710 ) | ( ~n13668 & n19548 ) | ( n17710 & n19548 ) ;
  assign n22508 = ( ~n9550 & n21081 ) | ( ~n9550 & n22507 ) | ( n21081 & n22507 ) ;
  assign n22511 = ( n5373 & n12015 ) | ( n5373 & n14960 ) | ( n12015 & n14960 ) ;
  assign n22509 = n16481 ^ n13491 ^ n3801 ;
  assign n22510 = ( n5615 & ~n18145 ) | ( n5615 & n22509 ) | ( ~n18145 & n22509 ) ;
  assign n22512 = n22511 ^ n22510 ^ n2246 ;
  assign n22513 = ( ~x32 & n10644 ) | ( ~x32 & n18778 ) | ( n10644 & n18778 ) ;
  assign n22514 = ( n6986 & n14177 ) | ( n6986 & n22513 ) | ( n14177 & n22513 ) ;
  assign n22518 = n21674 ^ n11494 ^ n8342 ;
  assign n22515 = ( n2746 & ~n5140 ) | ( n2746 & n8516 ) | ( ~n5140 & n8516 ) ;
  assign n22516 = n14529 ^ n4343 ^ n820 ;
  assign n22517 = ( n20289 & ~n22515 ) | ( n20289 & n22516 ) | ( ~n22515 & n22516 ) ;
  assign n22519 = n22518 ^ n22517 ^ n7999 ;
  assign n22520 = n22519 ^ n8590 ^ n7746 ;
  assign n22521 = ( n5455 & n9492 ) | ( n5455 & n18512 ) | ( n9492 & n18512 ) ;
  assign n22522 = ( n5195 & ~n8298 ) | ( n5195 & n17190 ) | ( ~n8298 & n17190 ) ;
  assign n22523 = ( n14357 & ~n19160 ) | ( n14357 & n22522 ) | ( ~n19160 & n22522 ) ;
  assign n22524 = n12404 ^ n5831 ^ n1416 ;
  assign n22525 = ( n18000 & ~n18193 ) | ( n18000 & n22524 ) | ( ~n18193 & n22524 ) ;
  assign n22526 = ( n2798 & ~n10994 ) | ( n2798 & n12312 ) | ( ~n10994 & n12312 ) ;
  assign n22527 = n22526 ^ n6868 ^ n1698 ;
  assign n22528 = ( ~n11574 & n14098 ) | ( ~n11574 & n22456 ) | ( n14098 & n22456 ) ;
  assign n22529 = ( n363 & n5514 ) | ( n363 & n13366 ) | ( n5514 & n13366 ) ;
  assign n22530 = n22529 ^ n8109 ^ n3929 ;
  assign n22531 = n22530 ^ n15131 ^ n4366 ;
  assign n22532 = n21475 ^ n20530 ^ n3786 ;
  assign n22533 = n22532 ^ n9991 ^ n7779 ;
  assign n22534 = ( ~n3159 & n7426 ) | ( ~n3159 & n21269 ) | ( n7426 & n21269 ) ;
  assign n22535 = ( n10045 & ~n17287 ) | ( n10045 & n22534 ) | ( ~n17287 & n22534 ) ;
  assign n22536 = ( n5983 & ~n20029 ) | ( n5983 & n21783 ) | ( ~n20029 & n21783 ) ;
  assign n22537 = ( n194 & n603 ) | ( n194 & ~n11408 ) | ( n603 & ~n11408 ) ;
  assign n22538 = n6817 ^ n1270 ^ x115 ;
  assign n22539 = n22538 ^ n17574 ^ n14906 ;
  assign n22540 = n5472 ^ n3150 ^ n1162 ;
  assign n22541 = ( n535 & ~n926 ) | ( n535 & n4264 ) | ( ~n926 & n4264 ) ;
  assign n22542 = ( ~n2019 & n12635 ) | ( ~n2019 & n22541 ) | ( n12635 & n22541 ) ;
  assign n22543 = ( n4103 & n22540 ) | ( n4103 & n22542 ) | ( n22540 & n22542 ) ;
  assign n22544 = ( ~n1453 & n2195 ) | ( ~n1453 & n16714 ) | ( n2195 & n16714 ) ;
  assign n22545 = ( n2020 & ~n4653 ) | ( n2020 & n17148 ) | ( ~n4653 & n17148 ) ;
  assign n22546 = ( n507 & n1552 ) | ( n507 & ~n7207 ) | ( n1552 & ~n7207 ) ;
  assign n22547 = n7633 ^ n2935 ^ x54 ;
  assign n22548 = ( n7223 & ~n13776 ) | ( n7223 & n22547 ) | ( ~n13776 & n22547 ) ;
  assign n22549 = ( n9991 & n22546 ) | ( n9991 & ~n22548 ) | ( n22546 & ~n22548 ) ;
  assign n22550 = ( n1865 & ~n2978 ) | ( n1865 & n21445 ) | ( ~n2978 & n21445 ) ;
  assign n22552 = ( n2769 & n16376 ) | ( n2769 & ~n18029 ) | ( n16376 & ~n18029 ) ;
  assign n22553 = ( ~n3187 & n4224 ) | ( ~n3187 & n22552 ) | ( n4224 & n22552 ) ;
  assign n22551 = ( n12752 & ~n16323 ) | ( n12752 & n18738 ) | ( ~n16323 & n18738 ) ;
  assign n22554 = n22553 ^ n22551 ^ n18346 ;
  assign n22555 = ( n8883 & n12557 ) | ( n8883 & ~n22554 ) | ( n12557 & ~n22554 ) ;
  assign n22556 = n16963 ^ n7416 ^ n5865 ;
  assign n22557 = ( n1606 & n9884 ) | ( n1606 & n14006 ) | ( n9884 & n14006 ) ;
  assign n22558 = n22557 ^ n18970 ^ n14218 ;
  assign n22559 = n16832 ^ n16216 ^ n15153 ;
  assign n22560 = ( n7729 & n13356 ) | ( n7729 & ~n22559 ) | ( n13356 & ~n22559 ) ;
  assign n22561 = n8658 ^ n5023 ^ n4679 ;
  assign n22562 = ( ~n10482 & n21686 ) | ( ~n10482 & n22561 ) | ( n21686 & n22561 ) ;
  assign n22563 = n15955 ^ n14553 ^ n5009 ;
  assign n22564 = ( ~n3690 & n13543 ) | ( ~n3690 & n20645 ) | ( n13543 & n20645 ) ;
  assign n22565 = ( ~n11889 & n22563 ) | ( ~n11889 & n22564 ) | ( n22563 & n22564 ) ;
  assign n22566 = ( ~n587 & n1566 ) | ( ~n587 & n4944 ) | ( n1566 & n4944 ) ;
  assign n22567 = ( n7955 & n9747 ) | ( n7955 & n22566 ) | ( n9747 & n22566 ) ;
  assign n22568 = ( n4821 & ~n14851 ) | ( n4821 & n17551 ) | ( ~n14851 & n17551 ) ;
  assign n22569 = ( n11927 & n22567 ) | ( n11927 & ~n22568 ) | ( n22567 & ~n22568 ) ;
  assign n22570 = n15655 ^ n7148 ^ n4864 ;
  assign n22571 = n22570 ^ n17310 ^ n13091 ;
  assign n22572 = ( n5996 & ~n16181 ) | ( n5996 & n22571 ) | ( ~n16181 & n22571 ) ;
  assign n22573 = n20657 ^ n17822 ^ n14392 ;
  assign n22574 = ( ~n4943 & n21060 ) | ( ~n4943 & n22573 ) | ( n21060 & n22573 ) ;
  assign n22575 = ( n10119 & ~n15009 ) | ( n10119 & n22574 ) | ( ~n15009 & n22574 ) ;
  assign n22576 = n19387 ^ n17376 ^ n13838 ;
  assign n22577 = n19694 ^ n11789 ^ n6937 ;
  assign n22578 = n22577 ^ n2665 ^ n345 ;
  assign n22579 = ( n9687 & ~n15765 ) | ( n9687 & n22578 ) | ( ~n15765 & n22578 ) ;
  assign n22580 = ( n1704 & ~n6740 ) | ( n1704 & n8342 ) | ( ~n6740 & n8342 ) ;
  assign n22581 = n22580 ^ n18069 ^ n4216 ;
  assign n22582 = n19144 ^ n7601 ^ n712 ;
  assign n22583 = ( ~n9884 & n10617 ) | ( ~n9884 & n15855 ) | ( n10617 & n15855 ) ;
  assign n22584 = ( n3773 & n22582 ) | ( n3773 & ~n22583 ) | ( n22582 & ~n22583 ) ;
  assign n22585 = n15812 ^ n14132 ^ n11904 ;
  assign n22586 = ( n7570 & n8817 ) | ( n7570 & ~n21219 ) | ( n8817 & ~n21219 ) ;
  assign n22587 = ( n15664 & n19573 ) | ( n15664 & ~n22586 ) | ( n19573 & ~n22586 ) ;
  assign n22588 = ( ~n4576 & n5185 ) | ( ~n4576 & n7838 ) | ( n5185 & n7838 ) ;
  assign n22589 = ( n12351 & n17674 ) | ( n12351 & n22588 ) | ( n17674 & n22588 ) ;
  assign n22590 = n21006 ^ n20642 ^ n18237 ;
  assign n22591 = ( n414 & n13886 ) | ( n414 & ~n15541 ) | ( n13886 & ~n15541 ) ;
  assign n22592 = n15730 ^ n9868 ^ n184 ;
  assign n22593 = ( n8444 & n18937 ) | ( n8444 & ~n22592 ) | ( n18937 & ~n22592 ) ;
  assign n22594 = ( n3446 & n6257 ) | ( n3446 & ~n17716 ) | ( n6257 & ~n17716 ) ;
  assign n22595 = n22594 ^ n21057 ^ n5185 ;
  assign n22596 = ( n2132 & ~n6066 ) | ( n2132 & n20314 ) | ( ~n6066 & n20314 ) ;
  assign n22597 = n21454 ^ n15954 ^ n3765 ;
  assign n22598 = ( ~n2170 & n4795 ) | ( ~n2170 & n6084 ) | ( n4795 & n6084 ) ;
  assign n22599 = n16390 ^ n13055 ^ n5904 ;
  assign n22600 = ( ~n10237 & n22598 ) | ( ~n10237 & n22599 ) | ( n22598 & n22599 ) ;
  assign n22601 = ( n1000 & n2731 ) | ( n1000 & ~n10352 ) | ( n2731 & ~n10352 ) ;
  assign n22602 = n22601 ^ n16595 ^ n7488 ;
  assign n22603 = ( n3966 & ~n5552 ) | ( n3966 & n9460 ) | ( ~n5552 & n9460 ) ;
  assign n22604 = n22603 ^ n4995 ^ n383 ;
  assign n22605 = ( n19143 & ~n22602 ) | ( n19143 & n22604 ) | ( ~n22602 & n22604 ) ;
  assign n22606 = n20948 ^ n19200 ^ n5474 ;
  assign n22607 = ( n6062 & n12071 ) | ( n6062 & ~n14699 ) | ( n12071 & ~n14699 ) ;
  assign n22608 = n22607 ^ n7924 ^ n7468 ;
  assign n22609 = n20757 ^ n13363 ^ n6465 ;
  assign n22610 = ( ~n825 & n3514 ) | ( ~n825 & n16335 ) | ( n3514 & n16335 ) ;
  assign n22611 = n22610 ^ n4940 ^ n1178 ;
  assign n22612 = n15955 ^ n13692 ^ n6798 ;
  assign n22613 = ( n2527 & n4930 ) | ( n2527 & ~n6405 ) | ( n4930 & ~n6405 ) ;
  assign n22614 = n22613 ^ n3484 ^ n2243 ;
  assign n22615 = ( n9636 & n11429 ) | ( n9636 & ~n22614 ) | ( n11429 & ~n22614 ) ;
  assign n22616 = n22615 ^ n19056 ^ n11985 ;
  assign n22617 = ( ~n2148 & n4457 ) | ( ~n2148 & n20285 ) | ( n4457 & n20285 ) ;
  assign n22618 = ( ~n11264 & n14660 ) | ( ~n11264 & n20010 ) | ( n14660 & n20010 ) ;
  assign n22619 = n11927 ^ n8062 ^ n1167 ;
  assign n22620 = n22619 ^ n16389 ^ n13523 ;
  assign n22621 = n22620 ^ n14058 ^ n9795 ;
  assign n22622 = n14581 ^ n11753 ^ n10994 ;
  assign n22623 = ( n5563 & n15861 ) | ( n5563 & ~n22622 ) | ( n15861 & ~n22622 ) ;
  assign n22624 = n22125 ^ n20907 ^ n982 ;
  assign n22625 = n22624 ^ n20208 ^ n5110 ;
  assign n22626 = ( n2143 & ~n9164 ) | ( n2143 & n9932 ) | ( ~n9164 & n9932 ) ;
  assign n22627 = ( ~n1911 & n10651 ) | ( ~n1911 & n12439 ) | ( n10651 & n12439 ) ;
  assign n22628 = ( ~n8723 & n16611 ) | ( ~n8723 & n21742 ) | ( n16611 & n21742 ) ;
  assign n22629 = n9991 ^ n5362 ^ n826 ;
  assign n22630 = n14923 ^ n5823 ^ n4508 ;
  assign n22631 = ( n8682 & n9163 ) | ( n8682 & ~n22630 ) | ( n9163 & ~n22630 ) ;
  assign n22632 = ( ~n13168 & n22629 ) | ( ~n13168 & n22631 ) | ( n22629 & n22631 ) ;
  assign n22633 = ( ~n20110 & n22628 ) | ( ~n20110 & n22632 ) | ( n22628 & n22632 ) ;
  assign n22634 = ( n1299 & n5683 ) | ( n1299 & ~n10213 ) | ( n5683 & ~n10213 ) ;
  assign n22635 = n22634 ^ n7175 ^ n4307 ;
  assign n22636 = n4419 ^ n450 ^ x118 ;
  assign n22637 = ( n2824 & n12854 ) | ( n2824 & ~n22636 ) | ( n12854 & ~n22636 ) ;
  assign n22638 = n22637 ^ n10251 ^ n8960 ;
  assign n22639 = ( ~n18630 & n20753 ) | ( ~n18630 & n22638 ) | ( n20753 & n22638 ) ;
  assign n22640 = n14520 ^ n2644 ^ n1320 ;
  assign n22641 = ( ~n4967 & n9890 ) | ( ~n4967 & n22640 ) | ( n9890 & n22640 ) ;
  assign n22642 = n13087 ^ n9897 ^ n9857 ;
  assign n22643 = ( ~n15876 & n22641 ) | ( ~n15876 & n22642 ) | ( n22641 & n22642 ) ;
  assign n22644 = ( n1053 & ~n2828 ) | ( n1053 & n4645 ) | ( ~n2828 & n4645 ) ;
  assign n22645 = n4897 ^ n4778 ^ n335 ;
  assign n22646 = ( n8666 & n22644 ) | ( n8666 & ~n22645 ) | ( n22644 & ~n22645 ) ;
  assign n22647 = ( ~n904 & n7020 ) | ( ~n904 & n13089 ) | ( n7020 & n13089 ) ;
  assign n22648 = ( n2388 & n22646 ) | ( n2388 & n22647 ) | ( n22646 & n22647 ) ;
  assign n22649 = ( n3682 & n5480 ) | ( n3682 & ~n8189 ) | ( n5480 & ~n8189 ) ;
  assign n22650 = n22649 ^ n20207 ^ n18244 ;
  assign n22651 = n22650 ^ n4859 ^ n3160 ;
  assign n22652 = ( n779 & ~n9567 ) | ( n779 & n18005 ) | ( ~n9567 & n18005 ) ;
  assign n22653 = n22652 ^ n13098 ^ n9068 ;
  assign n22654 = ( n2036 & n2124 ) | ( n2036 & ~n13533 ) | ( n2124 & ~n13533 ) ;
  assign n22655 = ( n8200 & ~n8974 ) | ( n8200 & n22654 ) | ( ~n8974 & n22654 ) ;
  assign n22657 = n16929 ^ n13579 ^ n10198 ;
  assign n22656 = n7176 ^ n4686 ^ n975 ;
  assign n22658 = n22657 ^ n22656 ^ n7678 ;
  assign n22659 = ( n8249 & ~n16751 ) | ( n8249 & n20927 ) | ( ~n16751 & n20927 ) ;
  assign n22660 = n14041 ^ n13491 ^ n6383 ;
  assign n22661 = n22660 ^ n19043 ^ n1496 ;
  assign n22662 = n20625 ^ n18410 ^ n5385 ;
  assign n22663 = n22662 ^ n20519 ^ n3249 ;
  assign n22664 = n18344 ^ n5920 ^ n2911 ;
  assign n22665 = ( n11079 & ~n22663 ) | ( n11079 & n22664 ) | ( ~n22663 & n22664 ) ;
  assign n22666 = ( n8333 & ~n10096 ) | ( n8333 & n12680 ) | ( ~n10096 & n12680 ) ;
  assign n22668 = ( n3714 & n6534 ) | ( n3714 & ~n19489 ) | ( n6534 & ~n19489 ) ;
  assign n22667 = n19406 ^ n17206 ^ n12070 ;
  assign n22669 = n22668 ^ n22667 ^ n9045 ;
  assign n22673 = n17106 ^ n3091 ^ n2440 ;
  assign n22674 = ( n3344 & ~n15740 ) | ( n3344 & n22673 ) | ( ~n15740 & n22673 ) ;
  assign n22671 = n16892 ^ n9314 ^ n4111 ;
  assign n22672 = n22671 ^ n22086 ^ n4610 ;
  assign n22670 = ( n5727 & ~n12545 ) | ( n5727 & n16965 ) | ( ~n12545 & n16965 ) ;
  assign n22675 = n22674 ^ n22672 ^ n22670 ;
  assign n22676 = ( n966 & ~n4508 ) | ( n966 & n21791 ) | ( ~n4508 & n21791 ) ;
  assign n22677 = ( ~n6609 & n14168 ) | ( ~n6609 & n15877 ) | ( n14168 & n15877 ) ;
  assign n22678 = ( n10058 & ~n21204 ) | ( n10058 & n22677 ) | ( ~n21204 & n22677 ) ;
  assign n22679 = n22678 ^ n14854 ^ n9907 ;
  assign n22680 = n22360 ^ n10103 ^ n5193 ;
  assign n22681 = n14278 ^ n9957 ^ n7357 ;
  assign n22682 = ( n7355 & n17291 ) | ( n7355 & n22681 ) | ( n17291 & n22681 ) ;
  assign n22683 = n22450 ^ n11869 ^ n8674 ;
  assign n22685 = n22634 ^ n14537 ^ n4876 ;
  assign n22686 = n10196 ^ n2512 ^ n2424 ;
  assign n22687 = n22686 ^ n9986 ^ n9623 ;
  assign n22688 = ( ~n4327 & n22685 ) | ( ~n4327 & n22687 ) | ( n22685 & n22687 ) ;
  assign n22684 = n14171 ^ n5664 ^ n130 ;
  assign n22689 = n22688 ^ n22684 ^ n2758 ;
  assign n22690 = ( n3552 & n12466 ) | ( n3552 & n22689 ) | ( n12466 & n22689 ) ;
  assign n22692 = ( ~n9062 & n10027 ) | ( ~n9062 & n13853 ) | ( n10027 & n13853 ) ;
  assign n22691 = n12162 ^ n11472 ^ n7374 ;
  assign n22693 = n22692 ^ n22691 ^ n7087 ;
  assign n22694 = n18073 ^ n7679 ^ n1465 ;
  assign n22695 = n20128 ^ n14069 ^ n4403 ;
  assign n22696 = n2598 ^ n1666 ^ n1328 ;
  assign n22697 = ( n5177 & n19681 ) | ( n5177 & ~n22696 ) | ( n19681 & ~n22696 ) ;
  assign n22698 = ( n158 & ~n2064 ) | ( n158 & n6487 ) | ( ~n2064 & n6487 ) ;
  assign n22699 = ( n7124 & ~n14301 ) | ( n7124 & n20149 ) | ( ~n14301 & n20149 ) ;
  assign n22700 = ( n3801 & n22698 ) | ( n3801 & n22699 ) | ( n22698 & n22699 ) ;
  assign n22701 = n22393 ^ n16292 ^ n10803 ;
  assign n22702 = ( ~n16950 & n19322 ) | ( ~n16950 & n19743 ) | ( n19322 & n19743 ) ;
  assign n22703 = ( n8831 & ~n21310 ) | ( n8831 & n22702 ) | ( ~n21310 & n22702 ) ;
  assign n22704 = ( ~n14265 & n18267 ) | ( ~n14265 & n21054 ) | ( n18267 & n21054 ) ;
  assign n22705 = n18358 ^ n1322 ^ n459 ;
  assign n22706 = n22570 ^ n5087 ^ n1672 ;
  assign n22707 = n21697 ^ n8214 ^ n5152 ;
  assign n22708 = n22707 ^ n5412 ^ n2509 ;
  assign n22709 = ( n728 & n22706 ) | ( n728 & ~n22708 ) | ( n22706 & ~n22708 ) ;
  assign n22711 = n18095 ^ n4030 ^ n2677 ;
  assign n22712 = n22711 ^ n11825 ^ n581 ;
  assign n22710 = ( n2028 & n13503 ) | ( n2028 & ~n18327 ) | ( n13503 & ~n18327 ) ;
  assign n22713 = n22712 ^ n22710 ^ n3002 ;
  assign n22714 = ( ~n11776 & n13463 ) | ( ~n11776 & n18157 ) | ( n13463 & n18157 ) ;
  assign n22715 = n11012 ^ n7803 ^ n5424 ;
  assign n22716 = n22715 ^ n8843 ^ n1874 ;
  assign n22717 = n13465 ^ n3344 ^ n1820 ;
  assign n22718 = n16959 ^ n10051 ^ n9107 ;
  assign n22719 = ( n7510 & n16415 ) | ( n7510 & n22718 ) | ( n16415 & n22718 ) ;
  assign n22720 = ( n3381 & ~n22717 ) | ( n3381 & n22719 ) | ( ~n22717 & n22719 ) ;
  assign n22721 = n22720 ^ n14714 ^ n9021 ;
  assign n22722 = n19725 ^ n19140 ^ n3406 ;
  assign n22723 = ( n2219 & n6005 ) | ( n2219 & n9364 ) | ( n6005 & n9364 ) ;
  assign n22724 = ( ~n6517 & n12254 ) | ( ~n6517 & n22723 ) | ( n12254 & n22723 ) ;
  assign n22725 = n22724 ^ n17770 ^ n4430 ;
  assign n22726 = n22725 ^ n16726 ^ n2713 ;
  assign n22727 = ( n21436 & n22722 ) | ( n21436 & n22726 ) | ( n22722 & n22726 ) ;
  assign n22728 = ( n844 & n6712 ) | ( n844 & n20334 ) | ( n6712 & n20334 ) ;
  assign n22729 = n22728 ^ n19362 ^ n6080 ;
  assign n22730 = ( n7419 & n7458 ) | ( n7419 & ~n10706 ) | ( n7458 & ~n10706 ) ;
  assign n22731 = n22730 ^ n19066 ^ n3282 ;
  assign n22732 = ( n1859 & n2296 ) | ( n1859 & ~n9032 ) | ( n2296 & ~n9032 ) ;
  assign n22733 = ( n9227 & n17122 ) | ( n9227 & n22732 ) | ( n17122 & n22732 ) ;
  assign n22734 = ( ~n19872 & n22731 ) | ( ~n19872 & n22733 ) | ( n22731 & n22733 ) ;
  assign n22735 = n18215 ^ n11202 ^ n3511 ;
  assign n22739 = n12995 ^ n8674 ^ n8494 ;
  assign n22740 = n22739 ^ n9420 ^ n1222 ;
  assign n22736 = n21661 ^ n13680 ^ n9399 ;
  assign n22737 = ( n9925 & ~n13178 ) | ( n9925 & n14972 ) | ( ~n13178 & n14972 ) ;
  assign n22738 = ( n11461 & n22736 ) | ( n11461 & n22737 ) | ( n22736 & n22737 ) ;
  assign n22741 = n22740 ^ n22738 ^ n10596 ;
  assign n22742 = ( n9980 & n15590 ) | ( n9980 & ~n19082 ) | ( n15590 & ~n19082 ) ;
  assign n22743 = n8201 ^ n6489 ^ n1657 ;
  assign n22744 = ( n10804 & ~n11052 ) | ( n10804 & n15213 ) | ( ~n11052 & n15213 ) ;
  assign n22747 = n15232 ^ n10863 ^ n1153 ;
  assign n22748 = n22747 ^ n8857 ^ n7391 ;
  assign n22745 = n6859 ^ n4029 ^ n2771 ;
  assign n22746 = n22745 ^ n1356 ^ n617 ;
  assign n22749 = n22748 ^ n22746 ^ n4403 ;
  assign n22750 = ( n7875 & n13221 ) | ( n7875 & n22749 ) | ( n13221 & n22749 ) ;
  assign n22751 = ( ~n3375 & n11326 ) | ( ~n3375 & n14573 ) | ( n11326 & n14573 ) ;
  assign n22752 = ( n2574 & n6448 ) | ( n2574 & n16772 ) | ( n6448 & n16772 ) ;
  assign n22753 = ( n22624 & n22751 ) | ( n22624 & n22752 ) | ( n22751 & n22752 ) ;
  assign n22754 = n13775 ^ n1872 ^ n1819 ;
  assign n22755 = n22754 ^ n8827 ^ n1067 ;
  assign n22756 = n14456 ^ n12037 ^ n7292 ;
  assign n22757 = n17203 ^ n12082 ^ n8588 ;
  assign n22758 = ( n2141 & n9496 ) | ( n2141 & n20184 ) | ( n9496 & n20184 ) ;
  assign n22759 = n22758 ^ n15172 ^ n461 ;
  assign n22760 = n22759 ^ n18160 ^ n11017 ;
  assign n22761 = n22760 ^ n19080 ^ n6744 ;
  assign n22762 = n10525 ^ n5189 ^ n4781 ;
  assign n22763 = n22762 ^ n14702 ^ n5984 ;
  assign n22764 = ( ~n10801 & n17644 ) | ( ~n10801 & n17982 ) | ( n17644 & n17982 ) ;
  assign n22765 = n22764 ^ n11364 ^ n10847 ;
  assign n22766 = ( n2160 & ~n5137 ) | ( n2160 & n11307 ) | ( ~n5137 & n11307 ) ;
  assign n22767 = n22766 ^ n8881 ^ n2147 ;
  assign n22768 = ( ~n5213 & n18327 ) | ( ~n5213 & n22767 ) | ( n18327 & n22767 ) ;
  assign n22774 = ( n3441 & n9412 ) | ( n3441 & n13689 ) | ( n9412 & n13689 ) ;
  assign n22773 = ( n6511 & n6805 ) | ( n6511 & n19385 ) | ( n6805 & n19385 ) ;
  assign n22770 = n20749 ^ n9956 ^ n4419 ;
  assign n22769 = ( n2229 & n5363 ) | ( n2229 & ~n13353 ) | ( n5363 & ~n13353 ) ;
  assign n22771 = n22770 ^ n22769 ^ n20778 ;
  assign n22772 = n22771 ^ n19069 ^ n15692 ;
  assign n22775 = n22774 ^ n22773 ^ n22772 ;
  assign n22776 = ( n13982 & n14037 ) | ( n13982 & ~n16003 ) | ( n14037 & ~n16003 ) ;
  assign n22777 = n22776 ^ n16803 ^ n9568 ;
  assign n22778 = n22634 ^ n21948 ^ n2353 ;
  assign n22779 = n22778 ^ n12349 ^ n10251 ;
  assign n22780 = ( n6024 & ~n18336 ) | ( n6024 & n22779 ) | ( ~n18336 & n22779 ) ;
  assign n22781 = ( n3100 & ~n6761 ) | ( n3100 & n12029 ) | ( ~n6761 & n12029 ) ;
  assign n22782 = ( n1260 & ~n2628 ) | ( n1260 & n3527 ) | ( ~n2628 & n3527 ) ;
  assign n22783 = n18250 ^ n12145 ^ n9568 ;
  assign n22784 = ( n5861 & ~n22782 ) | ( n5861 & n22783 ) | ( ~n22782 & n22783 ) ;
  assign n22785 = ( n19387 & n22781 ) | ( n19387 & ~n22784 ) | ( n22781 & ~n22784 ) ;
  assign n22786 = ( n1354 & n17710 ) | ( n1354 & n22785 ) | ( n17710 & n22785 ) ;
  assign n22787 = ( n7108 & ~n10023 ) | ( n7108 & n14596 ) | ( ~n10023 & n14596 ) ;
  assign n22788 = ( n428 & n2976 ) | ( n428 & ~n9325 ) | ( n2976 & ~n9325 ) ;
  assign n22789 = ( n8131 & n14351 ) | ( n8131 & n22788 ) | ( n14351 & n22788 ) ;
  assign n22790 = n15704 ^ n7148 ^ n5209 ;
  assign n22791 = n22790 ^ n17371 ^ n4677 ;
  assign n22792 = ( n3100 & n4412 ) | ( n3100 & ~n19704 ) | ( n4412 & ~n19704 ) ;
  assign n22793 = n20869 ^ n4101 ^ n2297 ;
  assign n22794 = ( ~n610 & n14044 ) | ( ~n610 & n22793 ) | ( n14044 & n22793 ) ;
  assign n22795 = ( ~n12565 & n22792 ) | ( ~n12565 & n22794 ) | ( n22792 & n22794 ) ;
  assign n22796 = n16193 ^ n9774 ^ n836 ;
  assign n22797 = n22796 ^ n15443 ^ n6755 ;
  assign n22798 = ( n3674 & ~n15542 ) | ( n3674 & n16464 ) | ( ~n15542 & n16464 ) ;
  assign n22800 = ( ~n192 & n6976 ) | ( ~n192 & n13398 ) | ( n6976 & n13398 ) ;
  assign n22799 = n15856 ^ n13479 ^ n6403 ;
  assign n22801 = n22800 ^ n22799 ^ n2942 ;
  assign n22802 = n11078 ^ n4219 ^ n696 ;
  assign n22803 = n22802 ^ n13358 ^ n7982 ;
  assign n22804 = ( ~n2765 & n15629 ) | ( ~n2765 & n18847 ) | ( n15629 & n18847 ) ;
  assign n22805 = n22804 ^ n17411 ^ n15898 ;
  assign n22806 = ( n1615 & n4128 ) | ( n1615 & n14437 ) | ( n4128 & n14437 ) ;
  assign n22807 = ( n1280 & n6285 ) | ( n1280 & ~n22806 ) | ( n6285 & ~n22806 ) ;
  assign n22808 = n15812 ^ n10970 ^ n4082 ;
  assign n22809 = n7083 ^ n1560 ^ n451 ;
  assign n22810 = n18135 ^ n7955 ^ n348 ;
  assign n22811 = ( n4214 & n4279 ) | ( n4214 & ~n15823 ) | ( n4279 & ~n15823 ) ;
  assign n22812 = n7728 ^ n7475 ^ n4011 ;
  assign n22813 = ( ~n2634 & n5397 ) | ( ~n2634 & n22812 ) | ( n5397 & n22812 ) ;
  assign n22814 = ( n8997 & n9443 ) | ( n8997 & n22813 ) | ( n9443 & n22813 ) ;
  assign n22815 = ( n1197 & n14793 ) | ( n1197 & n22814 ) | ( n14793 & n22814 ) ;
  assign n22819 = n19545 ^ n4820 ^ n1773 ;
  assign n22820 = ( n538 & ~n17490 ) | ( n538 & n22819 ) | ( ~n17490 & n22819 ) ;
  assign n22817 = ( n6923 & n11728 ) | ( n6923 & ~n16785 ) | ( n11728 & ~n16785 ) ;
  assign n22818 = n22817 ^ n15635 ^ n186 ;
  assign n22816 = n17076 ^ n8808 ^ n6994 ;
  assign n22821 = n22820 ^ n22818 ^ n22816 ;
  assign n22822 = ( ~n7397 & n16333 ) | ( ~n7397 & n22821 ) | ( n16333 & n22821 ) ;
  assign n22823 = n13634 ^ n4619 ^ n950 ;
  assign n22824 = ( n8371 & n18343 ) | ( n8371 & ~n22823 ) | ( n18343 & ~n22823 ) ;
  assign n22825 = ( n7018 & ~n13336 ) | ( n7018 & n15509 ) | ( ~n13336 & n15509 ) ;
  assign n22826 = n22825 ^ n12010 ^ n551 ;
  assign n22827 = n7928 ^ n4766 ^ n3148 ;
  assign n22828 = n18531 ^ n12859 ^ n2446 ;
  assign n22829 = ( ~n4204 & n22827 ) | ( ~n4204 & n22828 ) | ( n22827 & n22828 ) ;
  assign n22830 = n18166 ^ n9227 ^ n5488 ;
  assign n22831 = ( n7877 & n14041 ) | ( n7877 & ~n18149 ) | ( n14041 & ~n18149 ) ;
  assign n22832 = ( ~n3097 & n7325 ) | ( ~n3097 & n11041 ) | ( n7325 & n11041 ) ;
  assign n22833 = n6114 ^ n5727 ^ n3247 ;
  assign n22834 = ( n3972 & n6552 ) | ( n3972 & n7322 ) | ( n6552 & n7322 ) ;
  assign n22835 = n22834 ^ n13218 ^ n8252 ;
  assign n22836 = n22835 ^ n8650 ^ n7388 ;
  assign n22837 = ( n5860 & ~n16275 ) | ( n5860 & n22836 ) | ( ~n16275 & n22836 ) ;
  assign n22839 = ( n14808 & ~n18890 ) | ( n14808 & n21532 ) | ( ~n18890 & n21532 ) ;
  assign n22838 = n19604 ^ n18059 ^ n11415 ;
  assign n22840 = n22839 ^ n22838 ^ n12968 ;
  assign n22841 = n22840 ^ n4761 ^ n4469 ;
  assign n22842 = ( n1145 & ~n5982 ) | ( n1145 & n13215 ) | ( ~n5982 & n13215 ) ;
  assign n22843 = ( ~n6143 & n17833 ) | ( ~n6143 & n22842 ) | ( n17833 & n22842 ) ;
  assign n22844 = ( n5839 & ~n7359 ) | ( n5839 & n22843 ) | ( ~n7359 & n22843 ) ;
  assign n22845 = ( n13966 & n17934 ) | ( n13966 & n18366 ) | ( n17934 & n18366 ) ;
  assign n22846 = ( n5885 & ~n14284 ) | ( n5885 & n22540 ) | ( ~n14284 & n22540 ) ;
  assign n22847 = n16095 ^ n10281 ^ n6320 ;
  assign n22848 = ( n2694 & n6036 ) | ( n2694 & ~n22847 ) | ( n6036 & ~n22847 ) ;
  assign n22849 = ( n1553 & n8351 ) | ( n1553 & ~n10266 ) | ( n8351 & ~n10266 ) ;
  assign n22850 = ( n12106 & ~n20967 ) | ( n12106 & n22849 ) | ( ~n20967 & n22849 ) ;
  assign n22851 = n22850 ^ n9768 ^ n3393 ;
  assign n22852 = ( ~n2292 & n4122 ) | ( ~n2292 & n8953 ) | ( n4122 & n8953 ) ;
  assign n22853 = n9139 ^ n8728 ^ n2585 ;
  assign n22854 = ( n3790 & n22852 ) | ( n3790 & n22853 ) | ( n22852 & n22853 ) ;
  assign n22855 = ( n2186 & n7411 ) | ( n2186 & ~n21489 ) | ( n7411 & ~n21489 ) ;
  assign n22856 = ( n4882 & ~n11246 ) | ( n4882 & n12888 ) | ( ~n11246 & n12888 ) ;
  assign n22861 = ( n12289 & n16264 ) | ( n12289 & n21506 ) | ( n16264 & n21506 ) ;
  assign n22862 = ( n10603 & n11000 ) | ( n10603 & ~n22861 ) | ( n11000 & ~n22861 ) ;
  assign n22857 = n9905 ^ n7206 ^ n6645 ;
  assign n22858 = n22857 ^ n6377 ^ n5062 ;
  assign n22859 = n22858 ^ n6487 ^ n1406 ;
  assign n22860 = n22859 ^ n18765 ^ n1266 ;
  assign n22863 = n22862 ^ n22860 ^ n5963 ;
  assign n22864 = ( n1994 & n12876 ) | ( n1994 & ~n13651 ) | ( n12876 & ~n13651 ) ;
  assign n22865 = ( n3238 & n3695 ) | ( n3238 & ~n10660 ) | ( n3695 & ~n10660 ) ;
  assign n22866 = n22865 ^ n16329 ^ n5333 ;
  assign n22867 = n2450 ^ n660 ^ n186 ;
  assign n22868 = ( ~n8565 & n18754 ) | ( ~n8565 & n22867 ) | ( n18754 & n22867 ) ;
  assign n22869 = ( n10151 & n11364 ) | ( n10151 & ~n22868 ) | ( n11364 & ~n22868 ) ;
  assign n22870 = ( n2901 & ~n5105 ) | ( n2901 & n5958 ) | ( ~n5105 & n5958 ) ;
  assign n22871 = ( n11646 & n12318 ) | ( n11646 & ~n22870 ) | ( n12318 & ~n22870 ) ;
  assign n22872 = n22871 ^ n14438 ^ n11401 ;
  assign n22873 = ( ~n3697 & n15779 ) | ( ~n3697 & n22872 ) | ( n15779 & n22872 ) ;
  assign n22874 = ( n4172 & n20973 ) | ( n4172 & ~n22873 ) | ( n20973 & ~n22873 ) ;
  assign n22875 = ( n1860 & n21487 ) | ( n1860 & ~n21685 ) | ( n21487 & ~n21685 ) ;
  assign n22876 = ( n6564 & n16015 ) | ( n6564 & n22875 ) | ( n16015 & n22875 ) ;
  assign n22877 = ( n3230 & n10495 ) | ( n3230 & ~n15933 ) | ( n10495 & ~n15933 ) ;
  assign n22878 = n22877 ^ n7470 ^ n1404 ;
  assign n22879 = ( n6422 & ~n7231 ) | ( n6422 & n10403 ) | ( ~n7231 & n10403 ) ;
  assign n22880 = n22879 ^ n13478 ^ n12795 ;
  assign n22881 = ( n2294 & n3274 ) | ( n2294 & ~n5004 ) | ( n3274 & ~n5004 ) ;
  assign n22882 = ( n4885 & n12096 ) | ( n4885 & n22881 ) | ( n12096 & n22881 ) ;
  assign n22883 = ( n10237 & n11331 ) | ( n10237 & n14995 ) | ( n11331 & n14995 ) ;
  assign n22884 = n18722 ^ n9955 ^ n2797 ;
  assign n22885 = n19962 ^ n17488 ^ n11791 ;
  assign n22886 = ( n8932 & ~n18904 ) | ( n8932 & n19155 ) | ( ~n18904 & n19155 ) ;
  assign n22887 = ( ~n197 & n7763 ) | ( ~n197 & n11722 ) | ( n7763 & n11722 ) ;
  assign n22888 = ( n1079 & n15261 ) | ( n1079 & ~n22887 ) | ( n15261 & ~n22887 ) ;
  assign n22889 = ( n10050 & n11505 ) | ( n10050 & ~n22888 ) | ( n11505 & ~n22888 ) ;
  assign n22890 = ( ~n1128 & n4273 ) | ( ~n1128 & n5700 ) | ( n4273 & n5700 ) ;
  assign n22891 = n22890 ^ n22736 ^ n18650 ;
  assign n22892 = n22891 ^ n6210 ^ n531 ;
  assign n22893 = ( n2174 & n2359 ) | ( n2174 & ~n13990 ) | ( n2359 & ~n13990 ) ;
  assign n22894 = n22893 ^ n6514 ^ n4447 ;
  assign n22895 = ( n1337 & ~n2671 ) | ( n1337 & n22894 ) | ( ~n2671 & n22894 ) ;
  assign n22896 = n21699 ^ n12179 ^ n9434 ;
  assign n22897 = ( n8532 & n9586 ) | ( n8532 & ~n22896 ) | ( n9586 & ~n22896 ) ;
  assign n22898 = n4546 ^ n2752 ^ n1837 ;
  assign n22899 = n22898 ^ n4605 ^ n3367 ;
  assign n22900 = ( n2116 & ~n13599 ) | ( n2116 & n22899 ) | ( ~n13599 & n22899 ) ;
  assign n22901 = ( n14867 & n18271 ) | ( n14867 & ~n21225 ) | ( n18271 & ~n21225 ) ;
  assign n22902 = ( ~n6884 & n12062 ) | ( ~n6884 & n22548 ) | ( n12062 & n22548 ) ;
  assign n22903 = ( n412 & n16204 ) | ( n412 & ~n19467 ) | ( n16204 & ~n19467 ) ;
  assign n22904 = ( n10614 & ~n14979 ) | ( n10614 & n22903 ) | ( ~n14979 & n22903 ) ;
  assign n22907 = n18226 ^ n9523 ^ n5718 ;
  assign n22908 = ( n3154 & n12372 ) | ( n3154 & ~n22907 ) | ( n12372 & ~n22907 ) ;
  assign n22905 = n13912 ^ n6796 ^ n4614 ;
  assign n22906 = ( n10140 & n10294 ) | ( n10140 & n22905 ) | ( n10294 & n22905 ) ;
  assign n22909 = n22908 ^ n22906 ^ n13347 ;
  assign n22910 = n20616 ^ n10144 ^ n2333 ;
  assign n22911 = n22910 ^ n7488 ^ n3658 ;
  assign n22912 = ( n6624 & n18844 ) | ( n6624 & ~n22911 ) | ( n18844 & ~n22911 ) ;
  assign n22913 = ( n16736 & ~n22909 ) | ( n16736 & n22912 ) | ( ~n22909 & n22912 ) ;
  assign n22914 = ( n4520 & n4996 ) | ( n4520 & ~n5668 ) | ( n4996 & ~n5668 ) ;
  assign n22915 = ( n1372 & n16665 ) | ( n1372 & n22914 ) | ( n16665 & n22914 ) ;
  assign n22916 = ( n8625 & n11767 ) | ( n8625 & n22915 ) | ( n11767 & n22915 ) ;
  assign n22917 = n16006 ^ n8997 ^ n1491 ;
  assign n22918 = ( n2750 & n22916 ) | ( n2750 & ~n22917 ) | ( n22916 & ~n22917 ) ;
  assign n22919 = ( n148 & n1622 ) | ( n148 & n3737 ) | ( n1622 & n3737 ) ;
  assign n22920 = ( n3338 & n9418 ) | ( n3338 & ~n22919 ) | ( n9418 & ~n22919 ) ;
  assign n22921 = n22920 ^ n17305 ^ n1792 ;
  assign n22922 = ( ~n1270 & n2195 ) | ( ~n1270 & n6995 ) | ( n2195 & n6995 ) ;
  assign n22923 = n5899 ^ n440 ^ x119 ;
  assign n22924 = ( ~n441 & n2717 ) | ( ~n441 & n7151 ) | ( n2717 & n7151 ) ;
  assign n22925 = ( n977 & n1092 ) | ( n977 & n3937 ) | ( n1092 & n3937 ) ;
  assign n22926 = ( n15028 & n17027 ) | ( n15028 & ~n22925 ) | ( n17027 & ~n22925 ) ;
  assign n22927 = ( n3792 & n21544 ) | ( n3792 & n22926 ) | ( n21544 & n22926 ) ;
  assign n22928 = ( ~n4634 & n7071 ) | ( ~n4634 & n22927 ) | ( n7071 & n22927 ) ;
  assign n22929 = n5920 ^ n1961 ^ n1649 ;
  assign n22930 = ( n9728 & n15219 ) | ( n9728 & ~n20326 ) | ( n15219 & ~n20326 ) ;
  assign n22931 = ( ~n15435 & n21277 ) | ( ~n15435 & n22930 ) | ( n21277 & n22930 ) ;
  assign n22932 = ( n9419 & ~n11719 ) | ( n9419 & n16518 ) | ( ~n11719 & n16518 ) ;
  assign n22933 = n13571 ^ n1043 ^ n829 ;
  assign n22935 = n6771 ^ n2941 ^ n1530 ;
  assign n22934 = ( n3387 & n8026 ) | ( n3387 & ~n14471 ) | ( n8026 & ~n14471 ) ;
  assign n22936 = n22935 ^ n22934 ^ n11193 ;
  assign n22937 = ( n4342 & n11664 ) | ( n4342 & ~n16867 ) | ( n11664 & ~n16867 ) ;
  assign n22939 = n11486 ^ n2338 ^ n670 ;
  assign n22938 = n15772 ^ n611 ^ n231 ;
  assign n22940 = n22939 ^ n22938 ^ n3241 ;
  assign n22941 = n8051 ^ n2448 ^ n319 ;
  assign n22942 = n14094 ^ n6301 ^ n3644 ;
  assign n22943 = ( n20837 & ~n22941 ) | ( n20837 & n22942 ) | ( ~n22941 & n22942 ) ;
  assign n22949 = ( n465 & ~n1550 ) | ( n465 & n7954 ) | ( ~n1550 & n7954 ) ;
  assign n22950 = ( ~n8831 & n12816 ) | ( ~n8831 & n22949 ) | ( n12816 & n22949 ) ;
  assign n22944 = n8914 ^ n4173 ^ n1082 ;
  assign n22945 = n22944 ^ n16642 ^ n4786 ;
  assign n22946 = n21518 ^ n20520 ^ n16871 ;
  assign n22947 = ( ~n358 & n2394 ) | ( ~n358 & n22946 ) | ( n2394 & n22946 ) ;
  assign n22948 = ( n7875 & ~n22945 ) | ( n7875 & n22947 ) | ( ~n22945 & n22947 ) ;
  assign n22951 = n22950 ^ n22948 ^ n13538 ;
  assign n22952 = n18778 ^ n14220 ^ n9204 ;
  assign n22953 = n22503 ^ n21668 ^ n14591 ;
  assign n22954 = n19864 ^ n18936 ^ n16150 ;
  assign n22955 = ( n1559 & n3049 ) | ( n1559 & n5152 ) | ( n3049 & n5152 ) ;
  assign n22956 = ( n4197 & n10806 ) | ( n4197 & n22955 ) | ( n10806 & n22955 ) ;
  assign n22957 = ( ~n2232 & n21476 ) | ( ~n2232 & n22956 ) | ( n21476 & n22956 ) ;
  assign n22958 = n17306 ^ n10628 ^ n5542 ;
  assign n22959 = n6803 ^ n3963 ^ n3127 ;
  assign n22960 = n4001 ^ n1022 ^ n559 ;
  assign n22961 = n22960 ^ n9841 ^ n2205 ;
  assign n22962 = ( ~n10551 & n20031 ) | ( ~n10551 & n22961 ) | ( n20031 & n22961 ) ;
  assign n22963 = n22962 ^ n8058 ^ n793 ;
  assign n22964 = ( ~n3845 & n22959 ) | ( ~n3845 & n22963 ) | ( n22959 & n22963 ) ;
  assign n22965 = n18862 ^ n3381 ^ n1057 ;
  assign n22966 = n22965 ^ n11860 ^ n6081 ;
  assign n22967 = n19287 ^ n11586 ^ n1068 ;
  assign n22976 = n6954 ^ n4360 ^ n4221 ;
  assign n22973 = n10635 ^ n10324 ^ n9477 ;
  assign n22974 = n22973 ^ n12424 ^ n3708 ;
  assign n22971 = ( ~n1235 & n2583 ) | ( ~n1235 & n9881 ) | ( n2583 & n9881 ) ;
  assign n22972 = n22971 ^ n17943 ^ n1588 ;
  assign n22975 = n22974 ^ n22972 ^ n15470 ;
  assign n22968 = ( n2021 & n5081 ) | ( n2021 & ~n7067 ) | ( n5081 & ~n7067 ) ;
  assign n22969 = ( n4519 & n5603 ) | ( n4519 & ~n22968 ) | ( n5603 & ~n22968 ) ;
  assign n22970 = n22969 ^ n17100 ^ n5483 ;
  assign n22977 = n22976 ^ n22975 ^ n22970 ;
  assign n22978 = n18173 ^ n17136 ^ n15476 ;
  assign n22979 = ( n3157 & n5665 ) | ( n3157 & n20029 ) | ( n5665 & n20029 ) ;
  assign n22980 = n22979 ^ n22033 ^ n7520 ;
  assign n22981 = n13656 ^ n9422 ^ n680 ;
  assign n22982 = ( n19545 & ~n22980 ) | ( n19545 & n22981 ) | ( ~n22980 & n22981 ) ;
  assign n22983 = ( ~n1005 & n9151 ) | ( ~n1005 & n14707 ) | ( n9151 & n14707 ) ;
  assign n22984 = n21689 ^ n14374 ^ n568 ;
  assign n22985 = n20361 ^ n2187 ^ n1948 ;
  assign n22987 = ( n190 & n1597 ) | ( n190 & n2303 ) | ( n1597 & n2303 ) ;
  assign n22986 = n21318 ^ n18250 ^ n12040 ;
  assign n22988 = n22987 ^ n22986 ^ n3005 ;
  assign n22989 = ( n2875 & ~n9394 ) | ( n2875 & n15797 ) | ( ~n9394 & n15797 ) ;
  assign n22990 = ( ~n6195 & n7748 ) | ( ~n6195 & n13579 ) | ( n7748 & n13579 ) ;
  assign n22991 = n22990 ^ n10358 ^ n5439 ;
  assign n22992 = n18648 ^ n16927 ^ n10183 ;
  assign n22993 = n22992 ^ n22939 ^ n7214 ;
  assign n22994 = ( n1012 & ~n2079 ) | ( n1012 & n20893 ) | ( ~n2079 & n20893 ) ;
  assign n22995 = n11301 ^ n7523 ^ n1978 ;
  assign n22996 = ( n10787 & n12897 ) | ( n10787 & n16312 ) | ( n12897 & n16312 ) ;
  assign n22997 = ( ~n21677 & n22995 ) | ( ~n21677 & n22996 ) | ( n22995 & n22996 ) ;
  assign n22998 = n21229 ^ n8827 ^ n8755 ;
  assign n22999 = n22998 ^ n19669 ^ n19517 ;
  assign n23000 = n18829 ^ n14499 ^ n822 ;
  assign n23001 = n23000 ^ n12487 ^ n2389 ;
  assign n23002 = n23001 ^ n19684 ^ n6578 ;
  assign n23003 = n21971 ^ n10623 ^ n6883 ;
  assign n23004 = ( ~n5994 & n7832 ) | ( ~n5994 & n23003 ) | ( n7832 & n23003 ) ;
  assign n23005 = n21880 ^ n14181 ^ n8516 ;
  assign n23006 = n15592 ^ n10704 ^ n6082 ;
  assign n23007 = ( ~n3136 & n11098 ) | ( ~n3136 & n23006 ) | ( n11098 & n23006 ) ;
  assign n23008 = ( n3189 & n9558 ) | ( n3189 & ~n12734 ) | ( n9558 & ~n12734 ) ;
  assign n23009 = n23008 ^ n16988 ^ n12153 ;
  assign n23010 = ( n5997 & n6897 ) | ( n5997 & n14187 ) | ( n6897 & n14187 ) ;
  assign n23011 = ( n7170 & n10937 ) | ( n7170 & n23010 ) | ( n10937 & n23010 ) ;
  assign n23012 = n23011 ^ n14386 ^ n12139 ;
  assign n23013 = n23012 ^ n19548 ^ n5405 ;
  assign n23014 = n23013 ^ n1613 ^ n312 ;
  assign n23018 = ( ~n4298 & n4799 ) | ( ~n4298 & n5522 ) | ( n4799 & n5522 ) ;
  assign n23015 = n12651 ^ n9660 ^ n4051 ;
  assign n23016 = ( ~n1000 & n11716 ) | ( ~n1000 & n23015 ) | ( n11716 & n23015 ) ;
  assign n23017 = ( n10293 & ~n22315 ) | ( n10293 & n23016 ) | ( ~n22315 & n23016 ) ;
  assign n23019 = n23018 ^ n23017 ^ n6155 ;
  assign n23020 = n23019 ^ n10858 ^ n8950 ;
  assign n23021 = ( n7186 & n7670 ) | ( n7186 & ~n23020 ) | ( n7670 & ~n23020 ) ;
  assign n23024 = n7530 ^ n5269 ^ n2152 ;
  assign n23022 = n16332 ^ n6097 ^ n5938 ;
  assign n23023 = n23022 ^ n12416 ^ n2748 ;
  assign n23025 = n23024 ^ n23023 ^ n8460 ;
  assign n23026 = ( ~n2184 & n2739 ) | ( ~n2184 & n18193 ) | ( n2739 & n18193 ) ;
  assign n23027 = n23026 ^ n3932 ^ n746 ;
  assign n23028 = n10198 ^ n8148 ^ n2954 ;
  assign n23029 = n23028 ^ n4612 ^ n1804 ;
  assign n23030 = ( n4307 & n21081 ) | ( n4307 & n23029 ) | ( n21081 & n23029 ) ;
  assign n23031 = ( ~n2573 & n10464 ) | ( ~n2573 & n16774 ) | ( n10464 & n16774 ) ;
  assign n23032 = ( n18231 & n18745 ) | ( n18231 & n23031 ) | ( n18745 & n23031 ) ;
  assign n23033 = n23032 ^ n17108 ^ n8936 ;
  assign n23034 = n23033 ^ n18861 ^ n9869 ;
  assign n23036 = n12184 ^ n11503 ^ n5311 ;
  assign n23037 = ( ~n5095 & n10370 ) | ( ~n5095 & n22636 ) | ( n10370 & n22636 ) ;
  assign n23038 = ( ~n9903 & n23036 ) | ( ~n9903 & n23037 ) | ( n23036 & n23037 ) ;
  assign n23035 = n22939 ^ n21114 ^ n4251 ;
  assign n23039 = n23038 ^ n23035 ^ n16414 ;
  assign n23040 = n18224 ^ n2198 ^ n1265 ;
  assign n23042 = n9502 ^ n9064 ^ n996 ;
  assign n23041 = n21209 ^ n6698 ^ n3283 ;
  assign n23043 = n23042 ^ n23041 ^ n20875 ;
  assign n23044 = ( ~n13469 & n14472 ) | ( ~n13469 & n23043 ) | ( n14472 & n23043 ) ;
  assign n23045 = ( n1044 & n4387 ) | ( n1044 & n4840 ) | ( n4387 & n4840 ) ;
  assign n23046 = ( n1475 & ~n17240 ) | ( n1475 & n23045 ) | ( ~n17240 & n23045 ) ;
  assign n23047 = n16929 ^ n16824 ^ n4300 ;
  assign n23048 = n11373 ^ n10948 ^ n1241 ;
  assign n23049 = ( ~n3555 & n9103 ) | ( ~n3555 & n23048 ) | ( n9103 & n23048 ) ;
  assign n23050 = n23049 ^ n12820 ^ n8276 ;
  assign n23051 = ( n6278 & n7700 ) | ( n6278 & ~n10663 ) | ( n7700 & ~n10663 ) ;
  assign n23052 = ( n4154 & ~n9520 ) | ( n4154 & n13153 ) | ( ~n9520 & n13153 ) ;
  assign n23053 = ( n1330 & n23051 ) | ( n1330 & ~n23052 ) | ( n23051 & ~n23052 ) ;
  assign n23054 = ( n17851 & ~n23050 ) | ( n17851 & n23053 ) | ( ~n23050 & n23053 ) ;
  assign n23055 = ( ~n8769 & n9174 ) | ( ~n8769 & n10014 ) | ( n9174 & n10014 ) ;
  assign n23056 = ( n6975 & n15149 ) | ( n6975 & n23055 ) | ( n15149 & n23055 ) ;
  assign n23057 = n7493 ^ n4493 ^ n2926 ;
  assign n23058 = n23057 ^ n9757 ^ n6165 ;
  assign n23059 = ( n2583 & n2749 ) | ( n2583 & n14094 ) | ( n2749 & n14094 ) ;
  assign n23060 = ( n5823 & n8006 ) | ( n5823 & ~n23059 ) | ( n8006 & ~n23059 ) ;
  assign n23061 = ( n560 & ~n973 ) | ( n560 & n9587 ) | ( ~n973 & n9587 ) ;
  assign n23062 = ( n9959 & n12887 ) | ( n9959 & ~n23061 ) | ( n12887 & ~n23061 ) ;
  assign n23063 = ( n17053 & ~n23060 ) | ( n17053 & n23062 ) | ( ~n23060 & n23062 ) ;
  assign n23064 = ( n14734 & n23058 ) | ( n14734 & n23063 ) | ( n23058 & n23063 ) ;
  assign n23065 = ( n7273 & n15348 ) | ( n7273 & ~n22044 ) | ( n15348 & ~n22044 ) ;
  assign n23066 = n13631 ^ n6829 ^ n2694 ;
  assign n23067 = n23066 ^ n5871 ^ n5030 ;
  assign n23068 = n23067 ^ n20577 ^ n2383 ;
  assign n23069 = ( n4214 & n21655 ) | ( n4214 & ~n23068 ) | ( n21655 & ~n23068 ) ;
  assign n23070 = n14296 ^ n7646 ^ n3820 ;
  assign n23071 = n23070 ^ n18843 ^ n17080 ;
  assign n23072 = ( ~n4013 & n6335 ) | ( ~n4013 & n23071 ) | ( n6335 & n23071 ) ;
  assign n23073 = ( ~n2168 & n7729 ) | ( ~n2168 & n17597 ) | ( n7729 & n17597 ) ;
  assign n23074 = n23073 ^ n17062 ^ n247 ;
  assign n23075 = ( n1301 & n4766 ) | ( n1301 & ~n13614 ) | ( n4766 & ~n13614 ) ;
  assign n23076 = ( n1245 & ~n2574 ) | ( n1245 & n19938 ) | ( ~n2574 & n19938 ) ;
  assign n23077 = n23076 ^ n17941 ^ n12629 ;
  assign n23079 = n18570 ^ n4350 ^ n3535 ;
  assign n23080 = ( ~n3088 & n9600 ) | ( ~n3088 & n23079 ) | ( n9600 & n23079 ) ;
  assign n23078 = ( n572 & n16844 ) | ( n572 & n17740 ) | ( n16844 & n17740 ) ;
  assign n23081 = n23080 ^ n23078 ^ n12524 ;
  assign n23082 = n8984 ^ n1851 ^ n274 ;
  assign n23083 = ( n1531 & ~n8233 ) | ( n1531 & n23082 ) | ( ~n8233 & n23082 ) ;
  assign n23086 = ( n3943 & ~n6297 ) | ( n3943 & n14565 ) | ( ~n6297 & n14565 ) ;
  assign n23087 = n23086 ^ n14150 ^ n9637 ;
  assign n23088 = n23087 ^ n22250 ^ n5884 ;
  assign n23089 = n23088 ^ n9321 ^ n4799 ;
  assign n23084 = ( n6123 & ~n9855 ) | ( n6123 & n17470 ) | ( ~n9855 & n17470 ) ;
  assign n23085 = ( ~n8499 & n20132 ) | ( ~n8499 & n23084 ) | ( n20132 & n23084 ) ;
  assign n23090 = n23089 ^ n23085 ^ n1345 ;
  assign n23091 = ( n3055 & n4409 ) | ( n3055 & ~n5101 ) | ( n4409 & ~n5101 ) ;
  assign n23092 = ( ~n3576 & n17076 ) | ( ~n3576 & n23091 ) | ( n17076 & n23091 ) ;
  assign n23093 = ( ~n1275 & n6704 ) | ( ~n1275 & n23092 ) | ( n6704 & n23092 ) ;
  assign n23094 = ( n1805 & ~n8030 ) | ( n1805 & n15312 ) | ( ~n8030 & n15312 ) ;
  assign n23095 = n19885 ^ n13959 ^ n7945 ;
  assign n23096 = n23095 ^ n6515 ^ n2401 ;
  assign n23097 = n8760 ^ n1884 ^ n374 ;
  assign n23098 = n23097 ^ n13776 ^ n12195 ;
  assign n23099 = ( n1659 & n11043 ) | ( n1659 & n11457 ) | ( n11043 & n11457 ) ;
  assign n23100 = ( n296 & ~n11178 ) | ( n296 & n15697 ) | ( ~n11178 & n15697 ) ;
  assign n23101 = ( n2211 & n3935 ) | ( n2211 & ~n23100 ) | ( n3935 & ~n23100 ) ;
  assign n23102 = n17507 ^ n16207 ^ n2046 ;
  assign n23103 = n21848 ^ n9797 ^ n9273 ;
  assign n23104 = ( n13206 & n23102 ) | ( n13206 & ~n23103 ) | ( n23102 & ~n23103 ) ;
  assign n23105 = n11468 ^ n10146 ^ n9136 ;
  assign n23106 = n23105 ^ n6188 ^ n6045 ;
  assign n23107 = n9102 ^ n6880 ^ n6140 ;
  assign n23108 = ( n5920 & n6183 ) | ( n5920 & ~n23107 ) | ( n6183 & ~n23107 ) ;
  assign n23109 = n17648 ^ n8479 ^ n4508 ;
  assign n23110 = n20010 ^ n5472 ^ n3588 ;
  assign n23111 = ( n402 & n14542 ) | ( n402 & ~n23110 ) | ( n14542 & ~n23110 ) ;
  assign n23112 = n23111 ^ n9072 ^ n8407 ;
  assign n23113 = n4662 ^ n4455 ^ n4212 ;
  assign n23115 = ( n8768 & n11038 ) | ( n8768 & n15326 ) | ( n11038 & n15326 ) ;
  assign n23114 = n19083 ^ n14085 ^ x109 ;
  assign n23116 = n23115 ^ n23114 ^ n1397 ;
  assign n23117 = n17955 ^ n9921 ^ n9117 ;
  assign n23118 = n23117 ^ n22057 ^ n7595 ;
  assign n23119 = n6941 ^ n2854 ^ n1040 ;
  assign n23120 = ( n6817 & n15888 ) | ( n6817 & n18209 ) | ( n15888 & n18209 ) ;
  assign n23121 = ( n11684 & ~n23119 ) | ( n11684 & n23120 ) | ( ~n23119 & n23120 ) ;
  assign n23122 = n23121 ^ n17361 ^ n1535 ;
  assign n23123 = ( n1572 & n2230 ) | ( n1572 & n3736 ) | ( n2230 & n3736 ) ;
  assign n23124 = n7846 ^ n7266 ^ n5308 ;
  assign n23125 = n23124 ^ n10050 ^ n7722 ;
  assign n23126 = ( n5856 & ~n23123 ) | ( n5856 & n23125 ) | ( ~n23123 & n23125 ) ;
  assign n23127 = ( ~n8621 & n14463 ) | ( ~n8621 & n17659 ) | ( n14463 & n17659 ) ;
  assign n23128 = n23127 ^ n5605 ^ n3004 ;
  assign n23130 = ( n5197 & ~n11071 ) | ( n5197 & n14094 ) | ( ~n11071 & n14094 ) ;
  assign n23129 = n3317 ^ n1868 ^ n672 ;
  assign n23131 = n23130 ^ n23129 ^ n23042 ;
  assign n23132 = n23131 ^ n11299 ^ n9371 ;
  assign n23133 = ( n8179 & n11413 ) | ( n8179 & ~n16302 ) | ( n11413 & ~n16302 ) ;
  assign n23134 = ( n23128 & n23132 ) | ( n23128 & ~n23133 ) | ( n23132 & ~n23133 ) ;
  assign n23135 = ( n3656 & n8673 ) | ( n3656 & n12070 ) | ( n8673 & n12070 ) ;
  assign n23145 = ( n9911 & n13518 ) | ( n9911 & ~n16572 ) | ( n13518 & ~n16572 ) ;
  assign n23141 = n9642 ^ n2739 ^ n1577 ;
  assign n23142 = n23141 ^ n13682 ^ n8678 ;
  assign n23140 = n16840 ^ n5307 ^ n2287 ;
  assign n23136 = n8507 ^ n1058 ^ x39 ;
  assign n23137 = n20691 ^ n4184 ^ n1670 ;
  assign n23138 = ( ~n212 & n14631 ) | ( ~n212 & n23137 ) | ( n14631 & n23137 ) ;
  assign n23139 = ( n16691 & ~n23136 ) | ( n16691 & n23138 ) | ( ~n23136 & n23138 ) ;
  assign n23143 = n23142 ^ n23140 ^ n23139 ;
  assign n23144 = n23143 ^ n17075 ^ n15751 ;
  assign n23146 = n23145 ^ n23144 ^ n18012 ;
  assign n23147 = n22782 ^ n9885 ^ n669 ;
  assign n23153 = ( ~n4731 & n17703 ) | ( ~n4731 & n18205 ) | ( n17703 & n18205 ) ;
  assign n23150 = n22488 ^ n11228 ^ n415 ;
  assign n23151 = n23150 ^ n17796 ^ n16824 ;
  assign n23148 = n9053 ^ n5570 ^ n2401 ;
  assign n23149 = n23148 ^ n9584 ^ n1821 ;
  assign n23152 = n23151 ^ n23149 ^ n5157 ;
  assign n23154 = n23153 ^ n23152 ^ n17443 ;
  assign n23155 = ( ~n7817 & n15226 ) | ( ~n7817 & n21258 ) | ( n15226 & n21258 ) ;
  assign n23156 = ( ~x50 & n11588 ) | ( ~x50 & n23155 ) | ( n11588 & n23155 ) ;
  assign n23157 = ( n7798 & n10454 ) | ( n7798 & n16416 ) | ( n10454 & n16416 ) ;
  assign n23158 = n23157 ^ n19196 ^ n5645 ;
  assign n23160 = n12631 ^ n7531 ^ n7335 ;
  assign n23161 = n23160 ^ n13057 ^ n4399 ;
  assign n23159 = n18859 ^ n9075 ^ n3606 ;
  assign n23162 = n23161 ^ n23159 ^ n1428 ;
  assign n23163 = ( ~n539 & n6090 ) | ( ~n539 & n21798 ) | ( n6090 & n21798 ) ;
  assign n23164 = n18575 ^ n9124 ^ n218 ;
  assign n23165 = ( n8331 & n21854 ) | ( n8331 & n23164 ) | ( n21854 & n23164 ) ;
  assign n23166 = n12965 ^ n5808 ^ n5054 ;
  assign n23167 = ( n1989 & n6225 ) | ( n1989 & n13938 ) | ( n6225 & n13938 ) ;
  assign n23168 = n23167 ^ n20701 ^ n2769 ;
  assign n23172 = ( n5889 & n13780 ) | ( n5889 & n15377 ) | ( n13780 & n15377 ) ;
  assign n23169 = ( n7076 & n8489 ) | ( n7076 & ~n9443 ) | ( n8489 & ~n9443 ) ;
  assign n23170 = n23169 ^ n8502 ^ n554 ;
  assign n23171 = n23170 ^ n20916 ^ n2051 ;
  assign n23173 = n23172 ^ n23171 ^ n2293 ;
  assign n23174 = n19492 ^ n1216 ^ n324 ;
  assign n23175 = ( x91 & n23173 ) | ( x91 & n23174 ) | ( n23173 & n23174 ) ;
  assign n23176 = ( ~n832 & n4370 ) | ( ~n832 & n23175 ) | ( n4370 & n23175 ) ;
  assign n23177 = n9067 ^ n5616 ^ n3009 ;
  assign n23178 = n23177 ^ n21366 ^ n8674 ;
  assign n23179 = n17335 ^ n11956 ^ n4449 ;
  assign n23180 = ( ~n3929 & n15823 ) | ( ~n3929 & n16545 ) | ( n15823 & n16545 ) ;
  assign n23181 = n23180 ^ n21504 ^ n13220 ;
  assign n23182 = n11699 ^ n10001 ^ n4625 ;
  assign n23183 = ( n4901 & n18488 ) | ( n4901 & n23182 ) | ( n18488 & n23182 ) ;
  assign n23187 = n18699 ^ n11665 ^ n677 ;
  assign n23184 = n17955 ^ n14523 ^ n11574 ;
  assign n23185 = n14804 ^ n6639 ^ n2664 ;
  assign n23186 = ( ~n14501 & n23184 ) | ( ~n14501 & n23185 ) | ( n23184 & n23185 ) ;
  assign n23188 = n23187 ^ n23186 ^ n17383 ;
  assign n23189 = n19066 ^ n15854 ^ n9737 ;
  assign n23190 = ( n2375 & n9165 ) | ( n2375 & n23189 ) | ( n9165 & n23189 ) ;
  assign n23191 = ( x55 & n7272 ) | ( x55 & n14244 ) | ( n7272 & n14244 ) ;
  assign n23194 = n15904 ^ n14202 ^ n2303 ;
  assign n23195 = n18602 ^ n10874 ^ n2466 ;
  assign n23196 = n23195 ^ n16930 ^ n10452 ;
  assign n23197 = n23196 ^ n7270 ^ n1697 ;
  assign n23198 = ( n2695 & n23194 ) | ( n2695 & ~n23197 ) | ( n23194 & ~n23197 ) ;
  assign n23192 = ( n9175 & n17098 ) | ( n9175 & ~n21869 ) | ( n17098 & ~n21869 ) ;
  assign n23193 = ( n8441 & n21852 ) | ( n8441 & n23192 ) | ( n21852 & n23192 ) ;
  assign n23199 = n23198 ^ n23193 ^ n10004 ;
  assign n23200 = ( n1609 & ~n23191 ) | ( n1609 & n23199 ) | ( ~n23191 & n23199 ) ;
  assign n23201 = ( n7734 & n11563 ) | ( n7734 & n23200 ) | ( n11563 & n23200 ) ;
  assign n23202 = ( n1404 & n6947 ) | ( n1404 & n20556 ) | ( n6947 & n20556 ) ;
  assign n23203 = n18269 ^ n8105 ^ n911 ;
  assign n23204 = ( n1965 & n7853 ) | ( n1965 & ~n19671 ) | ( n7853 & ~n19671 ) ;
  assign n23205 = ( n3275 & ~n17501 ) | ( n3275 & n23204 ) | ( ~n17501 & n23204 ) ;
  assign n23206 = ( n10842 & ~n16860 ) | ( n10842 & n20488 ) | ( ~n16860 & n20488 ) ;
  assign n23207 = ( n8337 & ~n16865 ) | ( n8337 & n23206 ) | ( ~n16865 & n23206 ) ;
  assign n23208 = n23207 ^ n10339 ^ n3447 ;
  assign n23209 = n21767 ^ n12552 ^ n2914 ;
  assign n23210 = n15872 ^ n12781 ^ n1216 ;
  assign n23211 = n23210 ^ n8889 ^ n7261 ;
  assign n23212 = ( n3161 & ~n5254 ) | ( n3161 & n6586 ) | ( ~n5254 & n6586 ) ;
  assign n23213 = ( n3893 & n13132 ) | ( n3893 & ~n18970 ) | ( n13132 & ~n18970 ) ;
  assign n23214 = n23213 ^ n16606 ^ n14106 ;
  assign n23215 = n18368 ^ n8316 ^ n6376 ;
  assign n23216 = ( n409 & n11211 ) | ( n409 & n15574 ) | ( n11211 & n15574 ) ;
  assign n23217 = n23216 ^ n20854 ^ n20361 ;
  assign n23218 = n23217 ^ n2921 ^ n2307 ;
  assign n23219 = ( n2487 & n7983 ) | ( n2487 & ~n21492 ) | ( n7983 & ~n21492 ) ;
  assign n23220 = ( n7114 & ~n12407 ) | ( n7114 & n18899 ) | ( ~n12407 & n18899 ) ;
  assign n23221 = ( n15303 & n21373 ) | ( n15303 & ~n23220 ) | ( n21373 & ~n23220 ) ;
  assign n23222 = ( n4213 & n5763 ) | ( n4213 & n18948 ) | ( n5763 & n18948 ) ;
  assign n23223 = n23222 ^ n16585 ^ n9471 ;
  assign n23227 = ( n2502 & n3587 ) | ( n2502 & ~n5217 ) | ( n3587 & ~n5217 ) ;
  assign n23224 = n12918 ^ n2725 ^ n318 ;
  assign n23225 = n23224 ^ n12784 ^ n5298 ;
  assign n23226 = n23225 ^ n16963 ^ n16562 ;
  assign n23228 = n23227 ^ n23226 ^ n7022 ;
  assign n23229 = ( ~n4615 & n10590 ) | ( ~n4615 & n15946 ) | ( n10590 & n15946 ) ;
  assign n23230 = ( n12523 & n17115 ) | ( n12523 & ~n21316 ) | ( n17115 & ~n21316 ) ;
  assign n23231 = n19734 ^ n15169 ^ n10714 ;
  assign n23232 = n13067 ^ n12537 ^ n9666 ;
  assign n23233 = ( n1034 & ~n10788 ) | ( n1034 & n11084 ) | ( ~n10788 & n11084 ) ;
  assign n23234 = n20176 ^ n8318 ^ n8045 ;
  assign n23235 = ( n6084 & ~n23233 ) | ( n6084 & n23234 ) | ( ~n23233 & n23234 ) ;
  assign n23236 = ( n2383 & n8414 ) | ( n2383 & n14252 ) | ( n8414 & n14252 ) ;
  assign n23237 = n23236 ^ n14950 ^ n2089 ;
  assign n23238 = n19892 ^ n12935 ^ n7517 ;
  assign n23239 = ( n1602 & n2284 ) | ( n1602 & ~n21101 ) | ( n2284 & ~n21101 ) ;
  assign n23245 = ( ~n252 & n8955 ) | ( ~n252 & n19866 ) | ( n8955 & n19866 ) ;
  assign n23240 = n14878 ^ n13465 ^ n1485 ;
  assign n23241 = ( ~n5700 & n13894 ) | ( ~n5700 & n23240 ) | ( n13894 & n23240 ) ;
  assign n23242 = n9413 ^ n6928 ^ n4167 ;
  assign n23243 = ( ~n1855 & n18189 ) | ( ~n1855 & n23242 ) | ( n18189 & n23242 ) ;
  assign n23244 = ( n8244 & ~n23241 ) | ( n8244 & n23243 ) | ( ~n23241 & n23243 ) ;
  assign n23246 = n23245 ^ n23244 ^ n4768 ;
  assign n23247 = ( n983 & n16255 ) | ( n983 & n23246 ) | ( n16255 & n23246 ) ;
  assign n23248 = ( n814 & ~n23239 ) | ( n814 & n23247 ) | ( ~n23239 & n23247 ) ;
  assign n23249 = ( ~n14544 & n23238 ) | ( ~n14544 & n23248 ) | ( n23238 & n23248 ) ;
  assign n23253 = n22920 ^ n15886 ^ n636 ;
  assign n23250 = n10060 ^ n9204 ^ n295 ;
  assign n23251 = n23250 ^ n7066 ^ n966 ;
  assign n23252 = n23251 ^ n21799 ^ n1162 ;
  assign n23254 = n23253 ^ n23252 ^ n13380 ;
  assign n23255 = ( n2877 & n12349 ) | ( n2877 & ~n16314 ) | ( n12349 & ~n16314 ) ;
  assign n23256 = n23255 ^ n15900 ^ n3950 ;
  assign n23257 = n23256 ^ n19661 ^ n15175 ;
  assign n23258 = n23257 ^ n17773 ^ n13363 ;
  assign n23259 = ( n592 & ~n663 ) | ( n592 & n4556 ) | ( ~n663 & n4556 ) ;
  assign n23260 = n15261 ^ n14912 ^ n11319 ;
  assign n23261 = n23260 ^ n19681 ^ n265 ;
  assign n23262 = ( n16423 & n23259 ) | ( n16423 & ~n23261 ) | ( n23259 & ~n23261 ) ;
  assign n23263 = n11887 ^ n4866 ^ n279 ;
  assign n23264 = ( n18251 & n19813 ) | ( n18251 & ~n23263 ) | ( n19813 & ~n23263 ) ;
  assign n23266 = ( ~n2047 & n5739 ) | ( ~n2047 & n8680 ) | ( n5739 & n8680 ) ;
  assign n23265 = n17573 ^ n15956 ^ n7148 ;
  assign n23267 = n23266 ^ n23265 ^ n16127 ;
  assign n23268 = n8778 ^ n5193 ^ n4659 ;
  assign n23269 = ( n9444 & n12839 ) | ( n9444 & n23268 ) | ( n12839 & n23268 ) ;
  assign n23270 = n23269 ^ n5824 ^ n5344 ;
  assign n23272 = n23182 ^ n13026 ^ n3715 ;
  assign n23273 = ( ~n19066 & n19469 ) | ( ~n19066 & n23272 ) | ( n19469 & n23272 ) ;
  assign n23271 = ( n9750 & n12340 ) | ( n9750 & ~n13684 ) | ( n12340 & ~n13684 ) ;
  assign n23274 = n23273 ^ n23271 ^ n195 ;
  assign n23275 = ( n426 & ~n7897 ) | ( n426 & n9196 ) | ( ~n7897 & n9196 ) ;
  assign n23276 = ( n5545 & ~n7999 ) | ( n5545 & n23275 ) | ( ~n7999 & n23275 ) ;
  assign n23277 = n23276 ^ n10948 ^ n8207 ;
  assign n23278 = ( n3528 & ~n10614 ) | ( n3528 & n11134 ) | ( ~n10614 & n11134 ) ;
  assign n23279 = n23278 ^ n22987 ^ n15513 ;
  assign n23280 = n17056 ^ n12918 ^ n7095 ;
  assign n23281 = n23280 ^ n17829 ^ n8803 ;
  assign n23282 = n9942 ^ n8754 ^ n2032 ;
  assign n23283 = n23282 ^ n17496 ^ n6001 ;
  assign n23284 = n19970 ^ n5218 ^ n584 ;
  assign n23285 = ( n6417 & n13862 ) | ( n6417 & n16858 ) | ( n13862 & n16858 ) ;
  assign n23292 = ( n1703 & n8898 ) | ( n1703 & n14613 ) | ( n8898 & n14613 ) ;
  assign n23293 = n23292 ^ n17486 ^ n8773 ;
  assign n23291 = ( n7340 & n13344 ) | ( n7340 & n18605 ) | ( n13344 & n18605 ) ;
  assign n23286 = ( n6001 & n9131 ) | ( n6001 & ~n9681 ) | ( n9131 & ~n9681 ) ;
  assign n23288 = ( ~n1459 & n2968 ) | ( ~n1459 & n7537 ) | ( n2968 & n7537 ) ;
  assign n23287 = n10512 ^ n5613 ^ n285 ;
  assign n23289 = n23288 ^ n23287 ^ n21246 ;
  assign n23290 = ( n12817 & n23286 ) | ( n12817 & ~n23289 ) | ( n23286 & ~n23289 ) ;
  assign n23294 = n23293 ^ n23291 ^ n23290 ;
  assign n23295 = n15994 ^ n12287 ^ n8303 ;
  assign n23296 = ( n8463 & ~n9597 ) | ( n8463 & n9982 ) | ( ~n9597 & n9982 ) ;
  assign n23297 = ( n4385 & ~n5901 ) | ( n4385 & n23296 ) | ( ~n5901 & n23296 ) ;
  assign n23298 = ( n609 & n2637 ) | ( n609 & ~n9595 ) | ( n2637 & ~n9595 ) ;
  assign n23299 = n23298 ^ n5937 ^ n4259 ;
  assign n23300 = ( n165 & ~n3884 ) | ( n165 & n8448 ) | ( ~n3884 & n8448 ) ;
  assign n23301 = ( n18838 & ~n23299 ) | ( n18838 & n23300 ) | ( ~n23299 & n23300 ) ;
  assign n23302 = ( n472 & ~n3492 ) | ( n472 & n21095 ) | ( ~n3492 & n21095 ) ;
  assign n23303 = n22920 ^ n21624 ^ n11327 ;
  assign n23304 = ( n9386 & n18884 ) | ( n9386 & n23303 ) | ( n18884 & n23303 ) ;
  assign n23305 = n23304 ^ n20694 ^ n9811 ;
  assign n23306 = ( n7255 & n15508 ) | ( n7255 & ~n16078 ) | ( n15508 & ~n16078 ) ;
  assign n23307 = n11884 ^ n10320 ^ n7732 ;
  assign n23308 = n18801 ^ n2283 ^ n496 ;
  assign n23309 = ( ~n8792 & n8884 ) | ( ~n8792 & n23308 ) | ( n8884 & n23308 ) ;
  assign n23310 = n15903 ^ n6371 ^ n5105 ;
  assign n23311 = ( n8178 & n12342 ) | ( n8178 & ~n13218 ) | ( n12342 & ~n13218 ) ;
  assign n23313 = ( ~n2434 & n5287 ) | ( ~n2434 & n6136 ) | ( n5287 & n6136 ) ;
  assign n23314 = ( n4209 & n21101 ) | ( n4209 & n23313 ) | ( n21101 & n23313 ) ;
  assign n23312 = n13927 ^ n9442 ^ n9001 ;
  assign n23315 = n23314 ^ n23312 ^ n3860 ;
  assign n23316 = ( n9415 & ~n17618 ) | ( n9415 & n23315 ) | ( ~n17618 & n23315 ) ;
  assign n23317 = ( ~n23310 & n23311 ) | ( ~n23310 & n23316 ) | ( n23311 & n23316 ) ;
  assign n23318 = n22104 ^ n5694 ^ n3340 ;
  assign n23319 = n16055 ^ n12909 ^ n4492 ;
  assign n23321 = n10552 ^ n4664 ^ n2208 ;
  assign n23320 = ( n2285 & ~n12635 ) | ( n2285 & n14365 ) | ( ~n12635 & n14365 ) ;
  assign n23322 = n23321 ^ n23320 ^ n7843 ;
  assign n23323 = ( n225 & n1123 ) | ( n225 & ~n3049 ) | ( n1123 & ~n3049 ) ;
  assign n23324 = ( n15926 & n17976 ) | ( n15926 & n23323 ) | ( n17976 & n23323 ) ;
  assign n23325 = ( n13214 & n15040 ) | ( n13214 & n23324 ) | ( n15040 & n23324 ) ;
  assign n23326 = ( n1025 & n6023 ) | ( n1025 & ~n23325 ) | ( n6023 & ~n23325 ) ;
  assign n23327 = ( n21131 & n23322 ) | ( n21131 & n23326 ) | ( n23322 & n23326 ) ;
  assign n23328 = ( ~n2964 & n4892 ) | ( ~n2964 & n19939 ) | ( n4892 & n19939 ) ;
  assign n23329 = n7429 ^ n2969 ^ n2345 ;
  assign n23330 = n16572 ^ n7365 ^ n2156 ;
  assign n23331 = ( n3311 & n4703 ) | ( n3311 & ~n23330 ) | ( n4703 & ~n23330 ) ;
  assign n23332 = ( n19007 & n23329 ) | ( n19007 & ~n23331 ) | ( n23329 & ~n23331 ) ;
  assign n23336 = ( n802 & n8285 ) | ( n802 & n9518 ) | ( n8285 & n9518 ) ;
  assign n23333 = n7077 ^ n6711 ^ n5689 ;
  assign n23334 = n23333 ^ n20927 ^ n11415 ;
  assign n23335 = n23334 ^ n6009 ^ n1245 ;
  assign n23337 = n23336 ^ n23335 ^ n22677 ;
  assign n23342 = n14562 ^ n6817 ^ n5136 ;
  assign n23339 = ( ~x11 & n515 ) | ( ~x11 & n9366 ) | ( n515 & n9366 ) ;
  assign n23340 = ( ~n4347 & n6947 ) | ( ~n4347 & n23339 ) | ( n6947 & n23339 ) ;
  assign n23338 = n16398 ^ n13426 ^ n9750 ;
  assign n23341 = n23340 ^ n23338 ^ n7411 ;
  assign n23343 = n23342 ^ n23341 ^ n22642 ;
  assign n23344 = ( n11830 & ~n15742 ) | ( n11830 & n17325 ) | ( ~n15742 & n17325 ) ;
  assign n23345 = n4920 ^ n3478 ^ n429 ;
  assign n23346 = ( n13649 & n14981 ) | ( n13649 & ~n23345 ) | ( n14981 & ~n23345 ) ;
  assign n23349 = n14034 ^ n3007 ^ n2743 ;
  assign n23350 = n23349 ^ n13356 ^ n2219 ;
  assign n23348 = ( n4931 & n12784 ) | ( n4931 & ~n17176 ) | ( n12784 & ~n17176 ) ;
  assign n23347 = n12937 ^ n10482 ^ n2071 ;
  assign n23351 = n23350 ^ n23348 ^ n23347 ;
  assign n23352 = ( n2170 & n4794 ) | ( n2170 & ~n23351 ) | ( n4794 & ~n23351 ) ;
  assign n23353 = n20306 ^ n8986 ^ n571 ;
  assign n23357 = ( x68 & n7609 ) | ( x68 & ~n14584 ) | ( n7609 & ~n14584 ) ;
  assign n23356 = ( ~n2028 & n4680 ) | ( ~n2028 & n6397 ) | ( n4680 & n6397 ) ;
  assign n23354 = ( n7897 & n14750 ) | ( n7897 & n15553 ) | ( n14750 & n15553 ) ;
  assign n23355 = ( n2911 & n18262 ) | ( n2911 & n23354 ) | ( n18262 & n23354 ) ;
  assign n23358 = n23357 ^ n23356 ^ n23355 ;
  assign n23359 = n22052 ^ n2598 ^ n630 ;
  assign n23360 = n19815 ^ n9712 ^ n7009 ;
  assign n23361 = ( n20944 & n23359 ) | ( n20944 & ~n23360 ) | ( n23359 & ~n23360 ) ;
  assign n23362 = n17635 ^ n5293 ^ n563 ;
  assign n23363 = n22644 ^ n18496 ^ n13228 ;
  assign n23364 = ( n18498 & ~n23362 ) | ( n18498 & n23363 ) | ( ~n23362 & n23363 ) ;
  assign n23365 = n10447 ^ n8523 ^ n1997 ;
  assign n23366 = ( ~n13869 & n16633 ) | ( ~n13869 & n23365 ) | ( n16633 & n23365 ) ;
  assign n23367 = n22769 ^ n8697 ^ x29 ;
  assign n23368 = ( x46 & n13402 ) | ( x46 & n19372 ) | ( n13402 & n19372 ) ;
  assign n23369 = ( n645 & n7028 ) | ( n645 & ~n23368 ) | ( n7028 & ~n23368 ) ;
  assign n23370 = ( n1880 & n7607 ) | ( n1880 & ~n17213 ) | ( n7607 & ~n17213 ) ;
  assign n23371 = ( n868 & ~n9263 ) | ( n868 & n23370 ) | ( ~n9263 & n23370 ) ;
  assign n23372 = ( ~n2722 & n10764 ) | ( ~n2722 & n23371 ) | ( n10764 & n23371 ) ;
  assign n23373 = n14071 ^ n3248 ^ n1834 ;
  assign n23374 = ( n3571 & ~n6882 ) | ( n3571 & n23373 ) | ( ~n6882 & n23373 ) ;
  assign n23376 = n16240 ^ n5590 ^ n622 ;
  assign n23375 = n16370 ^ n15953 ^ n7836 ;
  assign n23377 = n23376 ^ n23375 ^ n19552 ;
  assign n23379 = ( n399 & n3821 ) | ( n399 & n13061 ) | ( n3821 & n13061 ) ;
  assign n23378 = n16366 ^ n12475 ^ n3191 ;
  assign n23380 = n23379 ^ n23378 ^ n22916 ;
  assign n23381 = n2202 ^ n1754 ^ n463 ;
  assign n23382 = n23381 ^ n19897 ^ n4450 ;
  assign n23383 = n15964 ^ n11707 ^ n9524 ;
  assign n23384 = n23383 ^ n13563 ^ n11452 ;
  assign n23385 = n8532 ^ n7136 ^ n3943 ;
  assign n23386 = ( n4689 & n14034 ) | ( n4689 & n19931 ) | ( n14034 & n19931 ) ;
  assign n23387 = n18499 ^ n12036 ^ n10152 ;
  assign n23388 = ( n15383 & n17930 ) | ( n15383 & ~n23387 ) | ( n17930 & ~n23387 ) ;
  assign n23389 = n23388 ^ n10836 ^ n2276 ;
  assign n23390 = ( n21147 & n22432 ) | ( n21147 & ~n23389 ) | ( n22432 & ~n23389 ) ;
  assign n23391 = n23390 ^ n11021 ^ n3688 ;
  assign n23396 = ( n2757 & n6792 ) | ( n2757 & ~n8087 ) | ( n6792 & ~n8087 ) ;
  assign n23394 = n7371 ^ n2886 ^ n627 ;
  assign n23395 = ( n6788 & n11098 ) | ( n6788 & n23394 ) | ( n11098 & n23394 ) ;
  assign n23392 = ( ~n839 & n2318 ) | ( ~n839 & n3304 ) | ( n2318 & n3304 ) ;
  assign n23393 = n23392 ^ n13523 ^ n12374 ;
  assign n23397 = n23396 ^ n23395 ^ n23393 ;
  assign n23398 = ( n15554 & n20136 ) | ( n15554 & n20620 ) | ( n20136 & n20620 ) ;
  assign n23399 = ( ~n1697 & n2946 ) | ( ~n1697 & n8555 ) | ( n2946 & n8555 ) ;
  assign n23400 = ( ~n793 & n7812 ) | ( ~n793 & n19631 ) | ( n7812 & n19631 ) ;
  assign n23401 = ( ~n1081 & n18116 ) | ( ~n1081 & n23400 ) | ( n18116 & n23400 ) ;
  assign n23402 = ( n14537 & ~n23399 ) | ( n14537 & n23401 ) | ( ~n23399 & n23401 ) ;
  assign n23403 = n15415 ^ n9768 ^ n6670 ;
  assign n23407 = ( n3019 & n7601 ) | ( n3019 & ~n13891 ) | ( n7601 & ~n13891 ) ;
  assign n23408 = ( ~n4114 & n5954 ) | ( ~n4114 & n23407 ) | ( n5954 & n23407 ) ;
  assign n23409 = n23408 ^ n5733 ^ n2748 ;
  assign n23404 = ( n4088 & n6166 ) | ( n4088 & ~n14534 ) | ( n6166 & ~n14534 ) ;
  assign n23405 = ( n394 & ~n17383 ) | ( n394 & n23404 ) | ( ~n17383 & n23404 ) ;
  assign n23406 = ( ~n4852 & n19863 ) | ( ~n4852 & n23405 ) | ( n19863 & n23405 ) ;
  assign n23410 = n23409 ^ n23406 ^ n10553 ;
  assign n23411 = ( n1120 & n5513 ) | ( n1120 & n17349 ) | ( n5513 & n17349 ) ;
  assign n23412 = n23411 ^ n13089 ^ n6822 ;
  assign n23413 = n17731 ^ n15979 ^ n3779 ;
  assign n23414 = ( ~n7556 & n9965 ) | ( ~n7556 & n21393 ) | ( n9965 & n21393 ) ;
  assign n23415 = ( n1162 & ~n4025 ) | ( n1162 & n13180 ) | ( ~n4025 & n13180 ) ;
  assign n23416 = n23415 ^ n13459 ^ n2164 ;
  assign n23417 = ( n423 & n8717 ) | ( n423 & ~n18120 ) | ( n8717 & ~n18120 ) ;
  assign n23423 = ( x12 & n1405 ) | ( x12 & n3614 ) | ( n1405 & n3614 ) ;
  assign n23424 = ( n3691 & n5402 ) | ( n3691 & n23423 ) | ( n5402 & n23423 ) ;
  assign n23421 = ( n305 & ~n1316 ) | ( n305 & n5312 ) | ( ~n1316 & n5312 ) ;
  assign n23419 = ( ~n1971 & n4936 ) | ( ~n1971 & n5076 ) | ( n4936 & n5076 ) ;
  assign n23418 = ( n4374 & n10320 ) | ( n4374 & n17744 ) | ( n10320 & n17744 ) ;
  assign n23420 = n23419 ^ n23418 ^ n20051 ;
  assign n23422 = n23421 ^ n23420 ^ n12835 ;
  assign n23425 = n23424 ^ n23422 ^ n20065 ;
  assign n23426 = ( n2329 & n11703 ) | ( n2329 & ~n21019 ) | ( n11703 & ~n21019 ) ;
  assign n23427 = ( n1357 & n21168 ) | ( n1357 & ~n23426 ) | ( n21168 & ~n23426 ) ;
  assign n23428 = n10554 ^ n4021 ^ n2606 ;
  assign n23429 = n23428 ^ n15869 ^ n2061 ;
  assign n23430 = n20071 ^ n17604 ^ n12147 ;
  assign n23431 = n10606 ^ n5151 ^ n2670 ;
  assign n23432 = n23431 ^ n16831 ^ n4724 ;
  assign n23433 = ( n3806 & ~n10499 ) | ( n3806 & n13114 ) | ( ~n10499 & n13114 ) ;
  assign n23434 = ( n1223 & ~n9194 ) | ( n1223 & n23433 ) | ( ~n9194 & n23433 ) ;
  assign n23435 = ( n14911 & n15172 ) | ( n14911 & n23434 ) | ( n15172 & n23434 ) ;
  assign n23436 = n23435 ^ n19493 ^ n12853 ;
  assign n23437 = n10450 ^ n4888 ^ n4254 ;
  assign n23439 = ( n8049 & n8566 ) | ( n8049 & n19347 ) | ( n8566 & n19347 ) ;
  assign n23438 = n16109 ^ n13612 ^ n7494 ;
  assign n23440 = n23439 ^ n23438 ^ n18489 ;
  assign n23441 = ( n1280 & n5937 ) | ( n1280 & n14945 ) | ( n5937 & n14945 ) ;
  assign n23442 = n23441 ^ n18298 ^ n12481 ;
  assign n23443 = ( n7225 & n11282 ) | ( n7225 & n11283 ) | ( n11282 & n11283 ) ;
  assign n23444 = n23443 ^ n19511 ^ n9990 ;
  assign n23445 = n23444 ^ n22376 ^ n4095 ;
  assign n23446 = n12396 ^ n10471 ^ n10023 ;
  assign n23447 = ( ~n738 & n6392 ) | ( ~n738 & n18778 ) | ( n6392 & n18778 ) ;
  assign n23448 = ( ~n1860 & n8664 ) | ( ~n1860 & n23447 ) | ( n8664 & n23447 ) ;
  assign n23449 = n22663 ^ n22602 ^ n9607 ;
  assign n23450 = ( n15097 & ~n23448 ) | ( n15097 & n23449 ) | ( ~n23448 & n23449 ) ;
  assign n23451 = n8242 ^ n4778 ^ n3098 ;
  assign n23452 = ( n1935 & n5513 ) | ( n1935 & ~n23451 ) | ( n5513 & ~n23451 ) ;
  assign n23453 = n11990 ^ n6063 ^ n4855 ;
  assign n23454 = ( n4012 & ~n5615 ) | ( n4012 & n23453 ) | ( ~n5615 & n23453 ) ;
  assign n23455 = ( n6698 & n23452 ) | ( n6698 & ~n23454 ) | ( n23452 & ~n23454 ) ;
  assign n23460 = n12130 ^ n9070 ^ n3902 ;
  assign n23457 = ( n3870 & n6107 ) | ( n3870 & ~n6450 ) | ( n6107 & ~n6450 ) ;
  assign n23458 = ( n1989 & ~n15653 ) | ( n1989 & n23457 ) | ( ~n15653 & n23457 ) ;
  assign n23456 = ( n10232 & n18090 ) | ( n10232 & ~n22812 ) | ( n18090 & ~n22812 ) ;
  assign n23459 = n23458 ^ n23456 ^ n9398 ;
  assign n23461 = n23460 ^ n23459 ^ n10687 ;
  assign n23462 = n19995 ^ n6433 ^ n1681 ;
  assign n23463 = n6075 ^ n5522 ^ n2280 ;
  assign n23464 = n23463 ^ n20030 ^ n10211 ;
  assign n23465 = n5696 ^ n4869 ^ n2868 ;
  assign n23466 = n23465 ^ n21537 ^ n15505 ;
  assign n23467 = ( n6351 & n23464 ) | ( n6351 & ~n23466 ) | ( n23464 & ~n23466 ) ;
  assign n23468 = ( n12559 & n14881 ) | ( n12559 & n23467 ) | ( n14881 & n23467 ) ;
  assign n23469 = ( n14320 & n21895 ) | ( n14320 & ~n23468 ) | ( n21895 & ~n23468 ) ;
  assign n23470 = n22868 ^ n5109 ^ n2664 ;
  assign n23471 = ( ~n23462 & n23469 ) | ( ~n23462 & n23470 ) | ( n23469 & n23470 ) ;
  assign n23472 = n11928 ^ n3000 ^ n527 ;
  assign n23473 = n23472 ^ n15452 ^ n6269 ;
  assign n23474 = n23473 ^ n16063 ^ n5830 ;
  assign n23475 = n23474 ^ n17062 ^ n11402 ;
  assign n23476 = ( n2801 & ~n7420 ) | ( n2801 & n11520 ) | ( ~n7420 & n11520 ) ;
  assign n23477 = n14819 ^ n12915 ^ n6586 ;
  assign n23478 = ( n738 & n2553 ) | ( n738 & n13218 ) | ( n2553 & n13218 ) ;
  assign n23479 = ( n12360 & n16617 ) | ( n12360 & ~n23478 ) | ( n16617 & ~n23478 ) ;
  assign n23480 = ( x0 & n5241 ) | ( x0 & ~n10165 ) | ( n5241 & ~n10165 ) ;
  assign n23481 = n11366 ^ n8825 ^ n5485 ;
  assign n23482 = n23481 ^ n2094 ^ n756 ;
  assign n23483 = n16822 ^ n13641 ^ n1587 ;
  assign n23484 = n11660 ^ n5125 ^ n910 ;
  assign n23485 = ( n7248 & n18441 ) | ( n7248 & n23484 ) | ( n18441 & n23484 ) ;
  assign n23486 = ( n22215 & n23483 ) | ( n22215 & ~n23485 ) | ( n23483 & ~n23485 ) ;
  assign n23487 = ( n4396 & n7386 ) | ( n4396 & n11725 ) | ( n7386 & n11725 ) ;
  assign n23488 = ( ~n4023 & n20790 ) | ( ~n4023 & n22262 ) | ( n20790 & n22262 ) ;
  assign n23489 = n13801 ^ n2584 ^ n1688 ;
  assign n23490 = ( n761 & ~n12132 ) | ( n761 & n23489 ) | ( ~n12132 & n23489 ) ;
  assign n23491 = n23490 ^ n2214 ^ x90 ;
  assign n23492 = ( n5574 & ~n8389 ) | ( n5574 & n12102 ) | ( ~n8389 & n12102 ) ;
  assign n23493 = ( n2221 & n3401 ) | ( n2221 & n23492 ) | ( n3401 & n23492 ) ;
  assign n23494 = n17883 ^ n3388 ^ x4 ;
  assign n23495 = ( n10534 & ~n20143 ) | ( n10534 & n23494 ) | ( ~n20143 & n23494 ) ;
  assign n23496 = n23495 ^ n14864 ^ n1624 ;
  assign n23499 = n17935 ^ n13465 ^ n7426 ;
  assign n23500 = ( n1515 & n4489 ) | ( n1515 & ~n23499 ) | ( n4489 & ~n23499 ) ;
  assign n23497 = n9754 ^ n8390 ^ n2448 ;
  assign n23498 = ( n9201 & n18541 ) | ( n9201 & ~n23497 ) | ( n18541 & ~n23497 ) ;
  assign n23501 = n23500 ^ n23498 ^ n8543 ;
  assign n23502 = ( ~n14612 & n16281 ) | ( ~n14612 & n18637 ) | ( n16281 & n18637 ) ;
  assign n23503 = ( n8113 & n17903 ) | ( n8113 & n23502 ) | ( n17903 & n23502 ) ;
  assign n23504 = n19803 ^ n11981 ^ n11410 ;
  assign n23506 = ( n2239 & n18339 ) | ( n2239 & n19227 ) | ( n18339 & n19227 ) ;
  assign n23505 = n10339 ^ n4087 ^ n3396 ;
  assign n23507 = n23506 ^ n23505 ^ n5468 ;
  assign n23508 = n21099 ^ n14392 ^ n6972 ;
  assign n23509 = ( n1516 & n13010 ) | ( n1516 & ~n18590 ) | ( n13010 & ~n18590 ) ;
  assign n23510 = n11737 ^ n8598 ^ n6725 ;
  assign n23511 = n23510 ^ n11599 ^ n158 ;
  assign n23512 = n23511 ^ n17322 ^ n4067 ;
  assign n23513 = n22946 ^ n7502 ^ n227 ;
  assign n23514 = ( n5079 & n6822 ) | ( n5079 & n6929 ) | ( n6822 & n6929 ) ;
  assign n23515 = ( n2160 & n2411 ) | ( n2160 & n5428 ) | ( n2411 & n5428 ) ;
  assign n23516 = n14804 ^ n10031 ^ n3239 ;
  assign n23517 = ( n2071 & n23515 ) | ( n2071 & ~n23516 ) | ( n23515 & ~n23516 ) ;
  assign n23518 = n8517 ^ n4312 ^ n1589 ;
  assign n23523 = ( n1565 & n2699 ) | ( n1565 & n3259 ) | ( n2699 & n3259 ) ;
  assign n23520 = ( n2290 & n3374 ) | ( n2290 & n10003 ) | ( n3374 & n10003 ) ;
  assign n23521 = ( n12137 & n12810 ) | ( n12137 & ~n20728 ) | ( n12810 & ~n20728 ) ;
  assign n23522 = ( n15188 & n23520 ) | ( n15188 & n23521 ) | ( n23520 & n23521 ) ;
  assign n23519 = ( n8415 & n10438 ) | ( n8415 & n12549 ) | ( n10438 & n12549 ) ;
  assign n23524 = n23523 ^ n23522 ^ n23519 ;
  assign n23525 = ( n9175 & n10231 ) | ( n9175 & ~n18637 ) | ( n10231 & ~n18637 ) ;
  assign n23526 = ( n1555 & ~n9169 ) | ( n1555 & n20451 ) | ( ~n9169 & n20451 ) ;
  assign n23527 = ( ~n3701 & n23525 ) | ( ~n3701 & n23526 ) | ( n23525 & n23526 ) ;
  assign n23528 = ( n3657 & n8318 ) | ( n3657 & ~n10463 ) | ( n8318 & ~n10463 ) ;
  assign n23529 = ( n1342 & n2464 ) | ( n1342 & n11280 ) | ( n2464 & n11280 ) ;
  assign n23530 = n12800 ^ n10781 ^ n3247 ;
  assign n23531 = n23530 ^ n19110 ^ n4227 ;
  assign n23532 = n23531 ^ n13831 ^ n3667 ;
  assign n23533 = ( n951 & ~n1763 ) | ( n951 & n11505 ) | ( ~n1763 & n11505 ) ;
  assign n23534 = n23533 ^ n18814 ^ n5350 ;
  assign n23535 = ( n1507 & ~n23532 ) | ( n1507 & n23534 ) | ( ~n23532 & n23534 ) ;
  assign n23537 = ( ~n11308 & n12357 ) | ( ~n11308 & n17245 ) | ( n12357 & n17245 ) ;
  assign n23536 = n23015 ^ n18090 ^ n10436 ;
  assign n23538 = n23537 ^ n23536 ^ n15548 ;
  assign n23539 = ( ~n365 & n4126 ) | ( ~n365 & n9060 ) | ( n4126 & n9060 ) ;
  assign n23540 = ( ~n11050 & n11290 ) | ( ~n11050 & n11449 ) | ( n11290 & n11449 ) ;
  assign n23541 = ( n3371 & n23539 ) | ( n3371 & n23540 ) | ( n23539 & n23540 ) ;
  assign n23542 = ( ~n4269 & n6333 ) | ( ~n4269 & n23541 ) | ( n6333 & n23541 ) ;
  assign n23543 = ( n2875 & n12712 ) | ( n2875 & n18655 ) | ( n12712 & n18655 ) ;
  assign n23544 = ( n1132 & n2609 ) | ( n1132 & ~n23543 ) | ( n2609 & ~n23543 ) ;
  assign n23545 = ( ~n3409 & n4732 ) | ( ~n3409 & n20019 ) | ( n4732 & n20019 ) ;
  assign n23546 = n23545 ^ n12566 ^ n2458 ;
  assign n23547 = ( n8447 & n13334 ) | ( n8447 & ~n14833 ) | ( n13334 & ~n14833 ) ;
  assign n23548 = n17056 ^ n13884 ^ n10013 ;
  assign n23549 = n7663 ^ n673 ^ n170 ;
  assign n23550 = ( n6412 & n9228 ) | ( n6412 & ~n23549 ) | ( n9228 & ~n23549 ) ;
  assign n23551 = n23550 ^ n23499 ^ n449 ;
  assign n23552 = ( ~n3675 & n4035 ) | ( ~n3675 & n15544 ) | ( n4035 & n15544 ) ;
  assign n23553 = n23552 ^ n20645 ^ n4804 ;
  assign n23554 = n19147 ^ n15806 ^ n1286 ;
  assign n23555 = n23554 ^ n19113 ^ n9794 ;
  assign n23556 = n15695 ^ n13109 ^ n9116 ;
  assign n23557 = n19350 ^ n7976 ^ n7681 ;
  assign n23558 = ( ~n2330 & n20263 ) | ( ~n2330 & n23557 ) | ( n20263 & n23557 ) ;
  assign n23559 = n23558 ^ n17226 ^ n12557 ;
  assign n23560 = n23559 ^ n6681 ^ n2923 ;
  assign n23563 = n8984 ^ n7701 ^ n4675 ;
  assign n23561 = ( ~n2632 & n10175 ) | ( ~n2632 & n20295 ) | ( n10175 & n20295 ) ;
  assign n23562 = n23561 ^ n8556 ^ n5745 ;
  assign n23564 = n23563 ^ n23562 ^ n14537 ;
  assign n23565 = ( ~n6484 & n7466 ) | ( ~n6484 & n23564 ) | ( n7466 & n23564 ) ;
  assign n23566 = n9501 ^ n5795 ^ n4107 ;
  assign n23567 = ( n5761 & n10124 ) | ( n5761 & ~n23566 ) | ( n10124 & ~n23566 ) ;
  assign n23569 = n5294 ^ n3549 ^ n1599 ;
  assign n23570 = ( n4109 & n7753 ) | ( n4109 & n23569 ) | ( n7753 & n23569 ) ;
  assign n23568 = n21800 ^ n15179 ^ n14146 ;
  assign n23571 = n23570 ^ n23568 ^ n11749 ;
  assign n23572 = ( n13233 & ~n20588 ) | ( n13233 & n22097 ) | ( ~n20588 & n22097 ) ;
  assign n23573 = ( n2459 & n15239 ) | ( n2459 & n23572 ) | ( n15239 & n23572 ) ;
  assign n23574 = n23573 ^ n6487 ^ n3829 ;
  assign n23575 = n12815 ^ n6322 ^ n3098 ;
  assign n23576 = ( ~n2516 & n6649 ) | ( ~n2516 & n23575 ) | ( n6649 & n23575 ) ;
  assign n23577 = n16942 ^ n13455 ^ n10371 ;
  assign n23578 = ( n9362 & n23576 ) | ( n9362 & ~n23577 ) | ( n23576 & ~n23577 ) ;
  assign n23579 = ( ~n1081 & n6303 ) | ( ~n1081 & n9884 ) | ( n6303 & n9884 ) ;
  assign n23580 = ( n1589 & ~n18201 ) | ( n1589 & n23579 ) | ( ~n18201 & n23579 ) ;
  assign n23581 = n23580 ^ n18959 ^ n1105 ;
  assign n23582 = n15825 ^ n8128 ^ n7121 ;
  assign n23583 = n23582 ^ n20558 ^ n936 ;
  assign n23584 = n15755 ^ n13903 ^ n7368 ;
  assign n23585 = n23584 ^ n20661 ^ n4775 ;
  assign n23587 = n6957 ^ n5510 ^ n3909 ;
  assign n23586 = n20255 ^ n10307 ^ n4237 ;
  assign n23588 = n23587 ^ n23586 ^ n14181 ;
  assign n23590 = n22433 ^ n11192 ^ n4256 ;
  assign n23589 = n20576 ^ n15431 ^ n9803 ;
  assign n23591 = n23590 ^ n23589 ^ n9528 ;
  assign n23592 = ( n996 & ~n1626 ) | ( n996 & n3033 ) | ( ~n1626 & n3033 ) ;
  assign n23593 = ( ~n2349 & n21586 ) | ( ~n2349 & n23592 ) | ( n21586 & n23592 ) ;
  assign n23594 = ( ~n2354 & n10297 ) | ( ~n2354 & n11411 ) | ( n10297 & n11411 ) ;
  assign n23596 = ( n358 & ~n1657 ) | ( n358 & n2295 ) | ( ~n1657 & n2295 ) ;
  assign n23595 = ( n2335 & n9598 ) | ( n2335 & ~n11125 ) | ( n9598 & ~n11125 ) ;
  assign n23597 = n23596 ^ n23595 ^ n7422 ;
  assign n23598 = n23597 ^ n3357 ^ n2919 ;
  assign n23599 = n16930 ^ n15411 ^ n12644 ;
  assign n23600 = n18631 ^ n8418 ^ n3900 ;
  assign n23601 = ( ~n23598 & n23599 ) | ( ~n23598 & n23600 ) | ( n23599 & n23600 ) ;
  assign n23602 = ( ~n3299 & n4408 ) | ( ~n3299 & n11415 ) | ( n4408 & n11415 ) ;
  assign n23603 = n23602 ^ n19127 ^ n9991 ;
  assign n23604 = ( n3285 & ~n9220 ) | ( n3285 & n17062 ) | ( ~n9220 & n17062 ) ;
  assign n23605 = n23604 ^ n10791 ^ n4253 ;
  assign n23606 = n23605 ^ n4795 ^ n286 ;
  assign n23607 = n4586 ^ n2512 ^ n251 ;
  assign n23608 = n23607 ^ n6928 ^ n2752 ;
  assign n23609 = ( ~n8477 & n12672 ) | ( ~n8477 & n23608 ) | ( n12672 & n23608 ) ;
  assign n23610 = n23609 ^ n23226 ^ n16809 ;
  assign n23611 = ( n6399 & n6651 ) | ( n6399 & ~n7197 ) | ( n6651 & ~n7197 ) ;
  assign n23612 = n23611 ^ n6327 ^ n3448 ;
  assign n23613 = n13078 ^ n12062 ^ n10602 ;
  assign n23614 = ( ~n4026 & n15693 ) | ( ~n4026 & n16059 ) | ( n15693 & n16059 ) ;
  assign n23615 = ( ~n1007 & n1741 ) | ( ~n1007 & n10039 ) | ( n1741 & n10039 ) ;
  assign n23616 = ( n4373 & ~n4777 ) | ( n4373 & n23615 ) | ( ~n4777 & n23615 ) ;
  assign n23619 = ( n3212 & n17720 ) | ( n3212 & n20596 ) | ( n17720 & n20596 ) ;
  assign n23617 = ( n9151 & n10410 ) | ( n9151 & ~n11258 ) | ( n10410 & ~n11258 ) ;
  assign n23618 = n23617 ^ n21585 ^ n2058 ;
  assign n23620 = n23619 ^ n23618 ^ n18062 ;
  assign n23622 = ( n2035 & n4981 ) | ( n2035 & n11156 ) | ( n4981 & n11156 ) ;
  assign n23621 = ( n1940 & ~n7416 ) | ( n1940 & n15864 ) | ( ~n7416 & n15864 ) ;
  assign n23623 = n23622 ^ n23621 ^ n11820 ;
  assign n23624 = n23623 ^ n10613 ^ n775 ;
  assign n23625 = ( n3522 & ~n4426 ) | ( n3522 & n8352 ) | ( ~n4426 & n8352 ) ;
  assign n23626 = ( n22934 & n23624 ) | ( n22934 & n23625 ) | ( n23624 & n23625 ) ;
  assign n23627 = n19539 ^ n13629 ^ n2368 ;
  assign n23631 = n14729 ^ n6915 ^ n6863 ;
  assign n23630 = n12394 ^ n10293 ^ n8115 ;
  assign n23628 = ( ~n809 & n11878 ) | ( ~n809 & n23453 ) | ( n11878 & n23453 ) ;
  assign n23629 = n23628 ^ n11010 ^ n360 ;
  assign n23632 = n23631 ^ n23630 ^ n23629 ;
  assign n23634 = ( n10468 & n11522 ) | ( n10468 & n13666 ) | ( n11522 & n13666 ) ;
  assign n23633 = n22908 ^ n20228 ^ n16398 ;
  assign n23635 = n23634 ^ n23633 ^ n2604 ;
  assign n23636 = n23635 ^ n15039 ^ n6776 ;
  assign n23637 = n18907 ^ n16356 ^ n8569 ;
  assign n23638 = n11237 ^ n7140 ^ n4375 ;
  assign n23639 = ( ~n11377 & n11881 ) | ( ~n11377 & n15775 ) | ( n11881 & n15775 ) ;
  assign n23640 = n13933 ^ n13455 ^ n5761 ;
  assign n23641 = ( n641 & n12494 ) | ( n641 & n18837 ) | ( n12494 & n18837 ) ;
  assign n23642 = ( ~n17400 & n23640 ) | ( ~n17400 & n23641 ) | ( n23640 & n23641 ) ;
  assign n23643 = n23642 ^ n14443 ^ n3326 ;
  assign n23644 = n10848 ^ n2445 ^ n944 ;
  assign n23645 = n23644 ^ n14311 ^ n7176 ;
  assign n23646 = ( ~n1254 & n4961 ) | ( ~n1254 & n13323 ) | ( n4961 & n13323 ) ;
  assign n23647 = ( n15069 & ~n20637 ) | ( n15069 & n23646 ) | ( ~n20637 & n23646 ) ;
  assign n23648 = n16610 ^ n4561 ^ n2325 ;
  assign n23649 = ( ~n264 & n4794 ) | ( ~n264 & n19359 ) | ( n4794 & n19359 ) ;
  assign n23650 = ( n1257 & n16081 ) | ( n1257 & ~n23649 ) | ( n16081 & ~n23649 ) ;
  assign n23651 = n19590 ^ n17668 ^ n1678 ;
  assign n23652 = ( n6634 & ~n13846 ) | ( n6634 & n23651 ) | ( ~n13846 & n23651 ) ;
  assign n23653 = ( n4398 & n8687 ) | ( n4398 & ~n11665 ) | ( n8687 & ~n11665 ) ;
  assign n23654 = ( ~n1272 & n8849 ) | ( ~n1272 & n9796 ) | ( n8849 & n9796 ) ;
  assign n23655 = ( ~n917 & n10066 ) | ( ~n917 & n23654 ) | ( n10066 & n23654 ) ;
  assign n23656 = ( n3045 & n5762 ) | ( n3045 & ~n18957 ) | ( n5762 & ~n18957 ) ;
  assign n23657 = ( n5017 & ~n7971 ) | ( n5017 & n17341 ) | ( ~n7971 & n17341 ) ;
  assign n23658 = ( n1106 & n7438 ) | ( n1106 & n15346 ) | ( n7438 & n15346 ) ;
  assign n23664 = n13850 ^ n10092 ^ n6121 ;
  assign n23662 = ( n3865 & n17952 ) | ( n3865 & n18337 ) | ( n17952 & n18337 ) ;
  assign n23660 = n14119 ^ n10519 ^ n7427 ;
  assign n23661 = ( n1437 & n4302 ) | ( n1437 & n23660 ) | ( n4302 & n23660 ) ;
  assign n23663 = n23662 ^ n23661 ^ n21125 ;
  assign n23659 = n6284 ^ n5720 ^ n1337 ;
  assign n23665 = n23664 ^ n23663 ^ n23659 ;
  assign n23666 = n9926 ^ n4155 ^ n2774 ;
  assign n23667 = ( n13951 & n15304 ) | ( n13951 & ~n23666 ) | ( n15304 & ~n23666 ) ;
  assign n23668 = n23667 ^ n22073 ^ n14673 ;
  assign n23670 = ( n4202 & n4577 ) | ( n4202 & ~n9072 ) | ( n4577 & ~n9072 ) ;
  assign n23669 = n18592 ^ n6709 ^ n923 ;
  assign n23671 = n23670 ^ n23669 ^ n2796 ;
  assign n23672 = n2580 ^ n492 ^ n351 ;
  assign n23673 = ( ~n6362 & n22812 ) | ( ~n6362 & n23672 ) | ( n22812 & n23672 ) ;
  assign n23674 = ( ~n5071 & n6005 ) | ( ~n5071 & n23673 ) | ( n6005 & n23673 ) ;
  assign n23675 = ( n4682 & ~n8396 ) | ( n4682 & n21162 ) | ( ~n8396 & n21162 ) ;
  assign n23676 = n23675 ^ n15509 ^ n852 ;
  assign n23677 = n13618 ^ n8557 ^ n7385 ;
  assign n23678 = n7558 ^ n2770 ^ n2562 ;
  assign n23679 = ( n22996 & n23677 ) | ( n22996 & ~n23678 ) | ( n23677 & ~n23678 ) ;
  assign n23680 = n15586 ^ n11513 ^ n10712 ;
  assign n23681 = n14186 ^ n12514 ^ n5730 ;
  assign n23682 = ( n10059 & n15734 ) | ( n10059 & n23681 ) | ( n15734 & n23681 ) ;
  assign n23683 = n15206 ^ n8285 ^ n3118 ;
  assign n23684 = ( ~n984 & n1254 ) | ( ~n984 & n10698 ) | ( n1254 & n10698 ) ;
  assign n23685 = n23684 ^ n12867 ^ n11081 ;
  assign n23690 = ( ~n4151 & n6553 ) | ( ~n4151 & n12456 ) | ( n6553 & n12456 ) ;
  assign n23691 = n23690 ^ n17838 ^ n9492 ;
  assign n23686 = n15341 ^ n15131 ^ n10694 ;
  assign n23687 = n23686 ^ n7966 ^ n6256 ;
  assign n23688 = n23687 ^ n6692 ^ n3059 ;
  assign n23689 = n23688 ^ n21814 ^ n3905 ;
  assign n23692 = n23691 ^ n23689 ^ n4445 ;
  assign n23693 = ( n2748 & n9567 ) | ( n2748 & ~n11468 ) | ( n9567 & ~n11468 ) ;
  assign n23694 = ( ~n4818 & n8194 ) | ( ~n4818 & n23693 ) | ( n8194 & n23693 ) ;
  assign n23695 = n23694 ^ n3448 ^ n2118 ;
  assign n23697 = ( n3096 & n15791 ) | ( n3096 & ~n23497 ) | ( n15791 & ~n23497 ) ;
  assign n23696 = ( ~n293 & n434 ) | ( ~n293 & n13083 ) | ( n434 & n13083 ) ;
  assign n23698 = n23697 ^ n23696 ^ n20901 ;
  assign n23699 = n23698 ^ n17592 ^ n15541 ;
  assign n23700 = ( n2195 & n8446 ) | ( n2195 & ~n23699 ) | ( n8446 & ~n23699 ) ;
  assign n23701 = n23700 ^ n21241 ^ n4556 ;
  assign n23702 = n20519 ^ n17537 ^ n16003 ;
  assign n23703 = ( n2387 & n9894 ) | ( n2387 & ~n16264 ) | ( n9894 & ~n16264 ) ;
  assign n23704 = ( n13828 & n19439 ) | ( n13828 & ~n23703 ) | ( n19439 & ~n23703 ) ;
  assign n23705 = ( n6366 & n8460 ) | ( n6366 & ~n23704 ) | ( n8460 & ~n23704 ) ;
  assign n23706 = ( n6439 & n9873 ) | ( n6439 & n23705 ) | ( n9873 & n23705 ) ;
  assign n23707 = n23706 ^ n7764 ^ n6058 ;
  assign n23708 = n12709 ^ n11350 ^ n8543 ;
  assign n23709 = n10397 ^ n6082 ^ n1697 ;
  assign n23710 = n23709 ^ n21976 ^ n7008 ;
  assign n23711 = n19995 ^ n19735 ^ n15540 ;
  assign n23712 = ( ~n4690 & n20121 ) | ( ~n4690 & n20715 ) | ( n20121 & n20715 ) ;
  assign n23713 = ( n5368 & n14928 ) | ( n5368 & ~n17668 ) | ( n14928 & ~n17668 ) ;
  assign n23714 = ( n1973 & n17297 ) | ( n1973 & ~n21041 ) | ( n17297 & ~n21041 ) ;
  assign n23715 = n13352 ^ n6288 ^ n2093 ;
  assign n23716 = n23715 ^ n19953 ^ n10515 ;
  assign n23718 = n11319 ^ n2553 ^ n1977 ;
  assign n23719 = n23718 ^ n21113 ^ n21028 ;
  assign n23717 = n8358 ^ n7999 ^ n4997 ;
  assign n23720 = n23719 ^ n23717 ^ n2626 ;
  assign n23721 = ( n15074 & ~n15718 ) | ( n15074 & n21162 ) | ( ~n15718 & n21162 ) ;
  assign n23722 = ( ~n13472 & n16871 ) | ( ~n13472 & n23721 ) | ( n16871 & n23721 ) ;
  assign n23723 = ( n3328 & n8773 ) | ( n3328 & ~n23722 ) | ( n8773 & ~n23722 ) ;
  assign n23724 = n17573 ^ n13882 ^ n7602 ;
  assign n23725 = ( n184 & n5125 ) | ( n184 & ~n15095 ) | ( n5125 & ~n15095 ) ;
  assign n23726 = ( n4957 & n22802 ) | ( n4957 & ~n23725 ) | ( n22802 & ~n23725 ) ;
  assign n23727 = ( ~n11228 & n23724 ) | ( ~n11228 & n23726 ) | ( n23724 & n23726 ) ;
  assign n23728 = n18503 ^ n5757 ^ n2304 ;
  assign n23729 = ( ~n267 & n12823 ) | ( ~n267 & n18399 ) | ( n12823 & n18399 ) ;
  assign n23730 = n23729 ^ n23354 ^ n6381 ;
  assign n23731 = ( ~n9550 & n10522 ) | ( ~n9550 & n16459 ) | ( n10522 & n16459 ) ;
  assign n23732 = ( n12197 & ~n23730 ) | ( n12197 & n23731 ) | ( ~n23730 & n23731 ) ;
  assign n23737 = n13938 ^ n8627 ^ n2675 ;
  assign n23738 = ( ~n5289 & n7784 ) | ( ~n5289 & n23737 ) | ( n7784 & n23737 ) ;
  assign n23739 = n23738 ^ n8267 ^ n5295 ;
  assign n23734 = ( n2023 & n6691 ) | ( n2023 & n11372 ) | ( n6691 & n11372 ) ;
  assign n23733 = n8467 ^ n2249 ^ n2184 ;
  assign n23735 = n23734 ^ n23733 ^ n2381 ;
  assign n23736 = n23735 ^ n17631 ^ n5622 ;
  assign n23740 = n23739 ^ n23736 ^ n11189 ;
  assign n23741 = ( n1403 & n1642 ) | ( n1403 & ~n11677 ) | ( n1642 & ~n11677 ) ;
  assign n23742 = n20627 ^ n10139 ^ n7688 ;
  assign n23743 = ( ~n782 & n23741 ) | ( ~n782 & n23742 ) | ( n23741 & n23742 ) ;
  assign n23744 = n23743 ^ n14716 ^ n9787 ;
  assign n23745 = ( n1331 & ~n13316 ) | ( n1331 & n14436 ) | ( ~n13316 & n14436 ) ;
  assign n23748 = n15865 ^ n4683 ^ n176 ;
  assign n23747 = n20218 ^ n14606 ^ n4293 ;
  assign n23749 = n23748 ^ n23747 ^ n14077 ;
  assign n23746 = n16071 ^ n13511 ^ n6244 ;
  assign n23750 = n23749 ^ n23746 ^ n20792 ;
  assign n23751 = n23750 ^ n16129 ^ n11043 ;
  assign n23752 = n23751 ^ n9920 ^ n6298 ;
  assign n23753 = ( n274 & n18752 ) | ( n274 & n21413 ) | ( n18752 & n21413 ) ;
  assign n23754 = ( n1073 & ~n19623 ) | ( n1073 & n23753 ) | ( ~n19623 & n23753 ) ;
  assign n23757 = n8345 ^ n6297 ^ n1139 ;
  assign n23758 = n23757 ^ n11450 ^ n545 ;
  assign n23755 = n11078 ^ n2904 ^ n557 ;
  assign n23756 = ( n3249 & n16113 ) | ( n3249 & n23755 ) | ( n16113 & n23755 ) ;
  assign n23759 = n23758 ^ n23756 ^ n3695 ;
  assign n23760 = n23759 ^ n22862 ^ n7598 ;
  assign n23761 = n17746 ^ n10063 ^ n1453 ;
  assign n23762 = ( n10958 & ~n11718 ) | ( n10958 & n23761 ) | ( ~n11718 & n23761 ) ;
  assign n23763 = ( n8477 & n10446 ) | ( n8477 & n22264 ) | ( n10446 & n22264 ) ;
  assign n23764 = n23763 ^ n15767 ^ n1896 ;
  assign n23765 = n7051 ^ n6991 ^ n6927 ;
  assign n23766 = n23765 ^ n14759 ^ n6463 ;
  assign n23767 = ( n19029 & n23764 ) | ( n19029 & n23766 ) | ( n23764 & n23766 ) ;
  assign n23768 = n8122 ^ n7871 ^ n7009 ;
  assign n23769 = ( n3704 & n9173 ) | ( n3704 & n23768 ) | ( n9173 & n23768 ) ;
  assign n23770 = n23769 ^ n20757 ^ n8064 ;
  assign n23771 = ( n6352 & n11660 ) | ( n6352 & ~n23770 ) | ( n11660 & ~n23770 ) ;
  assign n23772 = n15292 ^ n12709 ^ n1151 ;
  assign n23773 = ( n5020 & n7316 ) | ( n5020 & n7725 ) | ( n7316 & n7725 ) ;
  assign n23774 = n23773 ^ n20162 ^ n1359 ;
  assign n23775 = ( n5531 & n7216 ) | ( n5531 & n14201 ) | ( n7216 & n14201 ) ;
  assign n23776 = ( ~n6633 & n16394 ) | ( ~n6633 & n23775 ) | ( n16394 & n23775 ) ;
  assign n23777 = n23776 ^ n17047 ^ n4595 ;
  assign n23778 = ( n7015 & n13324 ) | ( n7015 & ~n20381 ) | ( n13324 & ~n20381 ) ;
  assign n23779 = n23778 ^ n11408 ^ n3835 ;
  assign n23780 = ( ~n5032 & n23777 ) | ( ~n5032 & n23779 ) | ( n23777 & n23779 ) ;
  assign n23781 = n16705 ^ n4696 ^ n1182 ;
  assign n23782 = n23781 ^ n18575 ^ n15900 ;
  assign n23783 = n10988 ^ n7030 ^ n6904 ;
  assign n23784 = n23783 ^ n14774 ^ n12037 ;
  assign n23785 = n23784 ^ n21153 ^ n3141 ;
  assign n23786 = n18251 ^ n11848 ^ n730 ;
  assign n23787 = n21123 ^ n20272 ^ n11364 ;
  assign n23788 = ( n17585 & ~n23786 ) | ( n17585 & n23787 ) | ( ~n23786 & n23787 ) ;
  assign n23789 = n12564 ^ n4571 ^ n4496 ;
  assign n23791 = n23419 ^ n794 ^ n413 ;
  assign n23790 = ( n2445 & ~n5324 ) | ( n2445 & n14618 ) | ( ~n5324 & n14618 ) ;
  assign n23792 = n23791 ^ n23790 ^ n5295 ;
  assign n23793 = n19869 ^ n19258 ^ n15683 ;
  assign n23794 = n14240 ^ n10679 ^ n9622 ;
  assign n23795 = ( n10309 & n23793 ) | ( n10309 & ~n23794 ) | ( n23793 & ~n23794 ) ;
  assign n23796 = n23795 ^ n12147 ^ n9419 ;
  assign n23797 = n15272 ^ n11250 ^ n6949 ;
  assign n23798 = n23797 ^ n16150 ^ n10609 ;
  assign n23799 = ( ~n4867 & n16868 ) | ( ~n4867 & n19125 ) | ( n16868 & n19125 ) ;
  assign n23800 = n23799 ^ n6009 ^ n2935 ;
  assign n23803 = n14516 ^ n3699 ^ n1292 ;
  assign n23801 = n14881 ^ n5486 ^ n1541 ;
  assign n23802 = n23801 ^ n21229 ^ n13413 ;
  assign n23804 = n23803 ^ n23802 ^ n2188 ;
  assign n23805 = n11150 ^ n9050 ^ n3306 ;
  assign n23806 = n23805 ^ n6673 ^ n2491 ;
  assign n23807 = n21717 ^ n15929 ^ n6940 ;
  assign n23809 = n17231 ^ n2726 ^ n827 ;
  assign n23810 = n23809 ^ n18591 ^ n6925 ;
  assign n23808 = n18306 ^ n7307 ^ n348 ;
  assign n23811 = n23810 ^ n23808 ^ n3812 ;
  assign n23812 = n19857 ^ n10189 ^ n7851 ;
  assign n23813 = n13426 ^ n755 ^ n290 ;
  assign n23814 = ( n5951 & ~n7501 ) | ( n5951 & n8977 ) | ( ~n7501 & n8977 ) ;
  assign n23815 = n20329 ^ n18786 ^ n18769 ;
  assign n23816 = ( n1795 & n2897 ) | ( n1795 & n5213 ) | ( n2897 & n5213 ) ;
  assign n23817 = ( n2469 & n13433 ) | ( n2469 & ~n23816 ) | ( n13433 & ~n23816 ) ;
  assign n23818 = n23817 ^ n10830 ^ n5462 ;
  assign n23819 = ( ~n15851 & n19426 ) | ( ~n15851 & n23818 ) | ( n19426 & n23818 ) ;
  assign n23820 = n16583 ^ n12177 ^ n11998 ;
  assign n23821 = n23820 ^ n17955 ^ n1945 ;
  assign n23822 = n23821 ^ n13577 ^ n9967 ;
  assign n23823 = ( n16238 & ~n23282 ) | ( n16238 & n23822 ) | ( ~n23282 & n23822 ) ;
  assign n23828 = n16150 ^ n9689 ^ n1040 ;
  assign n23829 = n4207 ^ n3667 ^ n1898 ;
  assign n23830 = ( n2449 & n6953 ) | ( n2449 & n23829 ) | ( n6953 & n23829 ) ;
  assign n23831 = ( n12896 & n23828 ) | ( n12896 & n23830 ) | ( n23828 & n23830 ) ;
  assign n23824 = ( n1636 & n7891 ) | ( n1636 & n16921 ) | ( n7891 & n16921 ) ;
  assign n23825 = ( n6124 & ~n15583 ) | ( n6124 & n23824 ) | ( ~n15583 & n23824 ) ;
  assign n23826 = ( ~n4713 & n11040 ) | ( ~n4713 & n17808 ) | ( n11040 & n17808 ) ;
  assign n23827 = ( n17914 & ~n23825 ) | ( n17914 & n23826 ) | ( ~n23825 & n23826 ) ;
  assign n23832 = n23831 ^ n23827 ^ n2786 ;
  assign n23833 = ( n4161 & ~n5999 ) | ( n4161 & n15236 ) | ( ~n5999 & n15236 ) ;
  assign n23834 = ( n6758 & ~n12749 ) | ( n6758 & n13649 ) | ( ~n12749 & n13649 ) ;
  assign n23835 = ( ~n3981 & n12763 ) | ( ~n3981 & n14200 ) | ( n12763 & n14200 ) ;
  assign n23836 = ( ~n5771 & n21460 ) | ( ~n5771 & n23835 ) | ( n21460 & n23835 ) ;
  assign n23837 = ( n3783 & ~n4189 ) | ( n3783 & n18725 ) | ( ~n4189 & n18725 ) ;
  assign n23838 = n23837 ^ n8555 ^ n1779 ;
  assign n23839 = ( n186 & ~n6742 ) | ( n186 & n16462 ) | ( ~n6742 & n16462 ) ;
  assign n23840 = n5284 ^ n5151 ^ n3414 ;
  assign n23841 = ( n916 & ~n7855 ) | ( n916 & n23840 ) | ( ~n7855 & n23840 ) ;
  assign n23842 = n23841 ^ n19209 ^ n1130 ;
  assign n23843 = ( n3141 & n5225 ) | ( n3141 & ~n23842 ) | ( n5225 & ~n23842 ) ;
  assign n23844 = ( n13030 & n23839 ) | ( n13030 & ~n23843 ) | ( n23839 & ~n23843 ) ;
  assign n23845 = n23563 ^ n23322 ^ n22526 ;
  assign n23846 = n15106 ^ n12966 ^ n11179 ;
  assign n23847 = n23846 ^ n14893 ^ n13618 ;
  assign n23848 = ( n8046 & n10506 ) | ( n8046 & n21250 ) | ( n10506 & n21250 ) ;
  assign n23849 = n23848 ^ n12160 ^ n8483 ;
  assign n23850 = ( n5123 & n9744 ) | ( n5123 & ~n23849 ) | ( n9744 & ~n23849 ) ;
  assign n23852 = n10626 ^ n10288 ^ n6941 ;
  assign n23851 = ( n9884 & n10441 ) | ( n9884 & ~n21087 ) | ( n10441 & ~n21087 ) ;
  assign n23853 = n23852 ^ n23851 ^ n12249 ;
  assign n23854 = ( n5406 & n7489 ) | ( n5406 & n8303 ) | ( n7489 & n8303 ) ;
  assign n23855 = ( n10241 & n10911 ) | ( n10241 & n22688 ) | ( n10911 & n22688 ) ;
  assign n23856 = ( n1748 & ~n23854 ) | ( n1748 & n23855 ) | ( ~n23854 & n23855 ) ;
  assign n23857 = n17273 ^ n6849 ^ n626 ;
  assign n23858 = ( n12536 & n14028 ) | ( n12536 & ~n17067 ) | ( n14028 & ~n17067 ) ;
  assign n23859 = n22728 ^ n18367 ^ n1121 ;
  assign n23860 = ( n3576 & n7699 ) | ( n3576 & ~n15333 ) | ( n7699 & ~n15333 ) ;
  assign n23861 = ( n508 & n20119 ) | ( n508 & n23860 ) | ( n20119 & n23860 ) ;
  assign n23862 = ( ~n14105 & n16292 ) | ( ~n14105 & n23861 ) | ( n16292 & n23861 ) ;
  assign n23863 = n22634 ^ n11470 ^ n4408 ;
  assign n23864 = n23863 ^ n16063 ^ n2957 ;
  assign n23865 = n12422 ^ n3332 ^ n2569 ;
  assign n23866 = n23865 ^ n20634 ^ n381 ;
  assign n23868 = n21117 ^ n5241 ^ n706 ;
  assign n23867 = n17793 ^ n12947 ^ n11087 ;
  assign n23869 = n23868 ^ n23867 ^ n7214 ;
  assign n23870 = ( ~n2965 & n3830 ) | ( ~n2965 & n4295 ) | ( n3830 & n4295 ) ;
  assign n23871 = n14224 ^ n5971 ^ n1592 ;
  assign n23872 = ( n6920 & ~n20331 ) | ( n6920 & n23871 ) | ( ~n20331 & n23871 ) ;
  assign n23878 = ( n1608 & n2408 ) | ( n1608 & ~n10969 ) | ( n2408 & ~n10969 ) ;
  assign n23877 = n14043 ^ n3797 ^ n2689 ;
  assign n23874 = ( n1204 & n3898 ) | ( n1204 & ~n11036 ) | ( n3898 & ~n11036 ) ;
  assign n23875 = ( n15261 & ~n22706 ) | ( n15261 & n23874 ) | ( ~n22706 & n23874 ) ;
  assign n23873 = ( n10074 & ~n11498 ) | ( n10074 & n14835 ) | ( ~n11498 & n14835 ) ;
  assign n23876 = n23875 ^ n23873 ^ n5862 ;
  assign n23879 = n23878 ^ n23877 ^ n23876 ;
  assign n23880 = ( ~n1171 & n5269 ) | ( ~n1171 & n8005 ) | ( n5269 & n8005 ) ;
  assign n23881 = n23880 ^ n18970 ^ n8990 ;
  assign n23882 = ( n6275 & ~n13465 ) | ( n6275 & n21519 ) | ( ~n13465 & n21519 ) ;
  assign n23883 = ( ~n22034 & n23881 ) | ( ~n22034 & n23882 ) | ( n23881 & n23882 ) ;
  assign n23884 = ( n1259 & n10726 ) | ( n1259 & n21982 ) | ( n10726 & n21982 ) ;
  assign n23885 = n23884 ^ n18135 ^ n292 ;
  assign n23886 = ( n4374 & ~n15504 ) | ( n4374 & n21274 ) | ( ~n15504 & n21274 ) ;
  assign n23887 = ( ~n3792 & n13859 ) | ( ~n3792 & n16397 ) | ( n13859 & n16397 ) ;
  assign n23888 = n23887 ^ n9907 ^ n3218 ;
  assign n23889 = ( ~n5623 & n10716 ) | ( ~n5623 & n23888 ) | ( n10716 & n23888 ) ;
  assign n23890 = n19562 ^ n10985 ^ n10342 ;
  assign n23891 = n10605 ^ n3812 ^ n970 ;
  assign n23892 = n23891 ^ n22111 ^ n20943 ;
  assign n23893 = ( ~n1272 & n3676 ) | ( ~n1272 & n14240 ) | ( n3676 & n14240 ) ;
  assign n23894 = ( n208 & n23892 ) | ( n208 & ~n23893 ) | ( n23892 & ~n23893 ) ;
  assign n23895 = ( n5583 & n8595 ) | ( n5583 & ~n13124 ) | ( n8595 & ~n13124 ) ;
  assign n23896 = n23895 ^ n19445 ^ n15154 ;
  assign n23897 = n12397 ^ n10683 ^ n3029 ;
  assign n23898 = ( ~n3335 & n18350 ) | ( ~n3335 & n19829 ) | ( n18350 & n19829 ) ;
  assign n23899 = ( n4120 & n7314 ) | ( n4120 & n11893 ) | ( n7314 & n11893 ) ;
  assign n23900 = n23899 ^ n21607 ^ n1885 ;
  assign n23901 = n17281 ^ n7522 ^ n6932 ;
  assign n23902 = n23901 ^ n6119 ^ n4742 ;
  assign n23903 = ( ~n10574 & n23900 ) | ( ~n10574 & n23902 ) | ( n23900 & n23902 ) ;
  assign n23904 = n14535 ^ n10132 ^ n5232 ;
  assign n23905 = ( ~n5945 & n23903 ) | ( ~n5945 & n23904 ) | ( n23903 & n23904 ) ;
  assign n23907 = n7746 ^ n6919 ^ n222 ;
  assign n23908 = n23907 ^ n17151 ^ n11066 ;
  assign n23906 = ( ~n4950 & n16064 ) | ( ~n4950 & n17961 ) | ( n16064 & n17961 ) ;
  assign n23909 = n23908 ^ n23906 ^ n8364 ;
  assign n23910 = ( n1903 & n16977 ) | ( n1903 & n23909 ) | ( n16977 & n23909 ) ;
  assign n23911 = n10601 ^ n5895 ^ n4253 ;
  assign n23912 = ( ~n18221 & n19078 ) | ( ~n18221 & n23495 ) | ( n19078 & n23495 ) ;
  assign n23913 = ( n2989 & ~n7557 ) | ( n2989 & n23912 ) | ( ~n7557 & n23912 ) ;
  assign n23914 = ( n16028 & n20322 ) | ( n16028 & ~n20709 ) | ( n20322 & ~n20709 ) ;
  assign n23915 = n12962 ^ n7010 ^ n4242 ;
  assign n23916 = n19111 ^ n7809 ^ n358 ;
  assign n23917 = ( ~n6098 & n18153 ) | ( ~n6098 & n23916 ) | ( n18153 & n23916 ) ;
  assign n23918 = ( n6738 & ~n17025 ) | ( n6738 & n23917 ) | ( ~n17025 & n23917 ) ;
  assign n23919 = n6414 ^ n6358 ^ n4865 ;
  assign n23920 = ( ~n7175 & n12333 ) | ( ~n7175 & n23919 ) | ( n12333 & n23919 ) ;
  assign n23921 = n23920 ^ n17993 ^ n3676 ;
  assign n23922 = n10715 ^ n9496 ^ n6823 ;
  assign n23923 = ( n1155 & ~n2827 ) | ( n1155 & n23068 ) | ( ~n2827 & n23068 ) ;
  assign n23924 = ( n532 & n19207 ) | ( n532 & n23923 ) | ( n19207 & n23923 ) ;
  assign n23925 = ( n627 & n23922 ) | ( n627 & ~n23924 ) | ( n23922 & ~n23924 ) ;
  assign n23926 = n6018 ^ n4162 ^ n3018 ;
  assign n23927 = ( n849 & n7955 ) | ( n849 & ~n23926 ) | ( n7955 & ~n23926 ) ;
  assign n23928 = n12587 ^ n8912 ^ n2177 ;
  assign n23929 = ( n3491 & ~n6867 ) | ( n3491 & n14366 ) | ( ~n6867 & n14366 ) ;
  assign n23930 = n16156 ^ n3921 ^ n1630 ;
  assign n23931 = ( ~n1368 & n1611 ) | ( ~n1368 & n20674 ) | ( n1611 & n20674 ) ;
  assign n23932 = n16722 ^ n13272 ^ n4215 ;
  assign n23933 = ( n7726 & n16730 ) | ( n7726 & ~n23390 ) | ( n16730 & ~n23390 ) ;
  assign n23934 = ( ~n16492 & n20085 ) | ( ~n16492 & n23933 ) | ( n20085 & n23933 ) ;
  assign n23935 = n20591 ^ n18539 ^ n16626 ;
  assign n23936 = n23935 ^ n12526 ^ n9572 ;
  assign n23938 = ( n256 & ~n1555 ) | ( n256 & n5854 ) | ( ~n1555 & n5854 ) ;
  assign n23939 = n20704 ^ n18600 ^ n3639 ;
  assign n23940 = ( n12743 & n23938 ) | ( n12743 & n23939 ) | ( n23938 & n23939 ) ;
  assign n23937 = ( n6780 & n21049 ) | ( n6780 & ~n23817 ) | ( n21049 & ~n23817 ) ;
  assign n23941 = n23940 ^ n23937 ^ n17365 ;
  assign n23942 = n15000 ^ n8214 ^ n1022 ;
  assign n23948 = ( n10111 & n11883 ) | ( n10111 & n15628 ) | ( n11883 & n15628 ) ;
  assign n23949 = ( n5470 & ~n23457 ) | ( n5470 & n23948 ) | ( ~n23457 & n23948 ) ;
  assign n23950 = ( n1554 & n15896 ) | ( n1554 & n23949 ) | ( n15896 & n23949 ) ;
  assign n23946 = n7793 ^ n2601 ^ n1392 ;
  assign n23947 = n23946 ^ n20189 ^ n9105 ;
  assign n23944 = ( n1406 & n3306 ) | ( n1406 & ~n5203 ) | ( n3306 & ~n5203 ) ;
  assign n23943 = ( n4678 & n15260 ) | ( n4678 & ~n17277 ) | ( n15260 & ~n17277 ) ;
  assign n23945 = n23944 ^ n23943 ^ n8303 ;
  assign n23951 = n23950 ^ n23947 ^ n23945 ;
  assign n23952 = n12115 ^ n3029 ^ n2837 ;
  assign n23953 = n6457 ^ n5190 ^ n2643 ;
  assign n23954 = n23953 ^ n13284 ^ n756 ;
  assign n23955 = ( ~n2821 & n11291 ) | ( ~n2821 & n23954 ) | ( n11291 & n23954 ) ;
  assign n23956 = n23955 ^ n19197 ^ n13946 ;
  assign n23957 = n23956 ^ n14981 ^ n8140 ;
  assign n23958 = ( n240 & n1360 ) | ( n240 & ~n23957 ) | ( n1360 & ~n23957 ) ;
  assign n23960 = ( ~n820 & n4193 ) | ( ~n820 & n10780 ) | ( n4193 & n10780 ) ;
  assign n23961 = n23960 ^ n5805 ^ n4108 ;
  assign n23959 = ( n2630 & ~n6070 ) | ( n2630 & n11351 ) | ( ~n6070 & n11351 ) ;
  assign n23962 = n23961 ^ n23959 ^ n11427 ;
  assign n23963 = ( n1627 & n4596 ) | ( n1627 & ~n23962 ) | ( n4596 & ~n23962 ) ;
  assign n23964 = n2414 ^ n2120 ^ n1929 ;
  assign n23966 = n17125 ^ n7317 ^ n6806 ;
  assign n23965 = n14026 ^ n8722 ^ n478 ;
  assign n23967 = n23966 ^ n23965 ^ n20893 ;
  assign n23968 = ( n8355 & n23964 ) | ( n8355 & n23967 ) | ( n23964 & n23967 ) ;
  assign n23969 = ( ~n14720 & n15642 ) | ( ~n14720 & n23263 ) | ( n15642 & n23263 ) ;
  assign n23970 = n22963 ^ n19545 ^ n19054 ;
  assign n23971 = ( n2848 & ~n3534 ) | ( n2848 & n22976 ) | ( ~n3534 & n22976 ) ;
  assign n23972 = n5476 ^ n2852 ^ n2127 ;
  assign n23973 = ( n23970 & ~n23971 ) | ( n23970 & n23972 ) | ( ~n23971 & n23972 ) ;
  assign n23974 = n23973 ^ n22034 ^ n18301 ;
  assign n23975 = n23974 ^ n8912 ^ n1193 ;
  assign n23978 = ( ~n735 & n4049 ) | ( ~n735 & n14216 ) | ( n4049 & n14216 ) ;
  assign n23976 = ( n1353 & n4027 ) | ( n1353 & n15853 ) | ( n4027 & n15853 ) ;
  assign n23977 = n23976 ^ n21754 ^ n9251 ;
  assign n23979 = n23978 ^ n23977 ^ n18559 ;
  assign n23980 = n16095 ^ n14577 ^ n7468 ;
  assign n23981 = n23980 ^ n17077 ^ n6670 ;
  assign n23982 = ( n5714 & n19940 ) | ( n5714 & ~n23981 ) | ( n19940 & ~n23981 ) ;
  assign n23983 = n12818 ^ n9725 ^ n4371 ;
  assign n23984 = ( n301 & n11786 ) | ( n301 & n23983 ) | ( n11786 & n23983 ) ;
  assign n23985 = ( n11488 & ~n12670 ) | ( n11488 & n23984 ) | ( ~n12670 & n23984 ) ;
  assign n23986 = ( n1083 & ~n12013 ) | ( n1083 & n12122 ) | ( ~n12013 & n12122 ) ;
  assign n23987 = n23986 ^ n4291 ^ n3678 ;
  assign n23988 = n23314 ^ n2624 ^ n319 ;
  assign n23989 = ( n3635 & n11143 ) | ( n3635 & ~n23988 ) | ( n11143 & ~n23988 ) ;
  assign n23990 = n13646 ^ n3305 ^ x76 ;
  assign n23991 = ( n9396 & ~n13778 ) | ( n9396 & n23990 ) | ( ~n13778 & n23990 ) ;
  assign n23992 = n22349 ^ n18322 ^ n6738 ;
  assign n23993 = n21393 ^ n17441 ^ n12312 ;
  assign n23994 = ( ~n8567 & n10149 ) | ( ~n8567 & n14819 ) | ( n10149 & n14819 ) ;
  assign n23995 = ( ~n515 & n3459 ) | ( ~n515 & n23994 ) | ( n3459 & n23994 ) ;
  assign n23996 = ( n2773 & n23993 ) | ( n2773 & n23995 ) | ( n23993 & n23995 ) ;
  assign n23997 = ( n2776 & n4988 ) | ( n2776 & n17945 ) | ( n4988 & n17945 ) ;
  assign n23998 = n23997 ^ n3587 ^ n1422 ;
  assign n23999 = ( n1181 & n5710 ) | ( n1181 & ~n11268 ) | ( n5710 & ~n11268 ) ;
  assign n24000 = n23999 ^ n22433 ^ n3579 ;
  assign n24001 = n22660 ^ n21585 ^ n16081 ;
  assign n24002 = n6890 ^ n6495 ^ n1931 ;
  assign n24003 = n24002 ^ n14248 ^ n1269 ;
  assign n24004 = n24003 ^ n5206 ^ n4899 ;
  assign n24005 = n24004 ^ n23144 ^ n5528 ;
  assign n24008 = n18753 ^ n12305 ^ n11088 ;
  assign n24006 = ( n3624 & n8159 ) | ( n3624 & n8875 ) | ( n8159 & n8875 ) ;
  assign n24007 = ( ~n12600 & n19402 ) | ( ~n12600 & n24006 ) | ( n19402 & n24006 ) ;
  assign n24009 = n24008 ^ n24007 ^ n18787 ;
  assign n24010 = n11871 ^ n4514 ^ n3878 ;
  assign n24011 = n24010 ^ n4553 ^ n1215 ;
  assign n24012 = ( n8767 & n13017 ) | ( n8767 & ~n15113 ) | ( n13017 & ~n15113 ) ;
  assign n24013 = n24012 ^ n21292 ^ n9415 ;
  assign n24014 = ( n2717 & n10009 ) | ( n2717 & ~n24013 ) | ( n10009 & ~n24013 ) ;
  assign n24015 = n24014 ^ n18660 ^ n9727 ;
  assign n24016 = ( n237 & n6057 ) | ( n237 & ~n7975 ) | ( n6057 & ~n7975 ) ;
  assign n24017 = n24016 ^ n4339 ^ n476 ;
  assign n24018 = n24017 ^ n16814 ^ n373 ;
  assign n24019 = n11071 ^ n8429 ^ n4783 ;
  assign n24020 = ( n1186 & n5959 ) | ( n1186 & n7891 ) | ( n5959 & n7891 ) ;
  assign n24021 = ( n19667 & ~n24019 ) | ( n19667 & n24020 ) | ( ~n24019 & n24020 ) ;
  assign n24022 = ( ~n4334 & n12560 ) | ( ~n4334 & n14595 ) | ( n12560 & n14595 ) ;
  assign n24023 = n24022 ^ n9499 ^ n4982 ;
  assign n24024 = n13510 ^ n12295 ^ n4135 ;
  assign n24025 = n17291 ^ n4551 ^ n1786 ;
  assign n24026 = n2885 ^ n1513 ^ n1410 ;
  assign n24027 = ( x102 & ~n5418 ) | ( x102 & n24026 ) | ( ~n5418 & n24026 ) ;
  assign n24029 = ( n2684 & ~n2818 ) | ( n2684 & n8100 ) | ( ~n2818 & n8100 ) ;
  assign n24030 = ( n12054 & n21304 ) | ( n12054 & n24029 ) | ( n21304 & n24029 ) ;
  assign n24028 = n7035 ^ n6183 ^ n643 ;
  assign n24031 = n24030 ^ n24028 ^ n16894 ;
  assign n24033 = ( ~n20242 & n20817 ) | ( ~n20242 & n21579 ) | ( n20817 & n21579 ) ;
  assign n24032 = ( ~n2539 & n7065 ) | ( ~n2539 & n20334 ) | ( n7065 & n20334 ) ;
  assign n24034 = n24033 ^ n24032 ^ n5071 ;
  assign n24038 = n7924 ^ n2229 ^ n325 ;
  assign n24036 = ( n259 & ~n3044 ) | ( n259 & n15102 ) | ( ~n3044 & n15102 ) ;
  assign n24037 = ( n4884 & n16710 ) | ( n4884 & ~n24036 ) | ( n16710 & ~n24036 ) ;
  assign n24039 = n24038 ^ n24037 ^ n9144 ;
  assign n24035 = ( n7552 & n8597 ) | ( n7552 & ~n13369 ) | ( n8597 & ~n13369 ) ;
  assign n24040 = n24039 ^ n24035 ^ n5566 ;
  assign n24041 = ( n4253 & n4510 ) | ( n4253 & ~n19650 ) | ( n4510 & ~n19650 ) ;
  assign n24042 = ( ~n895 & n21108 ) | ( ~n895 & n21242 ) | ( n21108 & n21242 ) ;
  assign n24043 = n24042 ^ n21359 ^ n19055 ;
  assign n24044 = n24043 ^ n21357 ^ x43 ;
  assign n24045 = ( n6805 & n6975 ) | ( n6805 & n21295 ) | ( n6975 & n21295 ) ;
  assign n24046 = n16821 ^ n4518 ^ n1786 ;
  assign n24047 = ( n3443 & ~n4509 ) | ( n3443 & n17289 ) | ( ~n4509 & n17289 ) ;
  assign n24048 = ( n21455 & n24046 ) | ( n21455 & n24047 ) | ( n24046 & n24047 ) ;
  assign n24049 = ( n4328 & ~n4598 ) | ( n4328 & n10570 ) | ( ~n4598 & n10570 ) ;
  assign n24050 = n16660 ^ n15328 ^ n7134 ;
  assign n24051 = ( ~n23586 & n24049 ) | ( ~n23586 & n24050 ) | ( n24049 & n24050 ) ;
  assign n24052 = ( n1025 & n4137 ) | ( n1025 & n18983 ) | ( n4137 & n18983 ) ;
  assign n24053 = ( n7485 & n8315 ) | ( n7485 & n9877 ) | ( n8315 & n9877 ) ;
  assign n24055 = ( n2696 & n12013 ) | ( n2696 & ~n12583 ) | ( n12013 & ~n12583 ) ;
  assign n24054 = n17022 ^ n9651 ^ n8892 ;
  assign n24056 = n24055 ^ n24054 ^ n3429 ;
  assign n24057 = ( ~n21714 & n24053 ) | ( ~n21714 & n24056 ) | ( n24053 & n24056 ) ;
  assign n24058 = n7497 ^ n5771 ^ n3023 ;
  assign n24059 = n24058 ^ n10856 ^ n10368 ;
  assign n24060 = n24059 ^ n11245 ^ n7962 ;
  assign n24061 = n24060 ^ n19747 ^ n5859 ;
  assign n24062 = n3551 ^ n3311 ^ n1638 ;
  assign n24063 = ( n1558 & ~n6573 ) | ( n1558 & n24062 ) | ( ~n6573 & n24062 ) ;
  assign n24064 = n17093 ^ n2691 ^ n679 ;
  assign n24065 = n24064 ^ n18894 ^ n1713 ;
  assign n24066 = ( n1792 & n9000 ) | ( n1792 & ~n20478 ) | ( n9000 & ~n20478 ) ;
  assign n24067 = n9161 ^ n6714 ^ n3565 ;
  assign n24068 = n24067 ^ n21476 ^ n16188 ;
  assign n24069 = n24068 ^ n18429 ^ n3238 ;
  assign n24070 = ( ~n9373 & n17104 ) | ( ~n9373 & n24069 ) | ( n17104 & n24069 ) ;
  assign n24071 = ( n9685 & n15355 ) | ( n9685 & n19905 ) | ( n15355 & n19905 ) ;
  assign n24072 = n24071 ^ n2287 ^ n1769 ;
  assign n24073 = ( x73 & n312 ) | ( x73 & ~n3183 ) | ( n312 & ~n3183 ) ;
  assign n24074 = ( n1641 & ~n9238 ) | ( n1641 & n24073 ) | ( ~n9238 & n24073 ) ;
  assign n24075 = n17093 ^ n13124 ^ n7797 ;
  assign n24076 = n24075 ^ n11172 ^ n5873 ;
  assign n24077 = n14932 ^ n4603 ^ n3278 ;
  assign n24078 = n24077 ^ n16689 ^ n8077 ;
  assign n24079 = n24078 ^ n20237 ^ n10202 ;
  assign n24080 = ( n1557 & ~n24076 ) | ( n1557 & n24079 ) | ( ~n24076 & n24079 ) ;
  assign n24081 = ( n16652 & ~n24074 ) | ( n16652 & n24080 ) | ( ~n24074 & n24080 ) ;
  assign n24082 = n6419 ^ n3404 ^ n2976 ;
  assign n24083 = ( n650 & n6283 ) | ( n650 & ~n19065 ) | ( n6283 & ~n19065 ) ;
  assign n24084 = ( ~n657 & n3184 ) | ( ~n657 & n20743 ) | ( n3184 & n20743 ) ;
  assign n24085 = ( n24082 & n24083 ) | ( n24082 & ~n24084 ) | ( n24083 & ~n24084 ) ;
  assign n24086 = ( n1020 & n3447 ) | ( n1020 & ~n19669 ) | ( n3447 & ~n19669 ) ;
  assign n24087 = ( ~n3656 & n4651 ) | ( ~n3656 & n24086 ) | ( n4651 & n24086 ) ;
  assign n24088 = ( x28 & ~n15708 ) | ( x28 & n24087 ) | ( ~n15708 & n24087 ) ;
  assign n24089 = ( ~n4378 & n10556 ) | ( ~n4378 & n24088 ) | ( n10556 & n24088 ) ;
  assign n24090 = ( n1985 & n4856 ) | ( n1985 & n13801 ) | ( n4856 & n13801 ) ;
  assign n24091 = ( n12121 & n14543 ) | ( n12121 & n24090 ) | ( n14543 & n24090 ) ;
  assign n24092 = ( n15379 & ~n20647 ) | ( n15379 & n22571 ) | ( ~n20647 & n22571 ) ;
  assign n24093 = ( n21548 & ~n24091 ) | ( n21548 & n24092 ) | ( ~n24091 & n24092 ) ;
  assign n24094 = n13334 ^ n11572 ^ n9938 ;
  assign n24095 = ( n502 & n8825 ) | ( n502 & ~n24094 ) | ( n8825 & ~n24094 ) ;
  assign n24096 = ( n9905 & n16352 ) | ( n9905 & ~n24095 ) | ( n16352 & ~n24095 ) ;
  assign n24097 = ( n5581 & n16917 ) | ( n5581 & ~n22737 ) | ( n16917 & ~n22737 ) ;
  assign n24098 = n7793 ^ n2580 ^ n2521 ;
  assign n24099 = ( n8990 & ~n24097 ) | ( n8990 & n24098 ) | ( ~n24097 & n24098 ) ;
  assign n24100 = ( ~n170 & n20468 ) | ( ~n170 & n24099 ) | ( n20468 & n24099 ) ;
  assign n24101 = ( n4486 & ~n6464 ) | ( n4486 & n14344 ) | ( ~n6464 & n14344 ) ;
  assign n24102 = ( n17580 & ~n21072 ) | ( n17580 & n24101 ) | ( ~n21072 & n24101 ) ;
  assign n24103 = n12742 ^ n12125 ^ n3203 ;
  assign n24104 = n24103 ^ n10659 ^ n8515 ;
  assign n24105 = n24104 ^ n973 ^ n539 ;
  assign n24106 = n23434 ^ n22223 ^ n11023 ;
  assign n24107 = ( n5495 & ~n16206 ) | ( n5495 & n23621 ) | ( ~n16206 & n23621 ) ;
  assign n24108 = ( ~n2388 & n24106 ) | ( ~n2388 & n24107 ) | ( n24106 & n24107 ) ;
  assign n24109 = ( n7672 & ~n10377 ) | ( n7672 & n14698 ) | ( ~n10377 & n14698 ) ;
  assign n24110 = n19304 ^ n14294 ^ n1787 ;
  assign n24111 = ( n21545 & n24109 ) | ( n21545 & n24110 ) | ( n24109 & n24110 ) ;
  assign n24112 = ( n1569 & ~n24108 ) | ( n1569 & n24111 ) | ( ~n24108 & n24111 ) ;
  assign n24113 = ( n2428 & ~n14273 ) | ( n2428 & n18765 ) | ( ~n14273 & n18765 ) ;
  assign n24114 = n24113 ^ n18300 ^ n13980 ;
  assign n24115 = n15046 ^ n3169 ^ x72 ;
  assign n24116 = ( n9170 & n15008 ) | ( n9170 & ~n24115 ) | ( n15008 & ~n24115 ) ;
  assign n24117 = n23031 ^ n10750 ^ n7818 ;
  assign n24118 = n22955 ^ n1744 ^ n256 ;
  assign n24119 = ( n4551 & ~n11155 ) | ( n4551 & n24118 ) | ( ~n11155 & n24118 ) ;
  assign n24120 = n10466 ^ n4052 ^ n3312 ;
  assign n24121 = ( x69 & n9826 ) | ( x69 & ~n24120 ) | ( n9826 & ~n24120 ) ;
  assign n24122 = n24121 ^ n18527 ^ n7525 ;
  assign n24123 = ( n12177 & n19849 ) | ( n12177 & ~n23497 ) | ( n19849 & ~n23497 ) ;
  assign n24124 = ( n3641 & ~n5675 ) | ( n3641 & n24123 ) | ( ~n5675 & n24123 ) ;
  assign n24125 = ( ~n2143 & n2943 ) | ( ~n2143 & n13063 ) | ( n2943 & n13063 ) ;
  assign n24126 = n21730 ^ n12660 ^ n2019 ;
  assign n24127 = ( n11084 & ~n22068 ) | ( n11084 & n24126 ) | ( ~n22068 & n24126 ) ;
  assign n24128 = ( n7987 & n24125 ) | ( n7987 & ~n24127 ) | ( n24125 & ~n24127 ) ;
  assign n24129 = n1883 ^ n1773 ^ n171 ;
  assign n24130 = ( n6301 & n16311 ) | ( n6301 & n24129 ) | ( n16311 & n24129 ) ;
  assign n24131 = ( n783 & n12877 ) | ( n783 & ~n14390 ) | ( n12877 & ~n14390 ) ;
  assign n24132 = ( n405 & ~n2096 ) | ( n405 & n4212 ) | ( ~n2096 & n4212 ) ;
  assign n24133 = ( n6959 & ~n13506 ) | ( n6959 & n24132 ) | ( ~n13506 & n24132 ) ;
  assign n24134 = ( ~n12379 & n13027 ) | ( ~n12379 & n19883 ) | ( n13027 & n19883 ) ;
  assign n24135 = n24134 ^ n19038 ^ n8678 ;
  assign n24136 = ( n346 & ~n3788 ) | ( n346 & n18526 ) | ( ~n3788 & n18526 ) ;
  assign n24137 = ( n15014 & n24135 ) | ( n15014 & n24136 ) | ( n24135 & n24136 ) ;
  assign n24138 = ( n451 & ~n3882 ) | ( n451 & n19246 ) | ( ~n3882 & n19246 ) ;
  assign n24139 = ( n9982 & ~n12386 ) | ( n9982 & n19830 ) | ( ~n12386 & n19830 ) ;
  assign n24140 = ( n2388 & ~n5632 ) | ( n2388 & n17442 ) | ( ~n5632 & n17442 ) ;
  assign n24141 = ( ~n788 & n10477 ) | ( ~n788 & n24140 ) | ( n10477 & n24140 ) ;
  assign n24142 = ( n13850 & ~n19218 ) | ( n13850 & n24141 ) | ( ~n19218 & n24141 ) ;
  assign n24143 = ( n11137 & ~n19916 ) | ( n11137 & n23784 ) | ( ~n19916 & n23784 ) ;
  assign n24144 = n4630 ^ n3278 ^ n696 ;
  assign n24145 = n17630 ^ n10863 ^ n945 ;
  assign n24146 = n24145 ^ n23148 ^ n160 ;
  assign n24147 = ( n1532 & n3742 ) | ( n1532 & ~n22171 ) | ( n3742 & ~n22171 ) ;
  assign n24148 = n19966 ^ n12937 ^ n2712 ;
  assign n24149 = ( n2577 & n4097 ) | ( n2577 & n13670 ) | ( n4097 & n13670 ) ;
  assign n24150 = ( n15617 & ~n19048 ) | ( n15617 & n24149 ) | ( ~n19048 & n24149 ) ;
  assign n24151 = n22467 ^ n21644 ^ n6045 ;
  assign n24152 = ( n21409 & n23172 ) | ( n21409 & n24151 ) | ( n23172 & n24151 ) ;
  assign n24153 = n21437 ^ n18602 ^ n5510 ;
  assign n24154 = ( n3272 & n8629 ) | ( n3272 & ~n11141 ) | ( n8629 & ~n11141 ) ;
  assign n24155 = n24154 ^ n19390 ^ n18961 ;
  assign n24156 = n18478 ^ n15115 ^ n13891 ;
  assign n24157 = ( n3250 & ~n19255 ) | ( n3250 & n24156 ) | ( ~n19255 & n24156 ) ;
  assign n24158 = ( n16633 & n24155 ) | ( n16633 & n24157 ) | ( n24155 & n24157 ) ;
  assign n24163 = ( n4682 & ~n7364 ) | ( n4682 & n17899 ) | ( ~n7364 & n17899 ) ;
  assign n24159 = n11769 ^ n11247 ^ n1141 ;
  assign n24160 = ( n6425 & ~n12528 ) | ( n6425 & n18986 ) | ( ~n12528 & n18986 ) ;
  assign n24161 = ( n4374 & ~n24159 ) | ( n4374 & n24160 ) | ( ~n24159 & n24160 ) ;
  assign n24162 = n24161 ^ n7130 ^ n6997 ;
  assign n24164 = n24163 ^ n24162 ^ n19227 ;
  assign n24165 = n24164 ^ n22186 ^ n15421 ;
  assign n24166 = ( n6280 & n7364 ) | ( n6280 & n13312 ) | ( n7364 & n13312 ) ;
  assign n24167 = n24166 ^ n20458 ^ n12756 ;
  assign n24168 = ( ~n5303 & n23768 ) | ( ~n5303 & n24167 ) | ( n23768 & n24167 ) ;
  assign n24169 = n18187 ^ n6015 ^ n5556 ;
  assign n24170 = n12225 ^ n9852 ^ n1756 ;
  assign n24171 = ( n9999 & n15076 ) | ( n9999 & n23686 ) | ( n15076 & n23686 ) ;
  assign n24172 = ( n3887 & n17403 ) | ( n3887 & ~n24171 ) | ( n17403 & ~n24171 ) ;
  assign n24173 = ( n8084 & ~n13132 ) | ( n8084 & n21007 ) | ( ~n13132 & n21007 ) ;
  assign n24174 = n24173 ^ n10803 ^ n2882 ;
  assign n24176 = ( n3783 & n5025 ) | ( n3783 & ~n19055 ) | ( n5025 & ~n19055 ) ;
  assign n24175 = ( n1352 & ~n21698 ) | ( n1352 & n22269 ) | ( ~n21698 & n22269 ) ;
  assign n24177 = n24176 ^ n24175 ^ n9480 ;
  assign n24178 = n17877 ^ n3717 ^ n256 ;
  assign n24179 = n24178 ^ n8889 ^ n593 ;
  assign n24180 = n20893 ^ n15045 ^ n2464 ;
  assign n24181 = n24180 ^ n11069 ^ n6645 ;
  assign n24182 = ( n421 & n19443 ) | ( n421 & n24181 ) | ( n19443 & n24181 ) ;
  assign n24183 = ( ~n15039 & n18336 ) | ( ~n15039 & n20096 ) | ( n18336 & n20096 ) ;
  assign n24184 = ( n12447 & n12497 ) | ( n12447 & ~n20160 ) | ( n12497 & ~n20160 ) ;
  assign n24185 = n21274 ^ n14369 ^ n11053 ;
  assign n24186 = n23408 ^ n8395 ^ n5512 ;
  assign n24187 = n8349 ^ n6615 ^ n2368 ;
  assign n24188 = n24187 ^ n20398 ^ n15724 ;
  assign n24190 = ( n5886 & n7379 ) | ( n5886 & n21831 ) | ( n7379 & n21831 ) ;
  assign n24189 = n18955 ^ n7715 ^ n6579 ;
  assign n24191 = n24190 ^ n24189 ^ n2539 ;
  assign n24192 = n11702 ^ n7794 ^ n6360 ;
  assign n24193 = n23691 ^ n20871 ^ n3493 ;
  assign n24194 = n24193 ^ n22224 ^ n3259 ;
  assign n24195 = ( n1306 & ~n7199 ) | ( n1306 & n12571 ) | ( ~n7199 & n12571 ) ;
  assign n24196 = ( ~n11923 & n23902 ) | ( ~n11923 & n24195 ) | ( n23902 & n24195 ) ;
  assign n24197 = ( ~n1198 & n6157 ) | ( ~n1198 & n8421 ) | ( n6157 & n8421 ) ;
  assign n24198 = n24197 ^ n10491 ^ n9081 ;
  assign n24199 = n6136 ^ n2678 ^ n2006 ;
  assign n24200 = ( ~n4213 & n24198 ) | ( ~n4213 & n24199 ) | ( n24198 & n24199 ) ;
  assign n24201 = ( n1940 & ~n13388 ) | ( n1940 & n18654 ) | ( ~n13388 & n18654 ) ;
  assign n24202 = ( n24196 & n24200 ) | ( n24196 & ~n24201 ) | ( n24200 & ~n24201 ) ;
  assign n24207 = n20454 ^ n5866 ^ n1532 ;
  assign n24205 = ( n2753 & ~n2860 ) | ( n2753 & n5336 ) | ( ~n2860 & n5336 ) ;
  assign n24203 = ( n2461 & ~n10731 ) | ( n2461 & n13277 ) | ( ~n10731 & n13277 ) ;
  assign n24204 = ( n9095 & ~n9421 ) | ( n9095 & n24203 ) | ( ~n9421 & n24203 ) ;
  assign n24206 = n24205 ^ n24204 ^ n20109 ;
  assign n24208 = n24207 ^ n24206 ^ n7378 ;
  assign n24209 = ( n9489 & n10596 ) | ( n9489 & n14031 ) | ( n10596 & n14031 ) ;
  assign n24210 = ( n10224 & n13939 ) | ( n10224 & n16063 ) | ( n13939 & n16063 ) ;
  assign n24211 = ( n14344 & ~n15346 ) | ( n14344 & n20301 ) | ( ~n15346 & n20301 ) ;
  assign n24212 = ( n1070 & ~n14660 ) | ( n1070 & n24211 ) | ( ~n14660 & n24211 ) ;
  assign n24213 = n8137 ^ n5406 ^ n1441 ;
  assign n24214 = n6270 ^ n2633 ^ n2017 ;
  assign n24215 = n24214 ^ n17483 ^ n752 ;
  assign n24216 = n24215 ^ n13366 ^ n13138 ;
  assign n24217 = ( n1627 & ~n3051 ) | ( n1627 & n24216 ) | ( ~n3051 & n24216 ) ;
  assign n24218 = ( n12355 & ~n24213 ) | ( n12355 & n24217 ) | ( ~n24213 & n24217 ) ;
  assign n24219 = ( n748 & n1922 ) | ( n748 & ~n2696 ) | ( n1922 & ~n2696 ) ;
  assign n24220 = n24219 ^ n12107 ^ n399 ;
  assign n24221 = ( n8012 & n13932 ) | ( n8012 & n16335 ) | ( n13932 & n16335 ) ;
  assign n24222 = n24221 ^ n11580 ^ n1212 ;
  assign n24223 = n24222 ^ n20208 ^ n19170 ;
  assign n24224 = ( n587 & ~n10248 ) | ( n587 & n23373 ) | ( ~n10248 & n23373 ) ;
  assign n24225 = n9718 ^ n6659 ^ n5491 ;
  assign n24226 = ( ~n16684 & n17399 ) | ( ~n16684 & n24225 ) | ( n17399 & n24225 ) ;
  assign n24227 = n18761 ^ n14922 ^ n10931 ;
  assign n24228 = ( ~n19249 & n20582 ) | ( ~n19249 & n23067 ) | ( n20582 & n23067 ) ;
  assign n24229 = ( ~n7724 & n7838 ) | ( ~n7724 & n16561 ) | ( n7838 & n16561 ) ;
  assign n24230 = n10468 ^ n3763 ^ n3357 ;
  assign n24233 = n11422 ^ n7958 ^ n7874 ;
  assign n24231 = n6735 ^ n3189 ^ n566 ;
  assign n24232 = ( n7558 & n24134 ) | ( n7558 & ~n24231 ) | ( n24134 & ~n24231 ) ;
  assign n24234 = n24233 ^ n24232 ^ n9549 ;
  assign n24235 = ( n6132 & n24230 ) | ( n6132 & ~n24234 ) | ( n24230 & ~n24234 ) ;
  assign n24236 = n11965 ^ n9459 ^ n6055 ;
  assign n24237 = n24236 ^ n4046 ^ n1002 ;
  assign n24238 = ( n601 & n1673 ) | ( n601 & n8490 ) | ( n1673 & n8490 ) ;
  assign n24239 = ( n14768 & n17186 ) | ( n14768 & ~n24238 ) | ( n17186 & ~n24238 ) ;
  assign n24240 = n16988 ^ n2462 ^ n600 ;
  assign n24241 = n24240 ^ n14790 ^ n3421 ;
  assign n24242 = ( n3582 & ~n13999 ) | ( n3582 & n24241 ) | ( ~n13999 & n24241 ) ;
  assign n24243 = ( n3795 & ~n10647 ) | ( n3795 & n24242 ) | ( ~n10647 & n24242 ) ;
  assign n24244 = ( ~n5254 & n7426 ) | ( ~n5254 & n19338 ) | ( n7426 & n19338 ) ;
  assign n24245 = ( ~n1369 & n2605 ) | ( ~n1369 & n24244 ) | ( n2605 & n24244 ) ;
  assign n24246 = n24245 ^ n13821 ^ n5105 ;
  assign n24247 = ( n1138 & ~n14872 ) | ( n1138 & n22906 ) | ( ~n14872 & n22906 ) ;
  assign n24248 = n16257 ^ n14558 ^ n1893 ;
  assign n24249 = ( n3814 & n4609 ) | ( n3814 & ~n24248 ) | ( n4609 & ~n24248 ) ;
  assign n24252 = n2590 ^ n1066 ^ n311 ;
  assign n24253 = ( ~n13379 & n14485 ) | ( ~n13379 & n24252 ) | ( n14485 & n24252 ) ;
  assign n24254 = n24253 ^ n7669 ^ n1308 ;
  assign n24251 = ( ~n5174 & n7750 ) | ( ~n5174 & n10224 ) | ( n7750 & n10224 ) ;
  assign n24255 = n24254 ^ n24251 ^ n1371 ;
  assign n24250 = ( ~n683 & n4066 ) | ( ~n683 & n15343 ) | ( n4066 & n15343 ) ;
  assign n24256 = n24255 ^ n24250 ^ n1575 ;
  assign n24257 = n17799 ^ n10426 ^ n6704 ;
  assign n24258 = ( n387 & ~n23389 ) | ( n387 & n24257 ) | ( ~n23389 & n24257 ) ;
  assign n24259 = ( ~n11806 & n14943 ) | ( ~n11806 & n24258 ) | ( n14943 & n24258 ) ;
  assign n24260 = ( n5390 & n10043 ) | ( n5390 & ~n22236 ) | ( n10043 & ~n22236 ) ;
  assign n24261 = ( n4993 & n5456 ) | ( n4993 & n24260 ) | ( n5456 & n24260 ) ;
  assign n24262 = n15424 ^ n9424 ^ n2269 ;
  assign n24263 = n24262 ^ n9277 ^ n5047 ;
  assign n24264 = n12326 ^ n4536 ^ n1523 ;
  assign n24265 = ( n155 & n3912 ) | ( n155 & n24264 ) | ( n3912 & n24264 ) ;
  assign n24266 = n6973 ^ n563 ^ x86 ;
  assign n24267 = n14714 ^ n10829 ^ n7491 ;
  assign n24271 = ( ~n188 & n862 ) | ( ~n188 & n21433 ) | ( n862 & n21433 ) ;
  assign n24268 = ( n10098 & n11571 ) | ( n10098 & ~n14169 ) | ( n11571 & ~n14169 ) ;
  assign n24269 = n24268 ^ n21628 ^ n8466 ;
  assign n24270 = ( ~x60 & n17092 ) | ( ~x60 & n24269 ) | ( n17092 & n24269 ) ;
  assign n24272 = n24271 ^ n24270 ^ n13891 ;
  assign n24273 = ( ~n3678 & n17498 ) | ( ~n3678 & n23962 ) | ( n17498 & n23962 ) ;
  assign n24274 = ( ~n4450 & n7042 ) | ( ~n4450 & n18894 ) | ( n7042 & n18894 ) ;
  assign n24275 = ( n2793 & n19527 ) | ( n2793 & n24274 ) | ( n19527 & n24274 ) ;
  assign n24276 = n16300 ^ n3196 ^ n1721 ;
  assign n24277 = ( n24273 & ~n24275 ) | ( n24273 & n24276 ) | ( ~n24275 & n24276 ) ;
  assign n24278 = ( n188 & ~n1076 ) | ( n188 & n17383 ) | ( ~n1076 & n17383 ) ;
  assign n24279 = ( n10583 & n14359 ) | ( n10583 & ~n21763 ) | ( n14359 & ~n21763 ) ;
  assign n24280 = n17597 ^ n7576 ^ n4416 ;
  assign n24281 = ( n4248 & ~n22766 ) | ( n4248 & n24280 ) | ( ~n22766 & n24280 ) ;
  assign n24282 = ( ~n314 & n4302 ) | ( ~n314 & n12421 ) | ( n4302 & n12421 ) ;
  assign n24283 = ( n3607 & n5718 ) | ( n3607 & n24282 ) | ( n5718 & n24282 ) ;
  assign n24284 = ( n7281 & n21618 ) | ( n7281 & ~n24283 ) | ( n21618 & ~n24283 ) ;
  assign n24285 = n19852 ^ n14997 ^ n5522 ;
  assign n24286 = ( n15232 & n24284 ) | ( n15232 & n24285 ) | ( n24284 & n24285 ) ;
  assign n24289 = ( n4179 & n6068 ) | ( n4179 & ~n7168 ) | ( n6068 & ~n7168 ) ;
  assign n24288 = ( n3381 & ~n7025 ) | ( n3381 & n11078 ) | ( ~n7025 & n11078 ) ;
  assign n24287 = n5406 ^ n5231 ^ n3961 ;
  assign n24290 = n24289 ^ n24288 ^ n24287 ;
  assign n24291 = ( ~n1741 & n2637 ) | ( ~n1741 & n7912 ) | ( n2637 & n7912 ) ;
  assign n24292 = ( n1142 & ~n16546 ) | ( n1142 & n24291 ) | ( ~n16546 & n24291 ) ;
  assign n24293 = ( n11380 & ~n16471 ) | ( n11380 & n24292 ) | ( ~n16471 & n24292 ) ;
  assign n24294 = ( n1133 & n7246 ) | ( n1133 & ~n23148 ) | ( n7246 & ~n23148 ) ;
  assign n24295 = n24294 ^ n19104 ^ n8818 ;
  assign n24296 = n24295 ^ n8089 ^ n3336 ;
  assign n24297 = n24296 ^ n15062 ^ n5558 ;
  assign n24298 = n24297 ^ n16436 ^ n9605 ;
  assign n24299 = n18527 ^ n6464 ^ n4455 ;
  assign n24300 = n24299 ^ n6850 ^ n3119 ;
  assign n24301 = ( ~n6699 & n15724 ) | ( ~n6699 & n24300 ) | ( n15724 & n24300 ) ;
  assign n24302 = ( n220 & n13221 ) | ( n220 & ~n17932 ) | ( n13221 & ~n17932 ) ;
  assign n24303 = n24302 ^ n23946 ^ n3618 ;
  assign n24304 = ( n2683 & n6788 ) | ( n2683 & ~n10401 ) | ( n6788 & ~n10401 ) ;
  assign n24305 = ( ~n7377 & n7940 ) | ( ~n7377 & n20231 ) | ( n7940 & n20231 ) ;
  assign n24306 = ( ~n12351 & n24304 ) | ( ~n12351 & n24305 ) | ( n24304 & n24305 ) ;
  assign n24307 = ( n652 & ~n3170 ) | ( n652 & n3648 ) | ( ~n3170 & n3648 ) ;
  assign n24308 = ( n929 & ~n10667 ) | ( n929 & n13198 ) | ( ~n10667 & n13198 ) ;
  assign n24309 = ( n12008 & n24307 ) | ( n12008 & ~n24308 ) | ( n24307 & ~n24308 ) ;
  assign n24310 = ( ~n8129 & n15792 ) | ( ~n8129 & n19377 ) | ( n15792 & n19377 ) ;
  assign n24311 = ( n11428 & n19343 ) | ( n11428 & n19631 ) | ( n19343 & n19631 ) ;
  assign n24312 = n4715 ^ n3389 ^ n3009 ;
  assign n24313 = ( ~n12916 & n21251 ) | ( ~n12916 & n24312 ) | ( n21251 & n24312 ) ;
  assign n24314 = ( n985 & n7347 ) | ( n985 & n24313 ) | ( n7347 & n24313 ) ;
  assign n24315 = ( x106 & n4641 ) | ( x106 & n22847 ) | ( n4641 & n22847 ) ;
  assign n24316 = n24315 ^ n14803 ^ n9162 ;
  assign n24317 = n24316 ^ n22827 ^ n14451 ;
  assign n24318 = ( ~n3497 & n6665 ) | ( ~n3497 & n13705 ) | ( n6665 & n13705 ) ;
  assign n24319 = n24318 ^ n18781 ^ n15353 ;
  assign n24320 = ( ~n243 & n3562 ) | ( ~n243 & n24319 ) | ( n3562 & n24319 ) ;
  assign n24321 = n24320 ^ n8378 ^ n5527 ;
  assign n24322 = n24321 ^ n18883 ^ n2176 ;
  assign n24323 = n21279 ^ n462 ^ n336 ;
  assign n24324 = n24323 ^ n23726 ^ n12570 ;
  assign n24325 = n24026 ^ n21174 ^ n10764 ;
  assign n24326 = ( ~n10038 & n12720 ) | ( ~n10038 & n20948 ) | ( n12720 & n20948 ) ;
  assign n24327 = n14061 ^ n11935 ^ n2196 ;
  assign n24328 = n8920 ^ n5846 ^ n3028 ;
  assign n24329 = n8554 ^ n3776 ^ n3641 ;
  assign n24330 = ( n403 & n3760 ) | ( n403 & n11313 ) | ( n3760 & n11313 ) ;
  assign n24331 = ( ~n3982 & n13715 ) | ( ~n3982 & n24330 ) | ( n13715 & n24330 ) ;
  assign n24332 = n20756 ^ n16531 ^ n11741 ;
  assign n24333 = n17305 ^ n13277 ^ n2378 ;
  assign n24334 = n20174 ^ n17098 ^ n1254 ;
  assign n24335 = n16693 ^ n12790 ^ n5674 ;
  assign n24336 = ( ~n6173 & n9004 ) | ( ~n6173 & n24335 ) | ( n9004 & n24335 ) ;
  assign n24337 = ( n17314 & ~n19079 ) | ( n17314 & n24336 ) | ( ~n19079 & n24336 ) ;
  assign n24338 = n20821 ^ n8771 ^ n1139 ;
  assign n24340 = ( x6 & n635 ) | ( x6 & n832 ) | ( n635 & n832 ) ;
  assign n24339 = ( n2906 & n5777 ) | ( n2906 & n12973 ) | ( n5777 & n12973 ) ;
  assign n24341 = n24340 ^ n24339 ^ n3441 ;
  assign n24342 = n12591 ^ n11051 ^ n3352 ;
  assign n24343 = ( ~n5105 & n5607 ) | ( ~n5105 & n13012 ) | ( n5607 & n13012 ) ;
  assign n24344 = n24343 ^ n16668 ^ n5313 ;
  assign n24345 = n24344 ^ n12131 ^ n1593 ;
  assign n24346 = n22050 ^ n9153 ^ n2022 ;
  assign n24348 = n22023 ^ n8823 ^ n1521 ;
  assign n24347 = ( ~n18264 & n20185 ) | ( ~n18264 & n20693 ) | ( n20185 & n20693 ) ;
  assign n24349 = n24348 ^ n24347 ^ n4553 ;
  assign n24350 = n9082 ^ n7443 ^ n2866 ;
  assign n24351 = ( n1105 & n2125 ) | ( n1105 & n10475 ) | ( n2125 & n10475 ) ;
  assign n24352 = n24351 ^ n20280 ^ n8783 ;
  assign n24353 = ( ~n7528 & n21165 ) | ( ~n7528 & n24352 ) | ( n21165 & n24352 ) ;
  assign n24354 = n7043 ^ n4422 ^ n1203 ;
  assign n24355 = n24354 ^ n16486 ^ n12942 ;
  assign n24356 = n24355 ^ n16264 ^ n4250 ;
  assign n24357 = ( ~n4449 & n8298 ) | ( ~n4449 & n13446 ) | ( n8298 & n13446 ) ;
  assign n24358 = ( n14052 & n24356 ) | ( n14052 & ~n24357 ) | ( n24356 & ~n24357 ) ;
  assign n24359 = ( ~n24350 & n24353 ) | ( ~n24350 & n24358 ) | ( n24353 & n24358 ) ;
  assign n24360 = ( n180 & n7019 ) | ( n180 & ~n8564 ) | ( n7019 & ~n8564 ) ;
  assign n24361 = n24360 ^ n14129 ^ n7023 ;
  assign n24362 = ( n1189 & n2487 ) | ( n1189 & ~n24361 ) | ( n2487 & ~n24361 ) ;
  assign n24363 = n24362 ^ n24240 ^ n2323 ;
  assign n24364 = ( ~n1865 & n5363 ) | ( ~n1865 & n24363 ) | ( n5363 & n24363 ) ;
  assign n24365 = ( n1306 & ~n8564 ) | ( n1306 & n24364 ) | ( ~n8564 & n24364 ) ;
  assign n24366 = ( n6025 & n7610 ) | ( n6025 & ~n8239 ) | ( n7610 & ~n8239 ) ;
  assign n24367 = ( n14230 & ~n15940 ) | ( n14230 & n24366 ) | ( ~n15940 & n24366 ) ;
  assign n24368 = ( n1186 & n2689 ) | ( n1186 & ~n5686 ) | ( n2689 & ~n5686 ) ;
  assign n24369 = n24368 ^ n14426 ^ n9160 ;
  assign n24370 = n16303 ^ n9009 ^ n5438 ;
  assign n24371 = n24370 ^ n18446 ^ n1229 ;
  assign n24372 = ( ~n12281 & n13430 ) | ( ~n12281 & n24371 ) | ( n13430 & n24371 ) ;
  assign n24373 = ( n13916 & n15184 ) | ( n13916 & ~n19072 ) | ( n15184 & ~n19072 ) ;
  assign n24374 = ( n2258 & n6196 ) | ( n2258 & n8088 ) | ( n6196 & n8088 ) ;
  assign n24375 = n24374 ^ n15034 ^ n4569 ;
  assign n24376 = n17635 ^ n8767 ^ n7962 ;
  assign n24378 = n3836 ^ n1066 ^ n295 ;
  assign n24377 = ( ~n848 & n11580 ) | ( ~n848 & n19524 ) | ( n11580 & n19524 ) ;
  assign n24379 = n24378 ^ n24377 ^ n23299 ;
  assign n24380 = n17969 ^ n7528 ^ n5190 ;
  assign n24381 = n24380 ^ n10586 ^ n7528 ;
  assign n24382 = ( ~n6191 & n16599 ) | ( ~n6191 & n24381 ) | ( n16599 & n24381 ) ;
  assign n24383 = ( n10255 & n12232 ) | ( n10255 & ~n16672 ) | ( n12232 & ~n16672 ) ;
  assign n24384 = n10827 ^ n9289 ^ n512 ;
  assign n24385 = n24384 ^ n19802 ^ n15537 ;
  assign n24386 = n10491 ^ n8555 ^ n2658 ;
  assign n24387 = ( n9056 & ~n11000 ) | ( n9056 & n24386 ) | ( ~n11000 & n24386 ) ;
  assign n24388 = ( ~n3055 & n11639 ) | ( ~n3055 & n24387 ) | ( n11639 & n24387 ) ;
  assign n24389 = ( n5541 & n15206 ) | ( n5541 & n24388 ) | ( n15206 & n24388 ) ;
  assign n24391 = n11791 ^ n2818 ^ n940 ;
  assign n24390 = n13055 ^ n10433 ^ n8484 ;
  assign n24392 = n24391 ^ n24390 ^ n2531 ;
  assign n24393 = n20027 ^ n4490 ^ n4466 ;
  assign n24394 = n10315 ^ n5390 ^ n1931 ;
  assign n24395 = n24394 ^ n23749 ^ n16943 ;
  assign n24399 = n9220 ^ n7509 ^ n5527 ;
  assign n24397 = ( ~n1065 & n1416 ) | ( ~n1065 & n10685 ) | ( n1416 & n10685 ) ;
  assign n24398 = n24397 ^ n23881 ^ n6889 ;
  assign n24396 = ( n2324 & n2901 ) | ( n2324 & ~n20733 ) | ( n2901 & ~n20733 ) ;
  assign n24400 = n24399 ^ n24398 ^ n24396 ;
  assign n24401 = n2749 ^ n2597 ^ n2516 ;
  assign n24402 = ( n2674 & ~n3579 ) | ( n2674 & n11933 ) | ( ~n3579 & n11933 ) ;
  assign n24403 = ( n9346 & ~n16268 ) | ( n9346 & n23966 ) | ( ~n16268 & n23966 ) ;
  assign n24404 = ( ~n2014 & n24402 ) | ( ~n2014 & n24403 ) | ( n24402 & n24403 ) ;
  assign n24405 = n20674 ^ n15818 ^ n4520 ;
  assign n24406 = n21974 ^ n6673 ^ n1052 ;
  assign n24407 = n16526 ^ n16075 ^ n6304 ;
  assign n24408 = ( n6393 & ~n7095 ) | ( n6393 & n16662 ) | ( ~n7095 & n16662 ) ;
  assign n24409 = n24408 ^ n19796 ^ n6926 ;
  assign n24410 = ( n10048 & ~n19382 ) | ( n10048 & n24409 ) | ( ~n19382 & n24409 ) ;
  assign n24412 = n16638 ^ n12536 ^ n3775 ;
  assign n24411 = ( ~n1176 & n1568 ) | ( ~n1176 & n19587 ) | ( n1568 & n19587 ) ;
  assign n24413 = n24412 ^ n24411 ^ n21440 ;
  assign n24414 = ( n5522 & n7443 ) | ( n5522 & ~n12135 ) | ( n7443 & ~n12135 ) ;
  assign n24415 = n14128 ^ n4452 ^ n4149 ;
  assign n24416 = ( n2894 & n9060 ) | ( n2894 & ~n17709 ) | ( n9060 & ~n17709 ) ;
  assign n24417 = ( n24414 & ~n24415 ) | ( n24414 & n24416 ) | ( ~n24415 & n24416 ) ;
  assign n24418 = n24417 ^ n9555 ^ n4484 ;
  assign n24419 = ( n9318 & n10282 ) | ( n9318 & ~n16205 ) | ( n10282 & ~n16205 ) ;
  assign n24420 = ( n3587 & ~n15067 ) | ( n3587 & n19276 ) | ( ~n15067 & n19276 ) ;
  assign n24421 = n24420 ^ n21879 ^ n593 ;
  assign n24422 = ( ~n2863 & n6629 ) | ( ~n2863 & n24421 ) | ( n6629 & n24421 ) ;
  assign n24425 = n15638 ^ n2011 ^ n1347 ;
  assign n24424 = n9520 ^ n4704 ^ n3441 ;
  assign n24423 = n23589 ^ n15296 ^ n1712 ;
  assign n24426 = n24425 ^ n24424 ^ n24423 ;
  assign n24427 = ( n261 & ~n13137 ) | ( n261 & n24426 ) | ( ~n13137 & n24426 ) ;
  assign n24428 = n9712 ^ n6746 ^ n3767 ;
  assign n24429 = ( ~n7517 & n9700 ) | ( ~n7517 & n24428 ) | ( n9700 & n24428 ) ;
  assign n24430 = n15320 ^ n13283 ^ n9766 ;
  assign n24431 = n24430 ^ n20591 ^ n11787 ;
  assign n24432 = ( ~n3280 & n24429 ) | ( ~n3280 & n24431 ) | ( n24429 & n24431 ) ;
  assign n24433 = n12100 ^ n9924 ^ n8915 ;
  assign n24434 = ( n7221 & n9089 ) | ( n7221 & n24433 ) | ( n9089 & n24433 ) ;
  assign n24436 = ( n1533 & n3529 ) | ( n1533 & ~n5185 ) | ( n3529 & ~n5185 ) ;
  assign n24437 = n24436 ^ n24361 ^ n22817 ;
  assign n24435 = ( ~n3303 & n4346 ) | ( ~n3303 & n14404 ) | ( n4346 & n14404 ) ;
  assign n24438 = n24437 ^ n24435 ^ n5463 ;
  assign n24439 = n16539 ^ n6235 ^ n3273 ;
  assign n24440 = ( n254 & ~n9411 ) | ( n254 & n24439 ) | ( ~n9411 & n24439 ) ;
  assign n24441 = ( ~n8915 & n9624 ) | ( ~n8915 & n24440 ) | ( n9624 & n24440 ) ;
  assign n24442 = ( n6617 & ~n15367 ) | ( n6617 & n19207 ) | ( ~n15367 & n19207 ) ;
  assign n24443 = ( ~n2862 & n7989 ) | ( ~n2862 & n10124 ) | ( n7989 & n10124 ) ;
  assign n24444 = n12190 ^ n11103 ^ n10419 ;
  assign n24445 = ( n9892 & n19010 ) | ( n9892 & ~n24444 ) | ( n19010 & ~n24444 ) ;
  assign n24446 = ( n1273 & n8583 ) | ( n1273 & ~n24445 ) | ( n8583 & ~n24445 ) ;
  assign n24447 = n14036 ^ n11225 ^ n2687 ;
  assign n24448 = ( ~n632 & n24446 ) | ( ~n632 & n24447 ) | ( n24446 & n24447 ) ;
  assign n24449 = ( n10695 & n13430 ) | ( n10695 & ~n23148 ) | ( n13430 & ~n23148 ) ;
  assign n24450 = n24449 ^ n8994 ^ n6632 ;
  assign n24451 = n24450 ^ n17530 ^ n16270 ;
  assign n24452 = ( n4422 & n5142 ) | ( n4422 & n15683 ) | ( n5142 & n15683 ) ;
  assign n24453 = n9774 ^ n1985 ^ n1798 ;
  assign n24454 = ( n4293 & ~n7979 ) | ( n4293 & n24453 ) | ( ~n7979 & n24453 ) ;
  assign n24455 = n11547 ^ n8970 ^ n6338 ;
  assign n24456 = ( ~n20000 & n23835 ) | ( ~n20000 & n24455 ) | ( n23835 & n24455 ) ;
  assign n24457 = n8441 ^ n3297 ^ n226 ;
  assign n24458 = ( n1786 & ~n3536 ) | ( n1786 & n24457 ) | ( ~n3536 & n24457 ) ;
  assign n24459 = ( n1396 & ~n8296 ) | ( n1396 & n14544 ) | ( ~n8296 & n14544 ) ;
  assign n24460 = ( n8271 & ~n24458 ) | ( n8271 & n24459 ) | ( ~n24458 & n24459 ) ;
  assign n24461 = n16814 ^ n10462 ^ n9424 ;
  assign n24462 = ( n2261 & n2947 ) | ( n2261 & n3210 ) | ( n2947 & n3210 ) ;
  assign n24463 = ( n11395 & n24461 ) | ( n11395 & n24462 ) | ( n24461 & n24462 ) ;
  assign n24464 = ( n2988 & n4040 ) | ( n2988 & n24463 ) | ( n4040 & n24463 ) ;
  assign n24465 = n13165 ^ n11670 ^ n4682 ;
  assign n24466 = ( n15191 & n20960 ) | ( n15191 & ~n24465 ) | ( n20960 & ~n24465 ) ;
  assign n24467 = ( n6590 & n10114 ) | ( n6590 & ~n10345 ) | ( n10114 & ~n10345 ) ;
  assign n24468 = ( n5873 & ~n9243 ) | ( n5873 & n14002 ) | ( ~n9243 & n14002 ) ;
  assign n24469 = n24468 ^ n17390 ^ n1730 ;
  assign n24470 = ( n15795 & ~n16438 ) | ( n15795 & n24469 ) | ( ~n16438 & n24469 ) ;
  assign n24471 = n24470 ^ n11141 ^ n3385 ;
  assign n24473 = n21372 ^ n18080 ^ n12308 ;
  assign n24474 = n24473 ^ n5315 ^ n3602 ;
  assign n24472 = n22460 ^ n18590 ^ n3070 ;
  assign n24475 = n24474 ^ n24472 ^ n16860 ;
  assign n24476 = ( n7323 & ~n11377 ) | ( n7323 & n16778 ) | ( ~n11377 & n16778 ) ;
  assign n24477 = n3763 ^ n1972 ^ n726 ;
  assign n24478 = n24477 ^ n8379 ^ n6274 ;
  assign n24479 = ( ~n11618 & n19162 ) | ( ~n11618 & n24478 ) | ( n19162 & n24478 ) ;
  assign n24480 = ( ~n5586 & n19342 ) | ( ~n5586 & n24479 ) | ( n19342 & n24479 ) ;
  assign n24481 = ( n6547 & n10737 ) | ( n6547 & ~n16911 ) | ( n10737 & ~n16911 ) ;
  assign n24482 = n9687 ^ n2539 ^ n1940 ;
  assign n24483 = n24482 ^ n15965 ^ n6488 ;
  assign n24484 = n18289 ^ n14605 ^ n6629 ;
  assign n24485 = ( n8067 & ~n14817 ) | ( n8067 & n24484 ) | ( ~n14817 & n24484 ) ;
  assign n24486 = ( n7614 & ~n17960 ) | ( n7614 & n18821 ) | ( ~n17960 & n18821 ) ;
  assign n24487 = n18103 ^ n11802 ^ n8119 ;
  assign n24488 = n14168 ^ n8610 ^ n3444 ;
  assign n24489 = n24488 ^ n6686 ^ n1246 ;
  assign n24490 = n24489 ^ n12218 ^ n4313 ;
  assign n24491 = ( n4555 & ~n10685 ) | ( n4555 & n16561 ) | ( ~n10685 & n16561 ) ;
  assign n24492 = ( ~n3046 & n15125 ) | ( ~n3046 & n24491 ) | ( n15125 & n24491 ) ;
  assign n24493 = ( n20051 & n24490 ) | ( n20051 & ~n24492 ) | ( n24490 & ~n24492 ) ;
  assign n24494 = n23289 ^ n18677 ^ n3746 ;
  assign n24495 = n17818 ^ n12939 ^ n4742 ;
  assign n24496 = n24495 ^ n840 ^ n479 ;
  assign n24497 = ( n17927 & n23060 ) | ( n17927 & n24496 ) | ( n23060 & n24496 ) ;
  assign n24498 = n24497 ^ n11569 ^ n3761 ;
  assign n24499 = n15481 ^ n11299 ^ n1388 ;
  assign n24500 = n24499 ^ n12480 ^ n9434 ;
  assign n24501 = ( n12218 & ~n18867 ) | ( n12218 & n19204 ) | ( ~n18867 & n19204 ) ;
  assign n24502 = ( n3163 & ~n8882 ) | ( n3163 & n24501 ) | ( ~n8882 & n24501 ) ;
  assign n24503 = ( ~n700 & n4385 ) | ( ~n700 & n14070 ) | ( n4385 & n14070 ) ;
  assign n24504 = n24503 ^ n20540 ^ n1682 ;
  assign n24505 = n24504 ^ n9583 ^ n7148 ;
  assign n24506 = n24505 ^ n4733 ^ n3588 ;
  assign n24507 = n13982 ^ n9007 ^ n5163 ;
  assign n24508 = ( n17976 & ~n18838 ) | ( n17976 & n24507 ) | ( ~n18838 & n24507 ) ;
  assign n24509 = n21530 ^ n19450 ^ n2024 ;
  assign n24510 = ( ~n13636 & n24508 ) | ( ~n13636 & n24509 ) | ( n24508 & n24509 ) ;
  assign n24511 = ( ~n2038 & n3381 ) | ( ~n2038 & n23341 ) | ( n3381 & n23341 ) ;
  assign n24512 = n22692 ^ n6767 ^ n4996 ;
  assign n24513 = ( n11670 & n13533 ) | ( n11670 & ~n18298 ) | ( n13533 & ~n18298 ) ;
  assign n24514 = n24513 ^ n8384 ^ n5226 ;
  assign n24515 = n12790 ^ n7570 ^ n7432 ;
  assign n24516 = ( n941 & n8069 ) | ( n941 & n24515 ) | ( n8069 & n24515 ) ;
  assign n24517 = ( n4864 & n15198 ) | ( n4864 & n18679 ) | ( n15198 & n18679 ) ;
  assign n24518 = ( n1877 & n24516 ) | ( n1877 & n24517 ) | ( n24516 & n24517 ) ;
  assign n24519 = n24518 ^ n23062 ^ n6254 ;
  assign n24520 = ( n186 & n1372 ) | ( n186 & ~n8629 ) | ( n1372 & ~n8629 ) ;
  assign n24521 = n24520 ^ n9131 ^ n8950 ;
  assign n24522 = n22437 ^ n10043 ^ n1201 ;
  assign n24523 = ( n17190 & n24521 ) | ( n17190 & n24522 ) | ( n24521 & n24522 ) ;
  assign n24524 = n18020 ^ n10131 ^ n9714 ;
  assign n24525 = n11940 ^ n7037 ^ n4298 ;
  assign n24526 = ( n8342 & ~n11284 ) | ( n8342 & n24525 ) | ( ~n11284 & n24525 ) ;
  assign n24527 = ( ~n714 & n4545 ) | ( ~n714 & n11571 ) | ( n4545 & n11571 ) ;
  assign n24528 = ( x24 & n22961 ) | ( x24 & ~n24527 ) | ( n22961 & ~n24527 ) ;
  assign n24529 = ( n3122 & n14753 ) | ( n3122 & n24528 ) | ( n14753 & n24528 ) ;
  assign n24530 = n24529 ^ n12383 ^ n8994 ;
  assign n24531 = n24297 ^ n14781 ^ n4169 ;
  assign n24532 = ( n3570 & n14810 ) | ( n3570 & n22285 ) | ( n14810 & n22285 ) ;
  assign n24533 = n20560 ^ n18776 ^ n11771 ;
  assign n24534 = n17199 ^ n7692 ^ n7603 ;
  assign n24535 = ( n7172 & n18766 ) | ( n7172 & ~n24534 ) | ( n18766 & ~n24534 ) ;
  assign n24536 = n10941 ^ n4855 ^ n1268 ;
  assign n24537 = n24536 ^ n5086 ^ n2527 ;
  assign n24538 = ( n5352 & n5470 ) | ( n5352 & n18335 ) | ( n5470 & n18335 ) ;
  assign n24539 = n24538 ^ n24289 ^ n5257 ;
  assign n24540 = ( n252 & n9573 ) | ( n252 & ~n18178 ) | ( n9573 & ~n18178 ) ;
  assign n24541 = ( ~n2913 & n4460 ) | ( ~n2913 & n24540 ) | ( n4460 & n24540 ) ;
  assign n24542 = n24541 ^ n16435 ^ n195 ;
  assign n24543 = n15541 ^ n3374 ^ n1593 ;
  assign n24544 = n20384 ^ n19246 ^ n10886 ;
  assign n24545 = n21784 ^ n21234 ^ n7840 ;
  assign n24546 = n20791 ^ n19325 ^ n16851 ;
  assign n24547 = ( n4103 & n18416 ) | ( n4103 & ~n19502 ) | ( n18416 & ~n19502 ) ;
  assign n24548 = ( n11135 & ~n24546 ) | ( n11135 & n24547 ) | ( ~n24546 & n24547 ) ;
  assign n24549 = n18263 ^ n3431 ^ x87 ;
  assign n24552 = ( n1853 & ~n19299 ) | ( n1853 & n22308 ) | ( ~n19299 & n22308 ) ;
  assign n24550 = ( n4887 & ~n6739 ) | ( n4887 & n10470 ) | ( ~n6739 & n10470 ) ;
  assign n24551 = ( n2795 & n9292 ) | ( n2795 & ~n24550 ) | ( n9292 & ~n24550 ) ;
  assign n24553 = n24552 ^ n24551 ^ n16720 ;
  assign n24555 = n8810 ^ n1075 ^ n445 ;
  assign n24556 = n24555 ^ n14575 ^ n1904 ;
  assign n24554 = ( n1733 & n4428 ) | ( n1733 & ~n14414 ) | ( n4428 & ~n14414 ) ;
  assign n24557 = n24556 ^ n24554 ^ n839 ;
  assign n24558 = n24557 ^ n2276 ^ n947 ;
  assign n24559 = ( n2661 & n9074 ) | ( n2661 & n24558 ) | ( n9074 & n24558 ) ;
  assign n24560 = n13811 ^ n13680 ^ n6815 ;
  assign n24561 = n24560 ^ n3802 ^ n3403 ;
  assign n24562 = n24561 ^ n11820 ^ n5503 ;
  assign n24563 = ( n4066 & ~n4327 ) | ( n4066 & n16803 ) | ( ~n4327 & n16803 ) ;
  assign n24566 = n19222 ^ n9386 ^ n3839 ;
  assign n24564 = ( ~n816 & n4225 ) | ( ~n816 & n5869 ) | ( n4225 & n5869 ) ;
  assign n24565 = ( n8962 & ~n12355 ) | ( n8962 & n24564 ) | ( ~n12355 & n24564 ) ;
  assign n24567 = n24566 ^ n24565 ^ n13925 ;
  assign n24568 = ( n12894 & ~n24563 ) | ( n12894 & n24567 ) | ( ~n24563 & n24567 ) ;
  assign n24570 = ( n4366 & n10714 ) | ( n4366 & n21461 ) | ( n10714 & n21461 ) ;
  assign n24569 = n9193 ^ n3242 ^ n783 ;
  assign n24571 = n24570 ^ n24569 ^ n19560 ;
  assign n24572 = n22434 ^ n17158 ^ n15017 ;
  assign n24573 = n24572 ^ n5567 ^ n2919 ;
  assign n24574 = n7453 ^ n3682 ^ n2325 ;
  assign n24575 = ( n4324 & n5750 ) | ( n4324 & n19047 ) | ( n5750 & n19047 ) ;
  assign n24578 = ( n2462 & n7357 ) | ( n2462 & ~n21316 ) | ( n7357 & ~n21316 ) ;
  assign n24576 = n15736 ^ n3215 ^ n2710 ;
  assign n24577 = n24576 ^ n19780 ^ n9911 ;
  assign n24579 = n24578 ^ n24577 ^ n617 ;
  assign n24580 = ( n1174 & ~n5880 ) | ( n1174 & n22738 ) | ( ~n5880 & n22738 ) ;
  assign n24581 = ( n9569 & n9880 ) | ( n9569 & ~n16485 ) | ( n9880 & ~n16485 ) ;
  assign n24582 = n24581 ^ n23868 ^ n17474 ;
  assign n24583 = ( n2695 & n16440 ) | ( n2695 & ~n17883 ) | ( n16440 & ~n17883 ) ;
  assign n24584 = n24583 ^ n3133 ^ n2827 ;
  assign n24585 = ( n3306 & n3893 ) | ( n3306 & ~n11963 ) | ( n3893 & ~n11963 ) ;
  assign n24586 = ( n5657 & n16453 ) | ( n5657 & n24585 ) | ( n16453 & n24585 ) ;
  assign n24587 = ( n587 & n24584 ) | ( n587 & ~n24586 ) | ( n24584 & ~n24586 ) ;
  assign n24588 = n16383 ^ n14485 ^ n4548 ;
  assign n24589 = ( n1669 & n5549 ) | ( n1669 & n20444 ) | ( n5549 & n20444 ) ;
  assign n24590 = ( n18591 & ~n23892 ) | ( n18591 & n24589 ) | ( ~n23892 & n24589 ) ;
  assign n24591 = n11728 ^ n9491 ^ n9203 ;
  assign n24592 = n24591 ^ n21686 ^ n7427 ;
  assign n24593 = n23275 ^ n23087 ^ n6861 ;
  assign n24594 = ( n870 & n2121 ) | ( n870 & ~n24593 ) | ( n2121 & ~n24593 ) ;
  assign n24595 = n9139 ^ n3965 ^ n1253 ;
  assign n24596 = ( n6819 & ~n20158 ) | ( n6819 & n21273 ) | ( ~n20158 & n21273 ) ;
  assign n24597 = n24252 ^ n6056 ^ n1967 ;
  assign n24598 = n24597 ^ n18994 ^ n18821 ;
  assign n24599 = n24598 ^ n24497 ^ n3036 ;
  assign n24600 = ( ~n5547 & n13481 ) | ( ~n5547 & n21296 ) | ( n13481 & n21296 ) ;
  assign n24601 = n17886 ^ n5059 ^ n2611 ;
  assign n24602 = ( ~n7577 & n23038 ) | ( ~n7577 & n24601 ) | ( n23038 & n24601 ) ;
  assign n24603 = n24602 ^ n19893 ^ n11343 ;
  assign n24604 = n16394 ^ n8353 ^ n5652 ;
  assign n24605 = n24604 ^ n21866 ^ n5467 ;
  assign n24606 = ( n4561 & n18166 ) | ( n4561 & ~n24605 ) | ( n18166 & ~n24605 ) ;
  assign n24607 = n6464 ^ n6443 ^ n3592 ;
  assign n24609 = n12077 ^ n11393 ^ n8842 ;
  assign n24608 = ( n7969 & n12345 ) | ( n7969 & n16204 ) | ( n12345 & n16204 ) ;
  assign n24610 = n24609 ^ n24608 ^ n12476 ;
  assign n24611 = ( ~n10866 & n24440 ) | ( ~n10866 & n24610 ) | ( n24440 & n24610 ) ;
  assign n24612 = ( ~n2220 & n24607 ) | ( ~n2220 & n24611 ) | ( n24607 & n24611 ) ;
  assign n24613 = ( n203 & ~n712 ) | ( n203 & n8152 ) | ( ~n712 & n8152 ) ;
  assign n24614 = n20479 ^ n13683 ^ n6117 ;
  assign n24615 = ( n5044 & n24613 ) | ( n5044 & ~n24614 ) | ( n24613 & ~n24614 ) ;
  assign n24616 = n10050 ^ n4938 ^ n4591 ;
  assign n24617 = n24616 ^ n10531 ^ n5633 ;
  assign n24618 = n24617 ^ n22422 ^ n5419 ;
  assign n24619 = n22636 ^ n10619 ^ n6986 ;
  assign n24620 = n24619 ^ n5045 ^ n1565 ;
  assign n24621 = ( ~n726 & n8266 ) | ( ~n726 & n16472 ) | ( n8266 & n16472 ) ;
  assign n24622 = n16968 ^ n6397 ^ n1002 ;
  assign n24623 = n24622 ^ n11084 ^ n8801 ;
  assign n24624 = n5715 ^ n5677 ^ n5549 ;
  assign n24625 = ( n559 & n11486 ) | ( n559 & ~n24624 ) | ( n11486 & ~n24624 ) ;
  assign n24626 = n8543 ^ n2721 ^ n1800 ;
  assign n24627 = n24626 ^ n14886 ^ n13627 ;
  assign n24630 = ( n3028 & n3397 ) | ( n3028 & n16757 ) | ( n3397 & n16757 ) ;
  assign n24629 = ( ~n561 & n14423 ) | ( ~n561 & n14673 ) | ( n14423 & n14673 ) ;
  assign n24628 = ( n3449 & n6898 ) | ( n3449 & n19112 ) | ( n6898 & n19112 ) ;
  assign n24631 = n24630 ^ n24629 ^ n24628 ;
  assign n24632 = ( n15097 & ~n24627 ) | ( n15097 & n24631 ) | ( ~n24627 & n24631 ) ;
  assign n24633 = ( n4940 & n5527 ) | ( n4940 & n18572 ) | ( n5527 & n18572 ) ;
  assign n24634 = n13135 ^ n7037 ^ n1803 ;
  assign n24635 = ( ~n3136 & n3905 ) | ( ~n3136 & n5172 ) | ( n3905 & n5172 ) ;
  assign n24636 = n11053 ^ n8773 ^ n3589 ;
  assign n24637 = ( ~n19126 & n24635 ) | ( ~n19126 & n24636 ) | ( n24635 & n24636 ) ;
  assign n24638 = n8768 ^ n4723 ^ n176 ;
  assign n24639 = ( n8075 & ~n11406 ) | ( n8075 & n12219 ) | ( ~n11406 & n12219 ) ;
  assign n24640 = ( ~n14710 & n17430 ) | ( ~n14710 & n24639 ) | ( n17430 & n24639 ) ;
  assign n24641 = ( ~n9785 & n24109 ) | ( ~n9785 & n24640 ) | ( n24109 & n24640 ) ;
  assign n24642 = n23625 ^ n23022 ^ n17937 ;
  assign n24643 = n17463 ^ n4110 ^ n3831 ;
  assign n24644 = ( n1562 & ~n1629 ) | ( n1562 & n14354 ) | ( ~n1629 & n14354 ) ;
  assign n24645 = ( n7882 & n24643 ) | ( n7882 & n24644 ) | ( n24643 & n24644 ) ;
  assign n24646 = ( ~n12485 & n21799 ) | ( ~n12485 & n24645 ) | ( n21799 & n24645 ) ;
  assign n24647 = ( ~n1416 & n5736 ) | ( ~n1416 & n8225 ) | ( n5736 & n8225 ) ;
  assign n24648 = n24647 ^ n24577 ^ n14630 ;
  assign n24649 = ( ~n3332 & n8367 ) | ( ~n3332 & n8438 ) | ( n8367 & n8438 ) ;
  assign n24650 = ( n4456 & ~n5965 ) | ( n4456 & n13910 ) | ( ~n5965 & n13910 ) ;
  assign n24651 = ( ~n5856 & n9032 ) | ( ~n5856 & n24650 ) | ( n9032 & n24650 ) ;
  assign n24652 = n24651 ^ n12216 ^ n3184 ;
  assign n24653 = ( ~n2180 & n8369 ) | ( ~n2180 & n8546 ) | ( n8369 & n8546 ) ;
  assign n24654 = n24653 ^ n16266 ^ n13885 ;
  assign n24655 = ( ~n6104 & n10363 ) | ( ~n6104 & n10800 ) | ( n10363 & n10800 ) ;
  assign n24656 = n24655 ^ n8032 ^ n2862 ;
  assign n24657 = n24656 ^ n4441 ^ n3321 ;
  assign n24658 = n14532 ^ n8859 ^ n7422 ;
  assign n24659 = n15437 ^ n11961 ^ n7490 ;
  assign n24660 = n24659 ^ n5953 ^ n1144 ;
  assign n24661 = ( n22081 & n24658 ) | ( n22081 & n24660 ) | ( n24658 & n24660 ) ;
  assign n24664 = n23558 ^ n14782 ^ n12062 ;
  assign n24662 = n5724 ^ n5248 ^ n4526 ;
  assign n24663 = n24662 ^ n13587 ^ n12576 ;
  assign n24665 = n24664 ^ n24663 ^ n9215 ;
  assign n24668 = ( n2110 & n2903 ) | ( n2110 & ~n9035 ) | ( n2903 & ~n9035 ) ;
  assign n24666 = n11036 ^ n9162 ^ n6296 ;
  assign n24667 = ( ~n9199 & n22934 ) | ( ~n9199 & n24666 ) | ( n22934 & n24666 ) ;
  assign n24669 = n24668 ^ n24667 ^ n24207 ;
  assign n24670 = n23469 ^ n20177 ^ n14801 ;
  assign n24671 = ( ~n2378 & n14370 ) | ( ~n2378 & n17430 ) | ( n14370 & n17430 ) ;
  assign n24672 = ( n165 & ~n23275 ) | ( n165 & n24671 ) | ( ~n23275 & n24671 ) ;
  assign n24673 = n22553 ^ n22360 ^ n16749 ;
  assign n24674 = ( n1316 & n2610 ) | ( n1316 & n21268 ) | ( n2610 & n21268 ) ;
  assign n24675 = ( n2110 & n4870 ) | ( n2110 & ~n12658 ) | ( n4870 & ~n12658 ) ;
  assign n24676 = ( n3592 & ~n18651 ) | ( n3592 & n24675 ) | ( ~n18651 & n24675 ) ;
  assign n24677 = n22802 ^ n22509 ^ n6240 ;
  assign n24678 = n4743 ^ n4019 ^ n1907 ;
  assign n24679 = ( ~n7801 & n11667 ) | ( ~n7801 & n19047 ) | ( n11667 & n19047 ) ;
  assign n24680 = n24679 ^ n22615 ^ n12008 ;
  assign n24682 = n7813 ^ n310 ^ x96 ;
  assign n24681 = ( n1888 & n15281 ) | ( n1888 & n20587 ) | ( n15281 & n20587 ) ;
  assign n24683 = n24682 ^ n24681 ^ n15476 ;
  assign n24684 = ( n171 & n1926 ) | ( n171 & ~n19358 ) | ( n1926 & ~n19358 ) ;
  assign n24685 = n24684 ^ n5093 ^ n3944 ;
  assign n24686 = n24685 ^ n21393 ^ n4065 ;
  assign n24687 = n13969 ^ n8988 ^ n6542 ;
  assign n24688 = n16897 ^ n16181 ^ n2252 ;
  assign n24689 = n24688 ^ n8154 ^ n1395 ;
  assign n24691 = ( ~n8768 & n10846 ) | ( ~n8768 & n15027 ) | ( n10846 & n15027 ) ;
  assign n24690 = ( n5023 & n6433 ) | ( n5023 & ~n18230 ) | ( n6433 & ~n18230 ) ;
  assign n24692 = n24691 ^ n24690 ^ n344 ;
  assign n24693 = n2732 ^ n1933 ^ n1730 ;
  assign n24694 = n24693 ^ n8959 ^ n1449 ;
  assign n24695 = ( ~n2629 & n13626 ) | ( ~n2629 & n16341 ) | ( n13626 & n16341 ) ;
  assign n24696 = ( ~n2541 & n10012 ) | ( ~n2541 & n11271 ) | ( n10012 & n11271 ) ;
  assign n24697 = ( ~n11626 & n17100 ) | ( ~n11626 & n20047 ) | ( n17100 & n20047 ) ;
  assign n24698 = ( n21537 & n24696 ) | ( n21537 & n24697 ) | ( n24696 & n24697 ) ;
  assign n24699 = ( n11677 & n12293 ) | ( n11677 & n24628 ) | ( n12293 & n24628 ) ;
  assign n24700 = n15489 ^ n11844 ^ n3828 ;
  assign n24701 = n11071 ^ n1847 ^ n1428 ;
  assign n24702 = ( n3132 & n6315 ) | ( n3132 & ~n24701 ) | ( n6315 & ~n24701 ) ;
  assign n24703 = ( n12583 & ~n23280 ) | ( n12583 & n24702 ) | ( ~n23280 & n24702 ) ;
  assign n24708 = n11011 ^ n6064 ^ n2578 ;
  assign n24706 = ( n2365 & n10338 ) | ( n2365 & n17982 ) | ( n10338 & n17982 ) ;
  assign n24707 = n24706 ^ n7241 ^ n6875 ;
  assign n24704 = n21743 ^ n16606 ^ n1557 ;
  assign n24705 = ( ~n4699 & n4937 ) | ( ~n4699 & n24704 ) | ( n4937 & n24704 ) ;
  assign n24709 = n24708 ^ n24707 ^ n24705 ;
  assign n24710 = n15486 ^ n8601 ^ n6297 ;
  assign n24711 = ( ~n14396 & n20977 ) | ( ~n14396 & n24710 ) | ( n20977 & n24710 ) ;
  assign n24712 = ( ~n6689 & n16534 ) | ( ~n6689 & n24711 ) | ( n16534 & n24711 ) ;
  assign n24713 = n22532 ^ n9021 ^ n313 ;
  assign n24716 = n17381 ^ n11370 ^ n3570 ;
  assign n24717 = n24716 ^ n12652 ^ n8418 ;
  assign n24718 = ( n6428 & n17479 ) | ( n6428 & n24717 ) | ( n17479 & n24717 ) ;
  assign n24714 = n14189 ^ n6411 ^ n3862 ;
  assign n24715 = n24714 ^ n1776 ^ n452 ;
  assign n24719 = n24718 ^ n24715 ^ n19818 ;
  assign n24720 = n20935 ^ n6263 ^ n4513 ;
  assign n24721 = ( n8062 & n12488 ) | ( n8062 & n16174 ) | ( n12488 & n16174 ) ;
  assign n24722 = ( n11684 & n24720 ) | ( n11684 & ~n24721 ) | ( n24720 & ~n24721 ) ;
  assign n24725 = ( ~n9043 & n10002 ) | ( ~n9043 & n11220 ) | ( n10002 & n11220 ) ;
  assign n24726 = n24725 ^ n10601 ^ n2200 ;
  assign n24723 = n7327 ^ n7043 ^ n4520 ;
  assign n24724 = ( n10004 & ~n18879 ) | ( n10004 & n24723 ) | ( ~n18879 & n24723 ) ;
  assign n24727 = n24726 ^ n24724 ^ n24219 ;
  assign n24728 = ( ~n1937 & n6915 ) | ( ~n1937 & n13904 ) | ( n6915 & n13904 ) ;
  assign n24733 = n11895 ^ n4968 ^ n1409 ;
  assign n24734 = n24733 ^ n10059 ^ n8366 ;
  assign n24729 = ( n4263 & n8331 ) | ( n4263 & n8966 ) | ( n8331 & n8966 ) ;
  assign n24730 = ( ~n5224 & n9441 ) | ( ~n5224 & n20627 ) | ( n9441 & n20627 ) ;
  assign n24731 = ( n16101 & ~n19796 ) | ( n16101 & n24730 ) | ( ~n19796 & n24730 ) ;
  assign n24732 = ( ~n2239 & n24729 ) | ( ~n2239 & n24731 ) | ( n24729 & n24731 ) ;
  assign n24735 = n24734 ^ n24732 ^ n4768 ;
  assign n24736 = ( ~n806 & n2233 ) | ( ~n806 & n3735 ) | ( n2233 & n3735 ) ;
  assign n24737 = ( n8460 & ~n22131 ) | ( n8460 & n23816 ) | ( ~n22131 & n23816 ) ;
  assign n24738 = ( n8070 & n24736 ) | ( n8070 & ~n24737 ) | ( n24736 & ~n24737 ) ;
  assign n24739 = ( ~n2293 & n17426 ) | ( ~n2293 & n24738 ) | ( n17426 & n24738 ) ;
  assign n24740 = n8735 ^ n6105 ^ n4899 ;
  assign n24741 = n24740 ^ n20030 ^ n7949 ;
  assign n24742 = n24162 ^ n15744 ^ n3022 ;
  assign n24743 = ( ~n2881 & n7615 ) | ( ~n2881 & n8842 ) | ( n7615 & n8842 ) ;
  assign n24744 = ( n6546 & n15873 ) | ( n6546 & n24743 ) | ( n15873 & n24743 ) ;
  assign n24745 = n24744 ^ n22325 ^ n14912 ;
  assign n24746 = ( n12366 & n14104 ) | ( n12366 & n14724 ) | ( n14104 & n14724 ) ;
  assign n24747 = ( n6108 & ~n17037 ) | ( n6108 & n24746 ) | ( ~n17037 & n24746 ) ;
  assign n24748 = ( n7206 & n10851 ) | ( n7206 & ~n23399 ) | ( n10851 & ~n23399 ) ;
  assign n24749 = n24748 ^ n7245 ^ n509 ;
  assign n24750 = ( ~n906 & n12491 ) | ( ~n906 & n21166 ) | ( n12491 & n21166 ) ;
  assign n24751 = ( ~n416 & n3550 ) | ( ~n416 & n24622 ) | ( n3550 & n24622 ) ;
  assign n24752 = n21299 ^ n14323 ^ n9099 ;
  assign n24753 = n20051 ^ n6240 ^ n734 ;
  assign n24754 = n12870 ^ n4973 ^ n1089 ;
  assign n24755 = ( n9679 & ~n24753 ) | ( n9679 & n24754 ) | ( ~n24753 & n24754 ) ;
  assign n24757 = ( n9402 & n20409 ) | ( n9402 & ~n22269 ) | ( n20409 & ~n22269 ) ;
  assign n24756 = n23693 ^ n20311 ^ n10714 ;
  assign n24758 = n24757 ^ n24756 ^ n11602 ;
  assign n24759 = ( n11574 & n15375 ) | ( n11574 & n19236 ) | ( n15375 & n19236 ) ;
  assign n24760 = n21213 ^ n3524 ^ n428 ;
  assign n24761 = ( n11700 & ~n18111 ) | ( n11700 & n21205 ) | ( ~n18111 & n21205 ) ;
  assign n24762 = ( ~n8301 & n11240 ) | ( ~n8301 & n24761 ) | ( n11240 & n24761 ) ;
  assign n24766 = ( ~n6077 & n6172 ) | ( ~n6077 & n23243 ) | ( n6172 & n23243 ) ;
  assign n24763 = n15082 ^ n2690 ^ n1420 ;
  assign n24764 = ( n13871 & n19705 ) | ( n13871 & n24763 ) | ( n19705 & n24763 ) ;
  assign n24765 = ( n4270 & ~n6576 ) | ( n4270 & n24764 ) | ( ~n6576 & n24764 ) ;
  assign n24767 = n24766 ^ n24765 ^ n4126 ;
  assign n24770 = ( n6284 & n18345 ) | ( n6284 & ~n22066 ) | ( n18345 & ~n22066 ) ;
  assign n24768 = ( ~n3003 & n21403 ) | ( ~n3003 & n24597 ) | ( n21403 & n24597 ) ;
  assign n24769 = ( n13714 & n15908 ) | ( n13714 & n24768 ) | ( n15908 & n24768 ) ;
  assign n24771 = n24770 ^ n24769 ^ n4269 ;
  assign n24772 = ( n354 & ~n3756 ) | ( n354 & n16025 ) | ( ~n3756 & n16025 ) ;
  assign n24773 = n9105 ^ n1505 ^ n742 ;
  assign n24774 = n24773 ^ n18289 ^ n8322 ;
  assign n24776 = n10671 ^ n8253 ^ n1229 ;
  assign n24775 = ( n7954 & n11488 ) | ( n7954 & n23830 ) | ( n11488 & n23830 ) ;
  assign n24777 = n24776 ^ n24775 ^ n10691 ;
  assign n24778 = n14969 ^ n5943 ^ n3999 ;
  assign n24779 = n7643 ^ n4184 ^ n3922 ;
  assign n24780 = ( n3890 & n9248 ) | ( n3890 & ~n24779 ) | ( n9248 & ~n24779 ) ;
  assign n24781 = ( n12640 & ~n24778 ) | ( n12640 & n24780 ) | ( ~n24778 & n24780 ) ;
  assign n24782 = n24781 ^ n17260 ^ n12878 ;
  assign n24783 = n2437 ^ n1413 ^ n1150 ;
  assign n24784 = n24783 ^ n13072 ^ n5282 ;
  assign n24785 = n24784 ^ n23024 ^ n22079 ;
  assign n24786 = n17645 ^ n15727 ^ n8559 ;
  assign n24787 = ( n7681 & ~n9938 ) | ( n7681 & n24786 ) | ( ~n9938 & n24786 ) ;
  assign n24790 = n12162 ^ n7761 ^ n4465 ;
  assign n24789 = ( n837 & n11783 ) | ( n837 & n18936 ) | ( n11783 & n18936 ) ;
  assign n24788 = ( n3595 & n6022 ) | ( n3595 & n19478 ) | ( n6022 & n19478 ) ;
  assign n24791 = n24790 ^ n24789 ^ n24788 ;
  assign n24792 = n6780 ^ n4709 ^ n1126 ;
  assign n24793 = ( ~n595 & n2681 ) | ( ~n595 & n24792 ) | ( n2681 & n24792 ) ;
  assign n24794 = n24793 ^ n17089 ^ n7350 ;
  assign n24795 = ( n10376 & n10804 ) | ( n10376 & n23622 ) | ( n10804 & n23622 ) ;
  assign n24796 = n24795 ^ n8361 ^ n6886 ;
  assign n24797 = ( ~n1836 & n9005 ) | ( ~n1836 & n10908 ) | ( n9005 & n10908 ) ;
  assign n24798 = n24797 ^ n13183 ^ n11395 ;
  assign n24799 = n24798 ^ n19107 ^ n762 ;
  assign n24800 = n2494 ^ n1998 ^ n238 ;
  assign n24801 = n24800 ^ n10745 ^ n4587 ;
  assign n24802 = ( n2001 & ~n3705 ) | ( n2001 & n24801 ) | ( ~n3705 & n24801 ) ;
  assign n24803 = n15168 ^ n5734 ^ n389 ;
  assign n24804 = ( n3450 & n12522 ) | ( n3450 & n20579 ) | ( n12522 & n20579 ) ;
  assign n24805 = ( x82 & n24803 ) | ( x82 & n24804 ) | ( n24803 & n24804 ) ;
  assign n24806 = ( n8161 & ~n8931 ) | ( n8161 & n24805 ) | ( ~n8931 & n24805 ) ;
  assign n24811 = n12358 ^ n11581 ^ n4813 ;
  assign n24812 = ( n7680 & n19610 ) | ( n7680 & ~n24811 ) | ( n19610 & ~n24811 ) ;
  assign n24813 = n24812 ^ n19164 ^ n4637 ;
  assign n24809 = n23887 ^ n4228 ^ n1631 ;
  assign n24807 = n8390 ^ n1588 ^ x118 ;
  assign n24808 = ( n7461 & n22140 ) | ( n7461 & n24807 ) | ( n22140 & n24807 ) ;
  assign n24810 = n24809 ^ n24808 ^ n8811 ;
  assign n24814 = n24813 ^ n24810 ^ n16603 ;
  assign n24815 = ( n24802 & n24806 ) | ( n24802 & n24814 ) | ( n24806 & n24814 ) ;
  assign n24816 = ( ~x3 & n866 ) | ( ~x3 & n2121 ) | ( n866 & n2121 ) ;
  assign n24817 = n24816 ^ n21449 ^ n379 ;
  assign n24818 = ( n16558 & n24536 ) | ( n16558 & ~n24817 ) | ( n24536 & ~n24817 ) ;
  assign n24819 = n17360 ^ n7428 ^ n142 ;
  assign n24820 = n11692 ^ n8387 ^ n4044 ;
  assign n24821 = ( ~n6365 & n24819 ) | ( ~n6365 & n24820 ) | ( n24819 & n24820 ) ;
  assign n24822 = n18036 ^ n15534 ^ n14673 ;
  assign n24823 = n18403 ^ n11429 ^ n11072 ;
  assign n24824 = n24823 ^ n24173 ^ n9942 ;
  assign n24825 = n24824 ^ n13891 ^ n4202 ;
  assign n24826 = ( n773 & ~n8480 ) | ( n773 & n14146 ) | ( ~n8480 & n14146 ) ;
  assign n24827 = ( n1384 & n3638 ) | ( n1384 & ~n24826 ) | ( n3638 & ~n24826 ) ;
  assign n24831 = n15933 ^ n6920 ^ n1692 ;
  assign n24832 = ( ~n4237 & n5280 ) | ( ~n4237 & n24831 ) | ( n5280 & n24831 ) ;
  assign n24829 = ( n12239 & ~n17434 ) | ( n12239 & n21701 ) | ( ~n17434 & n21701 ) ;
  assign n24828 = n4859 ^ n1240 ^ n1006 ;
  assign n24830 = n24829 ^ n24828 ^ n11010 ;
  assign n24833 = n24832 ^ n24830 ^ n3562 ;
  assign n24834 = ( ~n16829 & n22557 ) | ( ~n16829 & n24833 ) | ( n22557 & n24833 ) ;
  assign n24835 = n10744 ^ n5174 ^ n3782 ;
  assign n24836 = ( ~n3876 & n19379 ) | ( ~n3876 & n24835 ) | ( n19379 & n24835 ) ;
  assign n24837 = ( n3844 & n15551 ) | ( n3844 & n24836 ) | ( n15551 & n24836 ) ;
  assign n24838 = ( n320 & n6159 ) | ( n320 & ~n7641 ) | ( n6159 & ~n7641 ) ;
  assign n24839 = n24838 ^ n3529 ^ n334 ;
  assign n24840 = n24839 ^ n20271 ^ n8569 ;
  assign n24841 = ( n9182 & ~n13173 ) | ( n9182 & n15337 ) | ( ~n13173 & n15337 ) ;
  assign n24842 = n24841 ^ n11515 ^ n7206 ;
  assign n24843 = ( ~n7183 & n12390 ) | ( ~n7183 & n14591 ) | ( n12390 & n14591 ) ;
  assign n24844 = ( n683 & ~n12596 ) | ( n683 & n24843 ) | ( ~n12596 & n24843 ) ;
  assign n24845 = n16462 ^ n6844 ^ n3975 ;
  assign n24846 = ( n6713 & ~n9230 ) | ( n6713 & n21313 ) | ( ~n9230 & n21313 ) ;
  assign n24847 = n24846 ^ n11942 ^ n5612 ;
  assign n24848 = ( n4177 & ~n11455 ) | ( n4177 & n19669 ) | ( ~n11455 & n19669 ) ;
  assign n24849 = ( n2274 & n5175 ) | ( n2274 & ~n16583 ) | ( n5175 & ~n16583 ) ;
  assign n24850 = n15872 ^ n13057 ^ n2853 ;
  assign n24853 = ( n882 & n2234 ) | ( n882 & n11882 ) | ( n2234 & n11882 ) ;
  assign n24852 = n15385 ^ n14604 ^ n12860 ;
  assign n24851 = ( n5608 & n9087 ) | ( n5608 & n11945 ) | ( n9087 & n11945 ) ;
  assign n24854 = n24853 ^ n24852 ^ n24851 ;
  assign n24855 = n24854 ^ n14350 ^ n1588 ;
  assign n24856 = n14845 ^ n5166 ^ n2508 ;
  assign n24857 = n24856 ^ n23299 ^ n11182 ;
  assign n24858 = ( ~n7650 & n11429 ) | ( ~n7650 & n22324 ) | ( n11429 & n22324 ) ;
  assign n24859 = n22711 ^ n16667 ^ n5671 ;
  assign n24860 = ( ~n3162 & n24858 ) | ( ~n3162 & n24859 ) | ( n24858 & n24859 ) ;
  assign n24861 = ( n348 & n1334 ) | ( n348 & ~n3347 ) | ( n1334 & ~n3347 ) ;
  assign n24862 = ( n2594 & ~n7294 ) | ( n2594 & n17332 ) | ( ~n7294 & n17332 ) ;
  assign n24863 = ( n5542 & ~n10384 ) | ( n5542 & n23572 ) | ( ~n10384 & n23572 ) ;
  assign n24864 = ( n5989 & ~n21158 ) | ( n5989 & n24863 ) | ( ~n21158 & n24863 ) ;
  assign n24865 = ( n404 & ~n10679 ) | ( n404 & n22858 ) | ( ~n10679 & n22858 ) ;
  assign n24866 = n23481 ^ n4059 ^ n3733 ;
  assign n24867 = ( n8181 & n15899 ) | ( n8181 & ~n16864 ) | ( n15899 & ~n16864 ) ;
  assign n24868 = ( n18957 & ~n20032 ) | ( n18957 & n23204 ) | ( ~n20032 & n23204 ) ;
  assign n24869 = n9096 ^ n2725 ^ n2397 ;
  assign n24870 = ( ~n14517 & n24868 ) | ( ~n14517 & n24869 ) | ( n24868 & n24869 ) ;
  assign n24871 = ( n15415 & n24867 ) | ( n15415 & ~n24870 ) | ( n24867 & ~n24870 ) ;
  assign n24872 = n24640 ^ n14541 ^ n4486 ;
  assign n24873 = n12986 ^ n12061 ^ n4471 ;
  assign n24874 = n5574 ^ n3819 ^ x49 ;
  assign n24875 = n24874 ^ n23602 ^ n2741 ;
  assign n24876 = ( ~n6411 & n11542 ) | ( ~n6411 & n24875 ) | ( n11542 & n24875 ) ;
  assign n24877 = ( ~n4407 & n8393 ) | ( ~n4407 & n14674 ) | ( n8393 & n14674 ) ;
  assign n24878 = ( n14573 & n23053 ) | ( n14573 & n24877 ) | ( n23053 & n24877 ) ;
  assign n24879 = n21402 ^ n7340 ^ n6897 ;
  assign n24880 = n24879 ^ n19507 ^ n13414 ;
  assign n24881 = n21612 ^ n20707 ^ n7797 ;
  assign n24882 = n11935 ^ n8462 ^ n1298 ;
  assign n24883 = n24882 ^ n21519 ^ n11637 ;
  assign n24884 = n11013 ^ n1463 ^ n1344 ;
  assign n24885 = ( n836 & n8839 ) | ( n836 & ~n24884 ) | ( n8839 & ~n24884 ) ;
  assign n24886 = ( n11881 & n24883 ) | ( n11881 & n24885 ) | ( n24883 & n24885 ) ;
  assign n24887 = n19886 ^ n6520 ^ n5416 ;
  assign n24888 = n24887 ^ n20406 ^ n8327 ;
  assign n24889 = ( n3295 & n3455 ) | ( n3295 & n24888 ) | ( n3455 & n24888 ) ;
  assign n24890 = n11000 ^ n9478 ^ n9226 ;
  assign n24891 = ( n3271 & n5646 ) | ( n3271 & ~n11665 ) | ( n5646 & ~n11665 ) ;
  assign n24892 = ( n5624 & n13289 ) | ( n5624 & ~n24891 ) | ( n13289 & ~n24891 ) ;
  assign n24893 = ( ~n7934 & n10144 ) | ( ~n7934 & n16616 ) | ( n10144 & n16616 ) ;
  assign n24894 = n15737 ^ n13993 ^ n492 ;
  assign n24895 = n17392 ^ n5540 ^ n282 ;
  assign n24896 = n11932 ^ n10408 ^ n2125 ;
  assign n24897 = ( ~n18191 & n21875 ) | ( ~n18191 & n24896 ) | ( n21875 & n24896 ) ;
  assign n24898 = n24897 ^ n8770 ^ n1557 ;
  assign n24899 = ( n809 & n7566 ) | ( n809 & ~n22776 ) | ( n7566 & ~n22776 ) ;
  assign n24900 = n20020 ^ n19898 ^ n16349 ;
  assign n24901 = ( n1215 & ~n7716 ) | ( n1215 & n9365 ) | ( ~n7716 & n9365 ) ;
  assign n24902 = ( n24899 & ~n24900 ) | ( n24899 & n24901 ) | ( ~n24900 & n24901 ) ;
  assign n24903 = n7005 ^ n2569 ^ n700 ;
  assign n24904 = n24903 ^ n10926 ^ n1307 ;
  assign n24905 = n9591 ^ n5822 ^ n453 ;
  assign n24906 = ( n4382 & n17797 ) | ( n4382 & n24905 ) | ( n17797 & n24905 ) ;
  assign n24907 = ( n8886 & n19049 ) | ( n8886 & ~n19507 ) | ( n19049 & ~n19507 ) ;
  assign n24908 = n12458 ^ n11896 ^ n10040 ;
  assign n24909 = n23525 ^ n20199 ^ n10074 ;
  assign n24910 = ( n502 & ~n1214 ) | ( n502 & n13553 ) | ( ~n1214 & n13553 ) ;
  assign n24911 = ( n2935 & ~n9280 ) | ( n2935 & n24910 ) | ( ~n9280 & n24910 ) ;
  assign n24913 = n3689 ^ n3639 ^ n630 ;
  assign n24914 = ( n3653 & n7794 ) | ( n3653 & n24913 ) | ( n7794 & n24913 ) ;
  assign n24912 = n22559 ^ n14009 ^ n11081 ;
  assign n24915 = n24914 ^ n24912 ^ n16865 ;
  assign n24916 = ( n7881 & n10884 ) | ( n7881 & ~n22005 ) | ( n10884 & ~n22005 ) ;
  assign n24917 = n18019 ^ n12351 ^ n5309 ;
  assign n24918 = n20837 ^ n9228 ^ n8902 ;
  assign n24919 = ( n2814 & ~n3008 ) | ( n2814 & n14829 ) | ( ~n3008 & n14829 ) ;
  assign n24920 = n24919 ^ n10790 ^ n9830 ;
  assign n24921 = n10827 ^ n4853 ^ n2773 ;
  assign n24922 = n24921 ^ n10307 ^ n144 ;
  assign n24923 = ( n4739 & n8779 ) | ( n4739 & n24922 ) | ( n8779 & n24922 ) ;
  assign n24924 = n19781 ^ n4748 ^ n2034 ;
  assign n24925 = ( ~n1364 & n7643 ) | ( ~n1364 & n24924 ) | ( n7643 & n24924 ) ;
  assign n24926 = ( n2780 & n15228 ) | ( n2780 & ~n19353 ) | ( n15228 & ~n19353 ) ;
  assign n24927 = n20147 ^ n13009 ^ n8704 ;
  assign n24928 = ( n2181 & n24926 ) | ( n2181 & n24927 ) | ( n24926 & n24927 ) ;
  assign n24929 = n24928 ^ n21271 ^ n13062 ;
  assign n24931 = ( n169 & n594 ) | ( n169 & n1457 ) | ( n594 & n1457 ) ;
  assign n24930 = ( n5905 & n14891 ) | ( n5905 & n15443 ) | ( n14891 & n15443 ) ;
  assign n24932 = n24931 ^ n24930 ^ n15579 ;
  assign n24933 = ( n3847 & n14529 ) | ( n3847 & ~n21815 ) | ( n14529 & ~n21815 ) ;
  assign n24934 = n18617 ^ n17720 ^ n4863 ;
  assign n24935 = n24934 ^ n24145 ^ n6517 ;
  assign n24938 = n13150 ^ n4340 ^ x56 ;
  assign n24936 = ( n5959 & n6601 ) | ( n5959 & ~n10193 ) | ( n6601 & ~n10193 ) ;
  assign n24937 = n24936 ^ n11520 ^ n2027 ;
  assign n24939 = n24938 ^ n24937 ^ n14067 ;
  assign n24944 = n23755 ^ n19012 ^ n18205 ;
  assign n24941 = ( n720 & ~n4478 ) | ( n720 & n7842 ) | ( ~n4478 & n7842 ) ;
  assign n24942 = n24941 ^ n18423 ^ n14050 ;
  assign n24940 = ( ~n10238 & n10633 ) | ( ~n10238 & n13075 ) | ( n10633 & n13075 ) ;
  assign n24943 = n24942 ^ n24940 ^ n2761 ;
  assign n24945 = n24944 ^ n24943 ^ n3094 ;
  assign n24946 = ( n17460 & n19425 ) | ( n17460 & n22416 ) | ( n19425 & n22416 ) ;
  assign n24947 = n24946 ^ n11703 ^ n7982 ;
  assign n24948 = ( n181 & n6131 ) | ( n181 & n12682 ) | ( n6131 & n12682 ) ;
  assign n24949 = ( ~n502 & n4881 ) | ( ~n502 & n13728 ) | ( n4881 & n13728 ) ;
  assign n24950 = ( n18476 & ~n24948 ) | ( n18476 & n24949 ) | ( ~n24948 & n24949 ) ;
  assign n24951 = n24950 ^ n19445 ^ n2269 ;
  assign n24952 = ( n9219 & ~n15919 ) | ( n9219 & n24951 ) | ( ~n15919 & n24951 ) ;
  assign n24953 = ( ~n5944 & n11557 ) | ( ~n5944 & n16668 ) | ( n11557 & n16668 ) ;
  assign n24954 = ( ~n2164 & n9252 ) | ( ~n2164 & n20467 ) | ( n9252 & n20467 ) ;
  assign n24955 = ( n9820 & ~n24953 ) | ( n9820 & n24954 ) | ( ~n24953 & n24954 ) ;
  assign n24956 = ( ~n14179 & n21150 ) | ( ~n14179 & n22499 ) | ( n21150 & n22499 ) ;
  assign n24957 = ( ~n3917 & n24662 ) | ( ~n3917 & n24956 ) | ( n24662 & n24956 ) ;
  assign n24958 = n20795 ^ n17915 ^ n2138 ;
  assign n24959 = ( n21070 & ~n24708 ) | ( n21070 & n24958 ) | ( ~n24708 & n24958 ) ;
  assign n24960 = ( n15585 & ~n16284 ) | ( n15585 & n19888 ) | ( ~n16284 & n19888 ) ;
  assign n24961 = n13598 ^ n13334 ^ n11186 ;
  assign n24962 = n17648 ^ n15570 ^ n2803 ;
  assign n24963 = n24962 ^ n5685 ^ n5351 ;
  assign n24964 = ( n5805 & n17132 ) | ( n5805 & ~n23084 ) | ( n17132 & ~n23084 ) ;
  assign n24965 = n7890 ^ n2953 ^ n1704 ;
  assign n24966 = ( n10412 & n13287 ) | ( n10412 & n21398 ) | ( n13287 & n21398 ) ;
  assign n24971 = n11049 ^ n6849 ^ n6342 ;
  assign n24972 = ( n9469 & n13707 ) | ( n9469 & n24971 ) | ( n13707 & n24971 ) ;
  assign n24969 = n13089 ^ n7707 ^ n6150 ;
  assign n24970 = ( ~n970 & n12383 ) | ( ~n970 & n24969 ) | ( n12383 & n24969 ) ;
  assign n24967 = n21458 ^ n8016 ^ n5933 ;
  assign n24968 = n24967 ^ n22547 ^ n18348 ;
  assign n24973 = n24972 ^ n24970 ^ n24968 ;
  assign n24974 = ( n9531 & n11554 ) | ( n9531 & n13951 ) | ( n11554 & n13951 ) ;
  assign n24975 = n20013 ^ n6992 ^ n3688 ;
  assign n24976 = n24975 ^ n17464 ^ n8393 ;
  assign n24977 = n14664 ^ n10164 ^ n9304 ;
  assign n24978 = n24977 ^ n7985 ^ n4060 ;
  assign n24979 = n24978 ^ n11016 ^ x25 ;
  assign n24980 = ( n5713 & ~n17067 ) | ( n5713 & n21440 ) | ( ~n17067 & n21440 ) ;
  assign n24981 = n16042 ^ n10122 ^ n485 ;
  assign n24982 = ( n6289 & n8246 ) | ( n6289 & ~n20914 ) | ( n8246 & ~n20914 ) ;
  assign n24983 = n24982 ^ n16876 ^ n5159 ;
  assign n24984 = n22745 ^ n5805 ^ n1039 ;
  assign n24985 = ( ~n17613 & n20105 ) | ( ~n17613 & n21620 ) | ( n20105 & n21620 ) ;
  assign n24986 = ( n6360 & n7759 ) | ( n6360 & ~n14750 ) | ( n7759 & ~n14750 ) ;
  assign n24987 = n24798 ^ n18281 ^ n4996 ;
  assign n24988 = ( n12932 & ~n24986 ) | ( n12932 & n24987 ) | ( ~n24986 & n24987 ) ;
  assign n24991 = ( n1164 & n8962 ) | ( n1164 & n9412 ) | ( n8962 & n9412 ) ;
  assign n24989 = ( n4089 & ~n16076 ) | ( n4089 & n18744 ) | ( ~n16076 & n18744 ) ;
  assign n24990 = n24989 ^ n21644 ^ n1041 ;
  assign n24992 = n24991 ^ n24990 ^ n11584 ;
  assign n24993 = n24039 ^ n23787 ^ n3484 ;
  assign n24994 = ( ~n2562 & n10004 ) | ( ~n2562 & n15156 ) | ( n10004 & n15156 ) ;
  assign n24995 = n23543 ^ n22896 ^ n15975 ;
  assign n24996 = n10318 ^ n6196 ^ n4037 ;
  assign n24997 = ( n13629 & n15645 ) | ( n13629 & ~n24996 ) | ( n15645 & ~n24996 ) ;
  assign n24998 = n14714 ^ n8118 ^ n4593 ;
  assign n24999 = ( ~n587 & n23520 ) | ( ~n587 & n24998 ) | ( n23520 & n24998 ) ;
  assign n25000 = n20840 ^ n8389 ^ n7370 ;
  assign n25001 = n16657 ^ n14643 ^ n7761 ;
  assign n25002 = ( n982 & ~n11359 ) | ( n982 & n25001 ) | ( ~n11359 & n25001 ) ;
  assign n25003 = ( n4319 & ~n10060 ) | ( n4319 & n25002 ) | ( ~n10060 & n25002 ) ;
  assign n25004 = ( ~n4130 & n25000 ) | ( ~n4130 & n25003 ) | ( n25000 & n25003 ) ;
  assign n25007 = n11811 ^ n9009 ^ n2777 ;
  assign n25008 = n25007 ^ n16125 ^ n5982 ;
  assign n25006 = ( n2492 & ~n13761 ) | ( n2492 & n19638 ) | ( ~n13761 & n19638 ) ;
  assign n25005 = n22877 ^ n17596 ^ n16646 ;
  assign n25009 = n25008 ^ n25006 ^ n25005 ;
  assign n25010 = ( n1440 & ~n6232 ) | ( n1440 & n14889 ) | ( ~n6232 & n14889 ) ;
  assign n25011 = ( ~n11166 & n22363 ) | ( ~n11166 & n25010 ) | ( n22363 & n25010 ) ;
  assign n25012 = n25011 ^ n18542 ^ n1410 ;
  assign n25013 = n21723 ^ n18869 ^ n16780 ;
  assign n25014 = n18826 ^ n8583 ^ n5831 ;
  assign n25015 = ( n13283 & ~n16519 ) | ( n13283 & n25014 ) | ( ~n16519 & n25014 ) ;
  assign n25016 = n18217 ^ n1612 ^ n1603 ;
  assign n25017 = ( n4431 & n21994 ) | ( n4431 & n22853 ) | ( n21994 & n22853 ) ;
  assign n25018 = n19116 ^ n14852 ^ n6498 ;
  assign n25019 = ( n15023 & n16862 ) | ( n15023 & ~n23057 ) | ( n16862 & ~n23057 ) ;
  assign n25020 = ( n7302 & n16999 ) | ( n7302 & n19542 ) | ( n16999 & n19542 ) ;
  assign n25021 = ( x63 & n17383 ) | ( x63 & n25020 ) | ( n17383 & n25020 ) ;
  assign n25022 = ( n6406 & n6970 ) | ( n6406 & n18046 ) | ( n6970 & n18046 ) ;
  assign n25023 = ( ~n17110 & n19708 ) | ( ~n17110 & n25022 ) | ( n19708 & n25022 ) ;
  assign n25024 = n7204 ^ n6260 ^ n5260 ;
  assign n25025 = n25024 ^ n23536 ^ n16590 ;
  assign n25026 = n17511 ^ n15982 ^ n596 ;
  assign n25027 = n25026 ^ n9952 ^ n2892 ;
  assign n25028 = ( n2520 & ~n14016 ) | ( n2520 & n25027 ) | ( ~n14016 & n25027 ) ;
  assign n25029 = ( n1311 & ~n22796 ) | ( n1311 & n25028 ) | ( ~n22796 & n25028 ) ;
  assign n25030 = ( n3820 & ~n15420 ) | ( n3820 & n20104 ) | ( ~n15420 & n20104 ) ;
  assign n25035 = ( n3150 & ~n4515 ) | ( n3150 & n8341 ) | ( ~n4515 & n8341 ) ;
  assign n25036 = ( ~n17584 & n20016 ) | ( ~n17584 & n25035 ) | ( n20016 & n25035 ) ;
  assign n25031 = n19567 ^ n13511 ^ n1733 ;
  assign n25032 = ( n12847 & ~n24797 ) | ( n12847 & n25031 ) | ( ~n24797 & n25031 ) ;
  assign n25033 = n25032 ^ n5412 ^ x17 ;
  assign n25034 = ( n15554 & n19930 ) | ( n15554 & n25033 ) | ( n19930 & n25033 ) ;
  assign n25037 = n25036 ^ n25034 ^ n10363 ;
  assign n25038 = n15316 ^ n1762 ^ n997 ;
  assign n25039 = ( n7429 & n8306 ) | ( n7429 & n10958 ) | ( n8306 & n10958 ) ;
  assign n25040 = n25039 ^ n23573 ^ n9070 ;
  assign n25041 = n4903 ^ n2906 ^ n2673 ;
  assign n25042 = ( ~n957 & n6128 ) | ( ~n957 & n15054 ) | ( n6128 & n15054 ) ;
  assign n25043 = ( n13532 & ~n25041 ) | ( n13532 & n25042 ) | ( ~n25041 & n25042 ) ;
  assign n25044 = n19351 ^ n5161 ^ n2067 ;
  assign n25045 = ( n3650 & n9816 ) | ( n3650 & ~n25044 ) | ( n9816 & ~n25044 ) ;
  assign n25046 = ( n4319 & ~n8548 ) | ( n4319 & n25045 ) | ( ~n8548 & n25045 ) ;
  assign n25047 = n19410 ^ n6914 ^ n5699 ;
  assign n25048 = ( n6713 & n7481 ) | ( n6713 & n25047 ) | ( n7481 & n25047 ) ;
  assign n25049 = n25048 ^ n21165 ^ n3857 ;
  assign n25050 = ( n814 & n17545 ) | ( n814 & n22973 ) | ( n17545 & n22973 ) ;
  assign n25051 = ( n5195 & n15573 ) | ( n5195 & n25050 ) | ( n15573 & n25050 ) ;
  assign n25053 = ( n3989 & n4086 ) | ( n3989 & n24555 ) | ( n4086 & n24555 ) ;
  assign n25052 = n22672 ^ n6686 ^ n282 ;
  assign n25054 = n25053 ^ n25052 ^ n9956 ;
  assign n25055 = n19643 ^ n15278 ^ n6351 ;
  assign n25056 = n14127 ^ n1620 ^ n479 ;
  assign n25057 = ( n621 & n16284 ) | ( n621 & ~n25056 ) | ( n16284 & ~n25056 ) ;
  assign n25058 = ( n7145 & ~n8195 ) | ( n7145 & n11640 ) | ( ~n8195 & n11640 ) ;
  assign n25059 = n23000 ^ n14722 ^ n5928 ;
  assign n25060 = ( n7797 & n8299 ) | ( n7797 & ~n17158 ) | ( n8299 & ~n17158 ) ;
  assign n25061 = ( n10519 & n13021 ) | ( n10519 & n25060 ) | ( n13021 & n25060 ) ;
  assign n25062 = n19673 ^ n4352 ^ n3654 ;
  assign n25063 = ( n4577 & ~n10053 ) | ( n4577 & n25062 ) | ( ~n10053 & n25062 ) ;
  assign n25064 = n25063 ^ n24110 ^ n14094 ;
  assign n25065 = n25064 ^ n11099 ^ n6907 ;
  assign n25067 = n11441 ^ n6108 ^ n506 ;
  assign n25066 = ( ~n1786 & n9110 ) | ( ~n1786 & n15851 ) | ( n9110 & n15851 ) ;
  assign n25068 = n25067 ^ n25066 ^ n4919 ;
  assign n25071 = n9802 ^ n7340 ^ n1900 ;
  assign n25069 = n13140 ^ n6736 ^ n4003 ;
  assign n25070 = n25069 ^ n22614 ^ n11260 ;
  assign n25072 = n25071 ^ n25070 ^ n2607 ;
  assign n25073 = n12526 ^ n9561 ^ n5256 ;
  assign n25074 = ( n5174 & n12068 ) | ( n5174 & ~n15997 ) | ( n12068 & ~n15997 ) ;
  assign n25075 = ( n7303 & ~n25073 ) | ( n7303 & n25074 ) | ( ~n25073 & n25074 ) ;
  assign n25076 = ( n15281 & n25072 ) | ( n15281 & n25075 ) | ( n25072 & n25075 ) ;
  assign n25077 = n9281 ^ n2495 ^ n2238 ;
  assign n25078 = n19563 ^ n15940 ^ n4742 ;
  assign n25079 = n17871 ^ n6603 ^ n196 ;
  assign n25080 = ( ~n2352 & n13072 ) | ( ~n2352 & n14335 ) | ( n13072 & n14335 ) ;
  assign n25082 = n18595 ^ n7337 ^ n4868 ;
  assign n25083 = ( n18103 & n24658 ) | ( n18103 & n25082 ) | ( n24658 & n25082 ) ;
  assign n25081 = n20143 ^ n19415 ^ n2508 ;
  assign n25084 = n25083 ^ n25081 ^ n165 ;
  assign n25085 = n18995 ^ n14218 ^ n4454 ;
  assign n25086 = ( ~n3934 & n20579 ) | ( ~n3934 & n25085 ) | ( n20579 & n25085 ) ;
  assign n25087 = ( ~n11433 & n15245 ) | ( ~n11433 & n25086 ) | ( n15245 & n25086 ) ;
  assign n25088 = n23252 ^ n7457 ^ n2364 ;
  assign n25089 = n22240 ^ n19299 ^ n11927 ;
  assign n25090 = ( ~n1505 & n2165 ) | ( ~n1505 & n4272 ) | ( n2165 & n4272 ) ;
  assign n25091 = ( ~n5842 & n12610 ) | ( ~n5842 & n17835 ) | ( n12610 & n17835 ) ;
  assign n25095 = ( ~n1057 & n3101 ) | ( ~n1057 & n9526 ) | ( n3101 & n9526 ) ;
  assign n25092 = n15289 ^ n14110 ^ n1343 ;
  assign n25093 = ( n12193 & n21148 ) | ( n12193 & n25092 ) | ( n21148 & n25092 ) ;
  assign n25094 = ( n12444 & ~n20975 ) | ( n12444 & n25093 ) | ( ~n20975 & n25093 ) ;
  assign n25096 = n25095 ^ n25094 ^ n24557 ;
  assign n25097 = n10232 ^ n8919 ^ n913 ;
  assign n25098 = n25097 ^ n7686 ^ n2774 ;
  assign n25099 = ( ~n2972 & n22103 ) | ( ~n2972 & n25098 ) | ( n22103 & n25098 ) ;
  assign n25100 = n10974 ^ n8851 ^ n4706 ;
  assign n25101 = ( ~n429 & n8765 ) | ( ~n429 & n20125 ) | ( n8765 & n20125 ) ;
  assign n25102 = n25101 ^ n16190 ^ n8637 ;
  assign n25103 = n25102 ^ n13842 ^ n7435 ;
  assign n25104 = n19623 ^ n5959 ^ n4003 ;
  assign n25107 = ( ~n211 & n11392 ) | ( ~n211 & n24937 ) | ( n11392 & n24937 ) ;
  assign n25105 = n24491 ^ n5777 ^ n1163 ;
  assign n25106 = ( ~n6303 & n7095 ) | ( ~n6303 & n25105 ) | ( n7095 & n25105 ) ;
  assign n25108 = n25107 ^ n25106 ^ n7382 ;
  assign n25114 = ( n6102 & n10696 ) | ( n6102 & ~n16248 ) | ( n10696 & ~n16248 ) ;
  assign n25109 = n7041 ^ n5177 ^ n3559 ;
  assign n25110 = ( n4258 & n6999 ) | ( n4258 & ~n25109 ) | ( n6999 & ~n25109 ) ;
  assign n25111 = n4347 ^ n3656 ^ n702 ;
  assign n25112 = ( ~n17695 & n25110 ) | ( ~n17695 & n25111 ) | ( n25110 & n25111 ) ;
  assign n25113 = n25112 ^ n15846 ^ n13873 ;
  assign n25115 = n25114 ^ n25113 ^ n5945 ;
  assign n25116 = ( n7572 & n10297 ) | ( n7572 & n19298 ) | ( n10297 & n19298 ) ;
  assign n25117 = ( n13903 & ~n22169 ) | ( n13903 & n25116 ) | ( ~n22169 & n25116 ) ;
  assign n25118 = n21895 ^ n16744 ^ n10294 ;
  assign n25119 = ( n8615 & n13627 ) | ( n8615 & ~n25118 ) | ( n13627 & ~n25118 ) ;
  assign n25120 = n22318 ^ n18857 ^ n4199 ;
  assign n25121 = ( n764 & n3359 ) | ( n764 & ~n12680 ) | ( n3359 & ~n12680 ) ;
  assign n25122 = n8354 ^ n5997 ^ n5920 ;
  assign n25123 = n18948 ^ n11201 ^ n3630 ;
  assign n25124 = ( n5486 & n21321 ) | ( n5486 & ~n25123 ) | ( n21321 & ~n25123 ) ;
  assign n25126 = ( n7874 & n11791 ) | ( n7874 & ~n15437 ) | ( n11791 & ~n15437 ) ;
  assign n25125 = n24134 ^ n22684 ^ n9910 ;
  assign n25127 = n25126 ^ n25125 ^ n12683 ;
  assign n25128 = n20206 ^ n14351 ^ n1552 ;
  assign n25129 = ( n472 & n22247 ) | ( n472 & n23776 ) | ( n22247 & n23776 ) ;
  assign n25130 = ( n1647 & n1800 ) | ( n1647 & n12864 ) | ( n1800 & n12864 ) ;
  assign n25131 = n25130 ^ n19632 ^ n16571 ;
  assign n25132 = n24431 ^ n10698 ^ n706 ;
  assign n25133 = ( n4675 & n5087 ) | ( n4675 & n25132 ) | ( n5087 & n25132 ) ;
  assign n25134 = n25133 ^ n12911 ^ n9926 ;
  assign n25135 = n10638 ^ n8533 ^ n702 ;
  assign n25136 = ( n4769 & ~n14381 ) | ( n4769 & n16994 ) | ( ~n14381 & n16994 ) ;
  assign n25140 = ( n2066 & ~n3128 ) | ( n2066 & n5849 ) | ( ~n3128 & n5849 ) ;
  assign n25141 = ( n2380 & n2525 ) | ( n2380 & n25140 ) | ( n2525 & n25140 ) ;
  assign n25139 = ( n2077 & n4599 ) | ( n2077 & n12320 ) | ( n4599 & n12320 ) ;
  assign n25137 = ( n4027 & n6296 ) | ( n4027 & ~n21776 ) | ( n6296 & ~n21776 ) ;
  assign n25138 = n25137 ^ n13850 ^ n8918 ;
  assign n25142 = n25141 ^ n25139 ^ n25138 ;
  assign n25143 = n12771 ^ n10775 ^ n10183 ;
  assign n25144 = n25143 ^ n10257 ^ n829 ;
  assign n25145 = ( n15095 & n17831 ) | ( n15095 & ~n25144 ) | ( n17831 & ~n25144 ) ;
  assign n25146 = n17927 ^ n15248 ^ n7407 ;
  assign n25147 = ( ~n4937 & n9762 ) | ( ~n4937 & n25146 ) | ( n9762 & n25146 ) ;
  assign n25148 = ( n4174 & ~n11143 ) | ( n4174 & n25147 ) | ( ~n11143 & n25147 ) ;
  assign n25149 = ( n8537 & ~n23912 ) | ( n8537 & n25148 ) | ( ~n23912 & n25148 ) ;
  assign n25150 = ( n5101 & n15351 ) | ( n5101 & n24628 ) | ( n15351 & n24628 ) ;
  assign n25151 = n16628 ^ n7996 ^ n4360 ;
  assign n25152 = ( n1650 & ~n4904 ) | ( n1650 & n5635 ) | ( ~n4904 & n5635 ) ;
  assign n25153 = n25152 ^ n7110 ^ n6212 ;
  assign n25154 = n20479 ^ n13896 ^ n1785 ;
  assign n25155 = ( n10958 & ~n11136 ) | ( n10958 & n25154 ) | ( ~n11136 & n25154 ) ;
  assign n25156 = ( ~n14386 & n25153 ) | ( ~n14386 & n25155 ) | ( n25153 & n25155 ) ;
  assign n25157 = ( n7878 & ~n14788 ) | ( n7878 & n16466 ) | ( ~n14788 & n16466 ) ;
  assign n25158 = n23549 ^ n21248 ^ n6807 ;
  assign n25159 = n15899 ^ n8383 ^ n5918 ;
  assign n25160 = ( n1064 & n1125 ) | ( n1064 & ~n25159 ) | ( n1125 & ~n25159 ) ;
  assign n25161 = ( n7426 & n10038 ) | ( n7426 & ~n18858 ) | ( n10038 & ~n18858 ) ;
  assign n25162 = ( n10124 & n25160 ) | ( n10124 & ~n25161 ) | ( n25160 & ~n25161 ) ;
  assign n25163 = ( n3977 & n25158 ) | ( n3977 & n25162 ) | ( n25158 & n25162 ) ;
  assign n25164 = n25163 ^ n5095 ^ n3770 ;
  assign n25165 = ( n431 & ~n1729 ) | ( n431 & n9008 ) | ( ~n1729 & n9008 ) ;
  assign n25166 = n25165 ^ n20431 ^ n3774 ;
  assign n25167 = n5864 ^ n2695 ^ n2270 ;
  assign n25168 = n25167 ^ n2984 ^ n2665 ;
  assign n25169 = n16026 ^ n7312 ^ n1353 ;
  assign n25170 = n10351 ^ n7732 ^ n4908 ;
  assign n25171 = ( n2121 & n3077 ) | ( n2121 & n13646 ) | ( n3077 & n13646 ) ;
  assign n25172 = ( n911 & ~n11783 ) | ( n911 & n12581 ) | ( ~n11783 & n12581 ) ;
  assign n25173 = ( ~n9678 & n22941 ) | ( ~n9678 & n23121 ) | ( n22941 & n23121 ) ;
  assign n25174 = ( ~n21260 & n25172 ) | ( ~n21260 & n25173 ) | ( n25172 & n25173 ) ;
  assign n25182 = n18249 ^ n13887 ^ n6370 ;
  assign n25175 = n12763 ^ n6972 ^ n6760 ;
  assign n25179 = ( n15154 & n16941 ) | ( n15154 & ~n21814 ) | ( n16941 & ~n21814 ) ;
  assign n25176 = n12663 ^ n1620 ^ n604 ;
  assign n25177 = ( ~n15308 & n16718 ) | ( ~n15308 & n19186 ) | ( n16718 & n19186 ) ;
  assign n25178 = ( n9477 & ~n25176 ) | ( n9477 & n25177 ) | ( ~n25176 & n25177 ) ;
  assign n25180 = n25179 ^ n25178 ^ n164 ;
  assign n25181 = ( n3948 & ~n25175 ) | ( n3948 & n25180 ) | ( ~n25175 & n25180 ) ;
  assign n25183 = n25182 ^ n25181 ^ n11953 ;
  assign n25185 = ( n6323 & n10802 ) | ( n6323 & n17508 ) | ( n10802 & n17508 ) ;
  assign n25184 = n14585 ^ n4222 ^ n2111 ;
  assign n25186 = n25185 ^ n25184 ^ n12644 ;
  assign n25187 = n25186 ^ n17577 ^ n14529 ;
  assign n25188 = n23687 ^ n3340 ^ n3269 ;
  assign n25189 = n25188 ^ n23068 ^ n10071 ;
  assign n25190 = ( n1452 & n1861 ) | ( n1452 & ~n14909 ) | ( n1861 & ~n14909 ) ;
  assign n25191 = ( n5559 & n12624 ) | ( n5559 & n17582 ) | ( n12624 & n17582 ) ;
  assign n25192 = ( n7156 & n7607 ) | ( n7156 & ~n13004 ) | ( n7607 & ~n13004 ) ;
  assign n25197 = n18994 ^ n6278 ^ n3552 ;
  assign n25193 = ( ~n2525 & n5651 ) | ( ~n2525 & n21697 ) | ( n5651 & n21697 ) ;
  assign n25194 = ( n1971 & ~n5237 ) | ( n1971 & n25193 ) | ( ~n5237 & n25193 ) ;
  assign n25195 = n9972 ^ n7239 ^ n1360 ;
  assign n25196 = ( n8877 & ~n25194 ) | ( n8877 & n25195 ) | ( ~n25194 & n25195 ) ;
  assign n25198 = n25197 ^ n25196 ^ n23123 ;
  assign n25199 = ( n2230 & ~n9314 ) | ( n2230 & n22073 ) | ( ~n9314 & n22073 ) ;
  assign n25200 = n25199 ^ n18891 ^ n11534 ;
  assign n25201 = ( n8568 & n18425 ) | ( n8568 & ~n25200 ) | ( n18425 & ~n25200 ) ;
  assign n25202 = ( n10828 & n14996 ) | ( n10828 & ~n20109 ) | ( n14996 & ~n20109 ) ;
  assign n25203 = ( n9980 & n25201 ) | ( n9980 & ~n25202 ) | ( n25201 & ~n25202 ) ;
  assign n25204 = ( n6183 & n10545 ) | ( n6183 & n13286 ) | ( n10545 & n13286 ) ;
  assign n25205 = n17558 ^ n7000 ^ n6978 ;
  assign n25206 = ( ~n761 & n17980 ) | ( ~n761 & n25205 ) | ( n17980 & n25205 ) ;
  assign n25207 = n10926 ^ n1954 ^ n1880 ;
  assign n25208 = ( n14825 & n15064 ) | ( n14825 & n25207 ) | ( n15064 & n25207 ) ;
  assign n25215 = n13608 ^ n11939 ^ n7759 ;
  assign n25209 = ( ~n590 & n3554 ) | ( ~n590 & n12833 ) | ( n3554 & n12833 ) ;
  assign n25210 = ( n1981 & ~n2054 ) | ( n1981 & n4083 ) | ( ~n2054 & n4083 ) ;
  assign n25211 = ( n163 & n25209 ) | ( n163 & ~n25210 ) | ( n25209 & ~n25210 ) ;
  assign n25212 = n25211 ^ n21236 ^ n11171 ;
  assign n25213 = ( n5195 & n5802 ) | ( n5195 & ~n25212 ) | ( n5802 & ~n25212 ) ;
  assign n25214 = ( n6123 & ~n16015 ) | ( n6123 & n25213 ) | ( ~n16015 & n25213 ) ;
  assign n25216 = n25215 ^ n25214 ^ n21167 ;
  assign n25217 = ( n2660 & ~n18360 ) | ( n2660 & n19637 ) | ( ~n18360 & n19637 ) ;
  assign n25218 = n19679 ^ n17234 ^ n5856 ;
  assign n25220 = n7382 ^ n3492 ^ n3356 ;
  assign n25219 = ( ~n15453 & n16379 ) | ( ~n15453 & n19268 ) | ( n16379 & n19268 ) ;
  assign n25221 = n25220 ^ n25219 ^ n2746 ;
  assign n25222 = n25221 ^ n13185 ^ n12186 ;
  assign n25223 = ( n6315 & n6452 ) | ( n6315 & n9138 ) | ( n6452 & n9138 ) ;
  assign n25224 = ( n442 & ~n1106 ) | ( n442 & n2200 ) | ( ~n1106 & n2200 ) ;
  assign n25225 = n25224 ^ n19942 ^ n14620 ;
  assign n25226 = n4925 ^ n3090 ^ n1096 ;
  assign n25227 = ( n4235 & n14005 ) | ( n4235 & n25226 ) | ( n14005 & n25226 ) ;
  assign n25228 = n11338 ^ n7674 ^ n4526 ;
  assign n25229 = ( n5987 & n10454 ) | ( n5987 & n25228 ) | ( n10454 & n25228 ) ;
  assign n25230 = n14328 ^ n13695 ^ n374 ;
  assign n25231 = n25230 ^ n21262 ^ n6727 ;
  assign n25232 = ( n3654 & n15281 ) | ( n3654 & ~n15728 ) | ( n15281 & ~n15728 ) ;
  assign n25233 = ( n3518 & n15361 ) | ( n3518 & ~n25232 ) | ( n15361 & ~n25232 ) ;
  assign n25234 = n17467 ^ n11702 ^ n4870 ;
  assign n25235 = n23022 ^ n21160 ^ n12379 ;
  assign n25236 = n15668 ^ n14288 ^ n716 ;
  assign n25237 = ( n11488 & ~n19674 ) | ( n11488 & n25236 ) | ( ~n19674 & n25236 ) ;
  assign n25240 = ( ~n1209 & n5396 ) | ( ~n1209 & n9348 ) | ( n5396 & n9348 ) ;
  assign n25238 = ( n967 & n10630 ) | ( n967 & ~n20841 ) | ( n10630 & ~n20841 ) ;
  assign n25239 = ( ~n5723 & n12473 ) | ( ~n5723 & n25238 ) | ( n12473 & n25238 ) ;
  assign n25241 = n25240 ^ n25239 ^ n8691 ;
  assign n25242 = n25241 ^ n10539 ^ n1178 ;
  assign n25243 = n12190 ^ n9063 ^ n1832 ;
  assign n25244 = ( n334 & n6795 ) | ( n334 & n13739 ) | ( n6795 & n13739 ) ;
  assign n25245 = n25244 ^ n25139 ^ n14150 ;
  assign n25246 = ( ~n5734 & n6610 ) | ( ~n5734 & n21401 ) | ( n6610 & n21401 ) ;
  assign n25247 = n15149 ^ n8718 ^ n8690 ;
  assign n25248 = n25247 ^ n17566 ^ n5573 ;
  assign n25249 = ( n12433 & n25246 ) | ( n12433 & ~n25248 ) | ( n25246 & ~n25248 ) ;
  assign n25250 = ( n2856 & n9882 ) | ( n2856 & n17928 ) | ( n9882 & n17928 ) ;
  assign n25251 = ( n11134 & n12781 ) | ( n11134 & n21118 ) | ( n12781 & n21118 ) ;
  assign n25253 = ( n2085 & ~n3651 ) | ( n2085 & n4977 ) | ( ~n3651 & n4977 ) ;
  assign n25252 = ( ~n2082 & n10582 ) | ( ~n2082 & n18338 ) | ( n10582 & n18338 ) ;
  assign n25254 = n25253 ^ n25252 ^ n7820 ;
  assign n25255 = ( n6185 & ~n9725 ) | ( n6185 & n25254 ) | ( ~n9725 & n25254 ) ;
  assign n25256 = n25255 ^ n20086 ^ x14 ;
  assign n25258 = n11529 ^ n3968 ^ n242 ;
  assign n25259 = ( ~n740 & n20654 ) | ( ~n740 & n25258 ) | ( n20654 & n25258 ) ;
  assign n25257 = ( n1545 & ~n19394 ) | ( n1545 & n22068 ) | ( ~n19394 & n22068 ) ;
  assign n25260 = n25259 ^ n25257 ^ n285 ;
  assign n25261 = ( n6671 & n10018 ) | ( n6671 & ~n14516 ) | ( n10018 & ~n14516 ) ;
  assign n25264 = ( ~n4351 & n16492 ) | ( ~n4351 & n21209 ) | ( n16492 & n21209 ) ;
  assign n25262 = ( n4689 & n6768 ) | ( n4689 & n9586 ) | ( n6768 & n9586 ) ;
  assign n25263 = n25262 ^ n23449 ^ n21349 ;
  assign n25265 = n25264 ^ n25263 ^ n1178 ;
  assign n25266 = ( n15189 & n16252 ) | ( n15189 & ~n17055 ) | ( n16252 & ~n17055 ) ;
  assign n25267 = n9346 ^ n9304 ^ n8708 ;
  assign n25268 = n25267 ^ n13711 ^ n11356 ;
  assign n25269 = ( ~n23256 & n25069 ) | ( ~n23256 & n25268 ) | ( n25069 & n25268 ) ;
  assign n25270 = n22899 ^ n7419 ^ n2444 ;
  assign n25271 = n23895 ^ n21897 ^ n1005 ;
  assign n25272 = ( n7986 & ~n21271 ) | ( n7986 & n21550 ) | ( ~n21271 & n21550 ) ;
  assign n25273 = ( n866 & n3109 ) | ( n866 & ~n10619 ) | ( n3109 & ~n10619 ) ;
  assign n25274 = n25273 ^ n13874 ^ n4962 ;
  assign n25275 = ( n2785 & n10869 ) | ( n2785 & n14794 ) | ( n10869 & n14794 ) ;
  assign n25276 = ( ~n9139 & n23035 ) | ( ~n9139 & n25275 ) | ( n23035 & n25275 ) ;
  assign n25277 = n23849 ^ n12647 ^ n6442 ;
  assign n25278 = ( n5618 & ~n10065 ) | ( n5618 & n25026 ) | ( ~n10065 & n25026 ) ;
  assign n25279 = n2308 ^ n1852 ^ n459 ;
  assign n25280 = n13013 ^ n5146 ^ n4013 ;
  assign n25281 = n25280 ^ n17652 ^ n14420 ;
  assign n25282 = ( n702 & ~n25279 ) | ( n702 & n25281 ) | ( ~n25279 & n25281 ) ;
  assign n25283 = n14051 ^ n9438 ^ n7925 ;
  assign n25284 = ( n3048 & ~n10365 ) | ( n3048 & n25283 ) | ( ~n10365 & n25283 ) ;
  assign n25285 = ( ~n8846 & n20503 ) | ( ~n8846 & n23329 ) | ( n20503 & n23329 ) ;
  assign n25286 = ( n5610 & n23923 ) | ( n5610 & ~n25285 ) | ( n23923 & ~n25285 ) ;
  assign n25287 = n24874 ^ n14680 ^ n13846 ;
  assign n25288 = n25287 ^ n5312 ^ n775 ;
  assign n25289 = ( ~n25284 & n25286 ) | ( ~n25284 & n25288 ) | ( n25286 & n25288 ) ;
  assign n25290 = ( n7475 & n10249 ) | ( n7475 & n22671 ) | ( n10249 & n22671 ) ;
  assign n25291 = n25290 ^ n17817 ^ n7727 ;
  assign n25292 = n11148 ^ n8413 ^ n5604 ;
  assign n25293 = ( n14768 & n20390 ) | ( n14768 & ~n25292 ) | ( n20390 & ~n25292 ) ;
  assign n25294 = ( n747 & n16502 ) | ( n747 & ~n21346 ) | ( n16502 & ~n21346 ) ;
  assign n25295 = ( n2978 & n21783 ) | ( n2978 & ~n23182 ) | ( n21783 & ~n23182 ) ;
  assign n25296 = ( ~n8953 & n25294 ) | ( ~n8953 & n25295 ) | ( n25294 & n25295 ) ;
  assign n25297 = n23256 ^ n13866 ^ n9553 ;
  assign n25298 = n25297 ^ n16383 ^ n442 ;
  assign n25299 = n18809 ^ n10473 ^ n9235 ;
  assign n25300 = ( n25296 & ~n25298 ) | ( n25296 & n25299 ) | ( ~n25298 & n25299 ) ;
  assign n25301 = n16865 ^ n6739 ^ n1166 ;
  assign n25302 = ( ~n3865 & n5779 ) | ( ~n3865 & n19973 ) | ( n5779 & n19973 ) ;
  assign n25303 = ( n4245 & n10349 ) | ( n4245 & n25302 ) | ( n10349 & n25302 ) ;
  assign n25304 = ( n2020 & ~n7409 ) | ( n2020 & n18737 ) | ( ~n7409 & n18737 ) ;
  assign n25305 = n15168 ^ n10028 ^ n4990 ;
  assign n25306 = ( n5474 & n8026 ) | ( n5474 & ~n24784 ) | ( n8026 & ~n24784 ) ;
  assign n25307 = ( ~n4716 & n5466 ) | ( ~n4716 & n9270 ) | ( n5466 & n9270 ) ;
  assign n25308 = ( ~n1417 & n9787 ) | ( ~n1417 & n15642 ) | ( n9787 & n15642 ) ;
  assign n25309 = n25308 ^ n13470 ^ n4323 ;
  assign n25310 = ( ~n7851 & n16041 ) | ( ~n7851 & n22140 ) | ( n16041 & n22140 ) ;
  assign n25311 = ( ~n8432 & n9483 ) | ( ~n8432 & n12397 ) | ( n9483 & n12397 ) ;
  assign n25312 = ( n1178 & n5866 ) | ( n1178 & n25311 ) | ( n5866 & n25311 ) ;
  assign n25313 = n25312 ^ n10925 ^ n8332 ;
  assign n25314 = ( n12368 & n15272 ) | ( n12368 & ~n25313 ) | ( n15272 & ~n25313 ) ;
  assign n25315 = n25314 ^ n21829 ^ n3100 ;
  assign n25316 = ( n462 & ~n16174 ) | ( n462 & n17017 ) | ( ~n16174 & n17017 ) ;
  assign n25317 = n19018 ^ n7913 ^ n4338 ;
  assign n25318 = ( n5539 & ~n9051 ) | ( n5539 & n16757 ) | ( ~n9051 & n16757 ) ;
  assign n25319 = n7808 ^ n5587 ^ n3839 ;
  assign n25321 = ( ~n1288 & n11026 ) | ( ~n1288 & n16146 ) | ( n11026 & n16146 ) ;
  assign n25320 = ( n8950 & ~n15202 ) | ( n8950 & n23568 ) | ( ~n15202 & n23568 ) ;
  assign n25322 = n25321 ^ n25320 ^ n9503 ;
  assign n25323 = ( n7172 & n7949 ) | ( n7172 & n21274 ) | ( n7949 & n21274 ) ;
  assign n25324 = ( n762 & ~n6866 ) | ( n762 & n12625 ) | ( ~n6866 & n12625 ) ;
  assign n25325 = n25324 ^ n13474 ^ n1604 ;
  assign n25330 = n10735 ^ n10264 ^ n8217 ;
  assign n25326 = ( ~n3761 & n4425 ) | ( ~n3761 & n19266 ) | ( n4425 & n19266 ) ;
  assign n25327 = ( n2259 & n3080 ) | ( n2259 & ~n18862 ) | ( n3080 & ~n18862 ) ;
  assign n25328 = ( n6709 & n25326 ) | ( n6709 & ~n25327 ) | ( n25326 & ~n25327 ) ;
  assign n25329 = ( n359 & ~n9900 ) | ( n359 & n25328 ) | ( ~n9900 & n25328 ) ;
  assign n25331 = n25330 ^ n25329 ^ n13285 ;
  assign n25332 = ( n906 & ~n1082 ) | ( n906 & n8614 ) | ( ~n1082 & n8614 ) ;
  assign n25333 = n25332 ^ n17731 ^ n15878 ;
  assign n25334 = n25333 ^ n23874 ^ n5349 ;
  assign n25335 = ( n14191 & ~n15214 ) | ( n14191 & n24251 ) | ( ~n15214 & n24251 ) ;
  assign n25336 = ( n12885 & ~n17721 ) | ( n12885 & n18253 ) | ( ~n17721 & n18253 ) ;
  assign n25342 = n10961 ^ n5883 ^ n2465 ;
  assign n25337 = n5311 ^ n3382 ^ n1515 ;
  assign n25338 = ( ~n1345 & n3522 ) | ( ~n1345 & n25337 ) | ( n3522 & n25337 ) ;
  assign n25339 = n25338 ^ n7870 ^ n2957 ;
  assign n25340 = ( n15244 & n24688 ) | ( n15244 & n25339 ) | ( n24688 & n25339 ) ;
  assign n25341 = ( ~n625 & n10465 ) | ( ~n625 & n25340 ) | ( n10465 & n25340 ) ;
  assign n25343 = n25342 ^ n25341 ^ n3061 ;
  assign n25344 = n25343 ^ n17652 ^ n11829 ;
  assign n25345 = n19956 ^ n17513 ^ n10597 ;
  assign n25346 = n14062 ^ n10665 ^ n6933 ;
  assign n25347 = n25346 ^ n15113 ^ n5781 ;
  assign n25348 = ( n1642 & n13533 ) | ( n1642 & ~n14854 ) | ( n13533 & ~n14854 ) ;
  assign n25349 = ( n14779 & n23029 ) | ( n14779 & ~n25348 ) | ( n23029 & ~n25348 ) ;
  assign n25350 = n19815 ^ n18150 ^ n3403 ;
  assign n25351 = n13868 ^ n12585 ^ n4869 ;
  assign n25352 = n25351 ^ n23868 ^ n3494 ;
  assign n25353 = ( ~n1429 & n8616 ) | ( ~n1429 & n8647 ) | ( n8616 & n8647 ) ;
  assign n25354 = ( n2114 & n25109 ) | ( n2114 & ~n25353 ) | ( n25109 & ~n25353 ) ;
  assign n25355 = n25354 ^ n10806 ^ n1429 ;
  assign n25356 = ( n6281 & n10054 ) | ( n6281 & n25355 ) | ( n10054 & n25355 ) ;
  assign n25357 = ( n25350 & n25352 ) | ( n25350 & ~n25356 ) | ( n25352 & ~n25356 ) ;
  assign n25358 = n25357 ^ n8171 ^ n7574 ;
  assign n25359 = ( n10531 & ~n17486 ) | ( n10531 & n21996 ) | ( ~n17486 & n21996 ) ;
  assign n25360 = ( n4741 & ~n9150 ) | ( n4741 & n13598 ) | ( ~n9150 & n13598 ) ;
  assign n25363 = ( n1988 & n2095 ) | ( n1988 & ~n2803 ) | ( n2095 & ~n2803 ) ;
  assign n25361 = ( n3704 & n10071 ) | ( n3704 & n23734 ) | ( n10071 & n23734 ) ;
  assign n25362 = n25361 ^ n14016 ^ n13544 ;
  assign n25364 = n25363 ^ n25362 ^ n22249 ;
  assign n25365 = n18376 ^ n16419 ^ n15364 ;
  assign n25366 = n17026 ^ n14304 ^ n10671 ;
  assign n25367 = ( x44 & ~n1972 ) | ( x44 & n25366 ) | ( ~n1972 & n25366 ) ;
  assign n25368 = ( n4111 & n5193 ) | ( n4111 & ~n6168 ) | ( n5193 & ~n6168 ) ;
  assign n25369 = ( ~n7590 & n14990 ) | ( ~n7590 & n25368 ) | ( n14990 & n25368 ) ;
  assign n25370 = ( n15733 & n25137 ) | ( n15733 & ~n25369 ) | ( n25137 & ~n25369 ) ;
  assign n25371 = n15574 ^ n6491 ^ n736 ;
  assign n25372 = ( n1410 & n13211 ) | ( n1410 & ~n25371 ) | ( n13211 & ~n25371 ) ;
  assign n25373 = n25372 ^ n14035 ^ n11990 ;
  assign n25374 = ( n757 & ~n25370 ) | ( n757 & n25373 ) | ( ~n25370 & n25373 ) ;
  assign n25375 = ( ~n12733 & n25367 ) | ( ~n12733 & n25374 ) | ( n25367 & n25374 ) ;
  assign n25376 = ( x28 & ~n4907 ) | ( x28 & n5987 ) | ( ~n4907 & n5987 ) ;
  assign n25377 = n25376 ^ n7773 ^ n3318 ;
  assign n25378 = n25377 ^ n15727 ^ n9589 ;
  assign n25379 = n13041 ^ n11259 ^ n6979 ;
  assign n25380 = n25379 ^ n13737 ^ n1400 ;
  assign n25381 = n25380 ^ n13445 ^ n9420 ;
  assign n25382 = ( n396 & n25378 ) | ( n396 & ~n25381 ) | ( n25378 & ~n25381 ) ;
  assign n25383 = ( n6496 & n6624 ) | ( n6496 & ~n19087 ) | ( n6624 & ~n19087 ) ;
  assign n25384 = n22540 ^ n12523 ^ n1830 ;
  assign n25385 = n25384 ^ n6129 ^ n1652 ;
  assign n25386 = ( n6301 & ~n13408 ) | ( n6301 & n24941 ) | ( ~n13408 & n24941 ) ;
  assign n25387 = ( n5679 & ~n24049 ) | ( n5679 & n25386 ) | ( ~n24049 & n25386 ) ;
  assign n25388 = n12661 ^ n11013 ^ n431 ;
  assign n25389 = ( n6072 & n8449 ) | ( n6072 & n9155 ) | ( n8449 & n9155 ) ;
  assign n25390 = ( n4063 & n15341 ) | ( n4063 & ~n18453 ) | ( n15341 & ~n18453 ) ;
  assign n25391 = ( n2275 & n25389 ) | ( n2275 & n25390 ) | ( n25389 & n25390 ) ;
  assign n25392 = n25391 ^ n19246 ^ n6852 ;
  assign n25393 = ( n16530 & n25388 ) | ( n16530 & ~n25392 ) | ( n25388 & ~n25392 ) ;
  assign n25394 = ( n5042 & ~n17401 ) | ( n5042 & n17575 ) | ( ~n17401 & n17575 ) ;
  assign n25395 = ( n16574 & n18344 ) | ( n16574 & ~n19123 ) | ( n18344 & ~n19123 ) ;
  assign n25396 = ( n3340 & n6347 ) | ( n3340 & n22032 ) | ( n6347 & n22032 ) ;
  assign n25397 = ( n6901 & ~n10693 ) | ( n6901 & n25396 ) | ( ~n10693 & n25396 ) ;
  assign n25398 = n11990 ^ n8079 ^ n1156 ;
  assign n25399 = n25398 ^ n20510 ^ n812 ;
  assign n25400 = n7784 ^ n3142 ^ n2232 ;
  assign n25401 = n25400 ^ n7125 ^ n5151 ;
  assign n25402 = ( n18509 & ~n20681 ) | ( n18509 & n25401 ) | ( ~n20681 & n25401 ) ;
  assign n25403 = n23418 ^ n9194 ^ n5479 ;
  assign n25406 = ( n3061 & n13226 ) | ( n3061 & ~n25294 ) | ( n13226 & ~n25294 ) ;
  assign n25404 = n17799 ^ n9819 ^ n4819 ;
  assign n25405 = ( n15259 & n15383 ) | ( n15259 & ~n25404 ) | ( n15383 & ~n25404 ) ;
  assign n25407 = n25406 ^ n25405 ^ n11648 ;
  assign n25408 = ( n18018 & n25403 ) | ( n18018 & ~n25407 ) | ( n25403 & ~n25407 ) ;
  assign n25409 = n14096 ^ n13493 ^ n12046 ;
  assign n25410 = ( n6417 & ~n6586 ) | ( n6417 & n25409 ) | ( ~n6586 & n25409 ) ;
  assign n25411 = n13786 ^ n11749 ^ n1873 ;
  assign n25412 = n8413 ^ n6949 ^ n3166 ;
  assign n25413 = ( n12806 & ~n16504 ) | ( n12806 & n25412 ) | ( ~n16504 & n25412 ) ;
  assign n25414 = ( x26 & n3460 ) | ( x26 & n16303 ) | ( n3460 & n16303 ) ;
  assign n25415 = n25414 ^ n7343 ^ n6869 ;
  assign n25416 = ( n21124 & n24354 ) | ( n21124 & n25415 ) | ( n24354 & n25415 ) ;
  assign n25417 = n25416 ^ n12491 ^ n4378 ;
  assign n25418 = n20183 ^ n19892 ^ n14139 ;
  assign n25419 = ( n5777 & ~n13745 ) | ( n5777 & n25418 ) | ( ~n13745 & n25418 ) ;
  assign n25420 = ( n2629 & ~n15914 ) | ( n2629 & n24671 ) | ( ~n15914 & n24671 ) ;
  assign n25421 = ( n556 & n6262 ) | ( n556 & n24797 ) | ( n6262 & n24797 ) ;
  assign n25422 = ( n6886 & n11574 ) | ( n6886 & n17022 ) | ( n11574 & n17022 ) ;
  assign n25423 = ( n4314 & n19492 ) | ( n4314 & n25422 ) | ( n19492 & n25422 ) ;
  assign n25424 = n15883 ^ n1344 ^ n395 ;
  assign n25425 = ( n5545 & n7596 ) | ( n5545 & ~n25424 ) | ( n7596 & ~n25424 ) ;
  assign n25426 = n5663 ^ n2934 ^ n898 ;
  assign n25427 = n25426 ^ n7282 ^ n4401 ;
  assign n25428 = ( ~n280 & n1108 ) | ( ~n280 & n19352 ) | ( n1108 & n19352 ) ;
  assign n25429 = n25428 ^ n22455 ^ n17430 ;
  assign n25430 = ( n9221 & n25427 ) | ( n9221 & n25429 ) | ( n25427 & n25429 ) ;
  assign n25431 = ( ~n288 & n4530 ) | ( ~n288 & n11110 ) | ( n4530 & n11110 ) ;
  assign n25432 = n24214 ^ n21119 ^ n333 ;
  assign n25433 = ( n3229 & n25431 ) | ( n3229 & ~n25432 ) | ( n25431 & ~n25432 ) ;
  assign n25434 = ( n488 & n571 ) | ( n488 & n25433 ) | ( n571 & n25433 ) ;
  assign n25436 = n7071 ^ n452 ^ n245 ;
  assign n25435 = ( n10687 & n14874 ) | ( n10687 & ~n15104 ) | ( n14874 & ~n15104 ) ;
  assign n25437 = n25436 ^ n25435 ^ n14841 ;
  assign n25438 = ( n2948 & n7918 ) | ( n2948 & ~n9125 ) | ( n7918 & ~n9125 ) ;
  assign n25439 = n25438 ^ n18475 ^ n15949 ;
  assign n25440 = ( n4984 & ~n19820 ) | ( n4984 & n20791 ) | ( ~n19820 & n20791 ) ;
  assign n25441 = ( n704 & ~n23641 ) | ( n704 & n25440 ) | ( ~n23641 & n25440 ) ;
  assign n25442 = n19702 ^ n19302 ^ n15660 ;
  assign n25443 = ( n791 & n11298 ) | ( n791 & n15360 ) | ( n11298 & n15360 ) ;
  assign n25444 = ( n16667 & n19455 ) | ( n16667 & ~n25443 ) | ( n19455 & ~n25443 ) ;
  assign n25445 = ( n12542 & n25442 ) | ( n12542 & n25444 ) | ( n25442 & n25444 ) ;
  assign n25446 = n23563 ^ n18930 ^ n11155 ;
  assign n25447 = ( n2368 & n7908 ) | ( n2368 & ~n25446 ) | ( n7908 & ~n25446 ) ;
  assign n25448 = n25447 ^ n21645 ^ n10128 ;
  assign n25449 = n20197 ^ n16975 ^ n1606 ;
  assign n25450 = n23651 ^ n14965 ^ n2226 ;
  assign n25451 = n25450 ^ n16770 ^ n5666 ;
  assign n25452 = ( n3038 & n3502 ) | ( n3038 & n5334 ) | ( n3502 & n5334 ) ;
  assign n25453 = ( ~n1607 & n8381 ) | ( ~n1607 & n23169 ) | ( n8381 & n23169 ) ;
  assign n25454 = ( n3449 & ~n9137 ) | ( n3449 & n25453 ) | ( ~n9137 & n25453 ) ;
  assign n25455 = n23129 ^ n4665 ^ n3353 ;
  assign n25456 = ( n13223 & ~n14034 ) | ( n13223 & n25455 ) | ( ~n14034 & n25455 ) ;
  assign n25457 = ( n1115 & n9512 ) | ( n1115 & n11049 ) | ( n9512 & n11049 ) ;
  assign n25458 = ( n16606 & n24289 ) | ( n16606 & ~n25457 ) | ( n24289 & ~n25457 ) ;
  assign n25461 = n13757 ^ n2499 ^ n1715 ;
  assign n25459 = ( n2278 & ~n5666 ) | ( n2278 & n14663 ) | ( ~n5666 & n14663 ) ;
  assign n25460 = ( n8327 & n13262 ) | ( n8327 & n25459 ) | ( n13262 & n25459 ) ;
  assign n25462 = n25461 ^ n25460 ^ n6154 ;
  assign n25463 = n19428 ^ n10173 ^ n6629 ;
  assign n25464 = n25463 ^ n24828 ^ n6565 ;
  assign n25465 = n14952 ^ n13259 ^ n7054 ;
  assign n25466 = n25465 ^ n13506 ^ n11743 ;
  assign n25467 = ( ~n1402 & n11156 ) | ( ~n1402 & n19075 ) | ( n11156 & n19075 ) ;
  assign n25468 = ( n3854 & n14273 ) | ( n3854 & n25467 ) | ( n14273 & n25467 ) ;
  assign n25469 = n25468 ^ n7774 ^ n3858 ;
  assign n25470 = n16100 ^ n9660 ^ n5424 ;
  assign n25471 = n25470 ^ n19343 ^ n5040 ;
  assign n25472 = n4264 ^ n4028 ^ n672 ;
  assign n25473 = n25472 ^ n12397 ^ n4398 ;
  assign n25474 = n25473 ^ n2845 ^ n1571 ;
  assign n25475 = n25474 ^ n20119 ^ n10734 ;
  assign n25476 = n25475 ^ n14312 ^ n10182 ;
  assign n25477 = n15019 ^ n9933 ^ n5615 ;
  assign n25478 = n24408 ^ n18285 ^ n10217 ;
  assign n25479 = n25478 ^ n5946 ^ n1341 ;
  assign n25480 = n23561 ^ n3726 ^ n2794 ;
  assign n25481 = n8542 ^ n7368 ^ n2022 ;
  assign n25482 = n24203 ^ n22043 ^ n18263 ;
  assign n25483 = n25482 ^ n10657 ^ n5061 ;
  assign n25484 = ( n10717 & n12422 ) | ( n10717 & n25483 ) | ( n12422 & n25483 ) ;
  assign n25485 = ( n5694 & n10217 ) | ( n5694 & ~n25484 ) | ( n10217 & ~n25484 ) ;
  assign n25486 = ( n2200 & n14542 ) | ( n2200 & ~n24380 ) | ( n14542 & ~n24380 ) ;
  assign n25487 = ( n8890 & ~n9174 ) | ( n8890 & n25486 ) | ( ~n9174 & n25486 ) ;
  assign n25488 = ( ~n3603 & n21941 ) | ( ~n3603 & n25487 ) | ( n21941 & n25487 ) ;
  assign n25489 = ( n8395 & n9347 ) | ( n8395 & n19075 ) | ( n9347 & n19075 ) ;
  assign n25490 = ( ~n7085 & n12219 ) | ( ~n7085 & n16936 ) | ( n12219 & n16936 ) ;
  assign n25491 = n25490 ^ n7554 ^ n2189 ;
  assign n25492 = ( n1429 & n2294 ) | ( n1429 & n15549 ) | ( n2294 & n15549 ) ;
  assign n25493 = n25492 ^ n13897 ^ n9277 ;
  assign n25494 = n19731 ^ n17148 ^ n5144 ;
  assign n25495 = n25494 ^ n21138 ^ n9602 ;
  assign n25496 = n25495 ^ n19374 ^ n4960 ;
  assign n25497 = n24140 ^ n13134 ^ n8069 ;
  assign n25498 = ( ~n7436 & n7991 ) | ( ~n7436 & n21787 ) | ( n7991 & n21787 ) ;
  assign n25499 = n19162 ^ n8717 ^ n3204 ;
  assign n25500 = ( ~n2006 & n9800 ) | ( ~n2006 & n25499 ) | ( n9800 & n25499 ) ;
  assign n25501 = ( ~n9876 & n25498 ) | ( ~n9876 & n25500 ) | ( n25498 & n25500 ) ;
  assign n25502 = ( ~n3831 & n15998 ) | ( ~n3831 & n21530 ) | ( n15998 & n21530 ) ;
  assign n25503 = n5763 ^ n2233 ^ n1432 ;
  assign n25504 = ( n2333 & n25502 ) | ( n2333 & ~n25503 ) | ( n25502 & ~n25503 ) ;
  assign n25505 = n25504 ^ n16139 ^ n11940 ;
  assign n25506 = n25505 ^ n8230 ^ n7030 ;
  assign n25509 = ( n11026 & n12678 ) | ( n11026 & n14255 ) | ( n12678 & n14255 ) ;
  assign n25507 = ( ~n1748 & n9555 ) | ( ~n1748 & n12831 ) | ( n9555 & n12831 ) ;
  assign n25508 = ( n3914 & n23584 ) | ( n3914 & n25507 ) | ( n23584 & n25507 ) ;
  assign n25510 = n25509 ^ n25508 ^ n20975 ;
  assign n25511 = ( n1169 & n2273 ) | ( n1169 & n9841 ) | ( n2273 & n9841 ) ;
  assign n25512 = n25511 ^ n22406 ^ n7875 ;
  assign n25513 = n18252 ^ n5850 ^ n1213 ;
  assign n25518 = ( n2375 & n5829 ) | ( n2375 & n22273 ) | ( n5829 & n22273 ) ;
  assign n25519 = n25518 ^ n16650 ^ n867 ;
  assign n25516 = n12924 ^ n10136 ^ n1978 ;
  assign n25514 = n16303 ^ n5312 ^ n4542 ;
  assign n25515 = ( ~n1947 & n4364 ) | ( ~n1947 & n25514 ) | ( n4364 & n25514 ) ;
  assign n25517 = n25516 ^ n25515 ^ n12379 ;
  assign n25520 = n25519 ^ n25517 ^ n11414 ;
  assign n25521 = ( n16787 & n25513 ) | ( n16787 & ~n25520 ) | ( n25513 & ~n25520 ) ;
  assign n25522 = n25368 ^ n14996 ^ n9402 ;
  assign n25523 = ( n6359 & n12936 ) | ( n6359 & n25522 ) | ( n12936 & n25522 ) ;
  assign n25524 = ( n3811 & n15844 ) | ( n3811 & n25523 ) | ( n15844 & n25523 ) ;
  assign n25525 = ( n776 & ~n6384 ) | ( n776 & n20160 ) | ( ~n6384 & n20160 ) ;
  assign n25526 = n25525 ^ n16075 ^ n13534 ;
  assign n25527 = ( n8501 & n10430 ) | ( n8501 & n22406 ) | ( n10430 & n22406 ) ;
  assign n25528 = n24784 ^ n21768 ^ n6791 ;
  assign n25529 = ( n9500 & ~n16492 ) | ( n9500 & n21763 ) | ( ~n16492 & n21763 ) ;
  assign n25530 = ( n11779 & n16979 ) | ( n11779 & n25529 ) | ( n16979 & n25529 ) ;
  assign n25531 = ( n686 & n7067 ) | ( n686 & n12242 ) | ( n7067 & n12242 ) ;
  assign n25532 = ( n4367 & n20376 ) | ( n4367 & n25531 ) | ( n20376 & n25531 ) ;
  assign n25533 = n17140 ^ n2615 ^ n1540 ;
  assign n25534 = ( ~n224 & n2331 ) | ( ~n224 & n15537 ) | ( n2331 & n15537 ) ;
  assign n25535 = n25534 ^ n23322 ^ n20964 ;
  assign n25536 = n15672 ^ n8398 ^ n194 ;
  assign n25537 = n25536 ^ n17573 ^ n3317 ;
  assign n25539 = n10311 ^ n3978 ^ n1916 ;
  assign n25538 = n20924 ^ n15606 ^ n6717 ;
  assign n25540 = n25539 ^ n25538 ^ n10664 ;
  assign n25541 = ( ~n2064 & n10294 ) | ( ~n2064 & n15989 ) | ( n10294 & n15989 ) ;
  assign n25542 = ( n11599 & n15946 ) | ( n11599 & ~n16581 ) | ( n15946 & ~n16581 ) ;
  assign n25543 = n25542 ^ n16128 ^ n14662 ;
  assign n25544 = n23595 ^ n19660 ^ n3941 ;
  assign n25545 = n24198 ^ n17637 ^ n6635 ;
  assign n25547 = ( ~n756 & n7500 ) | ( ~n756 & n15998 ) | ( n7500 & n15998 ) ;
  assign n25546 = ( n5950 & n15094 ) | ( n5950 & n19613 ) | ( n15094 & n19613 ) ;
  assign n25548 = n25547 ^ n25546 ^ n22237 ;
  assign n25549 = ( ~n11334 & n21123 ) | ( ~n11334 & n22782 ) | ( n21123 & n22782 ) ;
  assign n25550 = n25549 ^ n21033 ^ n1843 ;
  assign n25551 = ( ~n7455 & n20543 ) | ( ~n7455 & n25550 ) | ( n20543 & n25550 ) ;
  assign n25552 = n14604 ^ n13422 ^ n194 ;
  assign n25553 = n25552 ^ n20163 ^ n7640 ;
  assign n25554 = n25553 ^ n13863 ^ n8044 ;
  assign n25555 = n25554 ^ n5737 ^ n489 ;
  assign n25556 = ( n6069 & ~n13338 ) | ( n6069 & n24987 ) | ( ~n13338 & n24987 ) ;
  assign n25557 = n20146 ^ n7445 ^ n1469 ;
  assign n25561 = ( n665 & n2067 ) | ( n665 & n16266 ) | ( n2067 & n16266 ) ;
  assign n25558 = n10038 ^ n1617 ^ n610 ;
  assign n25559 = n25558 ^ n6854 ^ n1017 ;
  assign n25560 = ( ~n18988 & n21146 ) | ( ~n18988 & n25559 ) | ( n21146 & n25559 ) ;
  assign n25562 = n25561 ^ n25560 ^ n14119 ;
  assign n25563 = ( n2188 & ~n9522 ) | ( n2188 & n14243 ) | ( ~n9522 & n14243 ) ;
  assign n25564 = ( n7607 & n16823 ) | ( n7607 & n25563 ) | ( n16823 & n25563 ) ;
  assign n25565 = n25564 ^ n19305 ^ n9038 ;
  assign n25568 = ( n3951 & n4756 ) | ( n3951 & n13996 ) | ( n4756 & n13996 ) ;
  assign n25569 = ( n158 & n23611 ) | ( n158 & n25568 ) | ( n23611 & n25568 ) ;
  assign n25570 = n25569 ^ n7001 ^ n5208 ;
  assign n25566 = ( n6507 & ~n9201 ) | ( n6507 & n23167 ) | ( ~n9201 & n23167 ) ;
  assign n25567 = n25566 ^ n19129 ^ n3776 ;
  assign n25571 = n25570 ^ n25567 ^ n5396 ;
  assign n25572 = n11967 ^ n6368 ^ n192 ;
  assign n25573 = n17425 ^ n14290 ^ n10781 ;
  assign n25574 = ( ~n16143 & n25572 ) | ( ~n16143 & n25573 ) | ( n25572 & n25573 ) ;
  assign n25575 = ( ~n13306 & n20903 ) | ( ~n13306 & n25574 ) | ( n20903 & n25574 ) ;
  assign n25576 = ( ~n10377 & n22168 ) | ( ~n10377 & n24921 ) | ( n22168 & n24921 ) ;
  assign n25577 = ( n4584 & n6548 ) | ( n4584 & n25576 ) | ( n6548 & n25576 ) ;
  assign n25578 = n25577 ^ n14815 ^ n9124 ;
  assign n25579 = n25578 ^ n8968 ^ n2642 ;
  assign n25580 = n19848 ^ n19018 ^ n184 ;
  assign n25581 = ( n3064 & n12406 ) | ( n3064 & n13567 ) | ( n12406 & n13567 ) ;
  assign n25582 = ( ~n8432 & n25580 ) | ( ~n8432 & n25581 ) | ( n25580 & n25581 ) ;
  assign n25583 = ( n6169 & n13120 ) | ( n6169 & ~n25582 ) | ( n13120 & ~n25582 ) ;
  assign n25584 = ( n1277 & ~n7936 ) | ( n1277 & n14750 ) | ( ~n7936 & n14750 ) ;
  assign n25585 = ( n5713 & ~n6208 ) | ( n5713 & n25584 ) | ( ~n6208 & n25584 ) ;
  assign n25586 = n25585 ^ n2650 ^ n2497 ;
  assign n25587 = ( n9967 & n19640 ) | ( n9967 & n25586 ) | ( n19640 & n25586 ) ;
  assign n25588 = ( x58 & n8336 ) | ( x58 & ~n18366 ) | ( n8336 & ~n18366 ) ;
  assign n25591 = n22123 ^ n11485 ^ n8152 ;
  assign n25592 = ( n1270 & n10972 ) | ( n1270 & ~n25591 ) | ( n10972 & ~n25591 ) ;
  assign n25589 = n25552 ^ n20586 ^ n16828 ;
  assign n25590 = n25589 ^ n24030 ^ n3785 ;
  assign n25593 = n25592 ^ n25590 ^ n24425 ;
  assign n25594 = ( n5682 & n25588 ) | ( n5682 & ~n25593 ) | ( n25588 & ~n25593 ) ;
  assign n25595 = ( ~n607 & n722 ) | ( ~n607 & n6899 ) | ( n722 & n6899 ) ;
  assign n25596 = ( n3974 & n21210 ) | ( n3974 & ~n21651 ) | ( n21210 & ~n21651 ) ;
  assign n25597 = ( ~n13483 & n25595 ) | ( ~n13483 & n25596 ) | ( n25595 & n25596 ) ;
  assign n25598 = n25597 ^ n25472 ^ n19797 ;
  assign n25599 = ( n825 & ~n1535 ) | ( n825 & n2589 ) | ( ~n1535 & n2589 ) ;
  assign n25600 = ( n2943 & n21446 ) | ( n2943 & n25599 ) | ( n21446 & n25599 ) ;
  assign n25601 = ( n2978 & n6927 ) | ( n2978 & n20311 ) | ( n6927 & n20311 ) ;
  assign n25602 = n25601 ^ n19545 ^ n4195 ;
  assign n25603 = ( n2673 & n3045 ) | ( n2673 & n25602 ) | ( n3045 & n25602 ) ;
  assign n25604 = ( ~n704 & n7074 ) | ( ~n704 & n10792 ) | ( n7074 & n10792 ) ;
  assign n25605 = ( n4721 & n10018 ) | ( n4721 & ~n10562 ) | ( n10018 & ~n10562 ) ;
  assign n25606 = ( n4204 & ~n25604 ) | ( n4204 & n25605 ) | ( ~n25604 & n25605 ) ;
  assign n25607 = ( n12428 & n15139 ) | ( n12428 & ~n15437 ) | ( n15139 & ~n15437 ) ;
  assign n25608 = n9237 ^ n1854 ^ n420 ;
  assign n25609 = ( n1171 & ~n15541 ) | ( n1171 & n25608 ) | ( ~n15541 & n25608 ) ;
  assign n25610 = ( n4202 & n8522 ) | ( n4202 & ~n25609 ) | ( n8522 & ~n25609 ) ;
  assign n25611 = ( n4171 & n5853 ) | ( n4171 & n7922 ) | ( n5853 & n7922 ) ;
  assign n25612 = ( n1105 & n10157 ) | ( n1105 & ~n25611 ) | ( n10157 & ~n25611 ) ;
  assign n25613 = n25612 ^ n20818 ^ n3987 ;
  assign n25614 = n24073 ^ n1171 ^ n858 ;
  assign n25615 = ( n6831 & n9003 ) | ( n6831 & ~n25614 ) | ( n9003 & ~n25614 ) ;
  assign n25616 = ( n9827 & n12025 ) | ( n9827 & n14094 ) | ( n12025 & n14094 ) ;
  assign n25617 = ( ~n9909 & n19886 ) | ( ~n9909 & n25616 ) | ( n19886 & n25616 ) ;
  assign n25618 = ( n19907 & n23079 ) | ( n19907 & ~n25617 ) | ( n23079 & ~n25617 ) ;
  assign n25619 = ( n7729 & n8147 ) | ( n7729 & n15456 ) | ( n8147 & n15456 ) ;
  assign n25620 = ( n5511 & ~n8393 ) | ( n5511 & n25619 ) | ( ~n8393 & n25619 ) ;
  assign n25621 = ( n7318 & n17778 ) | ( n7318 & n25389 ) | ( n17778 & n25389 ) ;
  assign n25622 = ( ~n8192 & n24666 ) | ( ~n8192 & n25621 ) | ( n24666 & n25621 ) ;
  assign n25623 = n25622 ^ n12360 ^ n9213 ;
  assign n25624 = ( n3805 & n9120 ) | ( n3805 & n18340 ) | ( n9120 & n18340 ) ;
  assign n25625 = ( ~n1914 & n21914 ) | ( ~n1914 & n25624 ) | ( n21914 & n25624 ) ;
  assign n25626 = ( n7248 & ~n25623 ) | ( n7248 & n25625 ) | ( ~n25623 & n25625 ) ;
  assign n25627 = ( n10636 & n18192 ) | ( n10636 & ~n25241 ) | ( n18192 & ~n25241 ) ;
  assign n25628 = ( n5165 & n10314 ) | ( n5165 & n22266 ) | ( n10314 & n22266 ) ;
  assign n25629 = n25628 ^ n22615 ^ n2366 ;
  assign n25633 = n9112 ^ n2597 ^ n2282 ;
  assign n25632 = n18474 ^ n9091 ^ n1992 ;
  assign n25634 = n25633 ^ n25632 ^ n13025 ;
  assign n25630 = n10327 ^ n4549 ^ n4514 ;
  assign n25631 = n25630 ^ n18621 ^ n5170 ;
  assign n25635 = n25634 ^ n25631 ^ n801 ;
  assign n25636 = ( n15379 & n16692 ) | ( n15379 & n22827 ) | ( n16692 & n22827 ) ;
  assign n25637 = ( n13715 & ~n14523 ) | ( n13715 & n25636 ) | ( ~n14523 & n25636 ) ;
  assign n25638 = ( ~n6229 & n6244 ) | ( ~n6229 & n25637 ) | ( n6244 & n25637 ) ;
  assign n25641 = ( n4756 & n7636 ) | ( n4756 & ~n7699 ) | ( n7636 & ~n7699 ) ;
  assign n25639 = ( ~n1692 & n2461 ) | ( ~n1692 & n2624 ) | ( n2461 & n2624 ) ;
  assign n25640 = ( n1520 & n2320 ) | ( n1520 & n25639 ) | ( n2320 & n25639 ) ;
  assign n25642 = n25641 ^ n25640 ^ n14990 ;
  assign n25643 = n25642 ^ n7952 ^ n6416 ;
  assign n25644 = ( n3141 & n3181 ) | ( n3141 & ~n9931 ) | ( n3181 & ~n9931 ) ;
  assign n25646 = ( n8502 & n9137 ) | ( n8502 & n25473 ) | ( n9137 & n25473 ) ;
  assign n25645 = n14897 ^ n10913 ^ n5609 ;
  assign n25647 = n25646 ^ n25645 ^ n17136 ;
  assign n25648 = n25647 ^ n3477 ^ n853 ;
  assign n25649 = n12404 ^ n4782 ^ x72 ;
  assign n25650 = ( n11366 & n15558 ) | ( n11366 & n25649 ) | ( n15558 & n25649 ) ;
  assign n25651 = n14113 ^ n11530 ^ n5181 ;
  assign n25658 = ( n4416 & n10212 ) | ( n4416 & n20241 ) | ( n10212 & n20241 ) ;
  assign n25656 = ( x4 & n8641 ) | ( x4 & ~n18112 ) | ( n8641 & ~n18112 ) ;
  assign n25654 = ( n9322 & ~n15066 ) | ( n9322 & n22879 ) | ( ~n15066 & n22879 ) ;
  assign n25655 = ( n2805 & n5584 ) | ( n2805 & n25654 ) | ( n5584 & n25654 ) ;
  assign n25652 = n13185 ^ n4841 ^ n1026 ;
  assign n25653 = ( n16740 & n25220 ) | ( n16740 & ~n25652 ) | ( n25220 & ~n25652 ) ;
  assign n25657 = n25656 ^ n25655 ^ n25653 ;
  assign n25659 = n25658 ^ n25657 ^ n11344 ;
  assign n25660 = ( ~n9471 & n10108 ) | ( ~n9471 & n12754 ) | ( n10108 & n12754 ) ;
  assign n25661 = n13498 ^ n7495 ^ n7187 ;
  assign n25662 = n25661 ^ n19682 ^ n13904 ;
  assign n25663 = ( n4831 & ~n23621 ) | ( n4831 & n25662 ) | ( ~n23621 & n25662 ) ;
  assign n25664 = ( n5572 & n9370 ) | ( n5572 & n10176 ) | ( n9370 & n10176 ) ;
  assign n25665 = ( n8639 & n20901 ) | ( n8639 & ~n25664 ) | ( n20901 & ~n25664 ) ;
  assign n25666 = ( n6506 & ~n17756 ) | ( n6506 & n25665 ) | ( ~n17756 & n25665 ) ;
  assign n25667 = ( n1796 & n8486 ) | ( n1796 & n12971 ) | ( n8486 & n12971 ) ;
  assign n25668 = n25667 ^ n17473 ^ n5928 ;
  assign n25669 = n15933 ^ n9675 ^ n7380 ;
  assign n25670 = n25669 ^ n16482 ^ n15760 ;
  assign n25671 = ( n2378 & n6173 ) | ( n2378 & n14081 ) | ( n6173 & n14081 ) ;
  assign n25672 = n25671 ^ n5721 ^ n1957 ;
  assign n25673 = n23891 ^ n6033 ^ n5371 ;
  assign n25674 = n16923 ^ n16884 ^ n10891 ;
  assign n25675 = ( n450 & ~n2081 ) | ( n450 & n25674 ) | ( ~n2081 & n25674 ) ;
  assign n25676 = ( n7471 & n15930 ) | ( n7471 & n18229 ) | ( n15930 & n18229 ) ;
  assign n25677 = ( n2144 & ~n8680 ) | ( n2144 & n16718 ) | ( ~n8680 & n16718 ) ;
  assign n25678 = ( n164 & ~n2039 ) | ( n164 & n14297 ) | ( ~n2039 & n14297 ) ;
  assign n25679 = ( ~n5722 & n15067 ) | ( ~n5722 & n19725 ) | ( n15067 & n19725 ) ;
  assign n25680 = ( n2153 & n3163 ) | ( n2153 & n14042 ) | ( n3163 & n14042 ) ;
  assign n25681 = ( n7603 & ~n9281 ) | ( n7603 & n25680 ) | ( ~n9281 & n25680 ) ;
  assign n25682 = n7136 ^ n366 ^ n199 ;
  assign n25683 = ( n12115 & n17005 ) | ( n12115 & n25682 ) | ( n17005 & n25682 ) ;
  assign n25684 = n25683 ^ n23010 ^ n5978 ;
  assign n25685 = ( n5194 & n12721 ) | ( n5194 & ~n20448 ) | ( n12721 & ~n20448 ) ;
  assign n25686 = ( n9594 & n17724 ) | ( n9594 & n25685 ) | ( n17724 & n25685 ) ;
  assign n25687 = ( ~n6232 & n19574 ) | ( ~n6232 & n25686 ) | ( n19574 & n25686 ) ;
  assign n25688 = ( n19123 & ~n19651 ) | ( n19123 & n24171 ) | ( ~n19651 & n24171 ) ;
  assign n25689 = n7422 ^ n3083 ^ n1039 ;
  assign n25690 = n25689 ^ n13356 ^ n12846 ;
  assign n25691 = ( n20152 & n22225 ) | ( n20152 & ~n25690 ) | ( n22225 & ~n25690 ) ;
  assign n25692 = n19225 ^ n8513 ^ n485 ;
  assign n25693 = n25692 ^ n15930 ^ n6469 ;
  assign n25694 = ( n9193 & ~n9840 ) | ( n9193 & n25693 ) | ( ~n9840 & n25693 ) ;
  assign n25695 = ( x40 & ~n271 ) | ( x40 & n6521 ) | ( ~n271 & n6521 ) ;
  assign n25696 = ( n2691 & n9353 ) | ( n2691 & ~n25695 ) | ( n9353 & ~n25695 ) ;
  assign n25697 = n25696 ^ n21891 ^ n15483 ;
  assign n25706 = ( n4992 & ~n9538 ) | ( n4992 & n11364 ) | ( ~n9538 & n11364 ) ;
  assign n25704 = ( n4527 & ~n20357 ) | ( n4527 & n20454 ) | ( ~n20357 & n20454 ) ;
  assign n25705 = ( n5180 & n18047 ) | ( n5180 & ~n25704 ) | ( n18047 & ~n25704 ) ;
  assign n25698 = ( n2447 & n14446 ) | ( n2447 & ~n22782 ) | ( n14446 & ~n22782 ) ;
  assign n25699 = n16613 ^ n5439 ^ n4604 ;
  assign n25700 = n19886 ^ n17956 ^ n2201 ;
  assign n25701 = ( n5180 & n25699 ) | ( n5180 & ~n25700 ) | ( n25699 & ~n25700 ) ;
  assign n25702 = ( n4055 & n25698 ) | ( n4055 & ~n25701 ) | ( n25698 & ~n25701 ) ;
  assign n25703 = ( n10895 & n13336 ) | ( n10895 & n25702 ) | ( n13336 & n25702 ) ;
  assign n25707 = n25706 ^ n25705 ^ n25703 ;
  assign n25708 = ( n4576 & n6906 ) | ( n4576 & n9168 ) | ( n6906 & n9168 ) ;
  assign n25709 = n11926 ^ n8630 ^ n537 ;
  assign n25711 = n10837 ^ n7247 ^ n667 ;
  assign n25710 = n11077 ^ n9436 ^ n5816 ;
  assign n25712 = n25711 ^ n25710 ^ n23266 ;
  assign n25713 = ( n18710 & n25709 ) | ( n18710 & n25712 ) | ( n25709 & n25712 ) ;
  assign n25714 = ( n1614 & ~n7803 ) | ( n1614 & n11969 ) | ( ~n7803 & n11969 ) ;
  assign n25715 = ( n4095 & n8800 ) | ( n4095 & ~n25714 ) | ( n8800 & ~n25714 ) ;
  assign n25717 = n11648 ^ n9797 ^ n3218 ;
  assign n25718 = ( n10319 & n15991 ) | ( n10319 & n25717 ) | ( n15991 & n25717 ) ;
  assign n25716 = n25498 ^ n7877 ^ n6945 ;
  assign n25719 = n25718 ^ n25716 ^ n20893 ;
  assign n25720 = ( n2857 & ~n5533 ) | ( n2857 & n17775 ) | ( ~n5533 & n17775 ) ;
  assign n25721 = ( n1245 & n12835 ) | ( n1245 & n25720 ) | ( n12835 & n25720 ) ;
  assign n25722 = ( n6837 & ~n12400 ) | ( n6837 & n16635 ) | ( ~n12400 & n16635 ) ;
  assign n25723 = ( n4311 & n13449 ) | ( n4311 & n17789 ) | ( n13449 & n17789 ) ;
  assign n25724 = n25426 ^ n19821 ^ n12973 ;
  assign n25725 = ( n5794 & n8543 ) | ( n5794 & ~n20165 ) | ( n8543 & ~n20165 ) ;
  assign n25726 = ( n1263 & ~n25724 ) | ( n1263 & n25725 ) | ( ~n25724 & n25725 ) ;
  assign n25727 = n25726 ^ n15075 ^ n13198 ;
  assign n25728 = n25727 ^ n18602 ^ n15383 ;
  assign n25729 = n22722 ^ n17345 ^ n13145 ;
  assign n25730 = n25729 ^ n15412 ^ n10426 ;
  assign n25731 = ( n977 & n9146 ) | ( n977 & n13534 ) | ( n9146 & n13534 ) ;
  assign n25732 = ( ~n3357 & n8587 ) | ( ~n3357 & n12321 ) | ( n8587 & n12321 ) ;
  assign n25733 = ( ~n3624 & n5217 ) | ( ~n3624 & n10068 ) | ( n5217 & n10068 ) ;
  assign n25734 = n25733 ^ n24708 ^ n9319 ;
  assign n25735 = n4474 ^ n2130 ^ n931 ;
  assign n25737 = ( n953 & ~n3579 ) | ( n953 & n16975 ) | ( ~n3579 & n16975 ) ;
  assign n25738 = n25737 ^ n9184 ^ n5038 ;
  assign n25736 = ( n191 & n2391 ) | ( n191 & ~n17838 ) | ( n2391 & ~n17838 ) ;
  assign n25739 = n25738 ^ n25736 ^ n3296 ;
  assign n25740 = n21668 ^ n18123 ^ n12708 ;
  assign n25741 = ( n858 & n4867 ) | ( n858 & ~n19386 ) | ( n4867 & ~n19386 ) ;
  assign n25742 = ( n12837 & n24996 ) | ( n12837 & ~n25741 ) | ( n24996 & ~n25741 ) ;
  assign n25743 = n22541 ^ n22117 ^ n17672 ;
  assign n25744 = ( n3358 & n3822 ) | ( n3358 & ~n6081 ) | ( n3822 & ~n6081 ) ;
  assign n25745 = ( n1759 & ~n3368 ) | ( n1759 & n20207 ) | ( ~n3368 & n20207 ) ;
  assign n25746 = ( n3276 & ~n4592 ) | ( n3276 & n8042 ) | ( ~n4592 & n8042 ) ;
  assign n25747 = ( n8829 & ~n19634 ) | ( n8829 & n25746 ) | ( ~n19634 & n25746 ) ;
  assign n25748 = ( n1338 & ~n17578 ) | ( n1338 & n25747 ) | ( ~n17578 & n25747 ) ;
  assign n25749 = n25748 ^ n10054 ^ n928 ;
  assign n25750 = n21661 ^ n17323 ^ n4093 ;
  assign n25751 = ( ~n5975 & n6870 ) | ( ~n5975 & n7230 ) | ( n6870 & n7230 ) ;
  assign n25752 = ( n1462 & n8708 ) | ( n1462 & ~n25751 ) | ( n8708 & ~n25751 ) ;
  assign n25753 = ( n7070 & ~n25750 ) | ( n7070 & n25752 ) | ( ~n25750 & n25752 ) ;
  assign n25754 = n19735 ^ n13525 ^ n7839 ;
  assign n25755 = n25754 ^ n8135 ^ n2450 ;
  assign n25756 = ( ~n4360 & n17399 ) | ( ~n4360 & n25755 ) | ( n17399 & n25755 ) ;
  assign n25757 = n14273 ^ n14151 ^ n10734 ;
  assign n25758 = n20006 ^ n6221 ^ n2466 ;
  assign n25759 = ( n469 & ~n19613 ) | ( n469 & n25758 ) | ( ~n19613 & n25758 ) ;
  assign n25760 = ( n2941 & n5486 ) | ( n2941 & ~n7065 ) | ( n5486 & ~n7065 ) ;
  assign n25761 = n24931 ^ n1099 ^ n716 ;
  assign n25762 = ( n18269 & ~n19706 ) | ( n18269 & n25761 ) | ( ~n19706 & n25761 ) ;
  assign n25763 = n25194 ^ n18798 ^ n13106 ;
  assign n25764 = ( n3582 & ~n13951 ) | ( n3582 & n25763 ) | ( ~n13951 & n25763 ) ;
  assign n25765 = n14917 ^ n14327 ^ n9255 ;
  assign n25766 = n25765 ^ n15134 ^ n2826 ;
  assign n25767 = n16135 ^ n12261 ^ n181 ;
  assign n25768 = ( n8879 & ~n10946 ) | ( n8879 & n25767 ) | ( ~n10946 & n25767 ) ;
  assign n25769 = n25768 ^ n24875 ^ n10057 ;
  assign n25770 = n25769 ^ n6472 ^ n1101 ;
  assign n25772 = n19545 ^ n5661 ^ n5573 ;
  assign n25771 = n6034 ^ n4846 ^ n280 ;
  assign n25773 = n25772 ^ n25771 ^ n3686 ;
  assign n25774 = ( n23241 & ~n25727 ) | ( n23241 & n25773 ) | ( ~n25727 & n25773 ) ;
  assign n25775 = n23950 ^ n7281 ^ n2548 ;
  assign n25776 = ( n11953 & ~n12376 ) | ( n11953 & n13031 ) | ( ~n12376 & n13031 ) ;
  assign n25778 = n19161 ^ n17439 ^ n3717 ;
  assign n25777 = n11719 ^ n7701 ^ n3640 ;
  assign n25779 = n25778 ^ n25777 ^ n11201 ;
  assign n25780 = ( n5793 & ~n10152 ) | ( n5793 & n17474 ) | ( ~n10152 & n17474 ) ;
  assign n25781 = ( n1692 & n21258 ) | ( n1692 & n25780 ) | ( n21258 & n25780 ) ;
  assign n25782 = ( n4901 & ~n19133 ) | ( n4901 & n25781 ) | ( ~n19133 & n25781 ) ;
  assign n25783 = n25465 ^ n21956 ^ n12626 ;
  assign n25784 = n25783 ^ n6529 ^ n3565 ;
  assign n25785 = n8955 ^ n7811 ^ x11 ;
  assign n25786 = n25785 ^ n15708 ^ n8668 ;
  assign n25787 = ( n6400 & n6780 ) | ( n6400 & ~n11638 ) | ( n6780 & ~n11638 ) ;
  assign n25788 = ( n973 & ~n12211 ) | ( n973 & n25787 ) | ( ~n12211 & n25787 ) ;
  assign n25789 = n25788 ^ n22583 ^ n3660 ;
  assign n25790 = ( n14864 & n25786 ) | ( n14864 & n25789 ) | ( n25786 & n25789 ) ;
  assign n25791 = ( ~n12052 & n25784 ) | ( ~n12052 & n25790 ) | ( n25784 & n25790 ) ;
  assign n25792 = ( n2863 & n17474 ) | ( n2863 & ~n25714 ) | ( n17474 & ~n25714 ) ;
  assign n25793 = n20063 ^ n8780 ^ n660 ;
  assign n25794 = n10022 ^ n6890 ^ n5682 ;
  assign n25795 = ( n4299 & n6785 ) | ( n4299 & n10347 ) | ( n6785 & n10347 ) ;
  assign n25796 = ( n19452 & n25794 ) | ( n19452 & n25795 ) | ( n25794 & n25795 ) ;
  assign n25797 = ( ~n12156 & n16757 ) | ( ~n12156 & n17014 ) | ( n16757 & n17014 ) ;
  assign n25798 = ( n6997 & n22819 ) | ( n6997 & ~n25797 ) | ( n22819 & ~n25797 ) ;
  assign n25799 = n12040 ^ n8970 ^ n7542 ;
  assign n25800 = n23901 ^ n16225 ^ n343 ;
  assign n25801 = ( n19445 & ~n25799 ) | ( n19445 & n25800 ) | ( ~n25799 & n25800 ) ;
  assign n25802 = n12103 ^ n5632 ^ n1514 ;
  assign n25803 = ( n1529 & n4873 ) | ( n1529 & ~n17371 ) | ( n4873 & ~n17371 ) ;
  assign n25804 = n6772 ^ n4658 ^ n3798 ;
  assign n25805 = ( n7263 & ~n10233 ) | ( n7263 & n25804 ) | ( ~n10233 & n25804 ) ;
  assign n25806 = ( n16803 & ~n25803 ) | ( n16803 & n25805 ) | ( ~n25803 & n25805 ) ;
  assign n25807 = ( n6160 & n15802 ) | ( n6160 & n19280 ) | ( n15802 & n19280 ) ;
  assign n25808 = ( ~n7256 & n8705 ) | ( ~n7256 & n25807 ) | ( n8705 & n25807 ) ;
  assign n25809 = n14075 ^ n4531 ^ n2627 ;
  assign n25810 = n25809 ^ n22249 ^ n2926 ;
  assign n25811 = n11969 ^ n9185 ^ n4306 ;
  assign n25812 = ( ~n788 & n7595 ) | ( ~n788 & n15117 ) | ( n7595 & n15117 ) ;
  assign n25813 = ( ~n2074 & n25811 ) | ( ~n2074 & n25812 ) | ( n25811 & n25812 ) ;
  assign n25814 = n25813 ^ n4524 ^ n1458 ;
  assign n25815 = n18483 ^ n16661 ^ n3524 ;
  assign n25816 = ( ~n2104 & n2998 ) | ( ~n2104 & n25815 ) | ( n2998 & n25815 ) ;
  assign n25817 = ( ~n605 & n4224 ) | ( ~n605 & n10461 ) | ( n4224 & n10461 ) ;
  assign n25818 = n25817 ^ n19827 ^ n19360 ;
  assign n25819 = n12904 ^ n5439 ^ n392 ;
  assign n25820 = ( n337 & ~n2208 ) | ( n337 & n25819 ) | ( ~n2208 & n25819 ) ;
  assign n25821 = ( n14638 & n17429 ) | ( n14638 & ~n25820 ) | ( n17429 & ~n25820 ) ;
  assign n25822 = ( n5265 & n15501 ) | ( n5265 & n25821 ) | ( n15501 & n25821 ) ;
  assign n25823 = n11365 ^ n7153 ^ n3272 ;
  assign n25824 = n17408 ^ n11400 ^ n6795 ;
  assign n25825 = ( ~n8729 & n8852 ) | ( ~n8729 & n25824 ) | ( n8852 & n25824 ) ;
  assign n25826 = n12473 ^ n4264 ^ n1462 ;
  assign n25827 = ( n5441 & n18208 ) | ( n5441 & n25826 ) | ( n18208 & n25826 ) ;
  assign n25828 = n25827 ^ n14837 ^ n6649 ;
  assign n25829 = n2491 ^ n1809 ^ n618 ;
  assign n25830 = n25829 ^ n17620 ^ n10190 ;
  assign n25831 = ( n5102 & ~n19450 ) | ( n5102 & n25830 ) | ( ~n19450 & n25830 ) ;
  assign n25832 = ( n2250 & n9339 ) | ( n2250 & n20096 ) | ( n9339 & n20096 ) ;
  assign n25833 = ( n594 & ~n20591 ) | ( n594 & n22615 ) | ( ~n20591 & n22615 ) ;
  assign n25834 = n17148 ^ n1422 ^ x111 ;
  assign n25835 = ( ~n2491 & n11252 ) | ( ~n2491 & n25834 ) | ( n11252 & n25834 ) ;
  assign n25838 = n8593 ^ n7092 ^ n6505 ;
  assign n25839 = ( n7788 & n10300 ) | ( n7788 & n25838 ) | ( n10300 & n25838 ) ;
  assign n25840 = n25839 ^ n19587 ^ n9502 ;
  assign n25836 = ( n12147 & n12326 ) | ( n12147 & ~n16311 ) | ( n12326 & ~n16311 ) ;
  assign n25837 = ( n2585 & ~n19245 ) | ( n2585 & n25836 ) | ( ~n19245 & n25836 ) ;
  assign n25841 = n25840 ^ n25837 ^ n15115 ;
  assign n25842 = ( n3484 & n5784 ) | ( n3484 & n17584 ) | ( n5784 & n17584 ) ;
  assign n25843 = n25842 ^ n4753 ^ n3731 ;
  assign n25844 = ( n18770 & ~n24420 ) | ( n18770 & n25843 ) | ( ~n24420 & n25843 ) ;
  assign n25846 = ( n13094 & ~n13107 ) | ( n13094 & n13961 ) | ( ~n13107 & n13961 ) ;
  assign n25845 = ( n14858 & n22540 ) | ( n14858 & n23155 ) | ( n22540 & n23155 ) ;
  assign n25847 = n25846 ^ n25845 ^ n5034 ;
  assign n25848 = ( ~n6705 & n23912 ) | ( ~n6705 & n25692 ) | ( n23912 & n25692 ) ;
  assign n25849 = ( ~n1655 & n17371 ) | ( ~n1655 & n25848 ) | ( n17371 & n25848 ) ;
  assign n25850 = ( n15719 & n24853 ) | ( n15719 & ~n25849 ) | ( n24853 & ~n25849 ) ;
  assign n25851 = n17395 ^ n9400 ^ n7846 ;
  assign n25852 = n25851 ^ n17022 ^ n10396 ;
  assign n25853 = n25852 ^ n14981 ^ n6623 ;
  assign n25854 = n25853 ^ n9200 ^ x32 ;
  assign n25856 = ( n7175 & n14354 ) | ( n7175 & n23703 ) | ( n14354 & n23703 ) ;
  assign n25855 = n16163 ^ n15554 ^ n174 ;
  assign n25857 = n25856 ^ n25855 ^ n10745 ;
  assign n25858 = n25857 ^ n18621 ^ n17208 ;
  assign n25859 = ( n8943 & n21331 ) | ( n8943 & ~n25858 ) | ( n21331 & ~n25858 ) ;
  assign n25860 = ( n1833 & n2604 ) | ( n1833 & n17001 ) | ( n2604 & n17001 ) ;
  assign n25861 = ( n847 & n10108 ) | ( n847 & n25860 ) | ( n10108 & n25860 ) ;
  assign n25862 = ( ~n4866 & n17859 ) | ( ~n4866 & n19562 ) | ( n17859 & n19562 ) ;
  assign n25863 = ( ~n5880 & n11047 ) | ( ~n5880 & n25862 ) | ( n11047 & n25862 ) ;
  assign n25864 = n6316 ^ n4123 ^ n281 ;
  assign n25865 = ( n3047 & n9441 ) | ( n3047 & ~n25864 ) | ( n9441 & ~n25864 ) ;
  assign n25866 = ( n14163 & n17732 ) | ( n14163 & ~n24412 ) | ( n17732 & ~n24412 ) ;
  assign n25867 = n25866 ^ n21718 ^ n2973 ;
  assign n25868 = ( ~n7978 & n25865 ) | ( ~n7978 & n25867 ) | ( n25865 & n25867 ) ;
  assign n25869 = ( n15928 & ~n20962 ) | ( n15928 & n21026 ) | ( ~n20962 & n21026 ) ;
  assign n25870 = n3375 ^ n512 ^ n507 ;
  assign n25871 = n25870 ^ n23015 ^ n6595 ;
  assign n25872 = n25871 ^ n8919 ^ n5457 ;
  assign n25873 = ( n8487 & ~n9811 ) | ( n8487 & n15134 ) | ( ~n9811 & n15134 ) ;
  assign n25874 = ( n2530 & n11717 ) | ( n2530 & ~n18699 ) | ( n11717 & ~n18699 ) ;
  assign n25875 = ( n15854 & ~n16588 ) | ( n15854 & n18931 ) | ( ~n16588 & n18931 ) ;
  assign n25876 = ( ~n4025 & n7654 ) | ( ~n4025 & n25875 ) | ( n7654 & n25875 ) ;
  assign n25877 = n25876 ^ n9489 ^ n2753 ;
  assign n25878 = ( n4063 & n8452 ) | ( n4063 & n17822 ) | ( n8452 & n17822 ) ;
  assign n25879 = n25878 ^ n22199 ^ n15183 ;
  assign n25880 = ( n170 & n2092 ) | ( n170 & ~n25879 ) | ( n2092 & ~n25879 ) ;
  assign n25881 = n13340 ^ n12447 ^ n1906 ;
  assign n25882 = n25881 ^ n17206 ^ n13508 ;
  assign n25883 = ( n11026 & n11770 ) | ( n11026 & ~n24241 ) | ( n11770 & ~n24241 ) ;
  assign n25884 = n25883 ^ n20965 ^ n16226 ;
  assign n25885 = ( n12829 & n15046 ) | ( n12829 & n25884 ) | ( n15046 & n25884 ) ;
  assign n25886 = n15908 ^ n11655 ^ n5410 ;
  assign n25887 = n25886 ^ n10696 ^ n4343 ;
  assign n25888 = ( n9816 & n20172 ) | ( n9816 & n25238 ) | ( n20172 & n25238 ) ;
  assign n25889 = n25888 ^ n1861 ^ n1096 ;
  assign n25890 = n25889 ^ n2173 ^ n2037 ;
  assign n25891 = ( n12863 & n16127 ) | ( n12863 & ~n23878 ) | ( n16127 & ~n23878 ) ;
  assign n25892 = ( n263 & n3499 ) | ( n263 & ~n9850 ) | ( n3499 & ~n9850 ) ;
  assign n25893 = n25892 ^ n25252 ^ n3992 ;
  assign n25898 = n10423 ^ n9496 ^ n7421 ;
  assign n25896 = n19139 ^ n12338 ^ n4886 ;
  assign n25897 = n25896 ^ n17979 ^ n15815 ;
  assign n25894 = ( n6567 & n9991 ) | ( n6567 & n10373 ) | ( n9991 & n10373 ) ;
  assign n25895 = n25894 ^ n22469 ^ n22422 ;
  assign n25899 = n25898 ^ n25897 ^ n25895 ;
  assign n25900 = n13430 ^ n12874 ^ n8829 ;
  assign n25901 = n19848 ^ n12440 ^ n8509 ;
  assign n25902 = ( n4913 & n5327 ) | ( n4913 & ~n25901 ) | ( n5327 & ~n25901 ) ;
  assign n25903 = ( ~n11394 & n15289 ) | ( ~n11394 & n25902 ) | ( n15289 & n25902 ) ;
  assign n25904 = ( n12902 & n13171 ) | ( n12902 & n25903 ) | ( n13171 & n25903 ) ;
  assign n25905 = n25904 ^ n9243 ^ n1020 ;
  assign n25906 = n7019 ^ n3358 ^ n2293 ;
  assign n25907 = ( ~n8732 & n18981 ) | ( ~n8732 & n25906 ) | ( n18981 & n25906 ) ;
  assign n25908 = ( n16902 & n17403 ) | ( n16902 & ~n25907 ) | ( n17403 & ~n25907 ) ;
  assign n25911 = ( n2360 & n17486 ) | ( n2360 & n18334 ) | ( n17486 & n18334 ) ;
  assign n25909 = ( n1950 & n3610 ) | ( n1950 & ~n22754 ) | ( n3610 & ~n22754 ) ;
  assign n25910 = n25909 ^ n3498 ^ n1361 ;
  assign n25912 = n25911 ^ n25910 ^ n14553 ;
  assign n25913 = ( ~n1509 & n2027 ) | ( ~n1509 & n17802 ) | ( n2027 & n17802 ) ;
  assign n25914 = n25913 ^ n23935 ^ n3290 ;
  assign n25915 = n10605 ^ n9126 ^ n379 ;
  assign n25916 = ( n2361 & n3840 ) | ( n2361 & ~n10628 ) | ( n3840 & ~n10628 ) ;
  assign n25917 = n25916 ^ n15157 ^ n14234 ;
  assign n25918 = n23776 ^ n15157 ^ n14420 ;
  assign n25921 = ( n5282 & ~n8448 ) | ( n5282 & n8855 ) | ( ~n8448 & n8855 ) ;
  assign n25919 = n20741 ^ n18391 ^ n14443 ;
  assign n25920 = ( n15524 & n22417 ) | ( n15524 & ~n25919 ) | ( n22417 & ~n25919 ) ;
  assign n25922 = n25921 ^ n25920 ^ n24566 ;
  assign n25923 = ( n9087 & ~n13835 ) | ( n9087 & n17501 ) | ( ~n13835 & n17501 ) ;
  assign n25924 = ( n1788 & n24555 ) | ( n1788 & n25923 ) | ( n24555 & n25923 ) ;
  assign n25926 = n16554 ^ n9335 ^ n8152 ;
  assign n25925 = ( n6988 & n14366 ) | ( n6988 & ~n14528 ) | ( n14366 & ~n14528 ) ;
  assign n25927 = n25926 ^ n25925 ^ n25140 ;
  assign n25928 = ( n1423 & ~n8734 ) | ( n1423 & n25927 ) | ( ~n8734 & n25927 ) ;
  assign n25929 = n24356 ^ n4223 ^ n768 ;
  assign n25930 = ( n5020 & n16152 ) | ( n5020 & ~n23827 ) | ( n16152 & ~n23827 ) ;
  assign n25931 = ( n959 & n8385 ) | ( n959 & n19335 ) | ( n8385 & n19335 ) ;
  assign n25935 = ( n3885 & n14664 ) | ( n3885 & n20708 ) | ( n14664 & n20708 ) ;
  assign n25932 = n10470 ^ n10339 ^ n5509 ;
  assign n25933 = ( n154 & n4381 ) | ( n154 & ~n8856 ) | ( n4381 & ~n8856 ) ;
  assign n25934 = ( n5190 & ~n25932 ) | ( n5190 & n25933 ) | ( ~n25932 & n25933 ) ;
  assign n25936 = n25935 ^ n25934 ^ n1254 ;
  assign n25937 = ( n6592 & ~n14549 ) | ( n6592 & n25936 ) | ( ~n14549 & n25936 ) ;
  assign n25944 = ( n1309 & ~n3491 ) | ( n1309 & n16144 ) | ( ~n3491 & n16144 ) ;
  assign n25940 = n18226 ^ n12269 ^ n715 ;
  assign n25941 = ( ~n6753 & n8621 ) | ( ~n6753 & n25940 ) | ( n8621 & n25940 ) ;
  assign n25942 = ( n3237 & ~n3625 ) | ( n3237 & n25941 ) | ( ~n3625 & n25941 ) ;
  assign n25943 = ( n7515 & ~n23078 ) | ( n7515 & n25942 ) | ( ~n23078 & n25942 ) ;
  assign n25938 = n21261 ^ n12596 ^ n4468 ;
  assign n25939 = n25938 ^ n7194 ^ n7184 ;
  assign n25945 = n25944 ^ n25943 ^ n25939 ;
  assign n25946 = ( n2468 & ~n7256 ) | ( n2468 & n25945 ) | ( ~n7256 & n25945 ) ;
  assign n25947 = n23826 ^ n23609 ^ n6473 ;
  assign n25948 = n21814 ^ n20165 ^ n9344 ;
  assign n25949 = ( n9443 & ~n9785 ) | ( n9443 & n25948 ) | ( ~n9785 & n25948 ) ;
  assign n25950 = ( n19115 & ~n19566 ) | ( n19115 & n19929 ) | ( ~n19566 & n19929 ) ;
  assign n25951 = ( n315 & ~n16154 ) | ( n315 & n25950 ) | ( ~n16154 & n25950 ) ;
  assign n25955 = n14876 ^ n7171 ^ n1270 ;
  assign n25954 = n10926 ^ n7165 ^ n1714 ;
  assign n25952 = ( n259 & n3891 ) | ( n259 & n22032 ) | ( n3891 & n22032 ) ;
  assign n25953 = n25952 ^ n5386 ^ n3523 ;
  assign n25956 = n25955 ^ n25954 ^ n25953 ;
  assign n25957 = n23669 ^ n14138 ^ n1913 ;
  assign n25958 = ( n4156 & ~n12245 ) | ( n4156 & n25957 ) | ( ~n12245 & n25957 ) ;
  assign n25959 = n15069 ^ n14044 ^ n12746 ;
  assign n25960 = ( n4492 & n5958 ) | ( n4492 & ~n9548 ) | ( n5958 & ~n9548 ) ;
  assign n25961 = n20749 ^ n11871 ^ n2532 ;
  assign n25962 = ( ~n6448 & n25960 ) | ( ~n6448 & n25961 ) | ( n25960 & n25961 ) ;
  assign n25963 = ( n1672 & n3339 ) | ( n1672 & n25962 ) | ( n3339 & n25962 ) ;
  assign n25964 = n25795 ^ n16644 ^ n16169 ;
  assign n25965 = n25964 ^ n10340 ^ n7469 ;
  assign n25966 = ( n3762 & n22879 ) | ( n3762 & ~n23422 ) | ( n22879 & ~n23422 ) ;
  assign n25967 = n21806 ^ n8833 ^ x58 ;
  assign n25968 = n22106 ^ n7310 ^ n5975 ;
  assign n25969 = ( n11845 & ~n13701 ) | ( n11845 & n25968 ) | ( ~n13701 & n25968 ) ;
  assign n25970 = ( n10683 & ~n12167 ) | ( n10683 & n16186 ) | ( ~n12167 & n16186 ) ;
  assign n25971 = n25970 ^ n9043 ^ n5360 ;
  assign n25972 = n25008 ^ n14132 ^ n5166 ;
  assign n25973 = n14617 ^ n8060 ^ n8014 ;
  assign n25974 = ( n4003 & ~n22592 ) | ( n4003 & n25973 ) | ( ~n22592 & n25973 ) ;
  assign n25975 = ( n17063 & n21167 ) | ( n17063 & ~n24863 ) | ( n21167 & ~n24863 ) ;
  assign n25976 = n6527 ^ n4321 ^ n2189 ;
  assign n25977 = n12119 ^ n3857 ^ n1617 ;
  assign n25978 = ( ~n9829 & n23167 ) | ( ~n9829 & n25977 ) | ( n23167 & n25977 ) ;
  assign n25979 = n13671 ^ n8222 ^ n2894 ;
  assign n25980 = ( n23119 & n25179 ) | ( n23119 & n25979 ) | ( n25179 & n25979 ) ;
  assign n25981 = n8095 ^ n6656 ^ n1162 ;
  assign n25982 = ( n13663 & ~n18882 ) | ( n13663 & n25981 ) | ( ~n18882 & n25981 ) ;
  assign n25983 = ( n5981 & n8450 ) | ( n5981 & ~n12217 ) | ( n8450 & ~n12217 ) ;
  assign n25984 = ( n896 & n5476 ) | ( n896 & n25983 ) | ( n5476 & n25983 ) ;
  assign n25985 = ( n362 & ~n22073 ) | ( n362 & n25984 ) | ( ~n22073 & n25984 ) ;
  assign n25986 = ( ~n20419 & n25982 ) | ( ~n20419 & n25985 ) | ( n25982 & n25985 ) ;
  assign n25987 = ( n4236 & n8814 ) | ( n4236 & ~n17636 ) | ( n8814 & ~n17636 ) ;
  assign n25988 = n25987 ^ n16085 ^ n8025 ;
  assign n25990 = n10915 ^ n10397 ^ n9430 ;
  assign n25989 = n10714 ^ n9852 ^ n505 ;
  assign n25991 = n25990 ^ n25989 ^ n10458 ;
  assign n25992 = ( n10937 & n21114 ) | ( n10937 & n24003 ) | ( n21114 & n24003 ) ;
  assign n25993 = ( n8374 & n9492 ) | ( n8374 & ~n17435 ) | ( n9492 & ~n17435 ) ;
  assign n25994 = n23141 ^ n16247 ^ n1930 ;
  assign n25995 = ( n21044 & n25993 ) | ( n21044 & n25994 ) | ( n25993 & n25994 ) ;
  assign n25996 = ( n5380 & n10881 ) | ( n5380 & ~n14435 ) | ( n10881 & ~n14435 ) ;
  assign n25997 = ( n817 & n25995 ) | ( n817 & n25996 ) | ( n25995 & n25996 ) ;
  assign n25998 = ( n1923 & ~n7797 ) | ( n1923 & n8450 ) | ( ~n7797 & n8450 ) ;
  assign n25999 = ( ~n4910 & n6798 ) | ( ~n4910 & n14425 ) | ( n6798 & n14425 ) ;
  assign n26000 = n25999 ^ n13977 ^ n4001 ;
  assign n26001 = n26000 ^ n11430 ^ n7322 ;
  assign n26002 = ( n6619 & ~n9135 ) | ( n6619 & n16109 ) | ( ~n9135 & n16109 ) ;
  assign n26003 = ( n25998 & ~n26001 ) | ( n25998 & n26002 ) | ( ~n26001 & n26002 ) ;
  assign n26004 = ( n5634 & ~n7416 ) | ( n5634 & n21123 ) | ( ~n7416 & n21123 ) ;
  assign n26007 = n8770 ^ n6029 ^ n3119 ;
  assign n26005 = ( n1839 & n4351 ) | ( n1839 & n11856 ) | ( n4351 & n11856 ) ;
  assign n26006 = ( ~n1352 & n23523 ) | ( ~n1352 & n26005 ) | ( n23523 & n26005 ) ;
  assign n26008 = n26007 ^ n26006 ^ n4618 ;
  assign n26009 = n18890 ^ n10028 ^ n8779 ;
  assign n26010 = ( ~n5990 & n13653 ) | ( ~n5990 & n14164 ) | ( n13653 & n14164 ) ;
  assign n26011 = ( n2445 & ~n16993 ) | ( n2445 & n26010 ) | ( ~n16993 & n26010 ) ;
  assign n26012 = n16475 ^ n10371 ^ x117 ;
  assign n26013 = n22298 ^ n9778 ^ n4862 ;
  assign n26014 = n26013 ^ n8006 ^ n6547 ;
  assign n26015 = ( n12850 & n16524 ) | ( n12850 & n26014 ) | ( n16524 & n26014 ) ;
  assign n26016 = ( n19142 & ~n26012 ) | ( n19142 & n26015 ) | ( ~n26012 & n26015 ) ;
  assign n26017 = n11352 ^ n11119 ^ n5233 ;
  assign n26018 = ( ~n1344 & n8921 ) | ( ~n1344 & n26017 ) | ( n8921 & n26017 ) ;
  assign n26019 = n22959 ^ n22471 ^ n15265 ;
  assign n26020 = n26019 ^ n11119 ^ n7301 ;
  assign n26021 = ( n6693 & n26018 ) | ( n6693 & n26020 ) | ( n26018 & n26020 ) ;
  assign n26022 = ( ~n6553 & n22762 ) | ( ~n6553 & n26021 ) | ( n22762 & n26021 ) ;
  assign n26023 = n9117 ^ n5484 ^ n1950 ;
  assign n26024 = ( n11821 & n13229 ) | ( n11821 & ~n22104 ) | ( n13229 & ~n22104 ) ;
  assign n26025 = ( n7485 & ~n26023 ) | ( n7485 & n26024 ) | ( ~n26023 & n26024 ) ;
  assign n26026 = n9122 ^ n5126 ^ n2678 ;
  assign n26027 = n26026 ^ n12805 ^ n12773 ;
  assign n26028 = n26027 ^ n19355 ^ n19277 ;
  assign n26029 = ( n1783 & n12817 ) | ( n1783 & ~n17895 ) | ( n12817 & ~n17895 ) ;
  assign n26030 = ( n4431 & ~n10813 ) | ( n4431 & n26029 ) | ( ~n10813 & n26029 ) ;
  assign n26031 = ( n319 & n18632 ) | ( n319 & n19969 ) | ( n18632 & n19969 ) ;
  assign n26032 = n26031 ^ n7441 ^ n1023 ;
  assign n26033 = n15680 ^ n7699 ^ n1756 ;
  assign n26034 = n26033 ^ n14742 ^ n9047 ;
  assign n26035 = ( n13755 & n18180 ) | ( n13755 & n22334 ) | ( n18180 & n22334 ) ;
  assign n26036 = n26035 ^ n25622 ^ n11528 ;
  assign n26037 = n9882 ^ n6521 ^ n3412 ;
  assign n26038 = ( n1743 & ~n4150 ) | ( n1743 & n26037 ) | ( ~n4150 & n26037 ) ;
  assign n26039 = n26038 ^ n22238 ^ n8339 ;
  assign n26040 = ( n5236 & n26036 ) | ( n5236 & n26039 ) | ( n26036 & n26039 ) ;
  assign n26041 = n24012 ^ n6837 ^ n6034 ;
  assign n26042 = n13662 ^ n6842 ^ n3703 ;
  assign n26044 = n3372 ^ n2869 ^ n1180 ;
  assign n26045 = n26044 ^ n7738 ^ n4481 ;
  assign n26043 = ( ~x88 & n7576 ) | ( ~x88 & n9192 ) | ( n7576 & n9192 ) ;
  assign n26046 = n26045 ^ n26043 ^ n6979 ;
  assign n26047 = ( n26041 & n26042 ) | ( n26041 & ~n26046 ) | ( n26042 & ~n26046 ) ;
  assign n26048 = ( n2536 & n4775 ) | ( n2536 & n4910 ) | ( n4775 & n4910 ) ;
  assign n26049 = n26048 ^ n7456 ^ n1766 ;
  assign n26050 = n26049 ^ n9598 ^ n9065 ;
  assign n26051 = n26050 ^ n18061 ^ n11891 ;
  assign n26052 = ( n6156 & ~n10857 ) | ( n6156 & n25143 ) | ( ~n10857 & n25143 ) ;
  assign n26053 = n26052 ^ n6492 ^ n4487 ;
  assign n26054 = n9756 ^ n8229 ^ n3268 ;
  assign n26055 = n8842 ^ n8782 ^ n280 ;
  assign n26057 = n14095 ^ n12324 ^ n7544 ;
  assign n26056 = ( n600 & ~n2799 ) | ( n600 & n3423 ) | ( ~n2799 & n3423 ) ;
  assign n26058 = n26057 ^ n26056 ^ n3094 ;
  assign n26060 = n24781 ^ n13207 ^ n2573 ;
  assign n26061 = ( ~n1522 & n2083 ) | ( ~n1522 & n26060 ) | ( n2083 & n26060 ) ;
  assign n26062 = n26061 ^ n25041 ^ n11987 ;
  assign n26059 = n5594 ^ n5420 ^ n4282 ;
  assign n26063 = n26062 ^ n26059 ^ n301 ;
  assign n26064 = ( n5127 & n7902 ) | ( n5127 & n18256 ) | ( n7902 & n18256 ) ;
  assign n26065 = ( n6645 & n19832 ) | ( n6645 & n26064 ) | ( n19832 & n26064 ) ;
  assign n26066 = ( ~n6564 & n15209 ) | ( ~n6564 & n26065 ) | ( n15209 & n26065 ) ;
  assign n26067 = ( ~n4258 & n8376 ) | ( ~n4258 & n12082 ) | ( n8376 & n12082 ) ;
  assign n26068 = n23809 ^ n6537 ^ n6106 ;
  assign n26069 = ( n7210 & n16459 ) | ( n7210 & n26068 ) | ( n16459 & n26068 ) ;
  assign n26070 = ( n22297 & n26067 ) | ( n22297 & n26069 ) | ( n26067 & n26069 ) ;
  assign n26071 = ( n788 & n8906 ) | ( n788 & ~n26070 ) | ( n8906 & ~n26070 ) ;
  assign n26072 = n6379 ^ n2597 ^ n1456 ;
  assign n26076 = n18604 ^ n7998 ^ n7443 ;
  assign n26075 = n18106 ^ n8947 ^ n3926 ;
  assign n26077 = n26076 ^ n26075 ^ n5376 ;
  assign n26073 = ( n10753 & n15635 ) | ( n10753 & n16821 ) | ( n15635 & n16821 ) ;
  assign n26074 = ( n211 & n1010 ) | ( n211 & n26073 ) | ( n1010 & n26073 ) ;
  assign n26078 = n26077 ^ n26074 ^ n4132 ;
  assign n26079 = n9691 ^ n1848 ^ n625 ;
  assign n26080 = ( n16458 & n21210 ) | ( n16458 & ~n25568 ) | ( n21210 & ~n25568 ) ;
  assign n26081 = ( n3531 & n13009 ) | ( n3531 & ~n14760 ) | ( n13009 & ~n14760 ) ;
  assign n26082 = n26081 ^ n3624 ^ n369 ;
  assign n26083 = n20587 ^ n19951 ^ n15853 ;
  assign n26084 = n26083 ^ n24624 ^ n11707 ;
  assign n26085 = ( n9796 & n14459 ) | ( n9796 & ~n26084 ) | ( n14459 & ~n26084 ) ;
  assign n26086 = ( n5392 & n7093 ) | ( n5392 & n9203 ) | ( n7093 & n9203 ) ;
  assign n26087 = ( n2380 & n5180 ) | ( n2380 & n26086 ) | ( n5180 & n26086 ) ;
  assign n26088 = n26087 ^ n23978 ^ n21223 ;
  assign n26089 = ( n1635 & n10480 ) | ( n1635 & n26088 ) | ( n10480 & n26088 ) ;
  assign n26090 = n26089 ^ n5647 ^ n5217 ;
  assign n26091 = n7377 ^ n5376 ^ n1850 ;
  assign n26092 = ( n5225 & n6784 ) | ( n5225 & n26091 ) | ( n6784 & n26091 ) ;
  assign n26093 = n26092 ^ n2985 ^ n1611 ;
  assign n26094 = ( n6833 & ~n25205 ) | ( n6833 & n26093 ) | ( ~n25205 & n26093 ) ;
  assign n26095 = ( n8160 & n9633 ) | ( n8160 & ~n21963 ) | ( n9633 & ~n21963 ) ;
  assign n26096 = n26095 ^ n24399 ^ n14110 ;
  assign n26099 = n25472 ^ n15381 ^ n13658 ;
  assign n26097 = ( ~n5820 & n6860 ) | ( ~n5820 & n12038 ) | ( n6860 & n12038 ) ;
  assign n26098 = n26097 ^ n3945 ^ n3253 ;
  assign n26100 = n26099 ^ n26098 ^ n21397 ;
  assign n26101 = ( ~n4266 & n24071 ) | ( ~n4266 & n24829 ) | ( n24071 & n24829 ) ;
  assign n26102 = n2942 ^ n1810 ^ n534 ;
  assign n26103 = n26102 ^ n26000 ^ n12868 ;
  assign n26104 = n11829 ^ n7722 ^ n7570 ;
  assign n26105 = ( ~n6425 & n18350 ) | ( ~n6425 & n26104 ) | ( n18350 & n26104 ) ;
  assign n26106 = n20778 ^ n9472 ^ n1121 ;
  assign n26107 = n26106 ^ n16606 ^ n16218 ;
  assign n26108 = ( n19966 & ~n26105 ) | ( n19966 & n26107 ) | ( ~n26105 & n26107 ) ;
  assign n26109 = ( ~n6732 & n26103 ) | ( ~n6732 & n26108 ) | ( n26103 & n26108 ) ;
  assign n26110 = n16564 ^ n13961 ^ n5326 ;
  assign n26111 = n26110 ^ n5687 ^ n4907 ;
  assign n26112 = n14596 ^ n8304 ^ n5375 ;
  assign n26113 = n26112 ^ n24779 ^ n16077 ;
  assign n26114 = n12342 ^ n7046 ^ n3416 ;
  assign n26115 = n26114 ^ n3443 ^ n205 ;
  assign n26116 = n26115 ^ n8532 ^ n3779 ;
  assign n26117 = n26116 ^ n19911 ^ n5779 ;
  assign n26118 = n16516 ^ n7864 ^ n1022 ;
  assign n26119 = n26118 ^ n5884 ^ n3223 ;
  assign n26120 = ( n1776 & n12377 ) | ( n1776 & n26119 ) | ( n12377 & n26119 ) ;
  assign n26121 = ( n1346 & n6954 ) | ( n1346 & n10674 ) | ( n6954 & n10674 ) ;
  assign n26122 = n18232 ^ n6525 ^ n282 ;
  assign n26123 = n21581 ^ n10178 ^ n8670 ;
  assign n26124 = n19579 ^ n7346 ^ n3812 ;
  assign n26125 = ( n9816 & n21610 ) | ( n9816 & n26124 ) | ( n21610 & n26124 ) ;
  assign n26126 = ( x69 & ~n14121 ) | ( x69 & n26125 ) | ( ~n14121 & n26125 ) ;
  assign n26127 = ( n13720 & ~n26123 ) | ( n13720 & n26126 ) | ( ~n26123 & n26126 ) ;
  assign n26128 = ( n6346 & ~n26122 ) | ( n6346 & n26127 ) | ( ~n26122 & n26127 ) ;
  assign n26129 = ( x67 & n11464 ) | ( x67 & n18792 ) | ( n11464 & n18792 ) ;
  assign n26130 = n26129 ^ n17158 ^ n7798 ;
  assign n26131 = n26130 ^ n24851 ^ n7593 ;
  assign n26132 = n26131 ^ n4180 ^ x35 ;
  assign n26133 = n26132 ^ n5616 ^ n2690 ;
  assign n26134 = n6732 ^ n5007 ^ n4907 ;
  assign n26135 = n26134 ^ n10931 ^ n9543 ;
  assign n26136 = ( n747 & ~n2020 ) | ( n747 & n4483 ) | ( ~n2020 & n4483 ) ;
  assign n26137 = n26136 ^ n16525 ^ n10207 ;
  assign n26138 = ( ~n10442 & n11689 ) | ( ~n10442 & n21951 ) | ( n11689 & n21951 ) ;
  assign n26139 = ( n1356 & ~n13920 ) | ( n1356 & n26138 ) | ( ~n13920 & n26138 ) ;
  assign n26140 = n26139 ^ n14801 ^ n12197 ;
  assign n26141 = n20327 ^ n3442 ^ n349 ;
  assign n26142 = n22032 ^ n18458 ^ n6855 ;
  assign n26143 = ( n2998 & ~n4666 ) | ( n2998 & n5126 ) | ( ~n4666 & n5126 ) ;
  assign n26144 = n26143 ^ n17750 ^ n15550 ;
  assign n26145 = ( n13511 & n26142 ) | ( n13511 & n26144 ) | ( n26142 & n26144 ) ;
  assign n26146 = ( n283 & n13474 ) | ( n283 & n26145 ) | ( n13474 & n26145 ) ;
  assign n26147 = n22821 ^ n10193 ^ n6405 ;
  assign n26148 = ( n898 & n5787 ) | ( n898 & n8420 ) | ( n5787 & n8420 ) ;
  assign n26149 = ( n6699 & n8561 ) | ( n6699 & ~n18829 ) | ( n8561 & ~n18829 ) ;
  assign n26150 = n9970 ^ n7302 ^ n5470 ;
  assign n26151 = n14819 ^ n13068 ^ n1008 ;
  assign n26152 = n14902 ^ n9175 ^ n960 ;
  assign n26153 = n26152 ^ n6751 ^ n3048 ;
  assign n26154 = n16870 ^ n4753 ^ n4687 ;
  assign n26155 = ( n6106 & n7508 ) | ( n6106 & n8227 ) | ( n7508 & n8227 ) ;
  assign n26156 = n14637 ^ n13346 ^ n3378 ;
  assign n26157 = ( ~n2427 & n25741 ) | ( ~n2427 & n26156 ) | ( n25741 & n26156 ) ;
  assign n26158 = ( x19 & ~n1249 ) | ( x19 & n18858 ) | ( ~n1249 & n18858 ) ;
  assign n26159 = n23058 ^ n19757 ^ n9858 ;
  assign n26160 = n26159 ^ n5889 ^ x73 ;
  assign n26161 = ( n838 & n24780 ) | ( n838 & n26160 ) | ( n24780 & n26160 ) ;
  assign n26162 = ( n2995 & n4644 ) | ( n2995 & ~n11390 ) | ( n4644 & ~n11390 ) ;
  assign n26163 = ( ~n23378 & n24942 ) | ( ~n23378 & n26162 ) | ( n24942 & n26162 ) ;
  assign n26164 = ( n22551 & ~n23554 ) | ( n22551 & n25750 ) | ( ~n23554 & n25750 ) ;
  assign n26165 = ( n12331 & ~n24555 ) | ( n12331 & n26164 ) | ( ~n24555 & n26164 ) ;
  assign n26166 = n22075 ^ n9629 ^ n4303 ;
  assign n26167 = ( n5912 & n22049 ) | ( n5912 & n26166 ) | ( n22049 & n26166 ) ;
  assign n26168 = ( ~n8392 & n20566 ) | ( ~n8392 & n26167 ) | ( n20566 & n26167 ) ;
  assign n26169 = ( n17907 & n23893 ) | ( n17907 & n26168 ) | ( n23893 & n26168 ) ;
  assign n26170 = n8038 ^ n7424 ^ n2749 ;
  assign n26171 = n26170 ^ n16239 ^ n10603 ;
  assign n26172 = ( n3828 & n17366 ) | ( n3828 & ~n24302 ) | ( n17366 & ~n24302 ) ;
  assign n26173 = n26172 ^ n6127 ^ n898 ;
  assign n26174 = ( n11182 & ~n26171 ) | ( n11182 & n26173 ) | ( ~n26171 & n26173 ) ;
  assign n26175 = ( ~n15345 & n18638 ) | ( ~n15345 & n26007 ) | ( n18638 & n26007 ) ;
  assign n26176 = ( n4325 & n19659 ) | ( n4325 & ~n24007 ) | ( n19659 & ~n24007 ) ;
  assign n26177 = ( n6873 & ~n9226 ) | ( n6873 & n20488 ) | ( ~n9226 & n20488 ) ;
  assign n26178 = n26177 ^ n6747 ^ n3309 ;
  assign n26179 = ( n1620 & n10124 ) | ( n1620 & n26178 ) | ( n10124 & n26178 ) ;
  assign n26180 = ( n7015 & ~n15164 ) | ( n7015 & n26179 ) | ( ~n15164 & n26179 ) ;
  assign n26181 = n26180 ^ n12331 ^ n7940 ;
  assign n26182 = ( n1467 & n2353 ) | ( n1467 & ~n15685 ) | ( n2353 & ~n15685 ) ;
  assign n26183 = ( n2916 & ~n23420 ) | ( n2916 & n26182 ) | ( ~n23420 & n26182 ) ;
  assign n26184 = ( n16573 & n17495 ) | ( n16573 & ~n18134 ) | ( n17495 & ~n18134 ) ;
  assign n26185 = ( ~n537 & n19654 ) | ( ~n537 & n23266 ) | ( n19654 & n23266 ) ;
  assign n26186 = n5089 ^ n2977 ^ n1649 ;
  assign n26187 = n26186 ^ n20405 ^ n3610 ;
  assign n26188 = ( ~n11630 & n12792 ) | ( ~n11630 & n26159 ) | ( n12792 & n26159 ) ;
  assign n26189 = n24384 ^ n15205 ^ n12631 ;
  assign n26190 = ( n2751 & n3861 ) | ( n2751 & ~n20218 ) | ( n3861 & ~n20218 ) ;
  assign n26191 = ( n5969 & n8331 ) | ( n5969 & n26190 ) | ( n8331 & n26190 ) ;
  assign n26194 = ( n1071 & n2255 ) | ( n1071 & ~n3116 ) | ( n2255 & ~n3116 ) ;
  assign n26195 = ( n1213 & n5118 ) | ( n1213 & n26194 ) | ( n5118 & n26194 ) ;
  assign n26192 = ( ~n350 & n1280 ) | ( ~n350 & n7329 ) | ( n1280 & n7329 ) ;
  assign n26193 = ( n16204 & ~n19830 ) | ( n16204 & n26192 ) | ( ~n19830 & n26192 ) ;
  assign n26196 = n26195 ^ n26193 ^ n14535 ;
  assign n26197 = ( n1597 & n1652 ) | ( n1597 & ~n5795 ) | ( n1652 & ~n5795 ) ;
  assign n26198 = n26197 ^ n15440 ^ n2376 ;
  assign n26199 = n26198 ^ n15726 ^ n11618 ;
  assign n26200 = ( n1561 & ~n3694 ) | ( n1561 & n15277 ) | ( ~n3694 & n15277 ) ;
  assign n26201 = n26200 ^ n10559 ^ n5315 ;
  assign n26202 = n23308 ^ n12701 ^ n8332 ;
  assign n26203 = ( n1145 & n3159 ) | ( n1145 & n3267 ) | ( n3159 & n3267 ) ;
  assign n26204 = n26203 ^ n12730 ^ n6739 ;
  assign n26205 = n26204 ^ n13980 ^ n13270 ;
  assign n26206 = ( ~n1530 & n1561 ) | ( ~n1530 & n23124 ) | ( n1561 & n23124 ) ;
  assign n26207 = n23246 ^ n20546 ^ n2325 ;
  assign n26208 = n26207 ^ n25176 ^ n14896 ;
  assign n26209 = ( n1236 & n3634 ) | ( n1236 & ~n22106 ) | ( n3634 & ~n22106 ) ;
  assign n26210 = ( n14412 & n26194 ) | ( n14412 & n26209 ) | ( n26194 & n26209 ) ;
  assign n26211 = n13966 ^ n10119 ^ n726 ;
  assign n26212 = ( ~n884 & n2370 ) | ( ~n884 & n20840 ) | ( n2370 & n20840 ) ;
  assign n26213 = ( n6019 & n18735 ) | ( n6019 & n26212 ) | ( n18735 & n26212 ) ;
  assign n26214 = n26213 ^ n8075 ^ n7505 ;
  assign n26215 = ( ~n10198 & n14573 ) | ( ~n10198 & n18743 ) | ( n14573 & n18743 ) ;
  assign n26216 = n26215 ^ n17951 ^ n15291 ;
  assign n26217 = ( n25414 & n26214 ) | ( n25414 & ~n26216 ) | ( n26214 & ~n26216 ) ;
  assign n26218 = n25296 ^ n14730 ^ n5407 ;
  assign n26219 = n20288 ^ n14195 ^ n4828 ;
  assign n26220 = n26219 ^ n13708 ^ x89 ;
  assign n26221 = n26220 ^ n16352 ^ n11015 ;
  assign n26222 = ( ~n5874 & n6958 ) | ( ~n5874 & n26081 ) | ( n6958 & n26081 ) ;
  assign n26223 = n11220 ^ n5170 ^ n1867 ;
  assign n26224 = n26223 ^ n16312 ^ n7887 ;
  assign n26225 = n26224 ^ n17879 ^ n16785 ;
  assign n26226 = ( n8260 & ~n16291 ) | ( n8260 & n26225 ) | ( ~n16291 & n26225 ) ;
  assign n26227 = n15587 ^ n8885 ^ n1499 ;
  assign n26228 = ( n2714 & n22457 ) | ( n2714 & ~n26227 ) | ( n22457 & ~n26227 ) ;
  assign n26229 = n26228 ^ n22211 ^ n4741 ;
  assign n26230 = n23706 ^ n20462 ^ n3981 ;
  assign n26231 = n25925 ^ n3592 ^ n2728 ;
  assign n26232 = ( n2662 & n5946 ) | ( n2662 & n23299 ) | ( n5946 & n23299 ) ;
  assign n26233 = n16136 ^ n14312 ^ n12185 ;
  assign n26234 = ( n3462 & ~n18603 ) | ( n3462 & n22706 ) | ( ~n18603 & n22706 ) ;
  assign n26235 = ( n23474 & ~n24897 ) | ( n23474 & n26234 ) | ( ~n24897 & n26234 ) ;
  assign n26236 = ( n9321 & ~n10993 ) | ( n9321 & n18365 ) | ( ~n10993 & n18365 ) ;
  assign n26237 = ( ~n7254 & n15166 ) | ( ~n7254 & n26236 ) | ( n15166 & n26236 ) ;
  assign n26238 = n11207 ^ n10910 ^ n4130 ;
  assign n26239 = n26238 ^ n23661 ^ n1460 ;
  assign n26240 = ( n426 & ~n23721 ) | ( n426 & n26239 ) | ( ~n23721 & n26239 ) ;
  assign n26241 = ( ~n18012 & n26237 ) | ( ~n18012 & n26240 ) | ( n26237 & n26240 ) ;
  assign n26242 = ( n4300 & n15575 ) | ( n4300 & ~n17014 ) | ( n15575 & ~n17014 ) ;
  assign n26243 = ( n1911 & ~n6150 ) | ( n1911 & n26242 ) | ( ~n6150 & n26242 ) ;
  assign n26244 = ( ~n4873 & n16730 ) | ( ~n4873 & n26243 ) | ( n16730 & n26243 ) ;
  assign n26245 = n25851 ^ n4659 ^ n554 ;
  assign n26246 = ( n14890 & ~n22189 ) | ( n14890 & n26245 ) | ( ~n22189 & n26245 ) ;
  assign n26247 = ( ~n2596 & n21463 ) | ( ~n2596 & n26246 ) | ( n21463 & n26246 ) ;
  assign n26248 = n11754 ^ n6114 ^ n4734 ;
  assign n26249 = ( n556 & n5751 ) | ( n556 & ~n8725 ) | ( n5751 & ~n8725 ) ;
  assign n26250 = ( n7020 & n8545 ) | ( n7020 & n24711 ) | ( n8545 & n24711 ) ;
  assign n26251 = n26250 ^ n7575 ^ n610 ;
  assign n26252 = ( ~n4322 & n6237 ) | ( ~n4322 & n14815 ) | ( n6237 & n14815 ) ;
  assign n26253 = ( n1101 & ~n12859 ) | ( n1101 & n25821 ) | ( ~n12859 & n25821 ) ;
  assign n26254 = ( n2684 & n4800 ) | ( n2684 & ~n15884 ) | ( n4800 & ~n15884 ) ;
  assign n26255 = n26254 ^ n20749 ^ n4226 ;
  assign n26256 = ( ~n9257 & n9478 ) | ( ~n9257 & n15912 ) | ( n9478 & n15912 ) ;
  assign n26257 = ( n587 & ~n10581 ) | ( n587 & n17193 ) | ( ~n10581 & n17193 ) ;
  assign n26258 = n21763 ^ n11153 ^ n7225 ;
  assign n26259 = ( ~n2241 & n3619 ) | ( ~n2241 & n11200 ) | ( n3619 & n11200 ) ;
  assign n26262 = ( ~n2297 & n7181 ) | ( ~n2297 & n9132 ) | ( n7181 & n9132 ) ;
  assign n26260 = ( n321 & n8544 ) | ( n321 & ~n14823 ) | ( n8544 & ~n14823 ) ;
  assign n26261 = n26260 ^ n25443 ^ n18920 ;
  assign n26263 = n26262 ^ n26261 ^ n22095 ;
  assign n26264 = ( n20103 & n21449 ) | ( n20103 & n23018 ) | ( n21449 & n23018 ) ;
  assign n26265 = ( n3260 & ~n16632 ) | ( n3260 & n26264 ) | ( ~n16632 & n26264 ) ;
  assign n26266 = ( n2425 & n9148 ) | ( n2425 & n26265 ) | ( n9148 & n26265 ) ;
  assign n26267 = ( ~n2369 & n6952 ) | ( ~n2369 & n13409 ) | ( n6952 & n13409 ) ;
  assign n26268 = ( n456 & n25005 ) | ( n456 & n25239 ) | ( n25005 & n25239 ) ;
  assign n26269 = ( n3951 & n26267 ) | ( n3951 & n26268 ) | ( n26267 & n26268 ) ;
  assign n26271 = n20691 ^ n13191 ^ n4584 ;
  assign n26272 = n26271 ^ n10594 ^ n5900 ;
  assign n26270 = n26204 ^ n21648 ^ n675 ;
  assign n26273 = n26272 ^ n26270 ^ n9051 ;
  assign n26274 = ( n1745 & n6550 ) | ( n1745 & n13638 ) | ( n6550 & n13638 ) ;
  assign n26275 = n26274 ^ n24347 ^ n17221 ;
  assign n26276 = ( n157 & n19656 ) | ( n157 & ~n20080 ) | ( n19656 & ~n20080 ) ;
  assign n26277 = n13344 ^ n7593 ^ n3440 ;
  assign n26278 = ( n586 & ~n8797 ) | ( n586 & n11369 ) | ( ~n8797 & n11369 ) ;
  assign n26279 = n26278 ^ n9687 ^ n6353 ;
  assign n26280 = ( ~n7670 & n13389 ) | ( ~n7670 & n21104 ) | ( n13389 & n21104 ) ;
  assign n26281 = n26280 ^ n20207 ^ n664 ;
  assign n26282 = ( n6239 & n7655 ) | ( n6239 & n7991 ) | ( n7655 & n7991 ) ;
  assign n26283 = n15272 ^ n14939 ^ n4223 ;
  assign n26284 = ( n22804 & ~n26282 ) | ( n22804 & n26283 ) | ( ~n26282 & n26283 ) ;
  assign n26285 = ( n576 & n6154 ) | ( n576 & ~n14379 ) | ( n6154 & ~n14379 ) ;
  assign n26286 = ( n6161 & ~n9274 ) | ( n6161 & n18697 ) | ( ~n9274 & n18697 ) ;
  assign n26287 = n26286 ^ n21487 ^ n13236 ;
  assign n26288 = n10289 ^ n7447 ^ n6490 ;
  assign n26289 = ( ~n502 & n1283 ) | ( ~n502 & n15667 ) | ( n1283 & n15667 ) ;
  assign n26290 = n26289 ^ n25258 ^ n10149 ;
  assign n26291 = n18704 ^ n9050 ^ n7322 ;
  assign n26292 = n21799 ^ n16742 ^ n2083 ;
  assign n26293 = ( n23474 & n26291 ) | ( n23474 & ~n26292 ) | ( n26291 & ~n26292 ) ;
  assign n26294 = n20402 ^ n16912 ^ n6867 ;
  assign n26295 = ( n4497 & n15865 ) | ( n4497 & ~n17401 ) | ( n15865 & ~n17401 ) ;
  assign n26296 = n26295 ^ n25803 ^ n3263 ;
  assign n26297 = ( n3341 & ~n9780 ) | ( n3341 & n26296 ) | ( ~n9780 & n26296 ) ;
  assign n26298 = ( n3379 & ~n4512 ) | ( n3379 & n26297 ) | ( ~n4512 & n26297 ) ;
  assign n26299 = n17056 ^ n10773 ^ n4275 ;
  assign n26300 = n22908 ^ n16509 ^ n11134 ;
  assign n26301 = ( n3191 & n11678 ) | ( n3191 & n18676 ) | ( n11678 & n18676 ) ;
  assign n26302 = n26301 ^ n15917 ^ n14610 ;
  assign n26303 = ( n11196 & ~n12947 ) | ( n11196 & n21377 ) | ( ~n12947 & n21377 ) ;
  assign n26304 = ( ~n8749 & n9967 ) | ( ~n8749 & n26303 ) | ( n9967 & n26303 ) ;
  assign n26305 = n15894 ^ n6559 ^ n1572 ;
  assign n26306 = n7326 ^ n2069 ^ n1524 ;
  assign n26308 = ( n11407 & n14953 ) | ( n11407 & ~n24029 ) | ( n14953 & ~n24029 ) ;
  assign n26307 = ( n12668 & ~n16773 ) | ( n12668 & n17252 ) | ( ~n16773 & n17252 ) ;
  assign n26309 = n26308 ^ n26307 ^ n6501 ;
  assign n26310 = ( n2147 & n6069 ) | ( n2147 & ~n13671 ) | ( n6069 & ~n13671 ) ;
  assign n26311 = n26310 ^ n10423 ^ n10305 ;
  assign n26312 = n17999 ^ n11154 ^ n693 ;
  assign n26313 = ( ~n11702 & n26311 ) | ( ~n11702 & n26312 ) | ( n26311 & n26312 ) ;
  assign n26314 = ( ~n1753 & n5646 ) | ( ~n1753 & n8378 ) | ( n5646 & n8378 ) ;
  assign n26315 = ( n3209 & ~n11428 ) | ( n3209 & n16071 ) | ( ~n11428 & n16071 ) ;
  assign n26316 = n23566 ^ n15912 ^ n9676 ;
  assign n26323 = ( n4898 & n8113 ) | ( n4898 & ~n21828 ) | ( n8113 & ~n21828 ) ;
  assign n26319 = n19573 ^ n13016 ^ n2150 ;
  assign n26320 = ( n6324 & n7625 ) | ( n6324 & n26319 ) | ( n7625 & n26319 ) ;
  assign n26321 = n26320 ^ n18454 ^ n4658 ;
  assign n26322 = n26321 ^ n23828 ^ n14922 ;
  assign n26317 = ( n2595 & ~n9589 ) | ( n2595 & n10845 ) | ( ~n9589 & n10845 ) ;
  assign n26318 = n26317 ^ n8247 ^ n1259 ;
  assign n26324 = n26323 ^ n26322 ^ n26318 ;
  assign n26325 = ( ~n2631 & n8576 ) | ( ~n2631 & n13115 ) | ( n8576 & n13115 ) ;
  assign n26326 = n26325 ^ n8264 ^ n7935 ;
  assign n26327 = n6002 ^ n4132 ^ n4077 ;
  assign n26328 = n22264 ^ n7791 ^ n7368 ;
  assign n26329 = ( n10892 & ~n17481 ) | ( n10892 & n26328 ) | ( ~n17481 & n26328 ) ;
  assign n26330 = ( n8754 & ~n12421 ) | ( n8754 & n16306 ) | ( ~n12421 & n16306 ) ;
  assign n26331 = ( n17442 & ~n23315 ) | ( n17442 & n26330 ) | ( ~n23315 & n26330 ) ;
  assign n26332 = n26331 ^ n14618 ^ n12441 ;
  assign n26333 = ( ~n5064 & n9466 ) | ( ~n5064 & n12732 ) | ( n9466 & n12732 ) ;
  assign n26334 = ( n3095 & n5669 ) | ( n3095 & n7794 ) | ( n5669 & n7794 ) ;
  assign n26335 = n26334 ^ n13873 ^ n12321 ;
  assign n26336 = n25285 ^ n15754 ^ n5099 ;
  assign n26337 = ( n4396 & n13160 ) | ( n4396 & n23976 ) | ( n13160 & n23976 ) ;
  assign n26338 = ( n4413 & ~n7112 ) | ( n4413 & n7506 ) | ( ~n7112 & n7506 ) ;
  assign n26339 = n26338 ^ n18959 ^ n13932 ;
  assign n26340 = ( n1119 & ~n20523 ) | ( n1119 & n26339 ) | ( ~n20523 & n26339 ) ;
  assign n26341 = n17525 ^ n13485 ^ n10066 ;
  assign n26342 = ( n2837 & ~n3627 ) | ( n2837 & n13191 ) | ( ~n3627 & n13191 ) ;
  assign n26343 = ( n15616 & ~n19037 ) | ( n15616 & n26342 ) | ( ~n19037 & n26342 ) ;
  assign n26344 = ( ~n1449 & n26190 ) | ( ~n1449 & n26343 ) | ( n26190 & n26343 ) ;
  assign n26345 = n26344 ^ n21854 ^ n20980 ;
  assign n26346 = ( ~n5508 & n26341 ) | ( ~n5508 & n26345 ) | ( n26341 & n26345 ) ;
  assign n26347 = n12348 ^ n8139 ^ n2889 ;
  assign n26348 = n14659 ^ n12532 ^ n5460 ;
  assign n26349 = n23901 ^ n12577 ^ n3888 ;
  assign n26350 = ( n20845 & n26348 ) | ( n20845 & n26349 ) | ( n26348 & n26349 ) ;
  assign n26352 = n15594 ^ n13298 ^ n9776 ;
  assign n26351 = ( n2517 & n6087 ) | ( n2517 & ~n24459 ) | ( n6087 & ~n24459 ) ;
  assign n26353 = n26352 ^ n26351 ^ n10911 ;
  assign n26354 = ( n1286 & n17655 ) | ( n1286 & ~n19118 ) | ( n17655 & ~n19118 ) ;
  assign n26355 = n26354 ^ n23082 ^ n18066 ;
  assign n26356 = n12074 ^ n5363 ^ n1129 ;
  assign n26357 = n26356 ^ n13527 ^ n1400 ;
  assign n26358 = ( n2489 & n5048 ) | ( n2489 & n26357 ) | ( n5048 & n26357 ) ;
  assign n26360 = n13869 ^ n7549 ^ n1406 ;
  assign n26359 = n24101 ^ n16828 ^ x56 ;
  assign n26361 = n26360 ^ n26359 ^ n4843 ;
  assign n26362 = ( n424 & n9125 ) | ( n424 & n23684 ) | ( n9125 & n23684 ) ;
  assign n26363 = ( n1461 & ~n6835 ) | ( n1461 & n7999 ) | ( ~n6835 & n7999 ) ;
  assign n26364 = n26363 ^ n2590 ^ n1218 ;
  assign n26365 = ( n6148 & n7802 ) | ( n6148 & n13729 ) | ( n7802 & n13729 ) ;
  assign n26366 = ( n9574 & ~n26364 ) | ( n9574 & n26365 ) | ( ~n26364 & n26365 ) ;
  assign n26367 = ( n14716 & n16949 ) | ( n14716 & ~n23827 ) | ( n16949 & ~n23827 ) ;
  assign n26368 = ( n3211 & ~n5814 ) | ( n3211 & n15151 ) | ( ~n5814 & n15151 ) ;
  assign n26369 = n26368 ^ n26098 ^ n15691 ;
  assign n26370 = ( n14033 & ~n19951 ) | ( n14033 & n22131 ) | ( ~n19951 & n22131 ) ;
  assign n26371 = ( ~n1307 & n2819 ) | ( ~n1307 & n26370 ) | ( n2819 & n26370 ) ;
  assign n26372 = ( n4159 & ~n14707 ) | ( n4159 & n18744 ) | ( ~n14707 & n18744 ) ;
  assign n26373 = n26372 ^ n20128 ^ n9524 ;
  assign n26374 = ( ~n16226 & n25022 ) | ( ~n16226 & n26373 ) | ( n25022 & n26373 ) ;
  assign n26375 = ( ~n4927 & n7616 ) | ( ~n4927 & n19302 ) | ( n7616 & n19302 ) ;
  assign n26376 = n26375 ^ n7410 ^ n6685 ;
  assign n26377 = n21769 ^ n13661 ^ n2579 ;
  assign n26378 = n26377 ^ n4782 ^ n848 ;
  assign n26379 = n6365 ^ n5486 ^ n1927 ;
  assign n26380 = n26379 ^ n12229 ^ n3454 ;
  assign n26381 = n26380 ^ n14255 ^ n13379 ;
  assign n26382 = n26381 ^ n20274 ^ n12568 ;
  assign n26383 = n13243 ^ n5886 ^ n2232 ;
  assign n26384 = n20493 ^ n9011 ^ n4997 ;
  assign n26385 = ( ~n5684 & n8545 ) | ( ~n5684 & n9936 ) | ( n8545 & n9936 ) ;
  assign n26386 = n26385 ^ n18456 ^ n4631 ;
  assign n26387 = ( ~n6141 & n26384 ) | ( ~n6141 & n26386 ) | ( n26384 & n26386 ) ;
  assign n26388 = ( ~n3389 & n26383 ) | ( ~n3389 & n26387 ) | ( n26383 & n26387 ) ;
  assign n26389 = ( n7023 & ~n7761 ) | ( n7023 & n15510 ) | ( ~n7761 & n15510 ) ;
  assign n26390 = n26389 ^ n18845 ^ n15183 ;
  assign n26391 = ( n4315 & ~n4925 ) | ( n4315 & n22056 ) | ( ~n4925 & n22056 ) ;
  assign n26392 = n26391 ^ n6598 ^ x76 ;
  assign n26395 = n12100 ^ n7958 ^ n7277 ;
  assign n26393 = n9530 ^ n3041 ^ n476 ;
  assign n26394 = n26393 ^ n5826 ^ n2108 ;
  assign n26396 = n26395 ^ n26394 ^ n21798 ;
  assign n26399 = n20467 ^ n4328 ^ n4039 ;
  assign n26397 = n13647 ^ n3866 ^ n1495 ;
  assign n26398 = ( n8675 & ~n11898 ) | ( n8675 & n26397 ) | ( ~n11898 & n26397 ) ;
  assign n26400 = n26399 ^ n26398 ^ n3868 ;
  assign n26403 = n20186 ^ n14320 ^ n12949 ;
  assign n26404 = n26403 ^ n22101 ^ n1359 ;
  assign n26401 = n14243 ^ n3140 ^ n971 ;
  assign n26402 = ( ~n5280 & n14042 ) | ( ~n5280 & n26401 ) | ( n14042 & n26401 ) ;
  assign n26405 = n26404 ^ n26402 ^ n8375 ;
  assign n26406 = ( n2008 & ~n4638 ) | ( n2008 & n9502 ) | ( ~n4638 & n9502 ) ;
  assign n26407 = ( ~n13823 & n16386 ) | ( ~n13823 & n26406 ) | ( n16386 & n26406 ) ;
  assign n26408 = ( n17640 & n19901 ) | ( n17640 & n26407 ) | ( n19901 & n26407 ) ;
  assign n26409 = n14938 ^ n11851 ^ n1044 ;
  assign n26410 = ( n4091 & n7094 ) | ( n4091 & n26409 ) | ( n7094 & n26409 ) ;
  assign n26411 = n4043 ^ n3626 ^ n1106 ;
  assign n26412 = ( n7737 & ~n9477 ) | ( n7737 & n16069 ) | ( ~n9477 & n16069 ) ;
  assign n26413 = ( n4511 & n7987 ) | ( n4511 & ~n26412 ) | ( n7987 & ~n26412 ) ;
  assign n26414 = ( n7468 & n19600 ) | ( n7468 & n22238 ) | ( n19600 & n22238 ) ;
  assign n26416 = n25207 ^ n17928 ^ n792 ;
  assign n26415 = ( n17206 & n21609 ) | ( n17206 & ~n24563 ) | ( n21609 & ~n24563 ) ;
  assign n26417 = n26416 ^ n26415 ^ n15636 ;
  assign n26418 = ( n2732 & ~n12020 ) | ( n2732 & n12906 ) | ( ~n12020 & n12906 ) ;
  assign n26419 = n6464 ^ n2361 ^ n1673 ;
  assign n26420 = ( n10845 & n13100 ) | ( n10845 & n26419 ) | ( n13100 & n26419 ) ;
  assign n26422 = n2222 ^ n1824 ^ n782 ;
  assign n26421 = n12118 ^ n12083 ^ n2421 ;
  assign n26423 = n26422 ^ n26421 ^ n5946 ;
  assign n26424 = n26423 ^ n8141 ^ n7985 ;
  assign n26425 = n17857 ^ n13233 ^ n9006 ;
  assign n26427 = n20310 ^ n1243 ^ n1183 ;
  assign n26426 = n23690 ^ n4631 ^ n2621 ;
  assign n26428 = n26427 ^ n26426 ^ n6329 ;
  assign n26429 = ( n2118 & n4225 ) | ( n2118 & n6717 ) | ( n4225 & n6717 ) ;
  assign n26430 = n26429 ^ n22821 ^ n13904 ;
  assign n26431 = ( n426 & n1559 ) | ( n426 & n1589 ) | ( n1559 & n1589 ) ;
  assign n26432 = n26431 ^ n10764 ^ n867 ;
  assign n26433 = n26432 ^ n25932 ^ n6266 ;
  assign n26434 = ( n4003 & n10938 ) | ( n4003 & n26433 ) | ( n10938 & n26433 ) ;
  assign n26435 = ( n1231 & ~n9504 ) | ( n1231 & n14791 ) | ( ~n9504 & n14791 ) ;
  assign n26436 = ( n5422 & n7625 ) | ( n5422 & n10965 ) | ( n7625 & n10965 ) ;
  assign n26437 = n26436 ^ n18355 ^ n15636 ;
  assign n26439 = n18096 ^ n10560 ^ n3742 ;
  assign n26438 = n10693 ^ n2127 ^ n1085 ;
  assign n26440 = n26439 ^ n26438 ^ n11675 ;
  assign n26441 = ( n11362 & ~n13920 ) | ( n11362 & n15825 ) | ( ~n13920 & n15825 ) ;
  assign n26442 = n16308 ^ n4841 ^ n1052 ;
  assign n26443 = n26442 ^ n14566 ^ n13433 ;
  assign n26444 = n14288 ^ n9333 ^ n6757 ;
  assign n26445 = ( n18070 & n26443 ) | ( n18070 & n26444 ) | ( n26443 & n26444 ) ;
  assign n26446 = n11596 ^ n5174 ^ n4662 ;
  assign n26447 = n26446 ^ n22310 ^ n17200 ;
  assign n26448 = n18011 ^ n14262 ^ n6859 ;
  assign n26449 = ( n2694 & ~n9031 ) | ( n2694 & n26448 ) | ( ~n9031 & n26448 ) ;
  assign n26452 = ( x55 & ~n8759 ) | ( x55 & n10999 ) | ( ~n8759 & n10999 ) ;
  assign n26453 = n26452 ^ n13366 ^ n8631 ;
  assign n26454 = n26453 ^ n22687 ^ n6360 ;
  assign n26455 = n26454 ^ n14339 ^ n1643 ;
  assign n26450 = ( n9521 & n20391 ) | ( n9521 & n20614 ) | ( n20391 & n20614 ) ;
  assign n26451 = ( n12965 & ~n18696 ) | ( n12965 & n26450 ) | ( ~n18696 & n26450 ) ;
  assign n26456 = n26455 ^ n26451 ^ n3215 ;
  assign n26457 = n20347 ^ n4829 ^ n2718 ;
  assign n26458 = n10660 ^ n3836 ^ n1165 ;
  assign n26461 = ( n4253 & ~n5029 ) | ( n4253 & n19147 ) | ( ~n5029 & n19147 ) ;
  assign n26460 = ( n718 & n14288 ) | ( n718 & ~n16949 ) | ( n14288 & ~n16949 ) ;
  assign n26459 = ( n4046 & ~n16670 ) | ( n4046 & n23080 ) | ( ~n16670 & n23080 ) ;
  assign n26462 = n26461 ^ n26460 ^ n26459 ;
  assign n26463 = n24242 ^ n17831 ^ n339 ;
  assign n26464 = n8496 ^ n3130 ^ n1960 ;
  assign n26465 = ( n262 & n11136 ) | ( n262 & ~n26464 ) | ( n11136 & ~n26464 ) ;
  assign n26466 = n23141 ^ n19113 ^ n5212 ;
  assign n26467 = ( ~n16936 & n22419 ) | ( ~n16936 & n26466 ) | ( n22419 & n26466 ) ;
  assign n26468 = ( n3297 & n21307 ) | ( n3297 & ~n26467 ) | ( n21307 & ~n26467 ) ;
  assign n26469 = n26468 ^ n6271 ^ n4512 ;
  assign n26470 = ( n2323 & ~n14825 ) | ( n2323 & n14977 ) | ( ~n14825 & n14977 ) ;
  assign n26471 = n24221 ^ n14983 ^ n1223 ;
  assign n26472 = ( ~n22946 & n26470 ) | ( ~n22946 & n26471 ) | ( n26470 & n26471 ) ;
  assign n26473 = ( n4362 & n4585 ) | ( n4362 & ~n9886 ) | ( n4585 & ~n9886 ) ;
  assign n26474 = n20694 ^ n13655 ^ n9251 ;
  assign n26475 = ( n12447 & ~n26473 ) | ( n12447 & n26474 ) | ( ~n26473 & n26474 ) ;
  assign n26476 = n7561 ^ n293 ^ x72 ;
  assign n26477 = n26476 ^ n19778 ^ n7150 ;
  assign n26478 = n26477 ^ n18811 ^ n3178 ;
  assign n26479 = n22080 ^ n17115 ^ n6687 ;
  assign n26480 = n26479 ^ n8830 ^ n8286 ;
  assign n26481 = ( n11980 & n13245 ) | ( n11980 & ~n26480 ) | ( n13245 & ~n26480 ) ;
  assign n26482 = n25003 ^ n11958 ^ n1517 ;
  assign n26483 = n13690 ^ n11364 ^ n6136 ;
  assign n26484 = ( ~n3777 & n10199 ) | ( ~n3777 & n11663 ) | ( n10199 & n11663 ) ;
  assign n26485 = ( n12394 & ~n26483 ) | ( n12394 & n26484 ) | ( ~n26483 & n26484 ) ;
  assign n26486 = ( ~n10383 & n15498 ) | ( ~n10383 & n18409 ) | ( n15498 & n18409 ) ;
  assign n26487 = n12195 ^ n6472 ^ n2260 ;
  assign n26488 = ( n3875 & n6744 ) | ( n3875 & ~n15726 ) | ( n6744 & ~n15726 ) ;
  assign n26489 = n25777 ^ n19190 ^ n3906 ;
  assign n26490 = ( n6678 & n26488 ) | ( n6678 & n26489 ) | ( n26488 & n26489 ) ;
  assign n26493 = ( n3086 & n5342 ) | ( n3086 & ~n7861 ) | ( n5342 & ~n7861 ) ;
  assign n26491 = n10848 ^ n8943 ^ n2209 ;
  assign n26492 = ( n10803 & ~n14133 ) | ( n10803 & n26491 ) | ( ~n14133 & n26491 ) ;
  assign n26494 = n26493 ^ n26492 ^ n24197 ;
  assign n26495 = n26494 ^ n18211 ^ n5978 ;
  assign n26496 = n26495 ^ n22812 ^ n6766 ;
  assign n26497 = n18070 ^ n6340 ^ n5475 ;
  assign n26498 = n26497 ^ n21689 ^ n8047 ;
  assign n26499 = ( n7578 & n18960 ) | ( n7578 & n22944 ) | ( n18960 & n22944 ) ;
  assign n26500 = n26499 ^ n26265 ^ n5380 ;
  assign n26501 = n17039 ^ n12446 ^ n7607 ;
  assign n26502 = n16060 ^ n13751 ^ n4456 ;
  assign n26503 = ( n749 & n2669 ) | ( n749 & ~n5130 ) | ( n2669 & ~n5130 ) ;
  assign n26504 = ( n2758 & n10750 ) | ( n2758 & ~n26503 ) | ( n10750 & ~n26503 ) ;
  assign n26505 = ( n1855 & ~n3263 ) | ( n1855 & n25851 ) | ( ~n3263 & n25851 ) ;
  assign n26506 = ( ~n10124 & n13348 ) | ( ~n10124 & n26505 ) | ( n13348 & n26505 ) ;
  assign n26507 = ( n9391 & n14142 ) | ( n9391 & n26506 ) | ( n14142 & n26506 ) ;
  assign n26508 = ( n803 & n11000 ) | ( n803 & n14313 ) | ( n11000 & n14313 ) ;
  assign n26509 = ( n430 & ~n1381 ) | ( n430 & n4440 ) | ( ~n1381 & n4440 ) ;
  assign n26510 = n26509 ^ n12920 ^ n4751 ;
  assign n26511 = ( n2136 & n10855 ) | ( n2136 & n23329 ) | ( n10855 & n23329 ) ;
  assign n26512 = ( n433 & n6711 ) | ( n433 & ~n26511 ) | ( n6711 & ~n26511 ) ;
  assign n26513 = n22976 ^ n14939 ^ n1545 ;
  assign n26514 = n26513 ^ n4961 ^ n3268 ;
  assign n26515 = ( n10611 & n26512 ) | ( n10611 & n26514 ) | ( n26512 & n26514 ) ;
  assign n26516 = ( n2611 & n7613 ) | ( n2611 & n13371 ) | ( n7613 & n13371 ) ;
  assign n26517 = n8778 ^ n3180 ^ n1921 ;
  assign n26518 = n19094 ^ n4336 ^ n804 ;
  assign n26519 = ( ~n26516 & n26517 ) | ( ~n26516 & n26518 ) | ( n26517 & n26518 ) ;
  assign n26520 = ( n5191 & n8814 ) | ( n5191 & ~n25443 ) | ( n8814 & ~n25443 ) ;
  assign n26521 = ( ~n1577 & n10230 ) | ( ~n1577 & n26520 ) | ( n10230 & n26520 ) ;
  assign n26522 = n14140 ^ n8162 ^ n5282 ;
  assign n26523 = n21707 ^ n13655 ^ n5825 ;
  assign n26524 = ( ~n13897 & n23124 ) | ( ~n13897 & n26523 ) | ( n23124 & n26523 ) ;
  assign n26525 = ( ~n4814 & n18131 ) | ( ~n4814 & n23988 ) | ( n18131 & n23988 ) ;
  assign n26526 = ( n5500 & n19885 ) | ( n5500 & n22034 ) | ( n19885 & n22034 ) ;
  assign n26527 = ( ~n20447 & n21936 ) | ( ~n20447 & n23519 ) | ( n21936 & n23519 ) ;
  assign n26529 = ( ~n6137 & n12954 ) | ( ~n6137 & n14308 ) | ( n12954 & n14308 ) ;
  assign n26528 = n14906 ^ n5990 ^ n3555 ;
  assign n26530 = n26529 ^ n26528 ^ n17578 ;
  assign n26531 = ( ~n7188 & n12870 ) | ( ~n7188 & n20681 ) | ( n12870 & n20681 ) ;
  assign n26532 = ( n8226 & n20834 ) | ( n8226 & n26531 ) | ( n20834 & n26531 ) ;
  assign n26533 = ( n10732 & n11395 ) | ( n10732 & ~n22080 ) | ( n11395 & ~n22080 ) ;
  assign n26534 = ( n1789 & n3936 ) | ( n1789 & n26533 ) | ( n3936 & n26533 ) ;
  assign n26535 = ( ~n9583 & n10455 ) | ( ~n9583 & n21652 ) | ( n10455 & n21652 ) ;
  assign n26536 = n26535 ^ n17880 ^ n4450 ;
  assign n26543 = n9744 ^ n6426 ^ n2865 ;
  assign n26540 = ( ~n2171 & n2570 ) | ( ~n2171 & n9333 ) | ( n2570 & n9333 ) ;
  assign n26541 = n26540 ^ n3745 ^ n1068 ;
  assign n26539 = ( n6833 & ~n22941 ) | ( n6833 & n24896 ) | ( ~n22941 & n24896 ) ;
  assign n26542 = n26541 ^ n26539 ^ n853 ;
  assign n26544 = n26543 ^ n26542 ^ n11769 ;
  assign n26537 = ( n4323 & n9269 ) | ( n4323 & ~n16259 ) | ( n9269 & ~n16259 ) ;
  assign n26538 = n26537 ^ n23031 ^ n3438 ;
  assign n26545 = n26544 ^ n26538 ^ n11479 ;
  assign n26548 = ( n1043 & n5228 ) | ( n1043 & ~n13543 ) | ( n5228 & ~n13543 ) ;
  assign n26547 = ( ~n9073 & n14292 ) | ( ~n9073 & n15869 ) | ( n14292 & n15869 ) ;
  assign n26546 = ( n6442 & n9570 ) | ( n6442 & ~n18689 ) | ( n9570 & ~n18689 ) ;
  assign n26549 = n26548 ^ n26547 ^ n26546 ;
  assign n26550 = ( n172 & n13864 ) | ( n172 & n17744 ) | ( n13864 & n17744 ) ;
  assign n26551 = ( n654 & n2762 ) | ( n654 & n6165 ) | ( n2762 & n6165 ) ;
  assign n26552 = ( n8336 & ~n8675 ) | ( n8336 & n16495 ) | ( ~n8675 & n16495 ) ;
  assign n26553 = ( ~n706 & n9960 ) | ( ~n706 & n18824 ) | ( n9960 & n18824 ) ;
  assign n26554 = ( n1668 & ~n13115 ) | ( n1668 & n26553 ) | ( ~n13115 & n26553 ) ;
  assign n26555 = n14644 ^ n1264 ^ n201 ;
  assign n26556 = ( n12833 & n20906 ) | ( n12833 & ~n26555 ) | ( n20906 & ~n26555 ) ;
  assign n26557 = n22619 ^ n9983 ^ n5195 ;
  assign n26558 = ( n4884 & ~n12215 ) | ( n4884 & n26557 ) | ( ~n12215 & n26557 ) ;
  assign n26559 = n23755 ^ n12513 ^ n4461 ;
  assign n26560 = n22131 ^ n19911 ^ n442 ;
  assign n26561 = ( ~n6402 & n24036 ) | ( ~n6402 & n26560 ) | ( n24036 & n26560 ) ;
  assign n26562 = ( n4760 & ~n18219 ) | ( n4760 & n23060 ) | ( ~n18219 & n23060 ) ;
  assign n26563 = n25727 ^ n11583 ^ n11519 ;
  assign n26564 = ( n5921 & n7025 ) | ( n5921 & ~n11524 ) | ( n7025 & ~n11524 ) ;
  assign n26565 = n10298 ^ n9026 ^ x47 ;
  assign n26566 = ( n18637 & n23086 ) | ( n18637 & ~n26565 ) | ( n23086 & ~n26565 ) ;
  assign n26567 = ( n8818 & ~n17335 ) | ( n8818 & n23955 ) | ( ~n17335 & n23955 ) ;
  assign n26568 = ( n4433 & ~n23901 ) | ( n4433 & n26567 ) | ( ~n23901 & n26567 ) ;
  assign n26569 = ( n20162 & n25748 ) | ( n20162 & n26568 ) | ( n25748 & n26568 ) ;
  assign n26570 = ( n8923 & ~n10042 ) | ( n8923 & n26569 ) | ( ~n10042 & n26569 ) ;
  assign n26571 = n5538 ^ n2885 ^ n1817 ;
  assign n26572 = ( n5101 & n5962 ) | ( n5101 & ~n15135 ) | ( n5962 & ~n15135 ) ;
  assign n26573 = n17335 ^ n15474 ^ n3085 ;
  assign n26574 = ( n26571 & ~n26572 ) | ( n26571 & n26573 ) | ( ~n26572 & n26573 ) ;
  assign n26575 = n18951 ^ n10159 ^ n8079 ;
  assign n26576 = n26575 ^ n16778 ^ n14643 ;
  assign n26577 = ( n3437 & n5581 ) | ( n3437 & ~n26576 ) | ( n5581 & ~n26576 ) ;
  assign n26578 = n26577 ^ n22457 ^ n5653 ;
  assign n26579 = ( ~n1974 & n12586 ) | ( ~n1974 & n26578 ) | ( n12586 & n26578 ) ;
  assign n26580 = n24516 ^ n16635 ^ n7621 ;
  assign n26581 = ( n4651 & n7732 ) | ( n4651 & ~n26580 ) | ( n7732 & ~n26580 ) ;
  assign n26582 = n21955 ^ n6688 ^ n1341 ;
  assign n26586 = n19106 ^ n6410 ^ n5119 ;
  assign n26585 = ( ~n2000 & n7132 ) | ( ~n2000 & n13934 ) | ( n7132 & n13934 ) ;
  assign n26583 = ( n6573 & n7408 ) | ( n6573 & n8352 ) | ( n7408 & n8352 ) ;
  assign n26584 = ( n8660 & n18499 ) | ( n8660 & n26583 ) | ( n18499 & n26583 ) ;
  assign n26587 = n26586 ^ n26585 ^ n26584 ;
  assign n26588 = ( ~n3319 & n21283 ) | ( ~n3319 & n26587 ) | ( n21283 & n26587 ) ;
  assign n26589 = ( n2664 & n10418 ) | ( n2664 & n25586 ) | ( n10418 & n25586 ) ;
  assign n26590 = n22566 ^ n11843 ^ n1462 ;
  assign n26591 = n25560 ^ n12053 ^ n8117 ;
  assign n26592 = n7464 ^ n4496 ^ n2095 ;
  assign n26593 = ( n23826 & n26591 ) | ( n23826 & n26592 ) | ( n26591 & n26592 ) ;
  assign n26594 = n26568 ^ n23559 ^ n16238 ;
  assign n26595 = ( ~n496 & n2540 ) | ( ~n496 & n7875 ) | ( n2540 & n7875 ) ;
  assign n26596 = n20439 ^ n16735 ^ n4162 ;
  assign n26597 = n26596 ^ n16436 ^ n1638 ;
  assign n26598 = n22198 ^ n17530 ^ n10496 ;
  assign n26599 = ( n1634 & n2313 ) | ( n1634 & ~n9910 ) | ( n2313 & ~n9910 ) ;
  assign n26600 = ( n16202 & ~n24129 ) | ( n16202 & n26599 ) | ( ~n24129 & n26599 ) ;
  assign n26601 = n26600 ^ n24478 ^ n4397 ;
  assign n26602 = n26601 ^ n20402 ^ n15382 ;
  assign n26603 = ( n13330 & n13596 ) | ( n13330 & n21409 ) | ( n13596 & n21409 ) ;
  assign n26604 = ( n7219 & ~n12018 ) | ( n7219 & n26603 ) | ( ~n12018 & n26603 ) ;
  assign n26605 = ( n18746 & n23563 ) | ( n18746 & n26604 ) | ( n23563 & n26604 ) ;
  assign n26606 = ( n2048 & n13203 ) | ( n2048 & ~n25197 ) | ( n13203 & ~n25197 ) ;
  assign n26607 = n26606 ^ n6505 ^ n4576 ;
  assign n26608 = n16634 ^ n7517 ^ n2301 ;
  assign n26609 = ( ~n5802 & n14235 ) | ( ~n5802 & n15269 ) | ( n14235 & n15269 ) ;
  assign n26610 = n8161 ^ n5696 ^ n5361 ;
  assign n26611 = ( n9791 & n26573 ) | ( n9791 & n26610 ) | ( n26573 & n26610 ) ;
  assign n26612 = ( ~n11118 & n23835 ) | ( ~n11118 & n26611 ) | ( n23835 & n26611 ) ;
  assign n26613 = ( n5060 & ~n26609 ) | ( n5060 & n26612 ) | ( ~n26609 & n26612 ) ;
  assign n26614 = n15601 ^ n3684 ^ n3287 ;
  assign n26615 = ( n13781 & n15923 ) | ( n13781 & n26614 ) | ( n15923 & n26614 ) ;
  assign n26616 = ( n3771 & n7533 ) | ( n3771 & n23721 ) | ( n7533 & n23721 ) ;
  assign n26617 = ( n12256 & ~n13418 ) | ( n12256 & n14510 ) | ( ~n13418 & n14510 ) ;
  assign n26618 = n26617 ^ n22992 ^ n17241 ;
  assign n26619 = n26476 ^ n15398 ^ n2029 ;
  assign n26620 = n26619 ^ n22956 ^ n5280 ;
  assign n26621 = n19715 ^ n8634 ^ n4582 ;
  assign n26622 = ( n14422 & n24598 ) | ( n14422 & n26621 ) | ( n24598 & n26621 ) ;
  assign n26623 = n3219 ^ n3212 ^ n2212 ;
  assign n26624 = n26623 ^ n17335 ^ x42 ;
  assign n26625 = n13161 ^ n9936 ^ n7319 ;
  assign n26626 = ( n4855 & n5761 ) | ( n4855 & n12845 ) | ( n5761 & n12845 ) ;
  assign n26627 = ( n1294 & n11936 ) | ( n1294 & ~n20960 ) | ( n11936 & ~n20960 ) ;
  assign n26628 = ( n6691 & ~n10119 ) | ( n6691 & n26627 ) | ( ~n10119 & n26627 ) ;
  assign n26629 = n26026 ^ n12566 ^ n6971 ;
  assign n26630 = ( n8609 & n11663 ) | ( n8609 & n26629 ) | ( n11663 & n26629 ) ;
  assign n26633 = n10092 ^ n8007 ^ n860 ;
  assign n26634 = n26633 ^ n17939 ^ n381 ;
  assign n26631 = n22202 ^ n7006 ^ n3773 ;
  assign n26632 = ( n7112 & n12334 ) | ( n7112 & ~n26631 ) | ( n12334 & ~n26631 ) ;
  assign n26635 = n26634 ^ n26632 ^ n7603 ;
  assign n26636 = ( ~n350 & n12684 ) | ( ~n350 & n20997 ) | ( n12684 & n20997 ) ;
  assign n26637 = n8348 ^ n5193 ^ n1220 ;
  assign n26638 = n26637 ^ n19747 ^ n9469 ;
  assign n26639 = ( n13006 & n14043 ) | ( n13006 & n26638 ) | ( n14043 & n26638 ) ;
  assign n26640 = n11462 ^ n7600 ^ x14 ;
  assign n26641 = ( n14197 & ~n17231 ) | ( n14197 & n26640 ) | ( ~n17231 & n26640 ) ;
  assign n26642 = n16078 ^ n10543 ^ n2935 ;
  assign n26643 = ( ~n3103 & n11107 ) | ( ~n3103 & n24362 ) | ( n11107 & n24362 ) ;
  assign n26644 = ( ~n617 & n2817 ) | ( ~n617 & n26643 ) | ( n2817 & n26643 ) ;
  assign n26645 = ( ~n7149 & n26642 ) | ( ~n7149 & n26644 ) | ( n26642 & n26644 ) ;
  assign n26646 = n26645 ^ n22270 ^ n2838 ;
  assign n26647 = n26646 ^ n7863 ^ n3948 ;
  assign n26648 = ( n26639 & n26641 ) | ( n26639 & n26647 ) | ( n26641 & n26647 ) ;
  assign n26649 = n22968 ^ n19305 ^ n9983 ;
  assign n26650 = ( ~n2617 & n6458 ) | ( ~n2617 & n16687 ) | ( n6458 & n16687 ) ;
  assign n26651 = n26650 ^ n6892 ^ n6137 ;
  assign n26652 = ( n2146 & ~n23802 ) | ( n2146 & n26651 ) | ( ~n23802 & n26651 ) ;
  assign n26653 = ( n1986 & ~n8498 ) | ( n1986 & n14949 ) | ( ~n8498 & n14949 ) ;
  assign n26654 = ( ~n8090 & n10994 ) | ( ~n8090 & n26653 ) | ( n10994 & n26653 ) ;
  assign n26655 = n16329 ^ n8933 ^ n8135 ;
  assign n26656 = ( n276 & n6609 ) | ( n276 & ~n26655 ) | ( n6609 & ~n26655 ) ;
  assign n26657 = n17460 ^ n11019 ^ n6912 ;
  assign n26658 = n6440 ^ n4555 ^ n1915 ;
  assign n26659 = ( n18406 & n26657 ) | ( n18406 & n26658 ) | ( n26657 & n26658 ) ;
  assign n26660 = ( n1983 & n3877 ) | ( n1983 & n3985 ) | ( n3877 & n3985 ) ;
  assign n26661 = n26660 ^ n2745 ^ n2404 ;
  assign n26662 = n18069 ^ n7923 ^ n3394 ;
  assign n26663 = ( n4678 & ~n10471 ) | ( n4678 & n20903 ) | ( ~n10471 & n20903 ) ;
  assign n26664 = ( n1197 & n6277 ) | ( n1197 & n14554 ) | ( n6277 & n14554 ) ;
  assign n26665 = ( ~x18 & n620 ) | ( ~x18 & n10828 ) | ( n620 & n10828 ) ;
  assign n26666 = ( ~n854 & n3619 ) | ( ~n854 & n18314 ) | ( n3619 & n18314 ) ;
  assign n26667 = n26666 ^ n14513 ^ n5018 ;
  assign n26668 = n26667 ^ n18732 ^ n8411 ;
  assign n26669 = ( ~n22021 & n26665 ) | ( ~n22021 & n26668 ) | ( n26665 & n26668 ) ;
  assign n26670 = n21994 ^ n18869 ^ n4272 ;
  assign n26671 = ( n7561 & n23322 ) | ( n7561 & n26670 ) | ( n23322 & n26670 ) ;
  assign n26672 = ( n5900 & n7402 ) | ( n5900 & ~n14637 ) | ( n7402 & ~n14637 ) ;
  assign n26673 = ( n583 & n1952 ) | ( n583 & n21132 ) | ( n1952 & n21132 ) ;
  assign n26674 = n26673 ^ n23225 ^ n5943 ;
  assign n26675 = ( n1860 & n26672 ) | ( n1860 & n26674 ) | ( n26672 & n26674 ) ;
  assign n26676 = ( n7573 & ~n13152 ) | ( n7573 & n13553 ) | ( ~n13152 & n13553 ) ;
  assign n26677 = ( n20713 & ~n24565 ) | ( n20713 & n26676 ) | ( ~n24565 & n26676 ) ;
  assign n26678 = n9707 ^ n8160 ^ n971 ;
  assign n26679 = ( n7974 & n10821 ) | ( n7974 & ~n10882 ) | ( n10821 & ~n10882 ) ;
  assign n26680 = n26679 ^ n22908 ^ n3508 ;
  assign n26681 = n23829 ^ n22823 ^ n5577 ;
  assign n26682 = n13243 ^ n5330 ^ n4248 ;
  assign n26683 = ( n13005 & n24335 ) | ( n13005 & ~n26682 ) | ( n24335 & ~n26682 ) ;
  assign n26684 = ( ~n13379 & n18268 ) | ( ~n13379 & n25952 ) | ( n18268 & n25952 ) ;
  assign n26685 = ( n9031 & n14779 ) | ( n9031 & ~n26684 ) | ( n14779 & ~n26684 ) ;
  assign n26686 = ( n448 & n14928 ) | ( n448 & n26685 ) | ( n14928 & n26685 ) ;
  assign n26687 = ( n3531 & n9865 ) | ( n3531 & ~n22138 ) | ( n9865 & ~n22138 ) ;
  assign n26688 = ( ~n2090 & n4493 ) | ( ~n2090 & n7586 ) | ( n4493 & n7586 ) ;
  assign n26689 = ( ~n1240 & n3557 ) | ( ~n1240 & n25852 ) | ( n3557 & n25852 ) ;
  assign n26690 = ( n3614 & ~n8620 ) | ( n3614 & n21125 ) | ( ~n8620 & n21125 ) ;
  assign n26691 = n26690 ^ n20020 ^ n14882 ;
  assign n26692 = ( n10727 & n23157 ) | ( n10727 & ~n23359 ) | ( n23157 & ~n23359 ) ;
  assign n26693 = ( ~n2209 & n10068 ) | ( ~n2209 & n11045 ) | ( n10068 & n11045 ) ;
  assign n26694 = n26693 ^ n12518 ^ n7201 ;
  assign n26695 = ( n2975 & ~n4612 ) | ( n2975 & n26694 ) | ( ~n4612 & n26694 ) ;
  assign n26696 = ( n6343 & ~n6926 ) | ( n6343 & n10649 ) | ( ~n6926 & n10649 ) ;
  assign n26697 = n14602 ^ n3907 ^ n2253 ;
  assign n26698 = ( ~n6859 & n15179 ) | ( ~n6859 & n26697 ) | ( n15179 & n26697 ) ;
  assign n26699 = ( ~n2496 & n9285 ) | ( ~n2496 & n26118 ) | ( n9285 & n26118 ) ;
  assign n26700 = n26699 ^ n19115 ^ n6765 ;
  assign n26701 = ( ~n10666 & n26698 ) | ( ~n10666 & n26700 ) | ( n26698 & n26700 ) ;
  assign n26702 = n20478 ^ n7471 ^ n3031 ;
  assign n26703 = n26702 ^ n20416 ^ n4124 ;
  assign n26704 = ( n3502 & n3791 ) | ( n3502 & ~n15201 ) | ( n3791 & ~n15201 ) ;
  assign n26705 = n26704 ^ n7175 ^ n1289 ;
  assign n26706 = ( n3666 & n6569 ) | ( n3666 & ~n17876 ) | ( n6569 & ~n17876 ) ;
  assign n26707 = n26706 ^ n24380 ^ n9606 ;
  assign n26708 = n26707 ^ n23738 ^ n19202 ;
  assign n26709 = ( n6869 & ~n25807 ) | ( n6869 & n26708 ) | ( ~n25807 & n26708 ) ;
  assign n26710 = ( n2290 & ~n4511 ) | ( n2290 & n19788 ) | ( ~n4511 & n19788 ) ;
  assign n26711 = ( n5733 & ~n9711 ) | ( n5733 & n13935 ) | ( ~n9711 & n13935 ) ;
  assign n26712 = n26711 ^ n24216 ^ n533 ;
  assign n26713 = ( n2239 & n26710 ) | ( n2239 & ~n26712 ) | ( n26710 & ~n26712 ) ;
  assign n26714 = n26713 ^ n26658 ^ n454 ;
  assign n26715 = n26714 ^ n11689 ^ n6372 ;
  assign n26716 = ( n802 & ~n10427 ) | ( n802 & n15089 ) | ( ~n10427 & n15089 ) ;
  assign n26717 = n26716 ^ n16874 ^ n16488 ;
  assign n26719 = n22645 ^ n19431 ^ n1881 ;
  assign n26718 = n13468 ^ n12705 ^ n1946 ;
  assign n26720 = n26719 ^ n26718 ^ n11652 ;
  assign n26721 = ( n11568 & ~n12819 ) | ( n11568 & n14180 ) | ( ~n12819 & n14180 ) ;
  assign n26722 = ( n814 & n15487 ) | ( n814 & n26721 ) | ( n15487 & n26721 ) ;
  assign n26723 = n23786 ^ n22861 ^ n20801 ;
  assign n26724 = n11214 ^ n3213 ^ n322 ;
  assign n26725 = ( n4813 & ~n16460 ) | ( n4813 & n26724 ) | ( ~n16460 & n26724 ) ;
  assign n26726 = n26725 ^ n24748 ^ n11481 ;
  assign n26727 = n22495 ^ n10007 ^ n1461 ;
  assign n26728 = ( ~n1245 & n6856 ) | ( ~n1245 & n13411 ) | ( n6856 & n13411 ) ;
  assign n26729 = n26728 ^ n11101 ^ n817 ;
  assign n26730 = n26729 ^ n23280 ^ n15326 ;
  assign n26731 = ( n14109 & n21211 ) | ( n14109 & ~n23904 ) | ( n21211 & ~n23904 ) ;
  assign n26732 = ( n528 & n2829 ) | ( n528 & ~n13976 ) | ( n2829 & ~n13976 ) ;
  assign n26733 = ( ~n2948 & n5484 ) | ( ~n2948 & n13496 ) | ( n5484 & n13496 ) ;
  assign n26734 = n14501 ^ n8298 ^ n3221 ;
  assign n26735 = n26734 ^ n19638 ^ n19467 ;
  assign n26736 = n26735 ^ n23572 ^ n5833 ;
  assign n26737 = ( n2067 & n9923 ) | ( n2067 & ~n12926 ) | ( n9923 & ~n12926 ) ;
  assign n26738 = ( n1244 & ~n14931 ) | ( n1244 & n23473 ) | ( ~n14931 & n23473 ) ;
  assign n26739 = n17025 ^ n5569 ^ n3650 ;
  assign n26740 = ( ~n5944 & n13503 ) | ( ~n5944 & n16981 ) | ( n13503 & n16981 ) ;
  assign n26741 = ( n3219 & n6784 ) | ( n3219 & ~n10526 ) | ( n6784 & ~n10526 ) ;
  assign n26742 = ( ~n11329 & n15742 ) | ( ~n11329 & n26741 ) | ( n15742 & n26741 ) ;
  assign n26743 = n26742 ^ n21460 ^ n1612 ;
  assign n26744 = n4070 ^ n2937 ^ n1165 ;
  assign n26745 = n26744 ^ n12780 ^ n10550 ;
  assign n26746 = ( n8615 & ~n12992 ) | ( n8615 & n23349 ) | ( ~n12992 & n23349 ) ;
  assign n26747 = n10997 ^ n2061 ^ n357 ;
  assign n26748 = n26747 ^ n20683 ^ n7475 ;
  assign n26749 = n26748 ^ n22538 ^ n8176 ;
  assign n26750 = n6020 ^ n4955 ^ n1790 ;
  assign n26751 = ( n8309 & ~n9040 ) | ( n8309 & n26750 ) | ( ~n9040 & n26750 ) ;
  assign n26752 = n26751 ^ n23562 ^ n497 ;
  assign n26753 = ( ~n11777 & n25173 ) | ( ~n11777 & n25884 ) | ( n25173 & n25884 ) ;
  assign n26754 = n8339 ^ n5415 ^ n4680 ;
  assign n26755 = n16337 ^ n11872 ^ n1019 ;
  assign n26756 = ( n12184 & n12329 ) | ( n12184 & ~n17965 ) | ( n12329 & ~n17965 ) ;
  assign n26757 = ( ~n12805 & n24726 ) | ( ~n12805 & n26756 ) | ( n24726 & n26756 ) ;
  assign n26758 = ( n3178 & n12131 ) | ( n3178 & n21153 ) | ( n12131 & n21153 ) ;
  assign n26759 = n5580 ^ n4280 ^ n1573 ;
  assign n26760 = n26759 ^ n14142 ^ n11002 ;
  assign n26763 = ( n2386 & n2583 ) | ( n2386 & n18007 ) | ( n2583 & n18007 ) ;
  assign n26761 = ( ~n5945 & n8922 ) | ( ~n5945 & n11125 ) | ( n8922 & n11125 ) ;
  assign n26762 = ( n4989 & n11363 ) | ( n4989 & ~n26761 ) | ( n11363 & ~n26761 ) ;
  assign n26764 = n26763 ^ n26762 ^ n5889 ;
  assign n26765 = ( n1663 & ~n3433 ) | ( n1663 & n9966 ) | ( ~n3433 & n9966 ) ;
  assign n26766 = ( n732 & ~n7792 ) | ( n732 & n23058 ) | ( ~n7792 & n23058 ) ;
  assign n26767 = n26766 ^ n9843 ^ n3480 ;
  assign n26768 = ( n1354 & n5285 ) | ( n1354 & ~n8226 ) | ( n5285 & ~n8226 ) ;
  assign n26769 = ( ~n9626 & n15429 ) | ( ~n9626 & n25492 ) | ( n15429 & n25492 ) ;
  assign n26773 = n7020 ^ n3567 ^ n3229 ;
  assign n26771 = n23060 ^ n6835 ^ n6172 ;
  assign n26772 = n26771 ^ n14694 ^ n4869 ;
  assign n26770 = ( n17776 & n19857 ) | ( n17776 & n20733 ) | ( n19857 & n20733 ) ;
  assign n26774 = n26773 ^ n26772 ^ n26770 ;
  assign n26775 = n16613 ^ n10009 ^ n2481 ;
  assign n26776 = n26775 ^ n20919 ^ n15081 ;
  assign n26777 = n11250 ^ n8923 ^ n2102 ;
  assign n26778 = n26777 ^ n4366 ^ n1879 ;
  assign n26779 = ( ~n5549 & n23597 ) | ( ~n5549 & n26778 ) | ( n23597 & n26778 ) ;
  assign n26780 = ( n12585 & n19965 ) | ( n12585 & ~n26779 ) | ( n19965 & ~n26779 ) ;
  assign n26781 = ( ~n6897 & n9000 ) | ( ~n6897 & n10127 ) | ( n9000 & n10127 ) ;
  assign n26782 = ( n945 & n12485 ) | ( n945 & n26781 ) | ( n12485 & n26781 ) ;
  assign n26783 = n22696 ^ n12427 ^ n3970 ;
  assign n26784 = ( n534 & ~n11245 ) | ( n534 & n26783 ) | ( ~n11245 & n26783 ) ;
  assign n26785 = ( n16256 & ~n20695 ) | ( n16256 & n26784 ) | ( ~n20695 & n26784 ) ;
  assign n26786 = n22215 ^ n16752 ^ n1928 ;
  assign n26787 = n7273 ^ n5583 ^ n4376 ;
  assign n26788 = n10861 ^ n7831 ^ n6693 ;
  assign n26789 = ( n13980 & n24436 ) | ( n13980 & n26788 ) | ( n24436 & n26788 ) ;
  assign n26790 = ( ~n24199 & n26787 ) | ( ~n24199 & n26789 ) | ( n26787 & n26789 ) ;
  assign n26791 = ( ~n19307 & n26786 ) | ( ~n19307 & n26790 ) | ( n26786 & n26790 ) ;
  assign n26792 = ( n17221 & n19492 ) | ( n17221 & n26476 ) | ( n19492 & n26476 ) ;
  assign n26793 = ( n1193 & n3660 ) | ( n1193 & n13350 ) | ( n3660 & n13350 ) ;
  assign n26794 = n10484 ^ n6491 ^ n2614 ;
  assign n26795 = n26794 ^ n11466 ^ n7820 ;
  assign n26796 = n19226 ^ n10089 ^ n3542 ;
  assign n26799 = ( n1131 & ~n3295 ) | ( n1131 & n10430 ) | ( ~n3295 & n10430 ) ;
  assign n26797 = ( ~n202 & n2785 ) | ( ~n202 & n5835 ) | ( n2785 & n5835 ) ;
  assign n26798 = n26797 ^ n6282 ^ n5123 ;
  assign n26800 = n26799 ^ n26798 ^ n14331 ;
  assign n26801 = ( n8380 & n11898 ) | ( n8380 & n13764 ) | ( n11898 & n13764 ) ;
  assign n26802 = n5051 ^ n4261 ^ n2117 ;
  assign n26803 = ( n13801 & ~n23944 ) | ( n13801 & n26802 ) | ( ~n23944 & n26802 ) ;
  assign n26804 = n17956 ^ n9262 ^ n3702 ;
  assign n26805 = ( n5696 & n6444 ) | ( n5696 & n26804 ) | ( n6444 & n26804 ) ;
  assign n26806 = ( n7847 & n10659 ) | ( n7847 & ~n26805 ) | ( n10659 & ~n26805 ) ;
  assign n26807 = n26806 ^ n24166 ^ n9376 ;
  assign n26808 = ( n11568 & ~n12171 ) | ( n11568 & n26807 ) | ( ~n12171 & n26807 ) ;
  assign n26809 = n26808 ^ n25595 ^ n1012 ;
  assign n26810 = ( n3982 & n16676 ) | ( n3982 & ~n26809 ) | ( n16676 & ~n26809 ) ;
  assign n26812 = ( n5933 & ~n6195 ) | ( n5933 & n9524 ) | ( ~n6195 & n9524 ) ;
  assign n26811 = n9436 ^ n9186 ^ n7034 ;
  assign n26813 = n26812 ^ n26811 ^ n19936 ;
  assign n26814 = ( n574 & n4299 ) | ( n574 & ~n10588 ) | ( n4299 & ~n10588 ) ;
  assign n26815 = n26814 ^ n23947 ^ n2145 ;
  assign n26816 = n8690 ^ n5010 ^ n3714 ;
  assign n26817 = ( n5622 & n20174 ) | ( n5622 & ~n26816 ) | ( n20174 & ~n26816 ) ;
  assign n26818 = ( n12645 & n20832 ) | ( n12645 & n21766 ) | ( n20832 & n21766 ) ;
  assign n26819 = n26818 ^ n8387 ^ n3767 ;
  assign n26822 = n20091 ^ n17154 ^ n8739 ;
  assign n26820 = ( n3245 & n14618 ) | ( n3245 & n15881 ) | ( n14618 & n15881 ) ;
  assign n26821 = ( n2194 & n15528 ) | ( n2194 & n26820 ) | ( n15528 & n26820 ) ;
  assign n26823 = n26822 ^ n26821 ^ n22903 ;
  assign n26824 = n24036 ^ n15383 ^ n5143 ;
  assign n26825 = ( n7393 & n13490 ) | ( n7393 & n15640 ) | ( n13490 & n15640 ) ;
  assign n26826 = ( n10172 & ~n26824 ) | ( n10172 & n26825 ) | ( ~n26824 & n26825 ) ;
  assign n26827 = ( ~n1328 & n2247 ) | ( ~n1328 & n21070 ) | ( n2247 & n21070 ) ;
  assign n26828 = ( n5225 & n12186 ) | ( n5225 & n26827 ) | ( n12186 & n26827 ) ;
  assign n26829 = ( n4441 & n13161 ) | ( n4441 & ~n19453 ) | ( n13161 & ~n19453 ) ;
  assign n26830 = n26829 ^ n26029 ^ n939 ;
  assign n26831 = n19962 ^ n10072 ^ n1143 ;
  assign n26832 = n20479 ^ n17206 ^ n1809 ;
  assign n26833 = ( n3396 & n26831 ) | ( n3396 & n26832 ) | ( n26831 & n26832 ) ;
  assign n26834 = ( ~n8868 & n10745 ) | ( ~n8868 & n19797 ) | ( n10745 & n19797 ) ;
  assign n26835 = n26834 ^ n9624 ^ n1814 ;
  assign n26836 = ( n2355 & ~n4691 ) | ( n2355 & n10013 ) | ( ~n4691 & n10013 ) ;
  assign n26837 = n26836 ^ n21624 ^ x73 ;
  assign n26838 = n5006 ^ n3336 ^ n1431 ;
  assign n26840 = ( ~n11193 & n18527 ) | ( ~n11193 & n25952 ) | ( n18527 & n25952 ) ;
  assign n26839 = n18434 ^ n7143 ^ n6200 ;
  assign n26841 = n26840 ^ n26839 ^ n8434 ;
  assign n26842 = ( n25147 & n26838 ) | ( n25147 & n26841 ) | ( n26838 & n26841 ) ;
  assign n26843 = n24296 ^ n20103 ^ n3431 ;
  assign n26844 = ( n8194 & n9057 ) | ( n8194 & n14134 ) | ( n9057 & n14134 ) ;
  assign n26845 = n7326 ^ n1371 ^ n430 ;
  assign n26846 = ( n4109 & n6369 ) | ( n4109 & ~n10410 ) | ( n6369 & ~n10410 ) ;
  assign n26847 = ( ~n4346 & n26845 ) | ( ~n4346 & n26846 ) | ( n26845 & n26846 ) ;
  assign n26848 = ( n9733 & ~n9963 ) | ( n9733 & n26847 ) | ( ~n9963 & n26847 ) ;
  assign n26849 = n10464 ^ n10384 ^ n6649 ;
  assign n26850 = ( ~n4497 & n6426 ) | ( ~n4497 & n26849 ) | ( n6426 & n26849 ) ;
  assign n26851 = ( n8432 & ~n11705 ) | ( n8432 & n26850 ) | ( ~n11705 & n26850 ) ;
  assign n26852 = n12785 ^ n2494 ^ n2419 ;
  assign n26853 = ( n1492 & n7953 ) | ( n1492 & ~n26852 ) | ( n7953 & ~n26852 ) ;
  assign n26854 = ( n19572 & ~n19824 ) | ( n19572 & n20863 ) | ( ~n19824 & n20863 ) ;
  assign n26855 = n26854 ^ n20011 ^ n12723 ;
  assign n26856 = ( ~n8368 & n10811 ) | ( ~n8368 & n22163 ) | ( n10811 & n22163 ) ;
  assign n26857 = ( n9731 & ~n14535 ) | ( n9731 & n26856 ) | ( ~n14535 & n26856 ) ;
  assign n26859 = ( n2309 & ~n4101 ) | ( n2309 & n9336 ) | ( ~n4101 & n9336 ) ;
  assign n26858 = n25341 ^ n16912 ^ n7471 ;
  assign n26860 = n26859 ^ n26858 ^ n8294 ;
  assign n26861 = n26860 ^ n8025 ^ n524 ;
  assign n26862 = ( n2871 & n4238 ) | ( n2871 & n15308 ) | ( n4238 & n15308 ) ;
  assign n26863 = ( n2890 & n5627 ) | ( n2890 & ~n26862 ) | ( n5627 & ~n26862 ) ;
  assign n26864 = n11869 ^ n10663 ^ n7422 ;
  assign n26865 = n26864 ^ n14331 ^ n10741 ;
  assign n26866 = ( ~n391 & n5670 ) | ( ~n391 & n8858 ) | ( n5670 & n8858 ) ;
  assign n26867 = ( n3190 & n7447 ) | ( n3190 & n26866 ) | ( n7447 & n26866 ) ;
  assign n26868 = n26867 ^ n16276 ^ n2036 ;
  assign n26869 = n10940 ^ n4611 ^ n1432 ;
  assign n26870 = n26869 ^ n11004 ^ n3274 ;
  assign n26871 = ( n7741 & ~n21124 ) | ( n7741 & n21380 ) | ( ~n21124 & n21380 ) ;
  assign n26872 = ( n1470 & n9153 ) | ( n1470 & ~n26871 ) | ( n9153 & ~n26871 ) ;
  assign n26873 = ( ~n13851 & n26870 ) | ( ~n13851 & n26872 ) | ( n26870 & n26872 ) ;
  assign n26874 = ( ~n5166 & n9838 ) | ( ~n5166 & n11154 ) | ( n9838 & n11154 ) ;
  assign n26875 = n26874 ^ n13914 ^ n7472 ;
  assign n26876 = n26875 ^ n1334 ^ n1092 ;
  assign n26877 = ( n8334 & ~n13340 ) | ( n8334 & n26876 ) | ( ~n13340 & n26876 ) ;
  assign n26878 = n21670 ^ n9200 ^ n7280 ;
  assign n26879 = ( ~n6371 & n14641 ) | ( ~n6371 & n15924 ) | ( n14641 & n15924 ) ;
  assign n26880 = n26879 ^ n21589 ^ n3774 ;
  assign n26881 = ( n2508 & n9204 ) | ( n2508 & n10974 ) | ( n9204 & n10974 ) ;
  assign n26882 = n26881 ^ n24296 ^ n16789 ;
  assign n26883 = n9731 ^ n6176 ^ n277 ;
  assign n26884 = ( n4704 & n11970 ) | ( n4704 & ~n26883 ) | ( n11970 & ~n26883 ) ;
  assign n26885 = ( n6047 & n9894 ) | ( n6047 & ~n26884 ) | ( n9894 & ~n26884 ) ;
  assign n26886 = n21253 ^ n12279 ^ n1391 ;
  assign n26888 = n14901 ^ n9399 ^ n2414 ;
  assign n26889 = n16313 ^ n5741 ^ n3316 ;
  assign n26890 = ( n10549 & n26888 ) | ( n10549 & ~n26889 ) | ( n26888 & ~n26889 ) ;
  assign n26887 = n19272 ^ n12796 ^ n3299 ;
  assign n26891 = n26890 ^ n26887 ^ n6593 ;
  assign n26892 = n22740 ^ n10937 ^ n7869 ;
  assign n26893 = n13560 ^ n1174 ^ n381 ;
  assign n26894 = ( n8149 & n13521 ) | ( n8149 & n26893 ) | ( n13521 & n26893 ) ;
  assign n26895 = ( n7485 & ~n15062 ) | ( n7485 & n16586 ) | ( ~n15062 & n16586 ) ;
  assign n26896 = n10823 ^ n9936 ^ n2809 ;
  assign n26897 = ( n1345 & n5720 ) | ( n1345 & ~n8901 ) | ( n5720 & ~n8901 ) ;
  assign n26898 = n15614 ^ n11088 ^ n2190 ;
  assign n26899 = n26898 ^ n25292 ^ n3699 ;
  assign n26900 = n26899 ^ n16596 ^ n11380 ;
  assign n26904 = ( ~n6681 & n6738 ) | ( ~n6681 & n9109 ) | ( n6738 & n9109 ) ;
  assign n26905 = ( n7631 & ~n10843 ) | ( n7631 & n26904 ) | ( ~n10843 & n26904 ) ;
  assign n26901 = n25692 ^ n8542 ^ n5245 ;
  assign n26902 = ( n960 & ~n4653 ) | ( n960 & n26901 ) | ( ~n4653 & n26901 ) ;
  assign n26903 = n26902 ^ n23185 ^ n21071 ;
  assign n26906 = n26905 ^ n26903 ^ n1454 ;
  assign n26909 = ( ~n11001 & n15652 ) | ( ~n11001 & n16412 ) | ( n15652 & n16412 ) ;
  assign n26910 = n26909 ^ n12657 ^ n12112 ;
  assign n26907 = n19066 ^ n11672 ^ n9300 ;
  assign n26908 = ( n11383 & ~n12834 ) | ( n11383 & n26907 ) | ( ~n12834 & n26907 ) ;
  assign n26911 = n26910 ^ n26908 ^ n13887 ;
  assign n26912 = ( ~n1819 & n7725 ) | ( ~n1819 & n23363 ) | ( n7725 & n23363 ) ;
  assign n26913 = n23532 ^ n22195 ^ n17508 ;
  assign n26914 = n26913 ^ n22432 ^ n3060 ;
  assign n26915 = ( n13951 & n21498 ) | ( n13951 & n26660 ) | ( n21498 & n26660 ) ;
  assign n26916 = n18253 ^ n17593 ^ n7787 ;
  assign n26917 = ( n18146 & ~n18581 ) | ( n18146 & n24280 ) | ( ~n18581 & n24280 ) ;
  assign n26918 = n23022 ^ n18157 ^ n6408 ;
  assign n26920 = ( n1525 & ~n6362 ) | ( n1525 & n15201 ) | ( ~n6362 & n15201 ) ;
  assign n26919 = n20045 ^ n16726 ^ n8759 ;
  assign n26921 = n26920 ^ n26919 ^ n2425 ;
  assign n26922 = n13586 ^ n9568 ^ n1236 ;
  assign n26925 = ( n5855 & ~n5880 ) | ( n5855 & n9045 ) | ( ~n5880 & n9045 ) ;
  assign n26923 = ( n9166 & n9283 ) | ( n9166 & n13339 ) | ( n9283 & n13339 ) ;
  assign n26924 = n26923 ^ n9144 ^ n3885 ;
  assign n26926 = n26925 ^ n26924 ^ n9658 ;
  assign n26927 = ( n3627 & n11006 ) | ( n3627 & ~n26389 ) | ( n11006 & ~n26389 ) ;
  assign n26929 = n7613 ^ n7149 ^ n2924 ;
  assign n26928 = n23422 ^ n21102 ^ n6816 ;
  assign n26930 = n26929 ^ n26928 ^ n26180 ;
  assign n26931 = ( n1289 & n1389 ) | ( n1289 & n15378 ) | ( n1389 & n15378 ) ;
  assign n26932 = ( x64 & n14049 ) | ( x64 & n17093 ) | ( n14049 & n17093 ) ;
  assign n26933 = ( n11246 & ~n26931 ) | ( n11246 & n26932 ) | ( ~n26931 & n26932 ) ;
  assign n26934 = n7083 ^ n1889 ^ n327 ;
  assign n26935 = ( n7267 & ~n22286 ) | ( n7267 & n26934 ) | ( ~n22286 & n26934 ) ;
  assign n26936 = n20283 ^ n19659 ^ n1521 ;
  assign n26937 = ( ~n7866 & n18797 ) | ( ~n7866 & n26936 ) | ( n18797 & n26936 ) ;
  assign n26938 = ( n8950 & n12649 ) | ( n8950 & ~n26937 ) | ( n12649 & ~n26937 ) ;
  assign n26939 = n14837 ^ n11251 ^ n3730 ;
  assign n26940 = ( n12154 & ~n18408 ) | ( n12154 & n26939 ) | ( ~n18408 & n26939 ) ;
  assign n26941 = ( ~n12558 & n16439 ) | ( ~n12558 & n26940 ) | ( n16439 & n26940 ) ;
  assign n26942 = ( n7943 & ~n12131 ) | ( n7943 & n26941 ) | ( ~n12131 & n26941 ) ;
  assign n26943 = ( ~n7859 & n9572 ) | ( ~n7859 & n25353 ) | ( n9572 & n25353 ) ;
  assign n26944 = ( n622 & n7537 ) | ( n622 & n16487 ) | ( n7537 & n16487 ) ;
  assign n26945 = n15661 ^ n5884 ^ n3749 ;
  assign n26946 = n26945 ^ n19196 ^ n15706 ;
  assign n26947 = ( n1151 & ~n1967 ) | ( n1151 & n2090 ) | ( ~n1967 & n2090 ) ;
  assign n26948 = ( ~n7174 & n15465 ) | ( ~n7174 & n26947 ) | ( n15465 & n26947 ) ;
  assign n26949 = n26948 ^ n21384 ^ n15661 ;
  assign n26950 = n8162 ^ n5482 ^ n538 ;
  assign n26951 = ( ~n4732 & n26604 ) | ( ~n4732 & n26950 ) | ( n26604 & n26950 ) ;
  assign n26952 = n21116 ^ n7612 ^ n7059 ;
  assign n26953 = ( n17659 & n26629 ) | ( n17659 & ~n26952 ) | ( n26629 & ~n26952 ) ;
  assign n26954 = ( n2772 & ~n11886 ) | ( n2772 & n13437 ) | ( ~n11886 & n13437 ) ;
  assign n26955 = ( n9236 & ~n12609 ) | ( n9236 & n23775 ) | ( ~n12609 & n23775 ) ;
  assign n26956 = n16024 ^ n9499 ^ n5459 ;
  assign n26957 = ( n13735 & n26955 ) | ( n13735 & n26956 ) | ( n26955 & n26956 ) ;
  assign n26958 = ( ~n1758 & n10994 ) | ( ~n1758 & n26957 ) | ( n10994 & n26957 ) ;
  assign n26959 = ( n1095 & n15868 ) | ( n1095 & n23893 ) | ( n15868 & n23893 ) ;
  assign n26960 = ( n5303 & n8049 ) | ( n5303 & n13008 ) | ( n8049 & n13008 ) ;
  assign n26961 = n26960 ^ n22463 ^ n19172 ;
  assign n26962 = ( n17604 & n18836 ) | ( n17604 & n26961 ) | ( n18836 & n26961 ) ;
  assign n26963 = ( n19248 & n26959 ) | ( n19248 & ~n26962 ) | ( n26959 & ~n26962 ) ;
  assign n26964 = ( n3495 & n6162 ) | ( n3495 & n16740 ) | ( n6162 & n16740 ) ;
  assign n26965 = n26964 ^ n26704 ^ n8027 ;
  assign n26966 = n26092 ^ n19374 ^ n14933 ;
  assign n26967 = ( n6575 & n15075 ) | ( n6575 & n26966 ) | ( n15075 & n26966 ) ;
  assign n26968 = ( ~n5396 & n25795 ) | ( ~n5396 & n26839 ) | ( n25795 & n26839 ) ;
  assign n26969 = ( n8910 & n10819 ) | ( n8910 & ~n25418 ) | ( n10819 & ~n25418 ) ;
  assign n26970 = n26969 ^ n25716 ^ n10911 ;
  assign n26971 = ( ~n1915 & n18167 ) | ( ~n1915 & n26970 ) | ( n18167 & n26970 ) ;
  assign n26972 = ( n2099 & n4567 ) | ( n2099 & ~n7802 ) | ( n4567 & ~n7802 ) ;
  assign n26973 = ( n3140 & ~n13244 ) | ( n3140 & n20753 ) | ( ~n13244 & n20753 ) ;
  assign n26974 = ( n3047 & n9266 ) | ( n3047 & ~n12203 ) | ( n9266 & ~n12203 ) ;
  assign n26975 = ( ~n1808 & n10596 ) | ( ~n1808 & n26974 ) | ( n10596 & n26974 ) ;
  assign n26976 = n20977 ^ n18717 ^ n4691 ;
  assign n26977 = n4691 ^ n4414 ^ n1759 ;
  assign n26978 = n26977 ^ n24797 ^ n23881 ;
  assign n26979 = n25158 ^ n23990 ^ n12864 ;
  assign n26980 = ( n6178 & n8443 ) | ( n6178 & ~n11407 ) | ( n8443 & ~n11407 ) ;
  assign n26981 = n26980 ^ n25178 ^ n11586 ;
  assign n26982 = n26585 ^ n5574 ^ x108 ;
  assign n26983 = ( ~n9467 & n16876 ) | ( ~n9467 & n26982 ) | ( n16876 & n26982 ) ;
  assign n26984 = ( ~n3985 & n12306 ) | ( ~n3985 & n15477 ) | ( n12306 & n15477 ) ;
  assign n26985 = ( ~n10621 & n23576 ) | ( ~n10621 & n26984 ) | ( n23576 & n26984 ) ;
  assign n26986 = ( n4110 & ~n24900 ) | ( n4110 & n26985 ) | ( ~n24900 & n26985 ) ;
  assign n26988 = n23622 ^ n1444 ^ x95 ;
  assign n26987 = ( n1524 & ~n7206 ) | ( n1524 & n9651 ) | ( ~n7206 & n9651 ) ;
  assign n26989 = n26988 ^ n26987 ^ n10118 ;
  assign n26990 = n15687 ^ n12801 ^ n8697 ;
  assign n26991 = ( n1000 & n8106 ) | ( n1000 & ~n13008 ) | ( n8106 & ~n13008 ) ;
  assign n26992 = n26991 ^ n18997 ^ n235 ;
  assign n26993 = ( n2868 & ~n4346 ) | ( n2868 & n26992 ) | ( ~n4346 & n26992 ) ;
  assign n26994 = ( n1198 & n4524 ) | ( n1198 & ~n9085 ) | ( n4524 & ~n9085 ) ;
  assign n26995 = ( ~n1971 & n14334 ) | ( ~n1971 & n19955 ) | ( n14334 & n19955 ) ;
  assign n26996 = n26995 ^ n13896 ^ n858 ;
  assign n26997 = n26996 ^ n19108 ^ n4493 ;
  assign n26998 = ( n3890 & n8553 ) | ( n3890 & n14834 ) | ( n8553 & n14834 ) ;
  assign n26999 = ( n13730 & n15358 ) | ( n13730 & ~n26998 ) | ( n15358 & ~n26998 ) ;
  assign n27001 = ( ~n4003 & n4933 ) | ( ~n4003 & n6828 ) | ( n4933 & n6828 ) ;
  assign n27000 = ( n19137 & n19454 ) | ( n19137 & n24948 ) | ( n19454 & n24948 ) ;
  assign n27002 = n27001 ^ n27000 ^ n20013 ;
  assign n27003 = ( ~n903 & n6878 ) | ( ~n903 & n19883 ) | ( n6878 & n19883 ) ;
  assign n27004 = ( ~n1875 & n19964 ) | ( ~n1875 & n20503 ) | ( n19964 & n20503 ) ;
  assign n27005 = ( ~n2720 & n3493 ) | ( ~n2720 & n27004 ) | ( n3493 & n27004 ) ;
  assign n27006 = ( n7427 & n27003 ) | ( n7427 & ~n27005 ) | ( n27003 & ~n27005 ) ;
  assign n27007 = ( ~n608 & n8660 ) | ( ~n608 & n27006 ) | ( n8660 & n27006 ) ;
  assign n27008 = n8940 ^ n3462 ^ n1937 ;
  assign n27009 = n11589 ^ n5851 ^ n4152 ;
  assign n27010 = n27009 ^ n21060 ^ n20396 ;
  assign n27011 = n27010 ^ n22164 ^ n17486 ;
  assign n27013 = ( n4977 & n22023 ) | ( n4977 & ~n23435 ) | ( n22023 & ~n23435 ) ;
  assign n27012 = ( n510 & n2082 ) | ( n510 & ~n11950 ) | ( n2082 & ~n11950 ) ;
  assign n27014 = n27013 ^ n27012 ^ n5916 ;
  assign n27015 = n8515 ^ n6641 ^ n492 ;
  assign n27016 = n26116 ^ n23341 ^ n18845 ;
  assign n27017 = ( n8139 & n18105 ) | ( n8139 & ~n24874 ) | ( n18105 & ~n24874 ) ;
  assign n27018 = n22446 ^ n20148 ^ n9461 ;
  assign n27019 = ( n5127 & n10228 ) | ( n5127 & n14166 ) | ( n10228 & n14166 ) ;
  assign n27020 = ( n1077 & n4437 ) | ( n1077 & n27019 ) | ( n4437 & n27019 ) ;
  assign n27021 = ( ~n3953 & n9872 ) | ( ~n3953 & n27020 ) | ( n9872 & n27020 ) ;
  assign n27022 = n27021 ^ n22686 ^ n15625 ;
  assign n27023 = n23495 ^ n18779 ^ x60 ;
  assign n27024 = ( ~n3846 & n5662 ) | ( ~n3846 & n14067 ) | ( n5662 & n14067 ) ;
  assign n27025 = ( n499 & ~n8147 ) | ( n499 & n27024 ) | ( ~n8147 & n27024 ) ;
  assign n27026 = ( n12372 & n26012 ) | ( n12372 & ~n27025 ) | ( n26012 & ~n27025 ) ;
  assign n27027 = ( ~n1379 & n9458 ) | ( ~n1379 & n19802 ) | ( n9458 & n19802 ) ;
  assign n27028 = n19314 ^ n16067 ^ n4289 ;
  assign n27029 = ( n5196 & n16423 ) | ( n5196 & ~n27028 ) | ( n16423 & ~n27028 ) ;
  assign n27032 = n17126 ^ n12717 ^ n10849 ;
  assign n27030 = ( n225 & n4734 ) | ( n225 & n10007 ) | ( n4734 & n10007 ) ;
  assign n27031 = ( n3124 & ~n9213 ) | ( n3124 & n27030 ) | ( ~n9213 & n27030 ) ;
  assign n27033 = n27032 ^ n27031 ^ n3084 ;
  assign n27034 = n18988 ^ n14535 ^ n9467 ;
  assign n27035 = n27034 ^ n12407 ^ n11035 ;
  assign n27036 = ( n3984 & n6336 ) | ( n3984 & ~n7577 ) | ( n6336 & ~n7577 ) ;
  assign n27037 = ( n1803 & n3074 ) | ( n1803 & ~n27036 ) | ( n3074 & ~n27036 ) ;
  assign n27038 = n8396 ^ n8237 ^ n348 ;
  assign n27039 = ( ~n10701 & n27037 ) | ( ~n10701 & n27038 ) | ( n27037 & n27038 ) ;
  assign n27040 = ( n15269 & ~n18326 ) | ( n15269 & n27039 ) | ( ~n18326 & n27039 ) ;
  assign n27041 = n25350 ^ n15830 ^ n9117 ;
  assign n27042 = ( ~n1840 & n24788 ) | ( ~n1840 & n27041 ) | ( n24788 & n27041 ) ;
  assign n27043 = n10087 ^ n2043 ^ n564 ;
  assign n27044 = ( n19502 & ~n27042 ) | ( n19502 & n27043 ) | ( ~n27042 & n27043 ) ;
  assign n27045 = n23280 ^ n6356 ^ n2649 ;
  assign n27046 = ( n11697 & n12954 ) | ( n11697 & ~n20502 ) | ( n12954 & ~n20502 ) ;
  assign n27047 = n27046 ^ n26017 ^ n14676 ;
  assign n27048 = ( n10698 & n16844 ) | ( n10698 & n27047 ) | ( n16844 & n27047 ) ;
  assign n27049 = n17401 ^ n4814 ^ n2275 ;
  assign n27050 = ( ~n17269 & n26514 ) | ( ~n17269 & n27049 ) | ( n26514 & n27049 ) ;
  assign n27051 = n17708 ^ n7362 ^ n2268 ;
  assign n27052 = ( n12066 & ~n14688 ) | ( n12066 & n27051 ) | ( ~n14688 & n27051 ) ;
  assign n27053 = ( n2785 & ~n4686 ) | ( n2785 & n16280 ) | ( ~n4686 & n16280 ) ;
  assign n27054 = ( n19291 & ~n27052 ) | ( n19291 & n27053 ) | ( ~n27052 & n27053 ) ;
  assign n27055 = ( n8797 & n15979 ) | ( n8797 & n16798 ) | ( n15979 & n16798 ) ;
  assign n27056 = ( n2708 & n7532 ) | ( n2708 & n23428 ) | ( n7532 & n23428 ) ;
  assign n27057 = ( n7476 & n17139 ) | ( n7476 & n27056 ) | ( n17139 & n27056 ) ;
  assign n27058 = n19651 ^ n2242 ^ n2189 ;
  assign n27059 = ( n14215 & n27057 ) | ( n14215 & n27058 ) | ( n27057 & n27058 ) ;
  assign n27060 = ( n5114 & n16102 ) | ( n5114 & ~n27059 ) | ( n16102 & ~n27059 ) ;
  assign n27061 = ( n2341 & ~n16036 ) | ( n2341 & n19545 ) | ( ~n16036 & n19545 ) ;
  assign n27062 = n22223 ^ n6776 ^ n2075 ;
  assign n27063 = n27062 ^ n18072 ^ n1794 ;
  assign n27064 = ( ~n17250 & n27061 ) | ( ~n17250 & n27063 ) | ( n27061 & n27063 ) ;
  assign n27065 = n15484 ^ n15438 ^ n10631 ;
  assign n27066 = ( ~n8115 & n25902 ) | ( ~n8115 & n27065 ) | ( n25902 & n27065 ) ;
  assign n27067 = ( n3004 & n8562 ) | ( n3004 & n15119 ) | ( n8562 & n15119 ) ;
  assign n27068 = n27067 ^ n16438 ^ n7658 ;
  assign n27070 = n19857 ^ n18191 ^ n9291 ;
  assign n27071 = ( n12623 & n23602 ) | ( n12623 & n27070 ) | ( n23602 & n27070 ) ;
  assign n27069 = n20410 ^ n7035 ^ n6585 ;
  assign n27072 = n27071 ^ n27069 ^ n13948 ;
  assign n27073 = ( n5884 & n10640 ) | ( n5884 & n22031 ) | ( n10640 & n22031 ) ;
  assign n27074 = ( n18841 & n26670 ) | ( n18841 & n27073 ) | ( n26670 & n27073 ) ;
  assign n27075 = ( n4005 & ~n7835 ) | ( n4005 & n23753 ) | ( ~n7835 & n23753 ) ;
  assign n27076 = n7901 ^ n6904 ^ n3814 ;
  assign n27077 = ( n12358 & n12751 ) | ( n12358 & n17370 ) | ( n12751 & n17370 ) ;
  assign n27078 = ( n2088 & n27076 ) | ( n2088 & ~n27077 ) | ( n27076 & ~n27077 ) ;
  assign n27079 = ( n7232 & n11467 ) | ( n7232 & n24097 ) | ( n11467 & n24097 ) ;
  assign n27080 = ( n9746 & n24660 ) | ( n9746 & n27079 ) | ( n24660 & n27079 ) ;
  assign n27081 = ( n400 & ~n2055 ) | ( n400 & n5939 ) | ( ~n2055 & n5939 ) ;
  assign n27082 = n27081 ^ n4498 ^ n2840 ;
  assign n27083 = n8460 ^ n6804 ^ n3316 ;
  assign n27084 = n18676 ^ n5363 ^ x16 ;
  assign n27085 = ( ~n379 & n3606 ) | ( ~n379 & n6367 ) | ( n3606 & n6367 ) ;
  assign n27086 = n27085 ^ n9937 ^ n3854 ;
  assign n27087 = n11952 ^ n10954 ^ n1722 ;
  assign n27088 = ( n7282 & n10572 ) | ( n7282 & ~n27087 ) | ( n10572 & ~n27087 ) ;
  assign n27089 = ( n1891 & n3367 ) | ( n1891 & ~n5546 ) | ( n3367 & ~n5546 ) ;
  assign n27090 = n27089 ^ n11071 ^ n1515 ;
  assign n27091 = ( n5989 & n27088 ) | ( n5989 & n27090 ) | ( n27088 & n27090 ) ;
  assign n27092 = n22200 ^ n4430 ^ n2210 ;
  assign n27093 = n19338 ^ n15659 ^ n12880 ;
  assign n27094 = ( n1665 & n8398 ) | ( n1665 & ~n15773 ) | ( n8398 & ~n15773 ) ;
  assign n27095 = ( n4793 & ~n8160 ) | ( n4793 & n27094 ) | ( ~n8160 & n27094 ) ;
  assign n27096 = ( n702 & ~n2127 ) | ( n702 & n21293 ) | ( ~n2127 & n21293 ) ;
  assign n27097 = n27096 ^ n25337 ^ n19996 ;
  assign n27098 = n27097 ^ n19425 ^ n1804 ;
  assign n27099 = n27098 ^ n15161 ^ n2773 ;
  assign n27100 = n19620 ^ n10629 ^ n9796 ;
  assign n27101 = ( n14339 & n19502 ) | ( n14339 & ~n27100 ) | ( n19502 & ~n27100 ) ;
  assign n27102 = ( ~n4113 & n24556 ) | ( ~n4113 & n27101 ) | ( n24556 & n27101 ) ;
  assign n27103 = n16787 ^ n13194 ^ n10790 ;
  assign n27104 = ( ~n3718 & n5248 ) | ( ~n3718 & n6345 ) | ( n5248 & n6345 ) ;
  assign n27105 = ( ~n5372 & n8802 ) | ( ~n5372 & n13749 ) | ( n8802 & n13749 ) ;
  assign n27106 = ( n5860 & n16860 ) | ( n5860 & ~n27105 ) | ( n16860 & ~n27105 ) ;
  assign n27107 = n21387 ^ n20943 ^ n19510 ;
  assign n27108 = ( ~n14714 & n20028 ) | ( ~n14714 & n25778 ) | ( n20028 & n25778 ) ;
  assign n27109 = ( ~n6547 & n16043 ) | ( ~n6547 & n27108 ) | ( n16043 & n27108 ) ;
  assign n27110 = ( n14978 & ~n18446 ) | ( n14978 & n20298 ) | ( ~n18446 & n20298 ) ;
  assign n27111 = n27110 ^ n13887 ^ n11732 ;
  assign n27112 = ( n1179 & n2343 ) | ( n1179 & n19501 ) | ( n2343 & n19501 ) ;
  assign n27113 = ( n4828 & n10880 ) | ( n4828 & ~n25916 ) | ( n10880 & ~n25916 ) ;
  assign n27114 = ( n3484 & ~n18572 ) | ( n3484 & n27113 ) | ( ~n18572 & n27113 ) ;
  assign n27115 = ( n5264 & ~n18041 ) | ( n5264 & n27114 ) | ( ~n18041 & n27114 ) ;
  assign n27116 = ( ~n5362 & n10709 ) | ( ~n5362 & n27115 ) | ( n10709 & n27115 ) ;
  assign n27117 = ( n2034 & n6942 ) | ( n2034 & ~n20496 ) | ( n6942 & ~n20496 ) ;
  assign n27118 = ( n805 & n2802 ) | ( n805 & n14354 ) | ( n2802 & n14354 ) ;
  assign n27119 = ( n846 & n23060 ) | ( n846 & n25110 ) | ( n23060 & n25110 ) ;
  assign n27120 = n7326 ^ n5968 ^ n1171 ;
  assign n27121 = n27120 ^ n22445 ^ n15004 ;
  assign n27122 = ( n24786 & ~n25671 ) | ( n24786 & n27121 ) | ( ~n25671 & n27121 ) ;
  assign n27123 = n24424 ^ n18902 ^ n3993 ;
  assign n27124 = n27123 ^ n17276 ^ n868 ;
  assign n27126 = n18316 ^ n11209 ^ n4398 ;
  assign n27125 = n16477 ^ n10561 ^ n7862 ;
  assign n27127 = n27126 ^ n27125 ^ n5449 ;
  assign n27128 = n8378 ^ n6856 ^ n3150 ;
  assign n27129 = ( n10182 & n12743 ) | ( n10182 & n27128 ) | ( n12743 & n27128 ) ;
  assign n27130 = ( n5459 & ~n5495 ) | ( n5459 & n14593 ) | ( ~n5495 & n14593 ) ;
  assign n27131 = ( n7818 & n27129 ) | ( n7818 & n27130 ) | ( n27129 & n27130 ) ;
  assign n27132 = ( n3858 & ~n9075 ) | ( n3858 & n13775 ) | ( ~n9075 & n13775 ) ;
  assign n27133 = ( n1872 & n15696 ) | ( n1872 & n16783 ) | ( n15696 & n16783 ) ;
  assign n27134 = ( ~n7074 & n17279 ) | ( ~n7074 & n27133 ) | ( n17279 & n27133 ) ;
  assign n27136 = ( n4115 & n5384 ) | ( n4115 & n8152 ) | ( n5384 & n8152 ) ;
  assign n27135 = n20627 ^ n17452 ^ n16906 ;
  assign n27137 = n27136 ^ n27135 ^ n23584 ;
  assign n27138 = n14645 ^ n12216 ^ n12123 ;
  assign n27139 = n27138 ^ n18446 ^ n136 ;
  assign n27140 = ( ~n8914 & n22620 ) | ( ~n8914 & n24655 ) | ( n22620 & n24655 ) ;
  assign n27141 = ( ~n5111 & n15391 ) | ( ~n5111 & n23981 ) | ( n15391 & n23981 ) ;
  assign n27142 = n23977 ^ n11010 ^ n7972 ;
  assign n27143 = ( ~n5472 & n13656 ) | ( ~n5472 & n13996 ) | ( n13656 & n13996 ) ;
  assign n27144 = n21413 ^ n13775 ^ n2348 ;
  assign n27145 = n16227 ^ n2812 ^ n2619 ;
  assign n27146 = ( n10844 & n11976 ) | ( n10844 & n27145 ) | ( n11976 & n27145 ) ;
  assign n27147 = n27146 ^ n11125 ^ n8713 ;
  assign n27148 = n10695 ^ n9430 ^ n4039 ;
  assign n27149 = n5684 ^ n5283 ^ n2204 ;
  assign n27150 = n17618 ^ n10106 ^ n944 ;
  assign n27153 = n20211 ^ n16650 ^ n7276 ;
  assign n27151 = ( n262 & n2231 ) | ( n262 & n22026 ) | ( n2231 & n22026 ) ;
  assign n27152 = n27151 ^ n22646 ^ n21210 ;
  assign n27154 = n27153 ^ n27152 ^ n24489 ;
  assign n27157 = ( ~n6830 & n13067 ) | ( ~n6830 & n20325 ) | ( n13067 & n20325 ) ;
  assign n27155 = ( ~n1954 & n5448 ) | ( ~n1954 & n9011 ) | ( n5448 & n9011 ) ;
  assign n27156 = n27155 ^ n14420 ^ n332 ;
  assign n27158 = n27157 ^ n27156 ^ n6901 ;
  assign n27159 = ( n738 & n17674 ) | ( n738 & n27158 ) | ( n17674 & n27158 ) ;
  assign n27160 = n27159 ^ n24058 ^ n7969 ;
  assign n27161 = ( n10350 & ~n13366 ) | ( n10350 & n24067 ) | ( ~n13366 & n24067 ) ;
  assign n27162 = n15045 ^ n9498 ^ n7713 ;
  assign n27163 = n27162 ^ n6918 ^ n2814 ;
  assign n27164 = ( n9179 & ~n10878 ) | ( n9179 & n23854 ) | ( ~n10878 & n23854 ) ;
  assign n27165 = ( n456 & n3034 ) | ( n456 & n13661 ) | ( n3034 & n13661 ) ;
  assign n27166 = ( ~n17316 & n27164 ) | ( ~n17316 & n27165 ) | ( n27164 & n27165 ) ;
  assign n27167 = ( ~n3601 & n12368 ) | ( ~n3601 & n21941 ) | ( n12368 & n21941 ) ;
  assign n27168 = n20478 ^ n6552 ^ n277 ;
  assign n27169 = ( n11204 & n27167 ) | ( n11204 & n27168 ) | ( n27167 & n27168 ) ;
  assign n27170 = ( n4558 & n7737 ) | ( n4558 & ~n23399 ) | ( n7737 & ~n23399 ) ;
  assign n27171 = ( n1900 & n5604 ) | ( n1900 & n27170 ) | ( n5604 & n27170 ) ;
  assign n27172 = n11556 ^ n8263 ^ n142 ;
  assign n27173 = ( n1558 & n5319 ) | ( n1558 & ~n12433 ) | ( n5319 & ~n12433 ) ;
  assign n27175 = ( n7904 & n15597 ) | ( n7904 & n25692 ) | ( n15597 & n25692 ) ;
  assign n27174 = n14771 ^ n9936 ^ n7595 ;
  assign n27176 = n27175 ^ n27174 ^ n21543 ;
  assign n27177 = n4479 ^ n1807 ^ n1061 ;
  assign n27178 = n27177 ^ n22613 ^ n14061 ;
  assign n27179 = ( n3681 & n4433 ) | ( n3681 & n6624 ) | ( n4433 & n6624 ) ;
  assign n27180 = n19570 ^ n14121 ^ n543 ;
  assign n27181 = ( n13511 & n17906 ) | ( n13511 & n19452 ) | ( n17906 & n19452 ) ;
  assign n27182 = n27181 ^ n6166 ^ n1311 ;
  assign n27183 = ( n13366 & n14144 ) | ( n13366 & n27182 ) | ( n14144 & n27182 ) ;
  assign n27184 = n27183 ^ n11319 ^ n1870 ;
  assign n27185 = ( n857 & ~n21091 ) | ( n857 & n23288 ) | ( ~n21091 & n23288 ) ;
  assign n27186 = n27185 ^ n20866 ^ n7472 ;
  assign n27187 = ( n11451 & n17366 ) | ( n11451 & ~n18371 ) | ( n17366 & ~n18371 ) ;
  assign n27188 = ( n10265 & n19383 ) | ( n10265 & n20989 ) | ( n19383 & n20989 ) ;
  assign n27189 = n16659 ^ n13808 ^ n7109 ;
  assign n27190 = n27189 ^ n22945 ^ n22183 ;
  assign n27193 = ( ~n1479 & n6009 ) | ( ~n1479 & n7951 ) | ( n6009 & n7951 ) ;
  assign n27192 = n23084 ^ n14349 ^ n1380 ;
  assign n27191 = ( n1783 & n7239 ) | ( n1783 & ~n12269 ) | ( n7239 & ~n12269 ) ;
  assign n27194 = n27193 ^ n27192 ^ n27191 ;
  assign n27195 = n7914 ^ n3636 ^ n1179 ;
  assign n27196 = ( n10586 & n10732 ) | ( n10586 & ~n18679 ) | ( n10732 & ~n18679 ) ;
  assign n27197 = ( n6103 & n13237 ) | ( n6103 & ~n27196 ) | ( n13237 & ~n27196 ) ;
  assign n27198 = n4774 ^ n4764 ^ n1875 ;
  assign n27199 = n21445 ^ n6271 ^ n3264 ;
  assign n27200 = ( n16403 & n23330 ) | ( n16403 & ~n27199 ) | ( n23330 & ~n27199 ) ;
  assign n27201 = ( n23439 & n27198 ) | ( n23439 & n27200 ) | ( n27198 & n27200 ) ;
  assign n27206 = ( n8811 & ~n15278 ) | ( n8811 & n15886 ) | ( ~n15278 & n15886 ) ;
  assign n27207 = n27206 ^ n23775 ^ n6235 ;
  assign n27205 = n21173 ^ n9869 ^ n8620 ;
  assign n27202 = n19060 ^ n6105 ^ n3864 ;
  assign n27203 = n27202 ^ n16229 ^ n14433 ;
  assign n27204 = ( n3593 & n11798 ) | ( n3593 & ~n27203 ) | ( n11798 & ~n27203 ) ;
  assign n27208 = n27207 ^ n27205 ^ n27204 ;
  assign n27209 = ( n17040 & ~n24733 ) | ( n17040 & n26156 ) | ( ~n24733 & n26156 ) ;
  assign n27210 = n19054 ^ n10989 ^ n5220 ;
  assign n27211 = n22240 ^ n21832 ^ n3126 ;
  assign n27212 = ( n19602 & ~n27210 ) | ( n19602 & n27211 ) | ( ~n27210 & n27211 ) ;
  assign n27213 = ( n8379 & n27209 ) | ( n8379 & n27212 ) | ( n27209 & n27212 ) ;
  assign n27217 = ( ~n1178 & n6099 ) | ( ~n1178 & n10611 ) | ( n6099 & n10611 ) ;
  assign n27215 = ( ~n876 & n5873 ) | ( ~n876 & n6776 ) | ( n5873 & n6776 ) ;
  assign n27214 = n12526 ^ n10850 ^ n2320 ;
  assign n27216 = n27215 ^ n27214 ^ n10690 ;
  assign n27218 = n27217 ^ n27216 ^ n10391 ;
  assign n27219 = ( n1318 & ~n2864 ) | ( n1318 & n3274 ) | ( ~n2864 & n3274 ) ;
  assign n27220 = ( ~n467 & n13648 ) | ( ~n467 & n19932 ) | ( n13648 & n19932 ) ;
  assign n27221 = ( n2830 & n6866 ) | ( n2830 & ~n9781 ) | ( n6866 & ~n9781 ) ;
  assign n27222 = n27221 ^ n12890 ^ n10298 ;
  assign n27223 = n17596 ^ n11990 ^ n7697 ;
  assign n27224 = ( ~n4488 & n5121 ) | ( ~n4488 & n5927 ) | ( n5121 & n5927 ) ;
  assign n27225 = n27224 ^ n27110 ^ n4484 ;
  assign n27226 = ( ~n636 & n16113 ) | ( ~n636 & n22321 ) | ( n16113 & n22321 ) ;
  assign n27227 = ( ~n1707 & n10161 ) | ( ~n1707 & n17855 ) | ( n10161 & n17855 ) ;
  assign n27228 = n27227 ^ n14860 ^ n4772 ;
  assign n27229 = ( x0 & ~n15672 ) | ( x0 & n27228 ) | ( ~n15672 & n27228 ) ;
  assign n27230 = ( ~n9078 & n22888 ) | ( ~n9078 & n24597 ) | ( n22888 & n24597 ) ;
  assign n27231 = n8798 ^ n6791 ^ n6417 ;
  assign n27232 = n27231 ^ n23473 ^ n16564 ;
  assign n27233 = n8801 ^ n5174 ^ n2044 ;
  assign n27234 = ( ~n2827 & n13422 ) | ( ~n2827 & n20376 ) | ( n13422 & n20376 ) ;
  assign n27235 = ( n4596 & ~n6189 ) | ( n4596 & n6754 ) | ( ~n6189 & n6754 ) ;
  assign n27236 = ( n4930 & n18473 ) | ( n4930 & n27235 ) | ( n18473 & n27235 ) ;
  assign n27237 = ( n19706 & n27234 ) | ( n19706 & ~n27236 ) | ( n27234 & ~n27236 ) ;
  assign n27238 = n18692 ^ n13315 ^ n9755 ;
  assign n27239 = n13848 ^ n11780 ^ n3638 ;
  assign n27240 = ( ~n24671 & n27238 ) | ( ~n24671 & n27239 ) | ( n27238 & n27239 ) ;
  assign n27241 = n27240 ^ n13449 ^ n10174 ;
  assign n27242 = ( n13923 & ~n18469 ) | ( n13923 & n21980 ) | ( ~n18469 & n21980 ) ;
  assign n27243 = n17466 ^ n13663 ^ n5034 ;
  assign n27244 = n17827 ^ n3107 ^ n260 ;
  assign n27245 = n27244 ^ n8200 ^ n242 ;
  assign n27246 = ( n22040 & n27243 ) | ( n22040 & ~n27245 ) | ( n27243 & ~n27245 ) ;
  assign n27247 = ( n1575 & ~n7301 ) | ( n1575 & n18434 ) | ( ~n7301 & n18434 ) ;
  assign n27248 = ( ~n22362 & n27246 ) | ( ~n22362 & n27247 ) | ( n27246 & n27247 ) ;
  assign n27249 = ( n949 & n7585 ) | ( n949 & ~n14114 ) | ( n7585 & ~n14114 ) ;
  assign n27250 = n19410 ^ n7976 ^ n3990 ;
  assign n27251 = ( n3514 & n12105 ) | ( n3514 & n27250 ) | ( n12105 & n27250 ) ;
  assign n27252 = ( n9716 & n27249 ) | ( n9716 & ~n27251 ) | ( n27249 & ~n27251 ) ;
  assign n27253 = ( n5286 & ~n10450 ) | ( n5286 & n27252 ) | ( ~n10450 & n27252 ) ;
  assign n27254 = ( n7357 & ~n8150 ) | ( n7357 & n17632 ) | ( ~n8150 & n17632 ) ;
  assign n27255 = ( n6036 & ~n9581 ) | ( n6036 & n15168 ) | ( ~n9581 & n15168 ) ;
  assign n27256 = ( n25568 & n27254 ) | ( n25568 & ~n27255 ) | ( n27254 & ~n27255 ) ;
  assign n27257 = ( ~n14545 & n26637 ) | ( ~n14545 & n27256 ) | ( n26637 & n27256 ) ;
  assign n27258 = ( n655 & n846 ) | ( n655 & n15250 ) | ( n846 & n15250 ) ;
  assign n27259 = n27258 ^ n15035 ^ n14675 ;
  assign n27260 = n19684 ^ n11327 ^ n4904 ;
  assign n27261 = ( ~n790 & n10320 ) | ( ~n790 & n20832 ) | ( n10320 & n20832 ) ;
  assign n27262 = ( n9972 & ~n11012 ) | ( n9972 & n16667 ) | ( ~n11012 & n16667 ) ;
  assign n27263 = ( ~n2673 & n13344 ) | ( ~n2673 & n27262 ) | ( n13344 & n27262 ) ;
  assign n27265 = n5183 ^ n788 ^ n622 ;
  assign n27264 = n4048 ^ n4034 ^ n635 ;
  assign n27266 = n27265 ^ n27264 ^ n11051 ;
  assign n27267 = n23704 ^ n17115 ^ n5587 ;
  assign n27268 = n27267 ^ n12295 ^ n7425 ;
  assign n27269 = ( n4503 & n8295 ) | ( n4503 & n8553 ) | ( n8295 & n8553 ) ;
  assign n27270 = ( n10057 & n27268 ) | ( n10057 & n27269 ) | ( n27268 & n27269 ) ;
  assign n27271 = ( ~n15159 & n20185 ) | ( ~n15159 & n22294 ) | ( n20185 & n22294 ) ;
  assign n27272 = ( n227 & ~n955 ) | ( n227 & n27271 ) | ( ~n955 & n27271 ) ;
  assign n27274 = ( n5435 & n10756 ) | ( n5435 & n10887 ) | ( n10756 & n10887 ) ;
  assign n27273 = n19510 ^ n18955 ^ n894 ;
  assign n27275 = n27274 ^ n27273 ^ n16635 ;
  assign n27276 = ( n8442 & n8445 ) | ( n8442 & n24053 ) | ( n8445 & n24053 ) ;
  assign n27277 = ( ~n152 & n11079 ) | ( ~n152 & n14707 ) | ( n11079 & n14707 ) ;
  assign n27278 = ( ~n20187 & n27276 ) | ( ~n20187 & n27277 ) | ( n27276 & n27277 ) ;
  assign n27279 = n19123 ^ n16665 ^ n7170 ;
  assign n27280 = n27279 ^ n20119 ^ n996 ;
  assign n27281 = n27280 ^ n20420 ^ n16516 ;
  assign n27282 = ( n7919 & n14244 ) | ( n7919 & ~n17818 ) | ( n14244 & ~n17818 ) ;
  assign n27283 = n25263 ^ n3698 ^ n1850 ;
  assign n27284 = n19471 ^ n17392 ^ n7352 ;
  assign n27285 = ( n4301 & ~n26070 ) | ( n4301 & n27284 ) | ( ~n26070 & n27284 ) ;
  assign n27286 = n8906 ^ n5092 ^ n4757 ;
  assign n27287 = ( ~n6380 & n9523 ) | ( ~n6380 & n13834 ) | ( n9523 & n13834 ) ;
  assign n27288 = ( n1682 & n10007 ) | ( n1682 & n15256 ) | ( n10007 & n15256 ) ;
  assign n27289 = ( n586 & ~n3671 ) | ( n586 & n25167 ) | ( ~n3671 & n25167 ) ;
  assign n27290 = n22360 ^ n15850 ^ n1157 ;
  assign n27291 = ( n4920 & ~n5541 ) | ( n4920 & n27290 ) | ( ~n5541 & n27290 ) ;
  assign n27292 = ( ~n7807 & n12008 ) | ( ~n7807 & n17795 ) | ( n12008 & n17795 ) ;
  assign n27293 = ( n16989 & n17215 ) | ( n16989 & ~n27292 ) | ( n17215 & ~n27292 ) ;
  assign n27294 = n24312 ^ n15121 ^ n3340 ;
  assign n27296 = n20146 ^ n9168 ^ n2837 ;
  assign n27295 = ( ~n1063 & n11773 ) | ( ~n1063 & n12524 ) | ( n11773 & n12524 ) ;
  assign n27297 = n27296 ^ n27295 ^ n4419 ;
  assign n27298 = ( n22399 & ~n27294 ) | ( n22399 & n27297 ) | ( ~n27294 & n27297 ) ;
  assign n27299 = n8161 ^ n3444 ^ n771 ;
  assign n27300 = ( n16521 & ~n22796 ) | ( n16521 & n27299 ) | ( ~n22796 & n27299 ) ;
  assign n27301 = n14171 ^ n13611 ^ n10946 ;
  assign n27302 = n1841 ^ n932 ^ n577 ;
  assign n27303 = ( n9811 & ~n16959 ) | ( n9811 & n27302 ) | ( ~n16959 & n27302 ) ;
  assign n27304 = ( n1664 & n2960 ) | ( n1664 & ~n9898 ) | ( n2960 & ~n9898 ) ;
  assign n27305 = n27304 ^ n15492 ^ n13116 ;
  assign n27306 = n27305 ^ n19312 ^ n14680 ;
  assign n27307 = ( n3952 & ~n21494 ) | ( n3952 & n22119 ) | ( ~n21494 & n22119 ) ;
  assign n27310 = ( n1979 & n8629 ) | ( n1979 & n18446 ) | ( n8629 & n18446 ) ;
  assign n27308 = ( n7510 & n7840 ) | ( n7510 & n13251 ) | ( n7840 & n13251 ) ;
  assign n27309 = ( n21067 & n23972 ) | ( n21067 & n27308 ) | ( n23972 & n27308 ) ;
  assign n27311 = n27310 ^ n27309 ^ n15054 ;
  assign n27312 = ( ~n12597 & n24626 ) | ( ~n12597 & n27311 ) | ( n24626 & n27311 ) ;
  assign n27313 = ( n17231 & ~n24971 ) | ( n17231 & n27037 ) | ( ~n24971 & n27037 ) ;
  assign n27314 = ( n3878 & n9583 ) | ( n3878 & ~n16083 ) | ( n9583 & ~n16083 ) ;
  assign n27315 = ( n1943 & n19978 ) | ( n1943 & ~n27314 ) | ( n19978 & ~n27314 ) ;
  assign n27316 = ( n2850 & n5654 ) | ( n2850 & n6432 ) | ( n5654 & n6432 ) ;
  assign n27317 = n26278 ^ n17903 ^ n6645 ;
  assign n27318 = ( n8838 & ~n27316 ) | ( n8838 & n27317 ) | ( ~n27316 & n27317 ) ;
  assign n27319 = ( ~n5660 & n7470 ) | ( ~n5660 & n7878 ) | ( n7470 & n7878 ) ;
  assign n27320 = ( n1034 & ~n5701 ) | ( n1034 & n16708 ) | ( ~n5701 & n16708 ) ;
  assign n27321 = n14852 ^ n11369 ^ n7316 ;
  assign n27322 = ( ~n7707 & n21953 ) | ( ~n7707 & n27321 ) | ( n21953 & n27321 ) ;
  assign n27323 = n25699 ^ n25116 ^ n15317 ;
  assign n27324 = n13373 ^ n9431 ^ n3152 ;
  assign n27325 = n27324 ^ n9466 ^ n3000 ;
  assign n27326 = ( n2972 & n3380 ) | ( n2972 & ~n27325 ) | ( n3380 & ~n27325 ) ;
  assign n27327 = ( n8445 & n9696 ) | ( n8445 & ~n19578 ) | ( n9696 & ~n19578 ) ;
  assign n27328 = ( n1702 & n11204 ) | ( n1702 & n27327 ) | ( n11204 & n27327 ) ;
  assign n27329 = n814 ^ n508 ^ x0 ;
  assign n27330 = ( n9020 & n10203 ) | ( n9020 & n23329 ) | ( n10203 & n23329 ) ;
  assign n27331 = n27330 ^ n14613 ^ n13280 ;
  assign n27332 = ( n9748 & ~n22432 ) | ( n9748 & n27331 ) | ( ~n22432 & n27331 ) ;
  assign n27333 = ( n3645 & ~n5225 ) | ( n3645 & n21148 ) | ( ~n5225 & n21148 ) ;
  assign n27334 = ( n274 & ~n14814 ) | ( n274 & n25321 ) | ( ~n14814 & n25321 ) ;
  assign n27335 = n25446 ^ n22409 ^ n11915 ;
  assign n27336 = ( n6839 & n6910 ) | ( n6839 & n27335 ) | ( n6910 & n27335 ) ;
  assign n27337 = ( ~n2583 & n18908 ) | ( ~n2583 & n27336 ) | ( n18908 & n27336 ) ;
  assign n27338 = n10971 ^ n8433 ^ n341 ;
  assign n27339 = n27338 ^ n16984 ^ n9475 ;
  assign n27340 = ( n2320 & n5302 ) | ( n2320 & n25576 ) | ( n5302 & n25576 ) ;
  assign n27341 = ( n1107 & n3575 ) | ( n1107 & ~n25024 ) | ( n3575 & ~n25024 ) ;
  assign n27342 = n24176 ^ n8259 ^ n7781 ;
  assign n27343 = n19226 ^ n11292 ^ n1966 ;
  assign n27344 = ( n12915 & n16238 ) | ( n12915 & n27343 ) | ( n16238 & n27343 ) ;
  assign n27345 = n26781 ^ n24354 ^ n22032 ;
  assign n27346 = ( n7140 & ~n9780 ) | ( n7140 & n27345 ) | ( ~n9780 & n27345 ) ;
  assign n27347 = ( ~n7791 & n16131 ) | ( ~n7791 & n20881 ) | ( n16131 & n20881 ) ;
  assign n27348 = n27347 ^ n25258 ^ n14876 ;
  assign n27349 = n23059 ^ n16155 ^ n10996 ;
  assign n27350 = ( n15320 & ~n17441 ) | ( n15320 & n19718 ) | ( ~n17441 & n19718 ) ;
  assign n27351 = ( n6645 & n8597 ) | ( n6645 & n17122 ) | ( n8597 & n17122 ) ;
  assign n27352 = n27351 ^ n6670 ^ n2153 ;
  assign n27353 = ( n15143 & n16421 ) | ( n15143 & ~n17372 ) | ( n16421 & ~n17372 ) ;
  assign n27354 = n8548 ^ n3904 ^ n3293 ;
  assign n27355 = ( n3029 & n4616 ) | ( n3029 & n9792 ) | ( n4616 & n9792 ) ;
  assign n27356 = n27355 ^ n19142 ^ n10212 ;
  assign n27357 = ( n5163 & ~n13488 ) | ( n5163 & n24162 ) | ( ~n13488 & n24162 ) ;
  assign n27362 = ( x65 & n942 ) | ( x65 & n971 ) | ( n942 & n971 ) ;
  assign n27359 = n7768 ^ n2568 ^ n1215 ;
  assign n27360 = n27359 ^ n23066 ^ n8600 ;
  assign n27358 = ( n6629 & n14300 ) | ( n6629 & n15045 ) | ( n14300 & n15045 ) ;
  assign n27361 = n27360 ^ n27358 ^ n4219 ;
  assign n27363 = n27362 ^ n27361 ^ n6845 ;
  assign n27364 = n16573 ^ n13365 ^ n10966 ;
  assign n27365 = n27364 ^ n10783 ^ n5100 ;
  assign n27366 = n27365 ^ n20358 ^ n11717 ;
  assign n27367 = ( n13893 & n15090 ) | ( n13893 & ~n20551 ) | ( n15090 & ~n20551 ) ;
  assign n27368 = ( n2472 & n13459 ) | ( n2472 & n27367 ) | ( n13459 & n27367 ) ;
  assign n27369 = ( n2814 & ~n10148 ) | ( n2814 & n10781 ) | ( ~n10148 & n10781 ) ;
  assign n27370 = n18685 ^ n6697 ^ n1862 ;
  assign n27371 = ( n1451 & n14067 ) | ( n1451 & n27370 ) | ( n14067 & n27370 ) ;
  assign n27372 = ( n5783 & n15906 ) | ( n5783 & ~n27371 ) | ( n15906 & ~n27371 ) ;
  assign n27373 = ( n387 & n11288 ) | ( n387 & n27372 ) | ( n11288 & n27372 ) ;
  assign n27374 = n9384 ^ n3464 ^ n1337 ;
  assign n27375 = ( n4407 & n15473 ) | ( n4407 & n16698 ) | ( n15473 & n16698 ) ;
  assign n27376 = ( n6784 & n9546 ) | ( n6784 & ~n10938 ) | ( n9546 & ~n10938 ) ;
  assign n27377 = n15238 ^ n12074 ^ n6346 ;
  assign n27378 = n10635 ^ n6798 ^ n5514 ;
  assign n27379 = ( n11598 & ~n23704 ) | ( n11598 & n27378 ) | ( ~n23704 & n27378 ) ;
  assign n27380 = ( n8844 & ~n17443 ) | ( n8844 & n19223 ) | ( ~n17443 & n19223 ) ;
  assign n27381 = n13714 ^ n3617 ^ n2417 ;
  assign n27382 = n27381 ^ n6997 ^ n4282 ;
  assign n27384 = n23944 ^ n22459 ^ n837 ;
  assign n27383 = ( n10695 & n17638 ) | ( n10695 & n20400 ) | ( n17638 & n20400 ) ;
  assign n27385 = n27384 ^ n27383 ^ n2056 ;
  assign n27387 = n12875 ^ n12386 ^ n2211 ;
  assign n27386 = n9894 ^ n3765 ^ n153 ;
  assign n27388 = n27387 ^ n27386 ^ n4154 ;
  assign n27389 = ( n5191 & n7207 ) | ( n5191 & ~n20645 ) | ( n7207 & ~n20645 ) ;
  assign n27390 = n27389 ^ n21102 ^ n2266 ;
  assign n27391 = n20833 ^ n5963 ^ n2850 ;
  assign n27392 = n10613 ^ n6520 ^ n4123 ;
  assign n27393 = ( n8520 & n27391 ) | ( n8520 & ~n27392 ) | ( n27391 & ~n27392 ) ;
  assign n27394 = n27393 ^ n16436 ^ n8724 ;
  assign n27395 = ( n6519 & ~n13367 ) | ( n6519 & n20983 ) | ( ~n13367 & n20983 ) ;
  assign n27396 = n23775 ^ n14806 ^ n5297 ;
  assign n27397 = ( ~n14759 & n22192 ) | ( ~n14759 & n23793 ) | ( n22192 & n23793 ) ;
  assign n27398 = ( n950 & n12107 ) | ( n950 & ~n19456 ) | ( n12107 & ~n19456 ) ;
  assign n27399 = n27398 ^ n11538 ^ n3977 ;
  assign n27400 = n27399 ^ n13531 ^ n11005 ;
  assign n27401 = n14982 ^ n12651 ^ n9144 ;
  assign n27402 = n27401 ^ n4394 ^ n2053 ;
  assign n27403 = n27402 ^ n14780 ^ n4687 ;
  assign n27404 = ( n548 & ~n14534 ) | ( n548 & n23950 ) | ( ~n14534 & n23950 ) ;
  assign n27405 = n12485 ^ n12002 ^ n11575 ;
  assign n27406 = ( n4622 & n15209 ) | ( n4622 & n26555 ) | ( n15209 & n26555 ) ;
  assign n27409 = n13174 ^ n10760 ^ n2795 ;
  assign n27407 = ( ~n265 & n7444 ) | ( ~n265 & n21444 ) | ( n7444 & n21444 ) ;
  assign n27408 = n27407 ^ n9179 ^ n597 ;
  assign n27410 = n27409 ^ n27408 ^ n21235 ;
  assign n27411 = ( n8389 & n12626 ) | ( n8389 & n18872 ) | ( n12626 & n18872 ) ;
  assign n27412 = n27411 ^ n18244 ^ n3910 ;
  assign n27413 = n18425 ^ n10329 ^ n2623 ;
  assign n27414 = ( ~n9771 & n13973 ) | ( ~n9771 & n18931 ) | ( n13973 & n18931 ) ;
  assign n27415 = ( ~n20153 & n20839 ) | ( ~n20153 & n27414 ) | ( n20839 & n27414 ) ;
  assign n27416 = ( n4079 & ~n27413 ) | ( n4079 & n27415 ) | ( ~n27413 & n27415 ) ;
  assign n27417 = ( n11267 & n12728 ) | ( n11267 & ~n16600 ) | ( n12728 & ~n16600 ) ;
  assign n27418 = n27417 ^ n5169 ^ n4595 ;
  assign n27419 = ( n2953 & n19701 ) | ( n2953 & ~n27418 ) | ( n19701 & ~n27418 ) ;
  assign n27420 = n17925 ^ n7119 ^ n610 ;
  assign n27421 = n13285 ^ n12100 ^ n2961 ;
  assign n27422 = n27421 ^ n26289 ^ n10545 ;
  assign n27423 = ( n5587 & n9591 ) | ( n5587 & ~n27422 ) | ( n9591 & ~n27422 ) ;
  assign n27424 = ( n3588 & n7919 ) | ( n3588 & ~n16596 ) | ( n7919 & ~n16596 ) ;
  assign n27425 = n27424 ^ n1031 ^ x83 ;
  assign n27426 = n27425 ^ n21964 ^ n15990 ;
  assign n27427 = ( n224 & n1899 ) | ( n224 & ~n18132 ) | ( n1899 & ~n18132 ) ;
  assign n27428 = n27427 ^ n19137 ^ n3775 ;
  assign n27430 = ( n5488 & n8372 ) | ( n5488 & ~n25829 ) | ( n8372 & ~n25829 ) ;
  assign n27429 = n23696 ^ n23050 ^ n11753 ;
  assign n27431 = n27430 ^ n27429 ^ n3469 ;
  assign n27432 = ( n2441 & ~n8330 ) | ( n2441 & n15521 ) | ( ~n8330 & n15521 ) ;
  assign n27433 = ( n8788 & n15709 ) | ( n8788 & n27432 ) | ( n15709 & n27432 ) ;
  assign n27434 = n27433 ^ n14136 ^ n9173 ;
  assign n27435 = n8268 ^ n7162 ^ n5844 ;
  assign n27436 = n27435 ^ n22029 ^ n16410 ;
  assign n27437 = ( ~n911 & n6664 ) | ( ~n911 & n27436 ) | ( n6664 & n27436 ) ;
  assign n27438 = n20363 ^ n16128 ^ n10673 ;
  assign n27439 = n27438 ^ n14020 ^ n1947 ;
  assign n27440 = n27439 ^ n21302 ^ n11875 ;
  assign n27444 = n8553 ^ n6631 ^ n3870 ;
  assign n27441 = ( n379 & n17082 ) | ( n379 & n23611 ) | ( n17082 & n23611 ) ;
  assign n27442 = n27441 ^ n11477 ^ n10532 ;
  assign n27443 = n27442 ^ n21059 ^ n6092 ;
  assign n27445 = n27444 ^ n27443 ^ n7858 ;
  assign n27446 = ( n1042 & n5291 ) | ( n1042 & n9093 ) | ( n5291 & n9093 ) ;
  assign n27447 = ( ~n2906 & n12958 ) | ( ~n2906 & n14687 ) | ( n12958 & n14687 ) ;
  assign n27448 = n8268 ^ n4993 ^ n1044 ;
  assign n27449 = n24546 ^ n23443 ^ n9519 ;
  assign n27450 = n20279 ^ n19752 ^ n3707 ;
  assign n27451 = ( n4862 & n6263 ) | ( n4862 & ~n27450 ) | ( n6263 & ~n27450 ) ;
  assign n27452 = ( n4850 & n24307 ) | ( n4850 & ~n27451 ) | ( n24307 & ~n27451 ) ;
  assign n27453 = n27452 ^ n23082 ^ n15398 ;
  assign n27454 = ( n2687 & ~n12087 ) | ( n2687 & n20771 ) | ( ~n12087 & n20771 ) ;
  assign n27456 = ( n144 & n3816 ) | ( n144 & n8743 ) | ( n3816 & n8743 ) ;
  assign n27455 = ( n10266 & ~n15490 ) | ( n10266 & n25631 ) | ( ~n15490 & n25631 ) ;
  assign n27457 = n27456 ^ n27455 ^ n25943 ;
  assign n27458 = n19583 ^ n13245 ^ n11318 ;
  assign n27459 = ( n4459 & n5867 ) | ( n4459 & n26637 ) | ( n5867 & n26637 ) ;
  assign n27460 = n27234 ^ n22557 ^ n14852 ;
  assign n27461 = n7380 ^ n4732 ^ n252 ;
  assign n27462 = n27461 ^ n12558 ^ n7164 ;
  assign n27463 = ( ~n637 & n8112 ) | ( ~n637 & n19029 ) | ( n8112 & n19029 ) ;
  assign n27464 = n20409 ^ n10790 ^ n8185 ;
  assign n27465 = n27464 ^ n22909 ^ n7150 ;
  assign n27466 = ( n4301 & n4868 ) | ( n4301 & ~n18148 ) | ( n4868 & ~n18148 ) ;
  assign n27467 = ( n4757 & n5436 ) | ( n4757 & ~n19985 ) | ( n5436 & ~n19985 ) ;
  assign n27468 = n26637 ^ n12251 ^ n11844 ;
  assign n27469 = ( n4623 & n11546 ) | ( n4623 & ~n27468 ) | ( n11546 & ~n27468 ) ;
  assign n27470 = n22511 ^ n10226 ^ n7640 ;
  assign n27471 = n14781 ^ n2766 ^ n939 ;
  assign n27472 = n27471 ^ n14707 ^ n10677 ;
  assign n27473 = ( n7471 & n8433 ) | ( n7471 & n24091 ) | ( n8433 & n24091 ) ;
  assign n27474 = ( ~n2502 & n5511 ) | ( ~n2502 & n27473 ) | ( n5511 & n27473 ) ;
  assign n27475 = ( n6427 & ~n15061 ) | ( n6427 & n16789 ) | ( ~n15061 & n16789 ) ;
  assign n27476 = ( n7094 & ~n9364 ) | ( n7094 & n27475 ) | ( ~n9364 & n27475 ) ;
  assign n27477 = n26307 ^ n10728 ^ n8799 ;
  assign n27478 = ( n1109 & n13400 ) | ( n1109 & ~n21811 ) | ( n13400 & ~n21811 ) ;
  assign n27479 = n15793 ^ n6704 ^ n3577 ;
  assign n27480 = n27479 ^ n26751 ^ n12190 ;
  assign n27481 = ( n5687 & n14331 ) | ( n5687 & n25623 ) | ( n14331 & n25623 ) ;
  assign n27482 = ( n1552 & ~n9391 ) | ( n1552 & n11840 ) | ( ~n9391 & n11840 ) ;
  assign n27483 = n27482 ^ n10623 ^ n3553 ;
  assign n27484 = n16411 ^ n15388 ^ n3068 ;
  assign n27485 = n11999 ^ n10306 ^ n10025 ;
  assign n27486 = ( n19211 & n27484 ) | ( n19211 & ~n27485 ) | ( n27484 & ~n27485 ) ;
  assign n27487 = ( ~n14255 & n18583 ) | ( ~n14255 & n27486 ) | ( n18583 & n27486 ) ;
  assign n27488 = n8439 ^ n8339 ^ n1763 ;
  assign n27489 = n23404 ^ n16072 ^ n11596 ;
  assign n27490 = ( n14177 & n16213 ) | ( n14177 & n27489 ) | ( n16213 & n27489 ) ;
  assign n27491 = ( ~n1090 & n5414 ) | ( ~n1090 & n10724 ) | ( n5414 & n10724 ) ;
  assign n27492 = ( ~n8570 & n17305 ) | ( ~n8570 & n27491 ) | ( n17305 & n27491 ) ;
  assign n27493 = ( ~n11844 & n22927 ) | ( ~n11844 & n23023 ) | ( n22927 & n23023 ) ;
  assign n27494 = n9684 ^ n7041 ^ n753 ;
  assign n27495 = n17187 ^ n7752 ^ n6288 ;
  assign n27496 = ( ~n18187 & n27494 ) | ( ~n18187 & n27495 ) | ( n27494 & n27495 ) ;
  assign n27497 = n27496 ^ n19100 ^ n10395 ;
  assign n27498 = n15612 ^ n6232 ^ n6202 ;
  assign n27499 = ( n9376 & ~n10275 ) | ( n9376 & n27498 ) | ( ~n10275 & n27498 ) ;
  assign n27500 = ( ~n4795 & n16515 ) | ( ~n4795 & n25685 ) | ( n16515 & n25685 ) ;
  assign n27501 = n9601 ^ n1773 ^ n1772 ;
  assign n27502 = n18242 ^ n14311 ^ n7248 ;
  assign n27503 = n27502 ^ n11352 ^ n1349 ;
  assign n27504 = n19579 ^ n11318 ^ n10431 ;
  assign n27505 = ( n6330 & ~n9047 ) | ( n6330 & n13538 ) | ( ~n9047 & n13538 ) ;
  assign n27506 = ( n16710 & n27504 ) | ( n16710 & n27505 ) | ( n27504 & n27505 ) ;
  assign n27507 = n25107 ^ n16336 ^ n10174 ;
  assign n27508 = ( n5858 & ~n8100 ) | ( n5858 & n27507 ) | ( ~n8100 & n27507 ) ;
  assign n27509 = n24517 ^ n14600 ^ n12307 ;
  assign n27510 = ( ~n6941 & n16207 ) | ( ~n6941 & n20235 ) | ( n16207 & n20235 ) ;
  assign n27511 = ( ~n2048 & n7945 ) | ( ~n2048 & n13774 ) | ( n7945 & n13774 ) ;
  assign n27512 = n27511 ^ n11447 ^ n2721 ;
  assign n27513 = ( n5851 & n10419 ) | ( n5851 & n20478 ) | ( n10419 & n20478 ) ;
  assign n27514 = n27513 ^ n25010 ^ n7301 ;
  assign n27515 = n18564 ^ n13868 ^ n5303 ;
  assign n27516 = ( n3893 & n16806 ) | ( n3893 & ~n27515 ) | ( n16806 & ~n27515 ) ;
  assign n27517 = n27516 ^ n20899 ^ n10230 ;
  assign n27518 = n27517 ^ n16388 ^ n5146 ;
  assign n27519 = ( n10808 & ~n14220 ) | ( n10808 & n24307 ) | ( ~n14220 & n24307 ) ;
  assign n27520 = ( n1016 & n17275 ) | ( n1016 & ~n26902 ) | ( n17275 & ~n26902 ) ;
  assign n27521 = ( n21336 & ~n23696 ) | ( n21336 & n27520 ) | ( ~n23696 & n27520 ) ;
  assign n27522 = n27521 ^ n20530 ^ n255 ;
  assign n27524 = ( n3501 & n7787 ) | ( n3501 & n26466 ) | ( n7787 & n26466 ) ;
  assign n27525 = ( n4144 & n15594 ) | ( n4144 & n23010 ) | ( n15594 & n23010 ) ;
  assign n27526 = ( n13400 & n27524 ) | ( n13400 & n27525 ) | ( n27524 & n27525 ) ;
  assign n27523 = n24189 ^ n6890 ^ n3577 ;
  assign n27527 = n27526 ^ n27523 ^ n8473 ;
  assign n27528 = n27527 ^ n12216 ^ n5485 ;
  assign n27530 = ( ~n2778 & n6368 ) | ( ~n2778 & n13419 ) | ( n6368 & n13419 ) ;
  assign n27529 = n24708 ^ n17137 ^ n2855 ;
  assign n27531 = n27530 ^ n27529 ^ n24149 ;
  assign n27532 = ( n11326 & n25736 ) | ( n11326 & n27531 ) | ( n25736 & n27531 ) ;
  assign n27533 = ( n841 & n4354 ) | ( n841 & n25083 ) | ( n4354 & n25083 ) ;
  assign n27534 = ( ~n5383 & n19916 ) | ( ~n5383 & n27533 ) | ( n19916 & n27533 ) ;
  assign n27535 = ( n2749 & n18924 ) | ( n2749 & n27534 ) | ( n18924 & n27534 ) ;
  assign n27536 = n15134 ^ n12091 ^ n6213 ;
  assign n27537 = ( n1091 & n8417 ) | ( n1091 & n19781 ) | ( n8417 & n19781 ) ;
  assign n27538 = n27537 ^ n25733 ^ n1441 ;
  assign n27539 = ( n6846 & n22939 ) | ( n6846 & ~n27538 ) | ( n22939 & ~n27538 ) ;
  assign n27541 = n12317 ^ n10837 ^ n1575 ;
  assign n27542 = ( ~n11616 & n20919 ) | ( ~n11616 & n27541 ) | ( n20919 & n27541 ) ;
  assign n27540 = n19953 ^ n17256 ^ n4308 ;
  assign n27543 = n27542 ^ n27540 ^ n8702 ;
  assign n27544 = n14664 ^ n5703 ^ n2459 ;
  assign n27545 = ( ~n13536 & n16815 ) | ( ~n13536 & n17144 ) | ( n16815 & n17144 ) ;
  assign n27546 = ( n608 & n1869 ) | ( n608 & n26505 ) | ( n1869 & n26505 ) ;
  assign n27547 = ( n7714 & ~n9163 ) | ( n7714 & n9831 ) | ( ~n9163 & n9831 ) ;
  assign n27548 = ( n282 & ~n615 ) | ( n282 & n2727 ) | ( ~n615 & n2727 ) ;
  assign n27549 = n27548 ^ n19179 ^ n1958 ;
  assign n27550 = ( n846 & n13932 ) | ( n846 & n27549 ) | ( n13932 & n27549 ) ;
  assign n27551 = ( n13872 & n17980 ) | ( n13872 & n27550 ) | ( n17980 & n27550 ) ;
  assign n27552 = ( n3374 & ~n9636 ) | ( n3374 & n19790 ) | ( ~n9636 & n19790 ) ;
  assign n27553 = n12867 ^ n11377 ^ n1109 ;
  assign n27554 = n27553 ^ n16819 ^ n14909 ;
  assign n27555 = n22840 ^ n12483 ^ n2126 ;
  assign n27556 = n27555 ^ n21416 ^ n14313 ;
  assign n27557 = n17395 ^ n11961 ^ n2966 ;
  assign n27558 = ( n4210 & ~n9149 ) | ( n4210 & n11428 ) | ( ~n9149 & n11428 ) ;
  assign n27559 = ( n2193 & n3985 ) | ( n2193 & n27558 ) | ( n3985 & n27558 ) ;
  assign n27560 = ( n871 & n4708 ) | ( n871 & ~n27559 ) | ( n4708 & ~n27559 ) ;
  assign n27561 = ( n9091 & n16129 ) | ( n9091 & n27560 ) | ( n16129 & n27560 ) ;
  assign n27562 = n27561 ^ n11071 ^ n9924 ;
  assign n27563 = n27562 ^ n22946 ^ n15895 ;
  assign n27564 = ( n1333 & ~n11311 ) | ( n1333 & n21974 ) | ( ~n11311 & n21974 ) ;
  assign n27565 = ( ~n12010 & n17595 ) | ( ~n12010 & n21941 ) | ( n17595 & n21941 ) ;
  assign n27566 = ( n906 & n7416 ) | ( n906 & ~n11154 ) | ( n7416 & ~n11154 ) ;
  assign n27567 = n27566 ^ n4354 ^ n3436 ;
  assign n27568 = n25195 ^ n10146 ^ n8524 ;
  assign n27569 = ( n13151 & n27567 ) | ( n13151 & ~n27568 ) | ( n27567 & ~n27568 ) ;
  assign n27570 = n27057 ^ n20265 ^ n2458 ;
  assign n27571 = n17674 ^ n3902 ^ n898 ;
  assign n27572 = n26118 ^ n19138 ^ n14536 ;
  assign n27573 = n27572 ^ n24435 ^ n23743 ;
  assign n27574 = n7613 ^ n7424 ^ n4943 ;
  assign n27575 = ( n4463 & ~n14380 ) | ( n4463 & n14848 ) | ( ~n14380 & n14848 ) ;
  assign n27576 = ( ~n7238 & n8601 ) | ( ~n7238 & n27575 ) | ( n8601 & n27575 ) ;
  assign n27577 = n19972 ^ n9050 ^ n2080 ;
  assign n27578 = ( ~n2050 & n14924 ) | ( ~n2050 & n18360 ) | ( n14924 & n18360 ) ;
  assign n27579 = ( ~n12546 & n27577 ) | ( ~n12546 & n27578 ) | ( n27577 & n27578 ) ;
  assign n27580 = n27579 ^ n16217 ^ n1841 ;
  assign n27581 = ( n2016 & n5478 ) | ( n2016 & n8333 ) | ( n5478 & n8333 ) ;
  assign n27582 = ( n331 & n2646 ) | ( n331 & n5331 ) | ( n2646 & n5331 ) ;
  assign n27583 = ( n1002 & n3812 ) | ( n1002 & n27582 ) | ( n3812 & n27582 ) ;
  assign n27584 = ( n19469 & n19714 ) | ( n19469 & ~n27583 ) | ( n19714 & ~n27583 ) ;
  assign n27585 = ( n15107 & n18837 ) | ( n15107 & n27146 ) | ( n18837 & n27146 ) ;
  assign n27586 = ( n13769 & n14744 ) | ( n13769 & ~n16401 ) | ( n14744 & ~n16401 ) ;
  assign n27587 = ( n6176 & ~n22081 ) | ( n6176 & n27586 ) | ( ~n22081 & n27586 ) ;
  assign n27588 = ( n3193 & ~n20193 ) | ( n3193 & n22825 ) | ( ~n20193 & n22825 ) ;
  assign n27589 = ( ~n519 & n11029 ) | ( ~n519 & n27588 ) | ( n11029 & n27588 ) ;
  assign n27590 = ( ~n3509 & n8727 ) | ( ~n3509 & n20599 ) | ( n8727 & n20599 ) ;
  assign n27591 = ( ~n12668 & n13347 ) | ( ~n12668 & n27590 ) | ( n13347 & n27590 ) ;
  assign n27592 = ( n11224 & ~n16311 ) | ( n11224 & n17549 ) | ( ~n16311 & n17549 ) ;
  assign n27593 = n25180 ^ n11515 ^ n6736 ;
  assign n27594 = ( n11969 & n26913 ) | ( n11969 & ~n27593 ) | ( n26913 & ~n27593 ) ;
  assign n27595 = n25591 ^ n10114 ^ n8348 ;
  assign n27596 = ( n3450 & ~n16475 ) | ( n3450 & n24507 ) | ( ~n16475 & n24507 ) ;
  assign n27597 = n27596 ^ n17683 ^ n9006 ;
  assign n27598 = ( n5536 & n27595 ) | ( n5536 & n27597 ) | ( n27595 & n27597 ) ;
  assign n27599 = ( n18550 & ~n20228 ) | ( n18550 & n27598 ) | ( ~n20228 & n27598 ) ;
  assign n27600 = n22526 ^ n15687 ^ n7725 ;
  assign n27601 = ( n2441 & ~n20303 ) | ( n2441 & n27600 ) | ( ~n20303 & n27600 ) ;
  assign n27602 = n27601 ^ n21532 ^ n7826 ;
  assign n27603 = n18596 ^ n9568 ^ n5933 ;
  assign n27604 = n27603 ^ n19179 ^ n7575 ;
  assign n27605 = ( ~n406 & n9506 ) | ( ~n406 & n17822 ) | ( n9506 & n17822 ) ;
  assign n27607 = ( n4383 & ~n5027 ) | ( n4383 & n5215 ) | ( ~n5027 & n5215 ) ;
  assign n27606 = n21888 ^ n16175 ^ n9589 ;
  assign n27608 = n27607 ^ n27606 ^ n23746 ;
  assign n27609 = ( ~n27604 & n27605 ) | ( ~n27604 & n27608 ) | ( n27605 & n27608 ) ;
  assign n27610 = n15534 ^ n15115 ^ n9638 ;
  assign n27611 = n27610 ^ n19613 ^ n7447 ;
  assign n27612 = ( n17632 & ~n17773 ) | ( n17632 & n27611 ) | ( ~n17773 & n27611 ) ;
  assign n27613 = n24718 ^ n9426 ^ n412 ;
  assign n27614 = n27613 ^ n18983 ^ n6930 ;
  assign n27615 = ( ~n26541 & n26601 ) | ( ~n26541 & n27614 ) | ( n26601 & n27614 ) ;
  assign n27616 = ( n8876 & ~n10882 ) | ( n8876 & n11916 ) | ( ~n10882 & n11916 ) ;
  assign n27619 = ( n3145 & ~n17479 ) | ( n3145 & n26242 ) | ( ~n17479 & n26242 ) ;
  assign n27617 = n10998 ^ n9080 ^ n3127 ;
  assign n27618 = n27617 ^ n8288 ^ n5325 ;
  assign n27620 = n27619 ^ n27618 ^ n20573 ;
  assign n27621 = n19512 ^ n10249 ^ n7947 ;
  assign n27622 = ( ~n5299 & n17341 ) | ( ~n5299 & n27621 ) | ( n17341 & n27621 ) ;
  assign n27623 = ( n879 & ~n19980 ) | ( n879 & n25148 ) | ( ~n19980 & n25148 ) ;
  assign n27624 = n18506 ^ n6928 ^ x12 ;
  assign n27625 = n9268 ^ n8913 ^ n5344 ;
  assign n27626 = ( ~n10504 & n19586 ) | ( ~n10504 & n24054 ) | ( n19586 & n24054 ) ;
  assign n27627 = ( ~n7131 & n9525 ) | ( ~n7131 & n27626 ) | ( n9525 & n27626 ) ;
  assign n27630 = n22842 ^ n10036 ^ n5106 ;
  assign n27628 = ( n3092 & ~n12688 ) | ( n3092 & n14204 ) | ( ~n12688 & n14204 ) ;
  assign n27629 = ( n13232 & ~n20539 ) | ( n13232 & n27628 ) | ( ~n20539 & n27628 ) ;
  assign n27631 = n27630 ^ n27629 ^ n17529 ;
  assign n27632 = n6247 ^ n4559 ^ n2379 ;
  assign n27633 = n27632 ^ n8126 ^ n2328 ;
  assign n27634 = n27633 ^ n23618 ^ n2259 ;
  assign n27635 = n25159 ^ n19278 ^ n2744 ;
  assign n27636 = ( ~n12064 & n21252 ) | ( ~n12064 & n27635 ) | ( n21252 & n27635 ) ;
  assign n27637 = n19211 ^ n13866 ^ n4271 ;
  assign n27638 = ( n7687 & n9176 ) | ( n7687 & n19714 ) | ( n9176 & n19714 ) ;
  assign n27640 = n9423 ^ n4381 ^ n2713 ;
  assign n27639 = ( n4976 & ~n22468 ) | ( n4976 & n27264 ) | ( ~n22468 & n27264 ) ;
  assign n27641 = n27640 ^ n27639 ^ n19330 ;
  assign n27644 = n16719 ^ n14508 ^ n2829 ;
  assign n27643 = n26845 ^ n22654 ^ n12388 ;
  assign n27642 = n12293 ^ n4247 ^ n3316 ;
  assign n27645 = n27644 ^ n27643 ^ n27642 ;
  assign n27646 = ( ~n1087 & n3414 ) | ( ~n1087 & n10301 ) | ( n3414 & n10301 ) ;
  assign n27647 = ( n138 & n14334 ) | ( n138 & n19764 ) | ( n14334 & n19764 ) ;
  assign n27648 = ( n4711 & n9704 ) | ( n4711 & n11154 ) | ( n9704 & n11154 ) ;
  assign n27649 = ( ~n9922 & n10442 ) | ( ~n9922 & n27648 ) | ( n10442 & n27648 ) ;
  assign n27650 = ( n1269 & n9418 ) | ( n1269 & ~n24835 ) | ( n9418 & ~n24835 ) ;
  assign n27651 = n22873 ^ n21600 ^ n13026 ;
  assign n27652 = ( n2627 & n7867 ) | ( n2627 & n17990 ) | ( n7867 & n17990 ) ;
  assign n27653 = ( n2080 & n6552 ) | ( n2080 & ~n27652 ) | ( n6552 & ~n27652 ) ;
  assign n27654 = n26404 ^ n6153 ^ n519 ;
  assign n27655 = ( n10003 & n15836 ) | ( n10003 & ~n27489 ) | ( n15836 & ~n27489 ) ;
  assign n27657 = ( n2570 & n19163 ) | ( n2570 & n19749 ) | ( n19163 & n19749 ) ;
  assign n27656 = n11427 ^ n8079 ^ n4048 ;
  assign n27658 = n27657 ^ n27656 ^ n26982 ;
  assign n27659 = ( n11384 & ~n12466 ) | ( n11384 & n27658 ) | ( ~n12466 & n27658 ) ;
  assign n27663 = n10660 ^ n7502 ^ n332 ;
  assign n27661 = n23549 ^ n16718 ^ n8386 ;
  assign n27662 = ( ~n3223 & n6963 ) | ( ~n3223 & n27661 ) | ( n6963 & n27661 ) ;
  assign n27660 = n18016 ^ n11153 ^ n7619 ;
  assign n27664 = n27663 ^ n27662 ^ n27660 ;
  assign n27665 = ( n5360 & ~n9352 ) | ( n5360 & n15222 ) | ( ~n9352 & n15222 ) ;
  assign n27666 = n27665 ^ n26067 ^ n3282 ;
  assign n27667 = n26516 ^ n7016 ^ n4136 ;
  assign n27668 = n6836 ^ n6830 ^ n1262 ;
  assign n27669 = ( n20962 & n25780 ) | ( n20962 & ~n27668 ) | ( n25780 & ~n27668 ) ;
  assign n27670 = ( n9993 & ~n27667 ) | ( n9993 & n27669 ) | ( ~n27667 & n27669 ) ;
  assign n27671 = n17830 ^ n3701 ^ n2224 ;
  assign n27672 = n27671 ^ n1838 ^ n1148 ;
  assign n27673 = ( ~n2896 & n16905 ) | ( ~n2896 & n27672 ) | ( n16905 & n27672 ) ;
  assign n27674 = ( n9811 & n19438 ) | ( n9811 & ~n21462 ) | ( n19438 & ~n21462 ) ;
  assign n27675 = ( n11377 & n23618 ) | ( n11377 & ~n27674 ) | ( n23618 & ~n27674 ) ;
  assign n27676 = ( n1623 & n6983 ) | ( n1623 & n21697 ) | ( n6983 & n21697 ) ;
  assign n27677 = ( n16197 & n24439 ) | ( n16197 & n27676 ) | ( n24439 & n27676 ) ;
  assign n27680 = ( ~x31 & n5916 ) | ( ~x31 & n15878 ) | ( n5916 & n15878 ) ;
  assign n27678 = n3722 ^ n2764 ^ n2525 ;
  assign n27679 = ( ~n7276 & n25866 ) | ( ~n7276 & n27678 ) | ( n25866 & n27678 ) ;
  assign n27681 = n27680 ^ n27679 ^ n4915 ;
  assign n27682 = ( n25177 & n27677 ) | ( n25177 & n27681 ) | ( n27677 & n27681 ) ;
  assign n27683 = ( n1900 & n6028 ) | ( n1900 & n13607 ) | ( n6028 & n13607 ) ;
  assign n27684 = ( n9728 & n13864 ) | ( n9728 & ~n20026 ) | ( n13864 & ~n20026 ) ;
  assign n27685 = n24684 ^ n10332 ^ n8019 ;
  assign n27686 = ( n19295 & ~n23329 ) | ( n19295 & n27685 ) | ( ~n23329 & n27685 ) ;
  assign n27687 = ( n18762 & ~n20074 ) | ( n18762 & n27686 ) | ( ~n20074 & n27686 ) ;
  assign n27688 = n25943 ^ n5305 ^ n4611 ;
  assign n27689 = ( n9340 & n15322 ) | ( n9340 & n23615 ) | ( n15322 & n23615 ) ;
  assign n27690 = n27689 ^ n15698 ^ n7063 ;
  assign n27691 = ( x31 & n301 ) | ( x31 & n2185 ) | ( n301 & n2185 ) ;
  assign n27692 = n27691 ^ n18725 ^ n8441 ;
  assign n27693 = n23980 ^ n22131 ^ n14016 ;
  assign n27694 = ( n1286 & n5939 ) | ( n1286 & n27693 ) | ( n5939 & n27693 ) ;
  assign n27695 = n17621 ^ n7106 ^ n6738 ;
  assign n27696 = ( n1539 & n15232 ) | ( n1539 & ~n27695 ) | ( n15232 & ~n27695 ) ;
  assign n27697 = ( ~n576 & n9986 ) | ( ~n576 & n27696 ) | ( n9986 & n27696 ) ;
  assign n27698 = ( ~n2399 & n2739 ) | ( ~n2399 & n27697 ) | ( n2739 & n27697 ) ;
  assign n27699 = n18844 ^ n14889 ^ n5364 ;
  assign n27700 = ( ~n3392 & n4843 ) | ( ~n3392 & n7594 ) | ( n4843 & n7594 ) ;
  assign n27701 = n27700 ^ n17298 ^ n6086 ;
  assign n27702 = ( n4205 & n11871 ) | ( n4205 & n15433 ) | ( n11871 & n15433 ) ;
  assign n27703 = ( n5471 & ~n7196 ) | ( n5471 & n10507 ) | ( ~n7196 & n10507 ) ;
  assign n27704 = ( n1683 & n26264 ) | ( n1683 & ~n27703 ) | ( n26264 & ~n27703 ) ;
  assign n27705 = n12221 ^ n10937 ^ n3369 ;
  assign n27706 = n27705 ^ n16901 ^ n5074 ;
  assign n27707 = ( n6520 & n13524 ) | ( n6520 & n27706 ) | ( n13524 & n27706 ) ;
  assign n27708 = ( ~n16348 & n19887 ) | ( ~n16348 & n27707 ) | ( n19887 & n27707 ) ;
  assign n27709 = n27708 ^ n23371 ^ n9360 ;
  assign n27710 = n27709 ^ n8542 ^ n2494 ;
  assign n27711 = ( n6102 & n15719 ) | ( n6102 & n19364 ) | ( n15719 & n19364 ) ;
  assign n27712 = n27711 ^ n25507 ^ n13872 ;
  assign n27713 = ( n938 & n11488 ) | ( n938 & ~n12196 ) | ( n11488 & ~n12196 ) ;
  assign n27714 = ( n8390 & n10599 ) | ( n8390 & n27713 ) | ( n10599 & n27713 ) ;
  assign n27715 = n8099 ^ n4131 ^ n488 ;
  assign n27716 = ( n7505 & n20510 ) | ( n7505 & ~n27715 ) | ( n20510 & ~n27715 ) ;
  assign n27717 = ( ~n7940 & n11997 ) | ( ~n7940 & n27716 ) | ( n11997 & n27716 ) ;
  assign n27718 = n12787 ^ n12748 ^ n3936 ;
  assign n27719 = ( ~n4479 & n11457 ) | ( ~n4479 & n26383 ) | ( n11457 & n26383 ) ;
  assign n27720 = n21170 ^ n7681 ^ n987 ;
  assign n27721 = ( ~n5474 & n7184 ) | ( ~n5474 & n26509 ) | ( n7184 & n26509 ) ;
  assign n27722 = ( n8246 & n14737 ) | ( n8246 & n27721 ) | ( n14737 & n27721 ) ;
  assign n27723 = n9991 ^ n5679 ^ n4215 ;
  assign n27724 = ( n2195 & ~n2529 ) | ( n2195 & n7252 ) | ( ~n2529 & n7252 ) ;
  assign n27725 = ( n1212 & n27723 ) | ( n1212 & ~n27724 ) | ( n27723 & ~n27724 ) ;
  assign n27726 = n27725 ^ n12854 ^ n4310 ;
  assign n27727 = ( n9181 & n10811 ) | ( n9181 & ~n27726 ) | ( n10811 & ~n27726 ) ;
  assign n27728 = ( n7675 & n10125 ) | ( n7675 & n16288 ) | ( n10125 & n16288 ) ;
  assign n27729 = n27728 ^ n27640 ^ n26890 ;
  assign n27730 = ( ~n2664 & n24928 ) | ( ~n2664 & n27729 ) | ( n24928 & n27729 ) ;
  assign n27733 = ( n10033 & n21790 ) | ( n10033 & ~n21832 ) | ( n21790 & ~n21832 ) ;
  assign n27734 = ( n2710 & n17804 ) | ( n2710 & n27733 ) | ( n17804 & n27733 ) ;
  assign n27735 = ( n11597 & n14688 ) | ( n11597 & ~n27734 ) | ( n14688 & ~n27734 ) ;
  assign n27731 = n26014 ^ n8073 ^ n3335 ;
  assign n27732 = n27731 ^ n18617 ^ n12955 ;
  assign n27736 = n27735 ^ n27732 ^ n24783 ;
  assign n27737 = n15039 ^ n10997 ^ x50 ;
  assign n27738 = n24551 ^ n15200 ^ n10298 ;
  assign n27739 = n16796 ^ n8856 ^ n2236 ;
  assign n27740 = n26744 ^ n13790 ^ n13409 ;
  assign n27741 = n27740 ^ n27156 ^ n23755 ;
  assign n27742 = n22148 ^ n19430 ^ n7995 ;
  assign n27743 = ( x54 & n9212 ) | ( x54 & n27742 ) | ( n9212 & n27742 ) ;
  assign n27744 = ( n1716 & n17525 ) | ( n1716 & ~n19680 ) | ( n17525 & ~n19680 ) ;
  assign n27745 = n27744 ^ n5133 ^ n2241 ;
  assign n27746 = n19982 ^ n12805 ^ n1254 ;
  assign n27747 = ( n797 & n13952 ) | ( n797 & ~n14714 ) | ( n13952 & ~n14714 ) ;
  assign n27748 = ( n13575 & n14290 ) | ( n13575 & ~n14371 ) | ( n14290 & ~n14371 ) ;
  assign n27749 = ( n7377 & n8383 ) | ( n7377 & n12511 ) | ( n8383 & n12511 ) ;
  assign n27750 = ( n3957 & n10606 ) | ( n3957 & n27749 ) | ( n10606 & n27749 ) ;
  assign n27751 = ( n182 & n6328 ) | ( n182 & ~n15534 ) | ( n6328 & ~n15534 ) ;
  assign n27752 = n26670 ^ n20284 ^ n6446 ;
  assign n27756 = ( n268 & n11498 ) | ( n268 & n15118 ) | ( n11498 & n15118 ) ;
  assign n27753 = ( n713 & n7864 ) | ( n713 & n13713 ) | ( n7864 & n13713 ) ;
  assign n27754 = ( n9131 & n10861 ) | ( n9131 & n17302 ) | ( n10861 & n17302 ) ;
  assign n27755 = ( n545 & n27753 ) | ( n545 & ~n27754 ) | ( n27753 & ~n27754 ) ;
  assign n27757 = n27756 ^ n27755 ^ n8332 ;
  assign n27758 = ( n16389 & n21693 ) | ( n16389 & ~n26162 ) | ( n21693 & ~n26162 ) ;
  assign n27759 = ( ~n14618 & n16423 ) | ( ~n14618 & n26729 ) | ( n16423 & n26729 ) ;
  assign n27760 = n15594 ^ n12426 ^ n4508 ;
  assign n27761 = ( ~n27758 & n27759 ) | ( ~n27758 & n27760 ) | ( n27759 & n27760 ) ;
  assign n27762 = n9073 ^ n5912 ^ n2384 ;
  assign n27763 = ( n366 & n22102 ) | ( n366 & n27762 ) | ( n22102 & n27762 ) ;
  assign n27766 = n11078 ^ n5588 ^ n2440 ;
  assign n27764 = n7826 ^ n2701 ^ n1904 ;
  assign n27765 = ( n176 & n9149 ) | ( n176 & n27764 ) | ( n9149 & n27764 ) ;
  assign n27767 = n27766 ^ n27765 ^ n7342 ;
  assign n27768 = ( ~n7620 & n10889 ) | ( ~n7620 & n17240 ) | ( n10889 & n17240 ) ;
  assign n27769 = ( ~n4722 & n8580 ) | ( ~n4722 & n11182 ) | ( n8580 & n11182 ) ;
  assign n27770 = n13081 ^ n9528 ^ x34 ;
  assign n27771 = n18731 ^ n14648 ^ n5939 ;
  assign n27772 = ( ~n20517 & n27770 ) | ( ~n20517 & n27771 ) | ( n27770 & n27771 ) ;
  assign n27773 = ( n12210 & ~n15279 ) | ( n12210 & n22193 ) | ( ~n15279 & n22193 ) ;
  assign n27774 = ( ~n11622 & n22446 ) | ( ~n11622 & n27773 ) | ( n22446 & n27773 ) ;
  assign n27775 = ( n8354 & n19691 ) | ( n8354 & n22038 ) | ( n19691 & n22038 ) ;
  assign n27783 = n22898 ^ n19127 ^ n11549 ;
  assign n27778 = ( n8207 & ~n17470 ) | ( n8207 & n26786 ) | ( ~n17470 & n26786 ) ;
  assign n27779 = n27778 ^ n7151 ^ n2988 ;
  assign n27780 = ( ~n8244 & n18038 ) | ( ~n8244 & n27779 ) | ( n18038 & n27779 ) ;
  assign n27776 = ( n2745 & ~n15953 ) | ( n2745 & n20748 ) | ( ~n15953 & n20748 ) ;
  assign n27777 = ( n13324 & n14445 ) | ( n13324 & n27776 ) | ( n14445 & n27776 ) ;
  assign n27781 = n27780 ^ n27777 ^ n8254 ;
  assign n27782 = n27781 ^ n12429 ^ n6220 ;
  assign n27784 = n27783 ^ n27782 ^ n24398 ;
  assign n27785 = n18014 ^ n8666 ^ n186 ;
  assign n27786 = ( n6518 & n11402 ) | ( n6518 & n13394 ) | ( n11402 & n13394 ) ;
  assign n27787 = n27786 ^ n4963 ^ n4703 ;
  assign n27788 = n27787 ^ n12163 ^ n11257 ;
  assign n27789 = ( ~n2822 & n18526 ) | ( ~n2822 & n27788 ) | ( n18526 & n27788 ) ;
  assign n27790 = ( n1596 & ~n12716 ) | ( n1596 & n21822 ) | ( ~n12716 & n21822 ) ;
  assign n27791 = ( n11493 & n21633 ) | ( n11493 & n26860 ) | ( n21633 & n26860 ) ;
  assign n27792 = n26617 ^ n9298 ^ n8986 ;
  assign n27793 = ( n516 & ~n13714 ) | ( n516 & n13928 ) | ( ~n13714 & n13928 ) ;
  assign n27794 = ( ~n6480 & n12811 ) | ( ~n6480 & n27793 ) | ( n12811 & n27793 ) ;
  assign n27795 = n27794 ^ n21714 ^ n16611 ;
  assign n27797 = ( n1473 & n9264 ) | ( n1473 & ~n16583 ) | ( n9264 & ~n16583 ) ;
  assign n27796 = n18565 ^ n17429 ^ n2810 ;
  assign n27798 = n27797 ^ n27796 ^ n12750 ;
  assign n27799 = ( n2998 & n5305 ) | ( n2998 & n21172 ) | ( n5305 & n21172 ) ;
  assign n27800 = n27799 ^ n25461 ^ n16055 ;
  assign n27801 = ( n19208 & ~n27798 ) | ( n19208 & n27800 ) | ( ~n27798 & n27800 ) ;
  assign n27802 = n27801 ^ n23017 ^ n1645 ;
  assign n27803 = n15499 ^ n6370 ^ n1224 ;
  assign n27804 = ( ~n3491 & n3860 ) | ( ~n3491 & n27803 ) | ( n3860 & n27803 ) ;
  assign n27805 = n15147 ^ n385 ^ n271 ;
  assign n27806 = ( n3940 & n17628 ) | ( n3940 & n21429 ) | ( n17628 & n21429 ) ;
  assign n27807 = n12748 ^ n5634 ^ n1188 ;
  assign n27808 = n27807 ^ n25178 ^ n11872 ;
  assign n27809 = ( n6308 & ~n25450 ) | ( n6308 & n26634 ) | ( ~n25450 & n26634 ) ;
  assign n27810 = n21616 ^ n13973 ^ n7992 ;
  assign n27812 = ( n4926 & n5228 ) | ( n4926 & n6914 ) | ( n5228 & n6914 ) ;
  assign n27811 = n22328 ^ n9500 ^ n1647 ;
  assign n27813 = n27812 ^ n27811 ^ n6872 ;
  assign n27814 = n27813 ^ n13389 ^ n2247 ;
  assign n27815 = n22213 ^ n2995 ^ n2530 ;
  assign n27816 = ( n8863 & ~n19232 ) | ( n8863 & n27815 ) | ( ~n19232 & n27815 ) ;
  assign n27817 = n5644 ^ n2495 ^ n605 ;
  assign n27818 = ( n7432 & n9764 ) | ( n7432 & n27817 ) | ( n9764 & n27817 ) ;
  assign n27819 = ( n3403 & n15439 ) | ( n3403 & ~n27818 ) | ( n15439 & ~n27818 ) ;
  assign n27820 = ( n5496 & n13598 ) | ( n5496 & ~n19248 ) | ( n13598 & ~n19248 ) ;
  assign n27821 = n27820 ^ n12652 ^ n1104 ;
  assign n27822 = n14755 ^ n10943 ^ n10089 ;
  assign n27823 = ( n589 & n1688 ) | ( n589 & ~n12888 ) | ( n1688 & ~n12888 ) ;
  assign n27824 = ( n764 & ~n2232 ) | ( n764 & n27823 ) | ( ~n2232 & n27823 ) ;
  assign n27825 = ( n11995 & ~n20618 ) | ( n11995 & n27824 ) | ( ~n20618 & n27824 ) ;
  assign n27826 = n27825 ^ n18136 ^ n6029 ;
  assign n27827 = n5973 ^ n3607 ^ n505 ;
  assign n27828 = ( n4828 & n4915 ) | ( n4828 & n27827 ) | ( n4915 & n27827 ) ;
  assign n27829 = ( n1341 & n2343 ) | ( n1341 & ~n27828 ) | ( n2343 & ~n27828 ) ;
  assign n27830 = n6837 ^ n545 ^ n180 ;
  assign n27831 = ( n2391 & n13546 ) | ( n2391 & n25207 ) | ( n13546 & n25207 ) ;
  assign n27832 = ( n8851 & ~n19495 ) | ( n8851 & n27831 ) | ( ~n19495 & n27831 ) ;
  assign n27833 = ( ~n4861 & n8823 ) | ( ~n4861 & n24198 ) | ( n8823 & n24198 ) ;
  assign n27834 = ( ~n361 & n21627 ) | ( ~n361 & n27833 ) | ( n21627 & n27833 ) ;
  assign n27835 = ( n3116 & n3930 ) | ( n3116 & ~n4059 ) | ( n3930 & ~n4059 ) ;
  assign n27836 = n27835 ^ n13365 ^ n6002 ;
  assign n27837 = n25716 ^ n7925 ^ n824 ;
  assign n27838 = ( n12754 & n16179 ) | ( n12754 & n25784 ) | ( n16179 & n25784 ) ;
  assign n27839 = ( n3203 & ~n23310 ) | ( n3203 & n27525 ) | ( ~n23310 & n27525 ) ;
  assign n27840 = n22469 ^ n5302 ^ n5016 ;
  assign n27843 = n15736 ^ n2560 ^ n1707 ;
  assign n27841 = n15169 ^ n8027 ^ n331 ;
  assign n27842 = n27841 ^ n24870 ^ n11862 ;
  assign n27844 = n27843 ^ n27842 ^ n20637 ;
  assign n27845 = ( n7022 & n16823 ) | ( n7022 & ~n19757 ) | ( n16823 & ~n19757 ) ;
  assign n27846 = n27845 ^ n11329 ^ n348 ;
  assign n27847 = ( x6 & ~n732 ) | ( x6 & n23463 ) | ( ~n732 & n23463 ) ;
  assign n27848 = n27847 ^ n12889 ^ n4689 ;
  assign n27852 = n25921 ^ n19634 ^ n12228 ;
  assign n27853 = n23035 ^ n13789 ^ n8860 ;
  assign n27854 = n27853 ^ n14714 ^ n11582 ;
  assign n27855 = ( ~n5116 & n14224 ) | ( ~n5116 & n24378 ) | ( n14224 & n24378 ) ;
  assign n27856 = n27855 ^ n6197 ^ n2084 ;
  assign n27857 = ( n27852 & n27854 ) | ( n27852 & n27856 ) | ( n27854 & n27856 ) ;
  assign n27850 = ( n1149 & ~n9691 ) | ( n1149 & n12932 ) | ( ~n9691 & n12932 ) ;
  assign n27849 = ( ~n6618 & n9918 ) | ( ~n6618 & n24187 ) | ( n9918 & n24187 ) ;
  assign n27851 = n27850 ^ n27849 ^ n22078 ;
  assign n27858 = n27857 ^ n27851 ^ n3242 ;
  assign n27859 = n25954 ^ n23058 ^ n3037 ;
  assign n27860 = n13324 ^ n7452 ^ n7349 ;
  assign n27861 = ( n9095 & ~n14508 ) | ( n9095 & n27860 ) | ( ~n14508 & n27860 ) ;
  assign n27862 = ( ~n8998 & n11529 ) | ( ~n8998 & n12275 ) | ( n11529 & n12275 ) ;
  assign n27863 = ( n14050 & ~n24398 ) | ( n14050 & n27862 ) | ( ~n24398 & n27862 ) ;
  assign n27864 = n17365 ^ n16328 ^ n6973 ;
  assign n27865 = ( n7195 & n8143 ) | ( n7195 & n11596 ) | ( n8143 & n11596 ) ;
  assign n27866 = n27865 ^ n19848 ^ n1342 ;
  assign n27867 = n22875 ^ n18623 ^ n10243 ;
  assign n27871 = n10763 ^ n9223 ^ n2563 ;
  assign n27869 = ( ~n327 & n7070 ) | ( ~n327 & n14109 ) | ( n7070 & n14109 ) ;
  assign n27870 = ( n7900 & n9053 ) | ( n7900 & n27869 ) | ( n9053 & n27869 ) ;
  assign n27872 = n27871 ^ n27870 ^ n14923 ;
  assign n27868 = ( n10735 & ~n11591 ) | ( n10735 & n11836 ) | ( ~n11591 & n11836 ) ;
  assign n27873 = n27872 ^ n27868 ^ n2973 ;
  assign n27874 = ( ~n8881 & n12789 ) | ( ~n8881 & n19126 ) | ( n12789 & n19126 ) ;
  assign n27875 = n27874 ^ n14960 ^ n14190 ;
  assign n27876 = n14460 ^ n4105 ^ x57 ;
  assign n27877 = n27876 ^ n18319 ^ n9054 ;
  assign n27878 = ( n503 & n21298 ) | ( n503 & ~n27877 ) | ( n21298 & ~n27877 ) ;
  assign n27879 = ( ~n13493 & n16239 ) | ( ~n13493 & n27878 ) | ( n16239 & n27878 ) ;
  assign n27880 = ( n10920 & n11990 ) | ( n10920 & n13468 ) | ( n11990 & n13468 ) ;
  assign n27881 = n19316 ^ n5538 ^ n938 ;
  assign n27882 = n27881 ^ n8360 ^ n8164 ;
  assign n27883 = n23349 ^ n9496 ^ n3977 ;
  assign n27884 = n27883 ^ n15553 ^ n10431 ;
  assign n27885 = ( ~n21258 & n27882 ) | ( ~n21258 & n27884 ) | ( n27882 & n27884 ) ;
  assign n27886 = n27371 ^ n23059 ^ n22817 ;
  assign n27887 = ( n912 & ~n19767 ) | ( n912 & n27886 ) | ( ~n19767 & n27886 ) ;
  assign n27888 = ( n5082 & n13269 ) | ( n5082 & ~n27887 ) | ( n13269 & ~n27887 ) ;
  assign n27889 = n27888 ^ n14133 ^ n8939 ;
  assign n27890 = n26619 ^ n26145 ^ n1147 ;
  assign n27891 = ( n1448 & n3422 ) | ( n1448 & n22938 ) | ( n3422 & n22938 ) ;
  assign n27892 = ( ~n4937 & n9788 ) | ( ~n4937 & n27891 ) | ( n9788 & n27891 ) ;
  assign n27893 = ( n10949 & n23984 ) | ( n10949 & n27892 ) | ( n23984 & n27892 ) ;
  assign n27894 = n27893 ^ n20689 ^ n15432 ;
  assign n27895 = ( n18365 & ~n20793 ) | ( n18365 & n26171 ) | ( ~n20793 & n26171 ) ;
  assign n27896 = n3296 ^ n1447 ^ n1248 ;
  assign n27897 = ( n7339 & ~n7945 ) | ( n7339 & n13104 ) | ( ~n7945 & n13104 ) ;
  assign n27898 = ( n17807 & ~n18264 ) | ( n17807 & n27897 ) | ( ~n18264 & n27897 ) ;
  assign n27899 = ( n5957 & ~n15437 ) | ( n5957 & n27898 ) | ( ~n15437 & n27898 ) ;
  assign n27900 = ( n14524 & n27896 ) | ( n14524 & n27899 ) | ( n27896 & n27899 ) ;
  assign n27901 = ( n821 & n6948 ) | ( n821 & ~n12102 ) | ( n6948 & ~n12102 ) ;
  assign n27902 = ( ~n1287 & n2131 ) | ( ~n1287 & n7890 ) | ( n2131 & n7890 ) ;
  assign n27903 = n27902 ^ n8173 ^ n510 ;
  assign n27904 = ( n8620 & n11536 ) | ( n8620 & n20463 ) | ( n11536 & n20463 ) ;
  assign n27905 = n27904 ^ n14850 ^ n8112 ;
  assign n27906 = n8222 ^ n1424 ^ n1392 ;
  assign n27909 = n9925 ^ n8438 ^ n7679 ;
  assign n27907 = ( n1804 & ~n7943 ) | ( n1804 & n17848 ) | ( ~n7943 & n17848 ) ;
  assign n27908 = n27907 ^ n12384 ^ n1307 ;
  assign n27910 = n27909 ^ n27908 ^ n22391 ;
  assign n27911 = ( ~n16733 & n27906 ) | ( ~n16733 & n27910 ) | ( n27906 & n27910 ) ;
  assign n27912 = ( n3969 & ~n15730 ) | ( n3969 & n18080 ) | ( ~n15730 & n18080 ) ;
  assign n27913 = n19530 ^ n7063 ^ n1462 ;
  assign n27914 = n27913 ^ n18264 ^ n4769 ;
  assign n27915 = n12256 ^ n9330 ^ n2476 ;
  assign n27916 = n16498 ^ n2923 ^ n1176 ;
  assign n27917 = n24088 ^ n20901 ^ n3517 ;
  assign n27918 = ( n12471 & ~n15671 ) | ( n12471 & n27917 ) | ( ~n15671 & n27917 ) ;
  assign n27919 = n19179 ^ n13163 ^ n9554 ;
  assign n27920 = n27919 ^ n7990 ^ n1735 ;
  assign n27921 = n27920 ^ n15399 ^ n8556 ;
  assign n27922 = ( ~n27916 & n27918 ) | ( ~n27916 & n27921 ) | ( n27918 & n27921 ) ;
  assign n27923 = ( n6063 & n7335 ) | ( n6063 & n9819 ) | ( n7335 & n9819 ) ;
  assign n27924 = ( n148 & n1847 ) | ( n148 & ~n6320 ) | ( n1847 & ~n6320 ) ;
  assign n27925 = ( ~n1841 & n27923 ) | ( ~n1841 & n27924 ) | ( n27923 & n27924 ) ;
  assign n27929 = ( x82 & n1252 ) | ( x82 & n13533 ) | ( n1252 & n13533 ) ;
  assign n27926 = n9704 ^ n7347 ^ n7108 ;
  assign n27927 = n17777 ^ n15223 ^ n2111 ;
  assign n27928 = ( n3764 & ~n27926 ) | ( n3764 & n27927 ) | ( ~n27926 & n27927 ) ;
  assign n27930 = n27929 ^ n27928 ^ n20505 ;
  assign n27931 = ( n8339 & ~n10429 ) | ( n8339 & n14899 ) | ( ~n10429 & n14899 ) ;
  assign n27932 = n14718 ^ n8257 ^ n6690 ;
  assign n27933 = n24970 ^ n9112 ^ n5703 ;
  assign n27934 = ( n4751 & n10658 ) | ( n4751 & ~n27933 ) | ( n10658 & ~n27933 ) ;
  assign n27935 = ( n5366 & ~n15438 ) | ( n5366 & n25830 ) | ( ~n15438 & n25830 ) ;
  assign n27936 = ( n8884 & n9815 ) | ( n8884 & n27935 ) | ( n9815 & n27935 ) ;
  assign n27937 = n27196 ^ n25500 ^ n21143 ;
  assign n27938 = n14641 ^ n7367 ^ n1135 ;
  assign n27939 = ( ~n933 & n4348 ) | ( ~n933 & n27938 ) | ( n4348 & n27938 ) ;
  assign n27940 = ( n5384 & ~n6121 ) | ( n5384 & n14091 ) | ( ~n6121 & n14091 ) ;
  assign n27941 = n27940 ^ n17307 ^ n7816 ;
  assign n27942 = ( ~n2255 & n5724 ) | ( ~n2255 & n5937 ) | ( n5724 & n5937 ) ;
  assign n27943 = n27942 ^ n6203 ^ n3044 ;
  assign n27944 = n27943 ^ n4182 ^ n992 ;
  assign n27945 = n21661 ^ n9715 ^ n5474 ;
  assign n27946 = n19791 ^ n12269 ^ n4098 ;
  assign n27947 = ( n657 & n7822 ) | ( n657 & n27946 ) | ( n7822 & n27946 ) ;
  assign n27949 = ( n4415 & n6818 ) | ( n4415 & n8938 ) | ( n6818 & n8938 ) ;
  assign n27948 = ( n2207 & n3204 ) | ( n2207 & n13814 ) | ( n3204 & n13814 ) ;
  assign n27950 = n27949 ^ n27948 ^ n1432 ;
  assign n27951 = ( ~n12148 & n12802 ) | ( ~n12148 & n17389 ) | ( n12802 & n17389 ) ;
  assign n27952 = ( n1183 & n15375 ) | ( n1183 & ~n20853 ) | ( n15375 & ~n20853 ) ;
  assign n27954 = ( ~n9054 & n10073 ) | ( ~n9054 & n16988 ) | ( n10073 & n16988 ) ;
  assign n27953 = n13734 ^ n12972 ^ n1377 ;
  assign n27955 = n27954 ^ n27953 ^ n2438 ;
  assign n27956 = n24807 ^ n18000 ^ n11824 ;
  assign n27957 = n24412 ^ n4460 ^ n4117 ;
  assign n27958 = n27957 ^ n21591 ^ n5238 ;
  assign n27959 = ( n12282 & n12654 ) | ( n12282 & ~n18094 ) | ( n12654 & ~n18094 ) ;
  assign n27960 = n24951 ^ n18457 ^ n446 ;
  assign n27961 = ( n1841 & n16442 ) | ( n1841 & n23359 ) | ( n16442 & n23359 ) ;
  assign n27962 = ( n5709 & ~n18948 ) | ( n5709 & n27961 ) | ( ~n18948 & n27961 ) ;
  assign n27963 = ( n2563 & n10498 ) | ( n2563 & n16855 ) | ( n10498 & n16855 ) ;
  assign n27964 = n27963 ^ n15236 ^ n13790 ;
  assign n27965 = ( n3629 & n6532 ) | ( n3629 & ~n27964 ) | ( n6532 & ~n27964 ) ;
  assign n27966 = ( ~n1041 & n5997 ) | ( ~n1041 & n27965 ) | ( n5997 & n27965 ) ;
  assign n27967 = n24737 ^ n8431 ^ n5360 ;
  assign n27968 = ( ~n4825 & n10021 ) | ( ~n4825 & n14311 ) | ( n10021 & n14311 ) ;
  assign n27969 = n27968 ^ n20106 ^ n15355 ;
  assign n27970 = ( ~n6901 & n11557 ) | ( ~n6901 & n19126 ) | ( n11557 & n19126 ) ;
  assign n27971 = n19118 ^ n4942 ^ n3875 ;
  assign n27972 = ( n9559 & n11035 ) | ( n9559 & ~n27971 ) | ( n11035 & ~n27971 ) ;
  assign n27973 = n20580 ^ n19482 ^ n19310 ;
  assign n27974 = n25436 ^ n3192 ^ x110 ;
  assign n27975 = n27974 ^ n11391 ^ n5908 ;
  assign n27976 = ( n18067 & n27973 ) | ( n18067 & ~n27975 ) | ( n27973 & ~n27975 ) ;
  assign n27977 = ( n10371 & ~n13296 ) | ( n10371 & n21146 ) | ( ~n13296 & n21146 ) ;
  assign n27978 = n27977 ^ n9700 ^ n7995 ;
  assign n27979 = ( n7807 & ~n10355 ) | ( n7807 & n27978 ) | ( ~n10355 & n27978 ) ;
  assign n27980 = n8451 ^ n6276 ^ n6041 ;
  assign n27981 = n27980 ^ n25034 ^ n11982 ;
  assign n27982 = ( n12895 & n18846 ) | ( n12895 & n19293 ) | ( n18846 & n19293 ) ;
  assign n27983 = n17804 ^ n7238 ^ x6 ;
  assign n27984 = ( n3650 & ~n11638 ) | ( n3650 & n27983 ) | ( ~n11638 & n27983 ) ;
  assign n27985 = n24555 ^ n16463 ^ n6117 ;
  assign n27986 = n27985 ^ n20062 ^ n15271 ;
  assign n27987 = ( n5257 & ~n27984 ) | ( n5257 & n27986 ) | ( ~n27984 & n27986 ) ;
  assign n27988 = n18038 ^ n14854 ^ n13506 ;
  assign n27991 = ( ~n11928 & n13543 ) | ( ~n11928 & n18002 ) | ( n13543 & n18002 ) ;
  assign n27989 = n21175 ^ n13134 ^ n5860 ;
  assign n27990 = n27989 ^ n17164 ^ x121 ;
  assign n27992 = n27991 ^ n27990 ^ n22101 ;
  assign n27993 = n12936 ^ n4311 ^ n3059 ;
  assign n27994 = ( ~n5061 & n16174 ) | ( ~n5061 & n22738 ) | ( n16174 & n22738 ) ;
  assign n27995 = n27994 ^ n4687 ^ n2009 ;
  assign n27998 = ( ~n6445 & n9377 ) | ( ~n6445 & n19701 ) | ( n9377 & n19701 ) ;
  assign n27996 = n9150 ^ n8137 ^ n5116 ;
  assign n27997 = n27996 ^ n14949 ^ n4666 ;
  assign n27999 = n27998 ^ n27997 ^ n3380 ;
  assign n28000 = n27999 ^ n10909 ^ n7380 ;
  assign n28001 = n19559 ^ n3343 ^ n2452 ;
  assign n28002 = n8470 ^ n5791 ^ n1846 ;
  assign n28003 = ( ~n4770 & n21210 ) | ( ~n4770 & n21768 ) | ( n21210 & n21768 ) ;
  assign n28004 = ( n26557 & n28002 ) | ( n26557 & ~n28003 ) | ( n28002 & ~n28003 ) ;
  assign n28005 = n7534 ^ n6598 ^ n2248 ;
  assign n28006 = ( n4088 & ~n14904 ) | ( n4088 & n28005 ) | ( ~n14904 & n28005 ) ;
  assign n28007 = n28006 ^ n14520 ^ n5132 ;
  assign n28008 = n28007 ^ n8132 ^ n2865 ;
  assign n28009 = n12992 ^ n9152 ^ n1740 ;
  assign n28010 = ( n15073 & n19113 ) | ( n15073 & n28009 ) | ( n19113 & n28009 ) ;
  assign n28011 = ( ~n2072 & n8434 ) | ( ~n2072 & n10220 ) | ( n8434 & n10220 ) ;
  assign n28013 = n24991 ^ n19022 ^ n2247 ;
  assign n28012 = ( n1777 & n10243 ) | ( n1777 & ~n15601 ) | ( n10243 & ~n15601 ) ;
  assign n28014 = n28013 ^ n28012 ^ n25273 ;
  assign n28015 = ( n11377 & n28011 ) | ( n11377 & n28014 ) | ( n28011 & n28014 ) ;
  assign n28016 = ( n1882 & ~n12934 ) | ( n1882 & n24643 ) | ( ~n12934 & n24643 ) ;
  assign n28017 = ( n1155 & n17709 ) | ( n1155 & n27849 ) | ( n17709 & n27849 ) ;
  assign n28019 = n24931 ^ n15927 ^ n2102 ;
  assign n28018 = n26567 ^ n8132 ^ n2255 ;
  assign n28020 = n28019 ^ n28018 ^ n6031 ;
  assign n28021 = n28020 ^ n27279 ^ n16289 ;
  assign n28022 = n24668 ^ n14191 ^ n6221 ;
  assign n28023 = ( n2519 & n11241 ) | ( n2519 & n21333 ) | ( n11241 & n21333 ) ;
  assign n28024 = ( n8629 & ~n26744 ) | ( n8629 & n28023 ) | ( ~n26744 & n28023 ) ;
  assign n28025 = ( n9316 & n13141 ) | ( n9316 & ~n14904 ) | ( n13141 & ~n14904 ) ;
  assign n28026 = n28025 ^ n25720 ^ n18159 ;
  assign n28027 = ( n5708 & n7099 ) | ( n5708 & ~n8536 ) | ( n7099 & ~n8536 ) ;
  assign n28028 = n14591 ^ n8003 ^ n7455 ;
  assign n28029 = n25888 ^ n7481 ^ n1706 ;
  assign n28030 = ( n20278 & n28028 ) | ( n20278 & ~n28029 ) | ( n28028 & ~n28029 ) ;
  assign n28031 = ( ~n17339 & n28027 ) | ( ~n17339 & n28030 ) | ( n28027 & n28030 ) ;
  assign n28032 = ( n1464 & ~n3067 ) | ( n1464 & n9772 ) | ( ~n3067 & n9772 ) ;
  assign n28033 = ( n25075 & n25407 ) | ( n25075 & ~n28032 ) | ( n25407 & ~n28032 ) ;
  assign n28034 = ( n5316 & n12342 ) | ( n5316 & ~n23552 ) | ( n12342 & ~n23552 ) ;
  assign n28035 = n12012 ^ n3035 ^ n2615 ;
  assign n28037 = n14505 ^ n6896 ^ n1840 ;
  assign n28036 = n9259 ^ n6604 ^ n3308 ;
  assign n28038 = n28037 ^ n28036 ^ n13139 ;
  assign n28039 = ( n10763 & n28035 ) | ( n10763 & ~n28038 ) | ( n28035 & ~n28038 ) ;
  assign n28040 = ( n12595 & n19979 ) | ( n12595 & ~n28039 ) | ( n19979 & ~n28039 ) ;
  assign n28041 = ( n1709 & n9615 ) | ( n1709 & n26452 ) | ( n9615 & n26452 ) ;
  assign n28042 = n28041 ^ n21770 ^ n6711 ;
  assign n28043 = n23459 ^ n20647 ^ n9241 ;
  assign n28044 = n26342 ^ n8005 ^ n5309 ;
  assign n28045 = n15555 ^ n6226 ^ n5157 ;
  assign n28046 = ( n13706 & ~n24846 ) | ( n13706 & n28045 ) | ( ~n24846 & n28045 ) ;
  assign n28047 = ( n22949 & ~n28044 ) | ( n22949 & n28046 ) | ( ~n28044 & n28046 ) ;
  assign n28048 = n8924 ^ n1265 ^ n220 ;
  assign n28049 = ( n1220 & n2874 ) | ( n1220 & n17907 ) | ( n2874 & n17907 ) ;
  assign n28050 = n28049 ^ n25275 ^ n3617 ;
  assign n28051 = ( ~n5668 & n28048 ) | ( ~n5668 & n28050 ) | ( n28048 & n28050 ) ;
  assign n28052 = ( n1370 & ~n6635 ) | ( n1370 & n10629 ) | ( ~n6635 & n10629 ) ;
  assign n28053 = ( ~n1850 & n8205 ) | ( ~n1850 & n18197 ) | ( n8205 & n18197 ) ;
  assign n28054 = ( n2691 & ~n28052 ) | ( n2691 & n28053 ) | ( ~n28052 & n28053 ) ;
  assign n28055 = n25440 ^ n16691 ^ n7924 ;
  assign n28056 = n25513 ^ n9127 ^ n6661 ;
  assign n28057 = n10927 ^ n7422 ^ n5796 ;
  assign n28058 = n7261 ^ n2881 ^ n913 ;
  assign n28059 = n28058 ^ n15580 ^ n14602 ;
  assign n28060 = ( n16553 & n28057 ) | ( n16553 & ~n28059 ) | ( n28057 & ~n28059 ) ;
  assign n28061 = n9544 ^ n9114 ^ n1795 ;
  assign n28062 = ( ~n22092 & n25247 ) | ( ~n22092 & n28061 ) | ( n25247 & n28061 ) ;
  assign n28063 = n26637 ^ n15028 ^ n11195 ;
  assign n28064 = n28063 ^ n28062 ^ n25147 ;
  assign n28065 = ( n23336 & ~n27560 ) | ( n23336 & n28064 ) | ( ~n27560 & n28064 ) ;
  assign n28066 = ( n3239 & ~n10434 ) | ( n3239 & n20420 ) | ( ~n10434 & n20420 ) ;
  assign n28067 = ( ~n28062 & n28065 ) | ( ~n28062 & n28066 ) | ( n28065 & n28066 ) ;
  assign n28068 = n21772 ^ n7523 ^ n6639 ;
  assign n28069 = n19128 ^ n14939 ^ n13205 ;
  assign n28070 = ( n16336 & n28068 ) | ( n16336 & ~n28069 ) | ( n28068 & ~n28069 ) ;
  assign n28071 = ( n15865 & n17549 ) | ( n15865 & n24617 ) | ( n17549 & n24617 ) ;
  assign n28072 = n22433 ^ n3473 ^ n2959 ;
  assign n28073 = n22647 ^ n14645 ^ n1343 ;
  assign n28074 = ( ~n530 & n4151 ) | ( ~n530 & n4515 ) | ( n4151 & n4515 ) ;
  assign n28075 = ( ~n9938 & n10502 ) | ( ~n9938 & n10870 ) | ( n10502 & n10870 ) ;
  assign n28076 = n28075 ^ n22022 ^ n9928 ;
  assign n28078 = n4466 ^ n3454 ^ n1767 ;
  assign n28077 = ( n2040 & n9203 ) | ( n2040 & ~n17421 ) | ( n9203 & ~n17421 ) ;
  assign n28079 = n28078 ^ n28077 ^ n11208 ;
  assign n28080 = n22319 ^ n17333 ^ n1068 ;
  assign n28081 = ( n571 & n638 ) | ( n571 & ~n15579 ) | ( n638 & ~n15579 ) ;
  assign n28082 = ( n5358 & n10563 ) | ( n5358 & n28081 ) | ( n10563 & n28081 ) ;
  assign n28083 = n26127 ^ n21369 ^ n18171 ;
  assign n28084 = n28083 ^ n12676 ^ n1919 ;
  assign n28085 = n12710 ^ n626 ^ x116 ;
  assign n28086 = ( ~n6324 & n10911 ) | ( ~n6324 & n28085 ) | ( n10911 & n28085 ) ;
  assign n28087 = ( ~n7874 & n10634 ) | ( ~n7874 & n28086 ) | ( n10634 & n28086 ) ;
  assign n28090 = n18152 ^ n15300 ^ n11042 ;
  assign n28088 = n21551 ^ n20321 ^ n10025 ;
  assign n28089 = n28088 ^ n10410 ^ n9089 ;
  assign n28091 = n28090 ^ n28089 ^ n26547 ;
  assign n28092 = n14031 ^ n13842 ^ n7939 ;
  assign n28093 = n28092 ^ n26339 ^ n12804 ;
  assign n28094 = ( n737 & ~n15272 ) | ( n737 & n19517 ) | ( ~n15272 & n19517 ) ;
  assign n28095 = n24833 ^ n23587 ^ n15337 ;
  assign n28096 = ( n8724 & ~n10480 ) | ( n8724 & n26143 ) | ( ~n10480 & n26143 ) ;
  assign n28097 = n25812 ^ n11433 ^ n2515 ;
  assign n28098 = ( n1098 & ~n13975 ) | ( n1098 & n28097 ) | ( ~n13975 & n28097 ) ;
  assign n28099 = n25378 ^ n13751 ^ n9106 ;
  assign n28100 = ( n12042 & n18498 ) | ( n12042 & n20728 ) | ( n18498 & n20728 ) ;
  assign n28101 = ( n18816 & ~n27129 ) | ( n18816 & n27409 ) | ( ~n27129 & n27409 ) ;
  assign n28102 = ( n4932 & ~n20984 ) | ( n4932 & n21181 ) | ( ~n20984 & n21181 ) ;
  assign n28103 = ( n1823 & ~n3027 ) | ( n1823 & n8159 ) | ( ~n3027 & n8159 ) ;
  assign n28104 = n16386 ^ n7649 ^ n1833 ;
  assign n28105 = n28104 ^ n12904 ^ n7486 ;
  assign n28106 = ( n188 & ~n5465 ) | ( n188 & n28105 ) | ( ~n5465 & n28105 ) ;
  assign n28107 = n28106 ^ n25178 ^ n8239 ;
  assign n28108 = ( n4539 & ~n8014 ) | ( n4539 & n11747 ) | ( ~n8014 & n11747 ) ;
  assign n28113 = n12518 ^ n9402 ^ n706 ;
  assign n28114 = ( n5610 & ~n10427 ) | ( n5610 & n28113 ) | ( ~n10427 & n28113 ) ;
  assign n28111 = n26007 ^ n10370 ^ n3984 ;
  assign n28112 = n28111 ^ n11652 ^ n8260 ;
  assign n28109 = n20790 ^ n7474 ^ n6701 ;
  assign n28110 = n28109 ^ n13063 ^ n5309 ;
  assign n28115 = n28114 ^ n28112 ^ n28110 ;
  assign n28116 = ( n6567 & n15575 ) | ( n6567 & ~n16583 ) | ( n15575 & ~n16583 ) ;
  assign n28117 = n20218 ^ n5034 ^ n3151 ;
  assign n28118 = ( n5237 & ~n15186 ) | ( n5237 & n28117 ) | ( ~n15186 & n28117 ) ;
  assign n28119 = ( n8032 & n8332 ) | ( n8032 & n24644 ) | ( n8332 & n24644 ) ;
  assign n28120 = ( n11281 & ~n14313 ) | ( n11281 & n27115 ) | ( ~n14313 & n27115 ) ;
  assign n28121 = n28120 ^ n9775 ^ n3737 ;
  assign n28122 = ( n4759 & ~n17901 ) | ( n4759 & n28121 ) | ( ~n17901 & n28121 ) ;
  assign n28123 = n28068 ^ n17809 ^ n13062 ;
  assign n28124 = ( n4574 & n10352 ) | ( n4574 & n28123 ) | ( n10352 & n28123 ) ;
  assign n28125 = ( n2233 & n20140 ) | ( n2233 & n22488 ) | ( n20140 & n22488 ) ;
  assign n28126 = n5403 ^ n3503 ^ n306 ;
  assign n28127 = ( n4518 & n8539 ) | ( n4518 & n28126 ) | ( n8539 & n28126 ) ;
  assign n28128 = ( ~n3394 & n28125 ) | ( ~n3394 & n28127 ) | ( n28125 & n28127 ) ;
  assign n28129 = ( n12800 & n15023 ) | ( n12800 & ~n19040 ) | ( n15023 & ~n19040 ) ;
  assign n28130 = ( n8432 & ~n18497 ) | ( n8432 & n28129 ) | ( ~n18497 & n28129 ) ;
  assign n28131 = n26317 ^ n11875 ^ n7008 ;
  assign n28132 = ( n13685 & n19245 ) | ( n13685 & n28131 ) | ( n19245 & n28131 ) ;
  assign n28133 = ( n6862 & n13402 ) | ( n6862 & ~n16407 ) | ( n13402 & ~n16407 ) ;
  assign n28134 = n28133 ^ n25982 ^ n2968 ;
  assign n28135 = ( n16816 & n19218 ) | ( n16816 & ~n28134 ) | ( n19218 & ~n28134 ) ;
  assign n28136 = ( ~n1778 & n6635 ) | ( ~n1778 & n20335 ) | ( n6635 & n20335 ) ;
  assign n28137 = n5103 ^ n638 ^ n286 ;
  assign n28138 = n24062 ^ n8280 ^ n531 ;
  assign n28139 = ( n276 & ~n21174 ) | ( n276 & n28138 ) | ( ~n21174 & n28138 ) ;
  assign n28140 = ( n28136 & n28137 ) | ( n28136 & ~n28139 ) | ( n28137 & ~n28139 ) ;
  assign n28141 = ( n1691 & n4410 ) | ( n1691 & n10624 ) | ( n4410 & n10624 ) ;
  assign n28142 = n7634 ^ n2641 ^ n380 ;
  assign n28143 = ( n27355 & ~n28141 ) | ( n27355 & n28142 ) | ( ~n28141 & n28142 ) ;
  assign n28144 = ( n3139 & ~n4992 ) | ( n3139 & n11706 ) | ( ~n4992 & n11706 ) ;
  assign n28145 = ( n1073 & ~n5990 ) | ( n1073 & n9542 ) | ( ~n5990 & n9542 ) ;
  assign n28146 = ( n15796 & n28144 ) | ( n15796 & ~n28145 ) | ( n28144 & ~n28145 ) ;
  assign n28147 = n28146 ^ n9907 ^ n4124 ;
  assign n28148 = ( n1280 & ~n7702 ) | ( n1280 & n14200 ) | ( ~n7702 & n14200 ) ;
  assign n28149 = ( n13510 & n28032 ) | ( n13510 & n28148 ) | ( n28032 & n28148 ) ;
  assign n28155 = ( n1786 & ~n11002 ) | ( n1786 & n12671 ) | ( ~n11002 & n12671 ) ;
  assign n28151 = ( n5241 & n9811 ) | ( n5241 & n16047 ) | ( n9811 & n16047 ) ;
  assign n28152 = n28151 ^ n21056 ^ n4070 ;
  assign n28150 = ( n6383 & n15083 ) | ( n6383 & n16078 ) | ( n15083 & n16078 ) ;
  assign n28153 = n28152 ^ n28150 ^ n2069 ;
  assign n28154 = n28153 ^ n25553 ^ n17743 ;
  assign n28156 = n28155 ^ n28154 ^ n14001 ;
  assign n28157 = ( n6897 & n22478 ) | ( n6897 & ~n22905 ) | ( n22478 & ~n22905 ) ;
  assign n28158 = n15494 ^ n10518 ^ n6714 ;
  assign n28159 = n28158 ^ n2388 ^ n485 ;
  assign n28160 = n25788 ^ n12214 ^ n6549 ;
  assign n28161 = n15381 ^ n12267 ^ x11 ;
  assign n28162 = ( n17180 & n18691 ) | ( n17180 & ~n28161 ) | ( n18691 & ~n28161 ) ;
  assign n28163 = ( n28159 & n28160 ) | ( n28159 & ~n28162 ) | ( n28160 & ~n28162 ) ;
  assign n28164 = n23678 ^ n9459 ^ n9109 ;
  assign n28165 = ( ~n2212 & n7265 ) | ( ~n2212 & n28164 ) | ( n7265 & n28164 ) ;
  assign n28166 = ( n10680 & n26531 ) | ( n10680 & n28165 ) | ( n26531 & n28165 ) ;
  assign n28167 = ( n545 & n7348 ) | ( n545 & n24816 ) | ( n7348 & n24816 ) ;
  assign n28168 = ( n10124 & n25513 ) | ( n10124 & n28167 ) | ( n25513 & n28167 ) ;
  assign n28169 = ( ~n3369 & n7615 ) | ( ~n3369 & n10212 ) | ( n7615 & n10212 ) ;
  assign n28170 = n28169 ^ n17925 ^ n8576 ;
  assign n28171 = n21296 ^ n6262 ^ n2923 ;
  assign n28172 = n20305 ^ n7199 ^ n2006 ;
  assign n28173 = ( n210 & n8544 ) | ( n210 & ~n27807 ) | ( n8544 & ~n27807 ) ;
  assign n28174 = n28173 ^ n17830 ^ n13332 ;
  assign n28175 = ( ~n1053 & n28172 ) | ( ~n1053 & n28174 ) | ( n28172 & n28174 ) ;
  assign n28176 = ( x24 & n5213 ) | ( x24 & n12587 ) | ( n5213 & n12587 ) ;
  assign n28177 = ( n7325 & n20301 ) | ( n7325 & n28176 ) | ( n20301 & n28176 ) ;
  assign n28178 = n28177 ^ n14128 ^ n6248 ;
  assign n28179 = n26786 ^ n10072 ^ x112 ;
  assign n28180 = n12324 ^ n8332 ^ n5646 ;
  assign n28181 = ( n5622 & n26693 ) | ( n5622 & n28180 ) | ( n26693 & n28180 ) ;
  assign n28182 = n24054 ^ n11396 ^ n6467 ;
  assign n28183 = n28182 ^ n17697 ^ n11373 ;
  assign n28184 = ( ~n11578 & n15499 ) | ( ~n11578 & n23867 ) | ( n15499 & n23867 ) ;
  assign n28185 = n25573 ^ n18269 ^ n11780 ;
  assign n28186 = n24765 ^ n17364 ^ n1586 ;
  assign n28187 = ( n8606 & n13715 ) | ( n8606 & n19673 ) | ( n13715 & n19673 ) ;
  assign n28188 = ( n1249 & n8647 ) | ( n1249 & ~n19165 ) | ( n8647 & ~n19165 ) ;
  assign n28189 = n28188 ^ n27943 ^ n15659 ;
  assign n28190 = ( n2955 & ~n9458 ) | ( n2955 & n12488 ) | ( ~n9458 & n12488 ) ;
  assign n28191 = n28190 ^ n24795 ^ n18970 ;
  assign n28193 = ( n3626 & ~n6999 ) | ( n3626 & n21514 ) | ( ~n6999 & n21514 ) ;
  assign n28192 = ( n5405 & n12495 ) | ( n5405 & ~n12588 ) | ( n12495 & ~n12588 ) ;
  assign n28194 = n28193 ^ n28192 ^ n8187 ;
  assign n28195 = ( n465 & ~n19033 ) | ( n465 & n24778 ) | ( ~n19033 & n24778 ) ;
  assign n28196 = n28195 ^ n19941 ^ n17773 ;
  assign n28199 = n9270 ^ n2765 ^ n1828 ;
  assign n28200 = ( n12142 & n22955 ) | ( n12142 & ~n28199 ) | ( n22955 & ~n28199 ) ;
  assign n28197 = n5844 ^ n4113 ^ n1689 ;
  assign n28198 = ( n8296 & n14985 ) | ( n8296 & n28197 ) | ( n14985 & n28197 ) ;
  assign n28201 = n28200 ^ n28198 ^ n18744 ;
  assign n28202 = ( n3508 & n6817 ) | ( n3508 & ~n7642 ) | ( n6817 & ~n7642 ) ;
  assign n28203 = n21873 ^ n5044 ^ n2215 ;
  assign n28204 = ( ~n23465 & n23877 ) | ( ~n23465 & n28203 ) | ( n23877 & n28203 ) ;
  assign n28205 = ( n12894 & n19314 ) | ( n12894 & n22233 ) | ( n19314 & n22233 ) ;
  assign n28206 = ( n9366 & n9865 ) | ( n9366 & ~n14243 ) | ( n9865 & ~n14243 ) ;
  assign n28207 = ( n2330 & n13439 ) | ( n2330 & ~n28206 ) | ( n13439 & ~n28206 ) ;
  assign n28208 = n20295 ^ n19739 ^ n18029 ;
  assign n28209 = ( n240 & n12016 ) | ( n240 & n28208 ) | ( n12016 & n28208 ) ;
  assign n28210 = ( n4616 & n11794 ) | ( n4616 & n14757 ) | ( n11794 & n14757 ) ;
  assign n28211 = ( n7289 & ~n26216 ) | ( n7289 & n26331 ) | ( ~n26216 & n26331 ) ;
  assign n28212 = ( n9620 & n19113 ) | ( n9620 & ~n24820 ) | ( n19113 & ~n24820 ) ;
  assign n28213 = ( n14439 & ~n23019 ) | ( n14439 & n23778 ) | ( ~n23019 & n23778 ) ;
  assign n28214 = n23691 ^ n4285 ^ n1935 ;
  assign n28215 = n20877 ^ n8933 ^ x74 ;
  assign n28216 = ( n15618 & n16519 ) | ( n15618 & ~n20515 ) | ( n16519 & ~n20515 ) ;
  assign n28217 = n28216 ^ n7044 ^ n3587 ;
  assign n28218 = ( n2137 & ~n3637 ) | ( n2137 & n6848 ) | ( ~n3637 & n6848 ) ;
  assign n28219 = n26018 ^ n22022 ^ n7794 ;
  assign n28220 = ( n5842 & ~n25355 ) | ( n5842 & n28219 ) | ( ~n25355 & n28219 ) ;
  assign n28221 = ( n11896 & ~n19106 ) | ( n11896 & n24555 ) | ( ~n19106 & n24555 ) ;
  assign n28222 = ( n17434 & ~n20569 ) | ( n17434 & n28221 ) | ( ~n20569 & n28221 ) ;
  assign n28223 = n28222 ^ n13515 ^ n12019 ;
  assign n28225 = n28177 ^ n5598 ^ n2158 ;
  assign n28224 = ( n5451 & n7597 ) | ( n5451 & ~n23123 ) | ( n7597 & ~n23123 ) ;
  assign n28226 = n28225 ^ n28224 ^ n9224 ;
  assign n28227 = n19362 ^ n13037 ^ n5731 ;
  assign n28228 = n14472 ^ n6733 ^ n319 ;
  assign n28229 = ( ~n5762 & n23860 ) | ( ~n5762 & n28228 ) | ( n23860 & n28228 ) ;
  assign n28230 = ( n7185 & n15923 ) | ( n7185 & ~n26446 ) | ( n15923 & ~n26446 ) ;
  assign n28231 = ( n7033 & n28229 ) | ( n7033 & ~n28230 ) | ( n28229 & ~n28230 ) ;
  assign n28233 = ( n7618 & ~n21436 ) | ( n7618 & n27524 ) | ( ~n21436 & n27524 ) ;
  assign n28234 = ( n3137 & n16834 ) | ( n3137 & ~n28233 ) | ( n16834 & ~n28233 ) ;
  assign n28235 = n28234 ^ n14338 ^ n399 ;
  assign n28232 = n11124 ^ n7384 ^ n1458 ;
  assign n28236 = n28235 ^ n28232 ^ n19574 ;
  assign n28237 = n13863 ^ n13732 ^ n7804 ;
  assign n28238 = ( n8775 & n14390 ) | ( n8775 & ~n28237 ) | ( n14390 & ~n28237 ) ;
  assign n28239 = n28238 ^ n8755 ^ n2186 ;
  assign n28240 = ( n21657 & n24077 ) | ( n21657 & ~n28239 ) | ( n24077 & ~n28239 ) ;
  assign n28241 = ( n1093 & ~n1214 ) | ( n1093 & n4410 ) | ( ~n1214 & n4410 ) ;
  assign n28242 = n16415 ^ n8848 ^ n260 ;
  assign n28243 = n23900 ^ n19669 ^ n19540 ;
  assign n28244 = ( n28241 & ~n28242 ) | ( n28241 & n28243 ) | ( ~n28242 & n28243 ) ;
  assign n28245 = n27705 ^ n10685 ^ n7574 ;
  assign n28246 = n12701 ^ n7549 ^ n6358 ;
  assign n28247 = ( ~n21397 & n23217 ) | ( ~n21397 & n28246 ) | ( n23217 & n28246 ) ;
  assign n28248 = n11084 ^ n6043 ^ n5965 ;
  assign n28249 = ( ~n9441 & n19209 ) | ( ~n9441 & n28248 ) | ( n19209 & n28248 ) ;
  assign n28250 = ( n5802 & n19444 ) | ( n5802 & n25361 ) | ( n19444 & n25361 ) ;
  assign n28251 = n19545 ^ n16964 ^ n7846 ;
  assign n28252 = ( ~n12293 & n22799 ) | ( ~n12293 & n28251 ) | ( n22799 & n28251 ) ;
  assign n28253 = n9853 ^ n6961 ^ n4348 ;
  assign n28254 = ( n217 & n7378 ) | ( n217 & ~n28253 ) | ( n7378 & ~n28253 ) ;
  assign n28255 = ( n1346 & n17153 ) | ( n1346 & ~n20815 ) | ( n17153 & ~n20815 ) ;
  assign n28256 = ( ~n7295 & n10390 ) | ( ~n7295 & n28255 ) | ( n10390 & n28255 ) ;
  assign n28257 = n28256 ^ n24028 ^ n3405 ;
  assign n28258 = n15321 ^ n7302 ^ n1203 ;
  assign n28259 = n28258 ^ n6323 ^ n3867 ;
  assign n28260 = n28259 ^ n27842 ^ n10581 ;
  assign n28261 = ( n1565 & ~n6325 ) | ( n1565 & n7274 ) | ( ~n6325 & n7274 ) ;
  assign n28262 = n28261 ^ n9059 ^ n361 ;
  assign n28263 = ( n12944 & n15219 ) | ( n12944 & ~n28262 ) | ( n15219 & ~n28262 ) ;
  assign n28266 = n19680 ^ n11998 ^ n625 ;
  assign n28264 = n13728 ^ n6265 ^ n1174 ;
  assign n28265 = n28264 ^ n19955 ^ n12511 ;
  assign n28267 = n28266 ^ n28265 ^ n5077 ;
  assign n28268 = ( n3678 & ~n19162 ) | ( n3678 & n23689 ) | ( ~n19162 & n23689 ) ;
  assign n28269 = n28268 ^ n26735 ^ n4901 ;
  assign n28270 = ( n2288 & ~n8779 ) | ( n2288 & n9630 ) | ( ~n8779 & n9630 ) ;
  assign n28271 = ( n7091 & n9777 ) | ( n7091 & ~n28270 ) | ( n9777 & ~n28270 ) ;
  assign n28272 = n28271 ^ n8805 ^ n2872 ;
  assign n28273 = ( n3240 & ~n11319 ) | ( n3240 & n28272 ) | ( ~n11319 & n28272 ) ;
  assign n28274 = ( n218 & n11501 ) | ( n218 & ~n18602 ) | ( n11501 & ~n18602 ) ;
  assign n28275 = ( ~n4192 & n23447 ) | ( ~n4192 & n28274 ) | ( n23447 & n28274 ) ;
  assign n28276 = ( n4072 & n11910 ) | ( n4072 & n28275 ) | ( n11910 & n28275 ) ;
  assign n28277 = n28276 ^ n23022 ^ n3666 ;
  assign n28278 = ( ~n8316 & n26093 ) | ( ~n8316 & n27652 ) | ( n26093 & n27652 ) ;
  assign n28279 = ( n7802 & n15946 ) | ( n7802 & ~n20063 ) | ( n15946 & ~n20063 ) ;
  assign n28280 = ( n4591 & n16763 ) | ( n4591 & ~n21752 ) | ( n16763 & ~n21752 ) ;
  assign n28282 = n18657 ^ n5388 ^ n3813 ;
  assign n28283 = n28282 ^ n15388 ^ n5838 ;
  assign n28281 = ( n3874 & n9567 ) | ( n3874 & ~n16870 ) | ( n9567 & ~n16870 ) ;
  assign n28284 = n28283 ^ n28281 ^ n6212 ;
  assign n28285 = ( n11378 & n14684 ) | ( n11378 & n21562 ) | ( n14684 & n21562 ) ;
  assign n28286 = n25373 ^ n11452 ^ n11450 ;
  assign n28287 = ( n2666 & n12907 ) | ( n2666 & ~n15074 ) | ( n12907 & ~n15074 ) ;
  assign n28288 = n6395 ^ n6243 ^ n4562 ;
  assign n28289 = ( n10032 & n20085 ) | ( n10032 & n28288 ) | ( n20085 & n28288 ) ;
  assign n28290 = ( ~n23977 & n28287 ) | ( ~n23977 & n28289 ) | ( n28287 & n28289 ) ;
  assign n28291 = ( ~n10849 & n13008 ) | ( ~n10849 & n23313 ) | ( n13008 & n23313 ) ;
  assign n28292 = n21941 ^ n11383 ^ n10831 ;
  assign n28293 = n28292 ^ n6299 ^ n3394 ;
  assign n28295 = ( ~n13984 & n15096 ) | ( ~n13984 & n17298 ) | ( n15096 & n17298 ) ;
  assign n28294 = ( n8778 & n18406 ) | ( n8778 & n25354 ) | ( n18406 & n25354 ) ;
  assign n28296 = n28295 ^ n28294 ^ n1689 ;
  assign n28297 = ( n10329 & n12769 ) | ( n10329 & n15480 ) | ( n12769 & n15480 ) ;
  assign n28298 = ( ~n742 & n1416 ) | ( ~n742 & n6776 ) | ( n1416 & n6776 ) ;
  assign n28299 = ( n1854 & ~n4536 ) | ( n1854 & n7543 ) | ( ~n4536 & n7543 ) ;
  assign n28300 = ( n316 & n1547 ) | ( n316 & n1639 ) | ( n1547 & n1639 ) ;
  assign n28301 = ( n12168 & n16081 ) | ( n12168 & ~n18820 ) | ( n16081 & ~n18820 ) ;
  assign n28302 = ( x41 & ~n10260 ) | ( x41 & n15422 ) | ( ~n10260 & n15422 ) ;
  assign n28303 = n28302 ^ n21508 ^ n21410 ;
  assign n28304 = ( n4170 & ~n27308 ) | ( n4170 & n28303 ) | ( ~n27308 & n28303 ) ;
  assign n28305 = n28304 ^ n25631 ^ n18173 ;
  assign n28306 = ( n2838 & n8435 ) | ( n2838 & ~n9075 ) | ( n8435 & ~n9075 ) ;
  assign n28307 = n28306 ^ n11418 ^ n7420 ;
  assign n28308 = ( n8167 & n9398 ) | ( n8167 & n28307 ) | ( n9398 & n28307 ) ;
  assign n28309 = n28308 ^ n6576 ^ n1012 ;
  assign n28310 = ( n855 & ~n10027 ) | ( n855 & n18244 ) | ( ~n10027 & n18244 ) ;
  assign n28311 = ( n2528 & ~n11552 ) | ( n2528 & n28310 ) | ( ~n11552 & n28310 ) ;
  assign n28312 = n20988 ^ n16232 ^ n10095 ;
  assign n28314 = ( ~n556 & n10174 ) | ( ~n556 & n14634 ) | ( n10174 & n14634 ) ;
  assign n28313 = n13049 ^ n12114 ^ n1167 ;
  assign n28315 = n28314 ^ n28313 ^ n5175 ;
  assign n28316 = n2301 ^ n1365 ^ n1350 ;
  assign n28317 = n28316 ^ n15677 ^ n14384 ;
  assign n28318 = n6191 ^ n3395 ^ n2405 ;
  assign n28319 = n28318 ^ n8567 ^ n5623 ;
  assign n28320 = n28319 ^ n24308 ^ n21481 ;
  assign n28321 = ( ~n624 & n3972 ) | ( ~n624 & n6966 ) | ( n3972 & n6966 ) ;
  assign n28322 = n28321 ^ n15013 ^ n441 ;
  assign n28323 = ( n11326 & ~n17616 ) | ( n11326 & n28322 ) | ( ~n17616 & n28322 ) ;
  assign n28324 = n28323 ^ n7031 ^ n6845 ;
  assign n28325 = n28323 ^ n19342 ^ n6964 ;
  assign n28326 = ( ~n667 & n12170 ) | ( ~n667 & n15094 ) | ( n12170 & n15094 ) ;
  assign n28327 = n28326 ^ n11800 ^ n3395 ;
  assign n28328 = ( ~n1044 & n8479 ) | ( ~n1044 & n15573 ) | ( n8479 & n15573 ) ;
  assign n28329 = n28328 ^ n19161 ^ n5732 ;
  assign n28330 = ( ~n7657 & n22426 ) | ( ~n7657 & n23045 ) | ( n22426 & n23045 ) ;
  assign n28331 = n21113 ^ n17294 ^ n1251 ;
  assign n28332 = ( n1025 & n11220 ) | ( n1025 & ~n15435 ) | ( n11220 & ~n15435 ) ;
  assign n28333 = n28332 ^ n26338 ^ n21393 ;
  assign n28334 = ( ~n9742 & n10242 ) | ( ~n9742 & n17441 ) | ( n10242 & n17441 ) ;
  assign n28335 = ( ~n4165 & n5555 ) | ( ~n4165 & n28334 ) | ( n5555 & n28334 ) ;
  assign n28336 = n3954 ^ n3747 ^ n2985 ;
  assign n28337 = ( n18349 & n21987 ) | ( n18349 & n28336 ) | ( n21987 & n28336 ) ;
  assign n28338 = n14636 ^ n8082 ^ n2710 ;
  assign n28339 = n10554 ^ n2442 ^ n988 ;
  assign n28340 = ( n5920 & n12016 ) | ( n5920 & ~n19980 ) | ( n12016 & ~n19980 ) ;
  assign n28341 = n22469 ^ n11692 ^ n2337 ;
  assign n28342 = ( n3910 & ~n11541 ) | ( n3910 & n16163 ) | ( ~n11541 & n16163 ) ;
  assign n28343 = ( n4332 & ~n8107 ) | ( n4332 & n28270 ) | ( ~n8107 & n28270 ) ;
  assign n28344 = n6299 ^ n2197 ^ n208 ;
  assign n28345 = n28344 ^ n22118 ^ n12728 ;
  assign n28346 = n17452 ^ n8247 ^ n5347 ;
  assign n28347 = n28346 ^ n24436 ^ n21071 ;
  assign n28348 = n28347 ^ n9862 ^ n2856 ;
  assign n28349 = n17155 ^ n13707 ^ n2289 ;
  assign n28350 = n19896 ^ n7660 ^ n7025 ;
  assign n28351 = n28350 ^ n25777 ^ n24584 ;
  assign n28352 = n28351 ^ n22245 ^ n15827 ;
  assign n28353 = n21603 ^ n17813 ^ n14673 ;
  assign n28354 = n18095 ^ n7538 ^ n6406 ;
  assign n28355 = n28354 ^ n27032 ^ n13798 ;
  assign n28356 = ( ~n379 & n9956 ) | ( ~n379 & n20276 ) | ( n9956 & n20276 ) ;
  assign n28357 = n28356 ^ n23243 ^ n3635 ;
  assign n28358 = n8077 ^ n5396 ^ n3883 ;
  assign n28359 = ( n4870 & n25639 ) | ( n4870 & ~n28358 ) | ( n25639 & ~n28358 ) ;
  assign n28360 = n8802 ^ n7204 ^ n3543 ;
  assign n28361 = n28360 ^ n8902 ^ n8427 ;
  assign n28362 = n12690 ^ n12574 ^ n398 ;
  assign n28363 = n12522 ^ n7178 ^ n1650 ;
  assign n28364 = n28363 ^ n15709 ^ n164 ;
  assign n28365 = ( n3245 & n7892 ) | ( n3245 & ~n14547 ) | ( n7892 & ~n14547 ) ;
  assign n28366 = n28365 ^ n10396 ^ n5575 ;
  assign n28367 = n28366 ^ n18030 ^ n11409 ;
  assign n28369 = n22050 ^ n20265 ^ n15989 ;
  assign n28370 = n28369 ^ n15789 ^ n10074 ;
  assign n28368 = n3299 ^ n1721 ^ n1337 ;
  assign n28371 = n28370 ^ n28368 ^ n25255 ;
  assign n28372 = n8952 ^ n1610 ^ n1003 ;
  assign n28373 = n28372 ^ n9458 ^ n4242 ;
  assign n28374 = n25447 ^ n19620 ^ n2676 ;
  assign n28375 = n28374 ^ n17829 ^ n13344 ;
  assign n28376 = n8587 ^ n7299 ^ n5500 ;
  assign n28377 = n21377 ^ n20011 ^ n10351 ;
  assign n28380 = n20689 ^ n15929 ^ n132 ;
  assign n28378 = ( ~n1865 & n4188 ) | ( ~n1865 & n15967 ) | ( n4188 & n15967 ) ;
  assign n28379 = n28378 ^ n8327 ^ n3724 ;
  assign n28381 = n28380 ^ n28379 ^ n5026 ;
  assign n28382 = ( n3452 & n20400 ) | ( n3452 & n20704 ) | ( n20400 & n20704 ) ;
  assign n28383 = ( ~n2410 & n13787 ) | ( ~n2410 & n22732 ) | ( n13787 & n22732 ) ;
  assign n28384 = ( n11395 & n12126 ) | ( n11395 & ~n28383 ) | ( n12126 & ~n28383 ) ;
  assign n28385 = n23457 ^ n11935 ^ n2155 ;
  assign n28386 = ( n17029 & n17629 ) | ( n17029 & n20809 ) | ( n17629 & n20809 ) ;
  assign n28387 = ( n22002 & ~n28385 ) | ( n22002 & n28386 ) | ( ~n28385 & n28386 ) ;
  assign n28388 = ( ~n4718 & n7559 ) | ( ~n4718 & n28387 ) | ( n7559 & n28387 ) ;
  assign n28389 = ( n1724 & ~n5435 ) | ( n1724 & n9443 ) | ( ~n5435 & n9443 ) ;
  assign n28390 = ( n3357 & n5074 ) | ( n3357 & ~n7966 ) | ( n5074 & ~n7966 ) ;
  assign n28391 = ( n264 & n1635 ) | ( n264 & n28390 ) | ( n1635 & n28390 ) ;
  assign n28392 = n28391 ^ n22788 ^ n9121 ;
  assign n28393 = ( n2673 & n2802 ) | ( n2673 & ~n21390 ) | ( n2802 & ~n21390 ) ;
  assign n28394 = ( n16817 & n20807 ) | ( n16817 & n28393 ) | ( n20807 & n28393 ) ;
  assign n28395 = n12895 ^ n7764 ^ n6698 ;
  assign n28396 = n14067 ^ n11445 ^ n9698 ;
  assign n28397 = n9376 ^ n6232 ^ n3892 ;
  assign n28398 = n28397 ^ n17430 ^ n3104 ;
  assign n28399 = ( n7992 & ~n14226 ) | ( n7992 & n19280 ) | ( ~n14226 & n19280 ) ;
  assign n28400 = ( n3940 & ~n6441 ) | ( n3940 & n25181 ) | ( ~n6441 & n25181 ) ;
  assign n28401 = n17784 ^ n13744 ^ n7648 ;
  assign n28402 = n19669 ^ n8327 ^ n677 ;
  assign n28403 = ( n4028 & ~n28401 ) | ( n4028 & n28402 ) | ( ~n28401 & n28402 ) ;
  assign n28404 = ( ~n1761 & n6703 ) | ( ~n1761 & n26627 ) | ( n6703 & n26627 ) ;
  assign n28405 = ( n7160 & n15967 ) | ( n7160 & ~n18127 ) | ( n15967 & ~n18127 ) ;
  assign n28406 = ( n7498 & n10963 ) | ( n7498 & n28405 ) | ( n10963 & n28405 ) ;
  assign n28407 = n28406 ^ n23396 ^ n20659 ;
  assign n28408 = ( n9623 & ~n14127 ) | ( n9623 & n22474 ) | ( ~n14127 & n22474 ) ;
  assign n28409 = n28408 ^ n3804 ^ n798 ;
  assign n28410 = n25371 ^ n14595 ^ n9292 ;
  assign n28411 = ( ~n270 & n10452 ) | ( ~n270 & n14872 ) | ( n10452 & n14872 ) ;
  assign n28412 = ( n19745 & n20487 ) | ( n19745 & n28411 ) | ( n20487 & n28411 ) ;
  assign n28413 = ( n12642 & n28410 ) | ( n12642 & n28412 ) | ( n28410 & n28412 ) ;
  assign n28415 = ( n1346 & n2411 ) | ( n1346 & ~n10422 ) | ( n2411 & ~n10422 ) ;
  assign n28414 = ( n642 & n13479 ) | ( n642 & ~n27731 ) | ( n13479 & ~n27731 ) ;
  assign n28416 = n28415 ^ n28414 ^ n16509 ;
  assign n28417 = ( ~n17039 & n22118 ) | ( ~n17039 & n22613 ) | ( n22118 & n22613 ) ;
  assign n28418 = n28417 ^ n12924 ^ n1550 ;
  assign n28419 = n28418 ^ n25888 ^ n3499 ;
  assign n28420 = n28419 ^ n23018 ^ n12925 ;
  assign n28421 = ( n2766 & n11496 ) | ( n2766 & ~n14128 ) | ( n11496 & ~n14128 ) ;
  assign n28422 = ( n3426 & n8244 ) | ( n3426 & n28421 ) | ( n8244 & n28421 ) ;
  assign n28423 = ( n1404 & n4307 ) | ( n1404 & n8374 ) | ( n4307 & n8374 ) ;
  assign n28424 = n28423 ^ n9183 ^ n4524 ;
  assign n28425 = n28424 ^ n25374 ^ n16923 ;
  assign n28426 = n28425 ^ n19513 ^ n3404 ;
  assign n28427 = ( n15002 & n24696 ) | ( n15002 & ~n28426 ) | ( n24696 & ~n28426 ) ;
  assign n28428 = ( n4095 & ~n15929 ) | ( n4095 & n16577 ) | ( ~n15929 & n16577 ) ;
  assign n28429 = n10419 ^ n5949 ^ n4207 ;
  assign n28430 = ( ~n9349 & n22960 ) | ( ~n9349 & n28429 ) | ( n22960 & n28429 ) ;
  assign n28431 = ( n3454 & n4030 ) | ( n3454 & ~n4199 ) | ( n4030 & ~n4199 ) ;
  assign n28432 = n28431 ^ n9828 ^ n6660 ;
  assign n28433 = ( n5112 & n12402 ) | ( n5112 & ~n15662 ) | ( n12402 & ~n15662 ) ;
  assign n28434 = n28433 ^ n19604 ^ n10700 ;
  assign n28435 = ( n481 & ~n21481 ) | ( n481 & n22104 ) | ( ~n21481 & n22104 ) ;
  assign n28436 = ( n17277 & n28434 ) | ( n17277 & n28435 ) | ( n28434 & n28435 ) ;
  assign n28439 = ( n2085 & n4796 ) | ( n2085 & n10779 ) | ( n4796 & n10779 ) ;
  assign n28440 = n28439 ^ n9850 ^ n1137 ;
  assign n28437 = n9564 ^ n9383 ^ n7485 ;
  assign n28438 = n28437 ^ n16562 ^ n1709 ;
  assign n28441 = n28440 ^ n28438 ^ n15909 ;
  assign n28442 = n17592 ^ n16853 ^ n14276 ;
  assign n28443 = ( n4113 & ~n9464 ) | ( n4113 & n28442 ) | ( ~n9464 & n28442 ) ;
  assign n28444 = n7820 ^ n6524 ^ n4077 ;
  assign n28445 = ( ~n2517 & n4004 ) | ( ~n2517 & n28444 ) | ( n4004 & n28444 ) ;
  assign n28446 = ( n4848 & n5091 ) | ( n4848 & ~n27606 ) | ( n5091 & ~n27606 ) ;
  assign n28447 = ( ~n3170 & n25767 ) | ( ~n3170 & n28446 ) | ( n25767 & n28446 ) ;
  assign n28451 = ( n20256 & n20557 ) | ( n20256 & ~n24273 ) | ( n20557 & ~n24273 ) ;
  assign n28448 = n15873 ^ n14886 ^ n2714 ;
  assign n28449 = ( n6631 & ~n12353 ) | ( n6631 & n28448 ) | ( ~n12353 & n28448 ) ;
  assign n28450 = n28449 ^ n19866 ^ n19139 ;
  assign n28452 = n28451 ^ n28450 ^ n9004 ;
  assign n28453 = n15359 ^ n10305 ^ n7597 ;
  assign n28454 = ( n1814 & n24232 ) | ( n1814 & n28453 ) | ( n24232 & n28453 ) ;
  assign n28455 = ( n7476 & ~n13425 ) | ( n7476 & n28454 ) | ( ~n13425 & n28454 ) ;
  assign n28456 = n22790 ^ n15740 ^ n15582 ;
  assign n28457 = n28456 ^ n12877 ^ n4485 ;
  assign n28458 = n12058 ^ n2418 ^ x111 ;
  assign n28459 = n27575 ^ n13821 ^ n2577 ;
  assign n28460 = n23447 ^ n11283 ^ n2061 ;
  assign n28461 = n28460 ^ n17812 ^ n16022 ;
  assign n28462 = ( n10643 & ~n13490 ) | ( n10643 & n21089 ) | ( ~n13490 & n21089 ) ;
  assign n28463 = ( n5016 & n16705 ) | ( n5016 & n20000 ) | ( n16705 & n20000 ) ;
  assign n28464 = n21175 ^ n10848 ^ n1877 ;
  assign n28465 = n28464 ^ n20114 ^ n17152 ;
  assign n28466 = n24859 ^ n22064 ^ n12126 ;
  assign n28467 = ( n3897 & ~n10174 ) | ( n3897 & n15844 ) | ( ~n10174 & n15844 ) ;
  assign n28468 = ( n6051 & n6502 ) | ( n6051 & n28467 ) | ( n6502 & n28467 ) ;
  assign n28469 = n28468 ^ n26852 ^ n4132 ;
  assign n28470 = ( ~n2798 & n6999 ) | ( ~n2798 & n28469 ) | ( n6999 & n28469 ) ;
  assign n28471 = n28470 ^ n23824 ^ n18570 ;
  assign n28472 = ( ~n2887 & n17037 ) | ( ~n2887 & n17434 ) | ( n17037 & n17434 ) ;
  assign n28473 = n28472 ^ n4167 ^ n3668 ;
  assign n28474 = ( n8502 & ~n22903 ) | ( n8502 & n22975 ) | ( ~n22903 & n22975 ) ;
  assign n28475 = ( ~n6540 & n12028 ) | ( ~n6540 & n22906 ) | ( n12028 & n22906 ) ;
  assign n28476 = n28475 ^ n13507 ^ n10744 ;
  assign n28477 = ( n1366 & n6090 ) | ( n1366 & n20634 ) | ( n6090 & n20634 ) ;
  assign n28478 = ( ~n9092 & n14024 ) | ( ~n9092 & n14369 ) | ( n14024 & n14369 ) ;
  assign n28479 = n15362 ^ n7817 ^ n5592 ;
  assign n28480 = ( n5521 & n28478 ) | ( n5521 & ~n28479 ) | ( n28478 & ~n28479 ) ;
  assign n28483 = n2279 ^ n1223 ^ x5 ;
  assign n28484 = ( n4995 & n20363 ) | ( n4995 & ~n28483 ) | ( n20363 & ~n28483 ) ;
  assign n28481 = n17822 ^ n15769 ^ n407 ;
  assign n28482 = n28481 ^ n22649 ^ n18211 ;
  assign n28485 = n28484 ^ n28482 ^ n13715 ;
  assign n28486 = ( n1078 & n19534 ) | ( n1078 & n20520 ) | ( n19534 & n20520 ) ;
  assign n28489 = n12461 ^ n8997 ^ n5583 ;
  assign n28487 = ( n11847 & n20526 ) | ( n11847 & ~n25729 ) | ( n20526 & ~n25729 ) ;
  assign n28488 = n28487 ^ n23127 ^ n19106 ;
  assign n28490 = n28489 ^ n28488 ^ n4473 ;
  assign n28491 = ( ~n12833 & n17083 ) | ( ~n12833 & n28490 ) | ( n17083 & n28490 ) ;
  assign n28494 = ( ~n5940 & n8604 ) | ( ~n5940 & n23874 ) | ( n8604 & n23874 ) ;
  assign n28492 = ( ~n971 & n1702 ) | ( ~n971 & n8698 ) | ( n1702 & n8698 ) ;
  assign n28493 = n28492 ^ n7512 ^ n637 ;
  assign n28495 = n28494 ^ n28493 ^ n11205 ;
  assign n28497 = ( n2737 & ~n2744 ) | ( n2737 & n3927 ) | ( ~n2744 & n3927 ) ;
  assign n28498 = ( ~n4499 & n5147 ) | ( ~n4499 & n28497 ) | ( n5147 & n28497 ) ;
  assign n28499 = ( n2574 & ~n27855 ) | ( n2574 & n28498 ) | ( ~n27855 & n28498 ) ;
  assign n28496 = ( x46 & n5299 ) | ( x46 & n12879 ) | ( n5299 & n12879 ) ;
  assign n28500 = n28499 ^ n28496 ^ n14637 ;
  assign n28501 = n20264 ^ n9162 ^ n5654 ;
  assign n28502 = ( n18318 & n25599 ) | ( n18318 & ~n28501 ) | ( n25599 & ~n28501 ) ;
  assign n28503 = ( n135 & n228 ) | ( n135 & ~n2353 ) | ( n228 & ~n2353 ) ;
  assign n28505 = ( n497 & n11182 ) | ( n497 & ~n13413 ) | ( n11182 & ~n13413 ) ;
  assign n28504 = n21905 ^ n12880 ^ n1640 ;
  assign n28506 = n28505 ^ n28504 ^ n8371 ;
  assign n28507 = ( ~n8095 & n10071 ) | ( ~n8095 & n28506 ) | ( n10071 & n28506 ) ;
  assign n28508 = n13191 ^ n11062 ^ n7276 ;
  assign n28509 = n28508 ^ n26599 ^ n13773 ;
  assign n28510 = n28509 ^ n27479 ^ n1580 ;
  assign n28511 = ( n5465 & n12559 ) | ( n5465 & ~n28510 ) | ( n12559 & ~n28510 ) ;
  assign n28512 = ( n6142 & ~n9080 ) | ( n6142 & n15186 ) | ( ~n9080 & n15186 ) ;
  assign n28513 = n28512 ^ n17622 ^ n6822 ;
  assign n28514 = n28513 ^ n11858 ^ n10574 ;
  assign n28515 = ( n3743 & ~n13675 ) | ( n3743 & n15153 ) | ( ~n13675 & n15153 ) ;
  assign n28516 = n6202 ^ n4163 ^ n3611 ;
  assign n28517 = n17786 ^ n2439 ^ n1105 ;
  assign n28518 = ( n9626 & n21146 ) | ( n9626 & n28517 ) | ( n21146 & n28517 ) ;
  assign n28519 = ( n28515 & ~n28516 ) | ( n28515 & n28518 ) | ( ~n28516 & n28518 ) ;
  assign n28520 = ( n3025 & n9062 ) | ( n3025 & ~n23452 ) | ( n9062 & ~n23452 ) ;
  assign n28521 = n28520 ^ n11290 ^ n7685 ;
  assign n28522 = n11998 ^ n8852 ^ n5567 ;
  assign n28523 = ( n144 & n5139 ) | ( n144 & ~n28522 ) | ( n5139 & ~n28522 ) ;
  assign n28524 = n14950 ^ n13789 ^ n565 ;
  assign n28525 = n28524 ^ n9271 ^ n2130 ;
  assign n28526 = ( n2880 & n26845 ) | ( n2880 & ~n28525 ) | ( n26845 & ~n28525 ) ;
  assign n28527 = ( n14819 & n28523 ) | ( n14819 & ~n28526 ) | ( n28523 & ~n28526 ) ;
  assign n28528 = n16417 ^ n10790 ^ n1497 ;
  assign n28529 = ( n4856 & n7866 ) | ( n4856 & n12028 ) | ( n7866 & n12028 ) ;
  assign n28530 = n19926 ^ n9056 ^ n6823 ;
  assign n28531 = ( n21954 & n27264 ) | ( n21954 & n28530 ) | ( n27264 & n28530 ) ;
  assign n28532 = ( n4637 & n5786 ) | ( n4637 & n11821 ) | ( n5786 & n11821 ) ;
  assign n28533 = ( ~n8675 & n15957 ) | ( ~n8675 & n28532 ) | ( n15957 & n28532 ) ;
  assign n28534 = ( n142 & ~n18196 ) | ( n142 & n28533 ) | ( ~n18196 & n28533 ) ;
  assign n28535 = ( n11447 & n22779 ) | ( n11447 & n23541 ) | ( n22779 & n23541 ) ;
  assign n28536 = n15383 ^ n12422 ^ n4111 ;
  assign n28537 = ( ~n4344 & n12919 ) | ( ~n4344 & n28536 ) | ( n12919 & n28536 ) ;
  assign n28538 = ( n8326 & ~n8855 ) | ( n8326 & n14960 ) | ( ~n8855 & n14960 ) ;
  assign n28539 = ( n8507 & n14811 ) | ( n8507 & ~n28538 ) | ( n14811 & ~n28538 ) ;
  assign n28540 = n28539 ^ n10106 ^ n5904 ;
  assign n28541 = n28540 ^ n14614 ^ n14058 ;
  assign n28542 = n28541 ^ n26538 ^ n11772 ;
  assign n28543 = n28366 ^ n9431 ^ n5840 ;
  assign n28546 = n23817 ^ n13813 ^ n13118 ;
  assign n28547 = n28546 ^ n12254 ^ n7621 ;
  assign n28544 = ( n2079 & n4162 ) | ( n2079 & n22213 ) | ( n4162 & n22213 ) ;
  assign n28545 = n28544 ^ n8747 ^ n1713 ;
  assign n28548 = n28547 ^ n28545 ^ n11477 ;
  assign n28549 = n28548 ^ n25979 ^ n23865 ;
  assign n28550 = n13255 ^ n12414 ^ n547 ;
  assign n28551 = ( n2687 & ~n7520 ) | ( n2687 & n28550 ) | ( ~n7520 & n28550 ) ;
  assign n28552 = n17121 ^ n14620 ^ n10058 ;
  assign n28553 = n28552 ^ n9570 ^ n2502 ;
  assign n28555 = n25095 ^ n19112 ^ n7994 ;
  assign n28554 = n13576 ^ n8029 ^ n6278 ;
  assign n28556 = n28555 ^ n28554 ^ n18346 ;
  assign n28557 = ( n3218 & ~n13340 ) | ( n3218 & n21571 ) | ( ~n13340 & n21571 ) ;
  assign n28558 = ( ~n8324 & n19180 ) | ( ~n8324 & n28557 ) | ( n19180 & n28557 ) ;
  assign n28559 = n22419 ^ n3996 ^ n2254 ;
  assign n28560 = ( n6977 & ~n26751 ) | ( n6977 & n28559 ) | ( ~n26751 & n28559 ) ;
  assign n28561 = n25827 ^ n23400 ^ n3161 ;
  assign n28562 = ( n1651 & n4153 ) | ( n1651 & ~n7215 ) | ( n4153 & ~n7215 ) ;
  assign n28563 = ( n293 & n2187 ) | ( n293 & ~n28562 ) | ( n2187 & ~n28562 ) ;
  assign n28564 = ( ~n21304 & n26643 ) | ( ~n21304 & n28563 ) | ( n26643 & n28563 ) ;
  assign n28565 = n28564 ^ n22288 ^ n2387 ;
  assign n28566 = n25351 ^ n14699 ^ n11998 ;
  assign n28567 = ( n869 & ~n6945 ) | ( n869 & n28566 ) | ( ~n6945 & n28566 ) ;
  assign n28568 = ( ~x82 & n8688 ) | ( ~x82 & n20817 ) | ( n8688 & n20817 ) ;
  assign n28569 = ( ~n4461 & n14686 ) | ( ~n4461 & n28568 ) | ( n14686 & n28568 ) ;
  assign n28570 = ( n4096 & n4287 ) | ( n4096 & n6085 ) | ( n4287 & n6085 ) ;
  assign n28571 = ( n11433 & n26988 ) | ( n11433 & ~n28570 ) | ( n26988 & ~n28570 ) ;
  assign n28572 = ( n10721 & n16553 ) | ( n10721 & ~n19164 ) | ( n16553 & ~n19164 ) ;
  assign n28573 = n26804 ^ n5654 ^ n424 ;
  assign n28574 = ( ~n9598 & n14494 ) | ( ~n9598 & n24126 ) | ( n14494 & n24126 ) ;
  assign n28575 = ( n390 & ~n5006 ) | ( n390 & n6994 ) | ( ~n5006 & n6994 ) ;
  assign n28576 = n28575 ^ n23863 ^ n22747 ;
  assign n28577 = n11266 ^ n6147 ^ n2629 ;
  assign n28578 = ( n18786 & ~n19562 ) | ( n18786 & n28577 ) | ( ~n19562 & n28577 ) ;
  assign n28579 = ( n747 & n6898 ) | ( n747 & n12355 ) | ( n6898 & n12355 ) ;
  assign n28580 = ( n979 & ~n23881 ) | ( n979 & n28579 ) | ( ~n23881 & n28579 ) ;
  assign n28581 = n28580 ^ n27211 ^ n15878 ;
  assign n28582 = ( n2362 & n18762 ) | ( n2362 & n23390 ) | ( n18762 & n23390 ) ;
  assign n28583 = ( n6796 & n7172 ) | ( n6796 & n9839 ) | ( n7172 & n9839 ) ;
  assign n28584 = ( n9432 & n14967 ) | ( n9432 & ~n22350 ) | ( n14967 & ~n22350 ) ;
  assign n28585 = ( ~n7183 & n8198 ) | ( ~n7183 & n18417 ) | ( n8198 & n18417 ) ;
  assign n28586 = n14276 ^ n10549 ^ n8203 ;
  assign n28587 = ( n1832 & n9829 ) | ( n1832 & n28586 ) | ( n9829 & n28586 ) ;
  assign n28588 = ( ~n3617 & n15736 ) | ( ~n3617 & n28587 ) | ( n15736 & n28587 ) ;
  assign n28589 = n21327 ^ n17787 ^ n13488 ;
  assign n28590 = n22788 ^ n10349 ^ n6141 ;
  assign n28591 = n22360 ^ n6618 ^ n2354 ;
  assign n28592 = ( n11702 & n13897 ) | ( n11702 & ~n25794 ) | ( n13897 & ~n25794 ) ;
  assign n28593 = ( ~n334 & n3315 ) | ( ~n334 & n28592 ) | ( n3315 & n28592 ) ;
  assign n28594 = n28593 ^ n15914 ^ n11175 ;
  assign n28595 = ( ~n28590 & n28591 ) | ( ~n28590 & n28594 ) | ( n28591 & n28594 ) ;
  assign n28596 = ( n455 & n3619 ) | ( n455 & ~n5092 ) | ( n3619 & ~n5092 ) ;
  assign n28597 = n28596 ^ n14422 ^ n2533 ;
  assign n28598 = n22516 ^ n14226 ^ n154 ;
  assign n28599 = n28598 ^ n15232 ^ n10567 ;
  assign n28600 = ( n2777 & n28597 ) | ( n2777 & n28599 ) | ( n28597 & n28599 ) ;
  assign n28601 = n28600 ^ n26840 ^ n11146 ;
  assign n28602 = ( n11016 & n12890 ) | ( n11016 & n28601 ) | ( n12890 & n28601 ) ;
  assign n28603 = ( n11457 & n19369 ) | ( n11457 & n23362 ) | ( n19369 & n23362 ) ;
  assign n28604 = n27558 ^ n11768 ^ n11699 ;
  assign n28605 = ( n2020 & ~n2681 ) | ( n2020 & n7520 ) | ( ~n2681 & n7520 ) ;
  assign n28606 = n28605 ^ n24386 ^ n15433 ;
  assign n28607 = ( ~n13565 & n15465 ) | ( ~n13565 & n28606 ) | ( n15465 & n28606 ) ;
  assign n28608 = n24260 ^ n11387 ^ n5675 ;
  assign n28609 = n17906 ^ n11564 ^ n3568 ;
  assign n28610 = ( n12317 & n15320 ) | ( n12317 & n22632 ) | ( n15320 & n22632 ) ;
  assign n28611 = ( ~n14695 & n15118 ) | ( ~n14695 & n17399 ) | ( n15118 & n17399 ) ;
  assign n28612 = n28611 ^ n21980 ^ n16828 ;
  assign n28613 = n28612 ^ n13396 ^ n3388 ;
  assign n28614 = n18989 ^ n9975 ^ n3088 ;
  assign n28615 = n28614 ^ n27424 ^ n8141 ;
  assign n28616 = ( n10114 & n18844 ) | ( n10114 & ~n26195 ) | ( n18844 & ~n26195 ) ;
  assign n28617 = ( n18134 & n18378 ) | ( n18134 & n25824 ) | ( n18378 & n25824 ) ;
  assign n28618 = n10879 ^ n8800 ^ n210 ;
  assign n28619 = n26182 ^ n14871 ^ n373 ;
  assign n28620 = ( ~n4525 & n6974 ) | ( ~n4525 & n8917 ) | ( n6974 & n8917 ) ;
  assign n28621 = n28620 ^ n13051 ^ n11958 ;
  assign n28622 = n16957 ^ n16923 ^ n7343 ;
  assign n28623 = ( n1876 & n9280 ) | ( n1876 & n28622 ) | ( n9280 & n28622 ) ;
  assign n28624 = ( n2463 & n6802 ) | ( n2463 & ~n25500 ) | ( n6802 & ~n25500 ) ;
  assign n28625 = ( n11501 & n20501 ) | ( n11501 & ~n27215 ) | ( n20501 & ~n27215 ) ;
  assign n28626 = ( n13774 & ~n21535 ) | ( n13774 & n28625 ) | ( ~n21535 & n28625 ) ;
  assign n28627 = ( ~n7381 & n8940 ) | ( ~n7381 & n28626 ) | ( n8940 & n28626 ) ;
  assign n28628 = n10217 ^ n4743 ^ n2947 ;
  assign n28629 = n28628 ^ n21167 ^ n16659 ;
  assign n28630 = ( ~n894 & n19123 ) | ( ~n894 & n26846 ) | ( n19123 & n26846 ) ;
  assign n28631 = n28630 ^ n25366 ^ n13201 ;
  assign n28632 = ( n195 & ~n17407 ) | ( n195 & n23552 ) | ( ~n17407 & n23552 ) ;
  assign n28634 = n14199 ^ n7383 ^ n1463 ;
  assign n28633 = ( n4408 & n5381 ) | ( n4408 & ~n11549 ) | ( n5381 & ~n11549 ) ;
  assign n28635 = n28634 ^ n28633 ^ n26179 ;
  assign n28636 = ( ~n10808 & n15144 ) | ( ~n10808 & n20044 ) | ( n15144 & n20044 ) ;
  assign n28637 = n25389 ^ n24340 ^ n1079 ;
  assign n28638 = ( n690 & n26798 ) | ( n690 & ~n28637 ) | ( n26798 & ~n28637 ) ;
  assign n28639 = n28638 ^ n14171 ^ n7747 ;
  assign n28640 = n28639 ^ n27916 ^ n14301 ;
  assign n28641 = ( n15910 & n28636 ) | ( n15910 & ~n28640 ) | ( n28636 & ~n28640 ) ;
  assign n28642 = ( ~n342 & n7679 ) | ( ~n342 & n17434 ) | ( n7679 & n17434 ) ;
  assign n28643 = n28642 ^ n22088 ^ n7198 ;
  assign n28645 = ( n778 & n9054 ) | ( n778 & n10555 ) | ( n9054 & n10555 ) ;
  assign n28644 = n24420 ^ n12536 ^ n10808 ;
  assign n28646 = n28645 ^ n28644 ^ x30 ;
  assign n28647 = n28646 ^ n18739 ^ n2130 ;
  assign n28648 = n13762 ^ n11859 ^ n753 ;
  assign n28649 = ( ~n6074 & n12270 ) | ( ~n6074 & n28648 ) | ( n12270 & n28648 ) ;
  assign n28650 = n8595 ^ n6474 ^ n580 ;
  assign n28651 = ( n5735 & n28649 ) | ( n5735 & ~n28650 ) | ( n28649 & ~n28650 ) ;
  assign n28652 = ( n3002 & ~n10735 ) | ( n3002 & n22086 ) | ( ~n10735 & n22086 ) ;
  assign n28653 = n24958 ^ n4583 ^ n4374 ;
  assign n28654 = n28653 ^ n15461 ^ n9191 ;
  assign n28655 = ( n4855 & ~n9549 ) | ( n4855 & n26470 ) | ( ~n9549 & n26470 ) ;
  assign n28656 = ( n2816 & n6266 ) | ( n2816 & ~n25153 ) | ( n6266 & ~n25153 ) ;
  assign n28657 = ( ~n3595 & n7201 ) | ( ~n3595 & n11634 ) | ( n7201 & n11634 ) ;
  assign n28659 = ( n737 & ~n2960 ) | ( n737 & n8116 ) | ( ~n2960 & n8116 ) ;
  assign n28658 = ( ~n3034 & n4259 ) | ( ~n3034 & n11675 ) | ( n4259 & n11675 ) ;
  assign n28660 = n28659 ^ n28658 ^ n18590 ;
  assign n28661 = ( n5322 & ~n5621 ) | ( n5322 & n5704 ) | ( ~n5621 & n5704 ) ;
  assign n28662 = n28661 ^ n27896 ^ n13249 ;
  assign n28663 = ( n8288 & n9215 ) | ( n8288 & ~n24264 ) | ( n9215 & ~n24264 ) ;
  assign n28664 = n7583 ^ n7037 ^ n1123 ;
  assign n28665 = ( ~n2428 & n14655 ) | ( ~n2428 & n22041 ) | ( n14655 & n22041 ) ;
  assign n28666 = n15242 ^ n9024 ^ n5755 ;
  assign n28667 = ( n5194 & n8763 ) | ( n5194 & n15317 ) | ( n8763 & n15317 ) ;
  assign n28668 = ( n159 & n3291 ) | ( n159 & n28667 ) | ( n3291 & n28667 ) ;
  assign n28669 = ( n19697 & n28666 ) | ( n19697 & n28668 ) | ( n28666 & n28668 ) ;
  assign n28670 = ( n8763 & ~n14092 ) | ( n8763 & n20674 ) | ( ~n14092 & n20674 ) ;
  assign n28671 = n28670 ^ n15098 ^ n6217 ;
  assign n28672 = ( n15742 & n17357 ) | ( n15742 & ~n27059 ) | ( n17357 & ~n27059 ) ;
  assign n28673 = ( ~n455 & n15120 ) | ( ~n455 & n23691 ) | ( n15120 & n23691 ) ;
  assign n28674 = ( ~n1679 & n18774 ) | ( ~n1679 & n28673 ) | ( n18774 & n28673 ) ;
  assign n28675 = n28674 ^ n10970 ^ n2126 ;
  assign n28676 = ( n6156 & n10495 ) | ( n6156 & n13852 ) | ( n10495 & n13852 ) ;
  assign n28677 = n28676 ^ n12204 ^ n1391 ;
  assign n28678 = ( n2937 & ~n23499 ) | ( n2937 & n28677 ) | ( ~n23499 & n28677 ) ;
  assign n28679 = n5787 ^ n1652 ^ n714 ;
  assign n28680 = n28679 ^ n21942 ^ n9806 ;
  assign n28681 = ( n4206 & n6486 ) | ( n4206 & ~n13197 ) | ( n6486 & ~n13197 ) ;
  assign n28682 = ( n414 & ~n15461 ) | ( n414 & n27968 ) | ( ~n15461 & n27968 ) ;
  assign n28683 = ( n20809 & n28681 ) | ( n20809 & n28682 ) | ( n28681 & n28682 ) ;
  assign n28684 = n28683 ^ n25138 ^ n10502 ;
  assign n28685 = ( n1549 & n15191 ) | ( n1549 & n16378 ) | ( n15191 & n16378 ) ;
  assign n28686 = ( n14116 & ~n19995 ) | ( n14116 & n20110 ) | ( ~n19995 & n20110 ) ;
  assign n28687 = n28686 ^ n18429 ^ n2241 ;
  assign n28688 = n19609 ^ n1242 ^ n876 ;
  assign n28689 = ( n20620 & ~n28687 ) | ( n20620 & n28688 ) | ( ~n28687 & n28688 ) ;
  assign n28690 = n28689 ^ n22887 ^ n15350 ;
  assign n28691 = n14950 ^ n4544 ^ n576 ;
  assign n28692 = ( n1911 & ~n4871 ) | ( n1911 & n21757 ) | ( ~n4871 & n21757 ) ;
  assign n28693 = n27909 ^ n23141 ^ n1448 ;
  assign n28694 = ( n2460 & n12603 ) | ( n2460 & ~n28693 ) | ( n12603 & ~n28693 ) ;
  assign n28695 = n19848 ^ n12961 ^ n5991 ;
  assign n28696 = ( ~n11011 & n28694 ) | ( ~n11011 & n28695 ) | ( n28694 & n28695 ) ;
  assign n28697 = ( ~n26674 & n28692 ) | ( ~n26674 & n28696 ) | ( n28692 & n28696 ) ;
  assign n28698 = ( n5164 & ~n5747 ) | ( n5164 & n11437 ) | ( ~n5747 & n11437 ) ;
  assign n28699 = ( n1566 & ~n7252 ) | ( n1566 & n17439 ) | ( ~n7252 & n17439 ) ;
  assign n28700 = ( ~n22360 & n28698 ) | ( ~n22360 & n28699 ) | ( n28698 & n28699 ) ;
  assign n28701 = n25875 ^ n21646 ^ n4066 ;
  assign n28702 = n13773 ^ n5053 ^ n4695 ;
  assign n28703 = n17248 ^ n17115 ^ n4170 ;
  assign n28704 = n17764 ^ n8163 ^ n1723 ;
  assign n28705 = ( n11765 & ~n19619 ) | ( n11765 & n26714 ) | ( ~n19619 & n26714 ) ;
  assign n28707 = n5732 ^ n3447 ^ n475 ;
  assign n28706 = n24478 ^ n13828 ^ n4995 ;
  assign n28708 = n28707 ^ n28706 ^ n3362 ;
  assign n28709 = n14237 ^ n8467 ^ n3434 ;
  assign n28710 = n9265 ^ n5681 ^ n4218 ;
  assign n28711 = ( n14107 & n25689 ) | ( n14107 & n28710 ) | ( n25689 & n28710 ) ;
  assign n28712 = n27096 ^ n20023 ^ n1261 ;
  assign n28713 = ( ~n1827 & n3722 ) | ( ~n1827 & n11703 ) | ( n3722 & n11703 ) ;
  assign n28714 = ( n19821 & ~n20599 ) | ( n19821 & n28713 ) | ( ~n20599 & n28713 ) ;
  assign n28716 = ( ~n2595 & n6014 ) | ( ~n2595 & n15439 ) | ( n6014 & n15439 ) ;
  assign n28717 = ( n1885 & ~n2758 ) | ( n1885 & n28716 ) | ( ~n2758 & n28716 ) ;
  assign n28715 = n26423 ^ n17398 ^ n8879 ;
  assign n28718 = n28717 ^ n28715 ^ n27907 ;
  assign n28719 = ( n13019 & n13183 ) | ( n13019 & n28718 ) | ( n13183 & n28718 ) ;
  assign n28720 = ( n2283 & ~n3932 ) | ( n2283 & n5135 ) | ( ~n3932 & n5135 ) ;
  assign n28721 = n28720 ^ n24013 ^ n3608 ;
  assign n28722 = n23335 ^ n11348 ^ n769 ;
  assign n28723 = ( n720 & n25720 ) | ( n720 & n28365 ) | ( n25720 & n28365 ) ;
  assign n28724 = ( n4209 & ~n6558 ) | ( n4209 & n13519 ) | ( ~n6558 & n13519 ) ;
  assign n28725 = ( n7851 & n13569 ) | ( n7851 & ~n13948 ) | ( n13569 & ~n13948 ) ;
  assign n28726 = n23192 ^ n13609 ^ n587 ;
  assign n28727 = ( n6082 & ~n15439 ) | ( n6082 & n28726 ) | ( ~n15439 & n28726 ) ;
  assign n28729 = n21450 ^ n18046 ^ n4016 ;
  assign n28728 = ( n19388 & n21465 ) | ( n19388 & ~n25712 ) | ( n21465 & ~n25712 ) ;
  assign n28730 = n28729 ^ n28728 ^ n25492 ;
  assign n28731 = ( ~x48 & n5016 ) | ( ~x48 & n5291 ) | ( n5016 & n5291 ) ;
  assign n28732 = ( ~n3103 & n4915 ) | ( ~n3103 & n28731 ) | ( n4915 & n28731 ) ;
  assign n28733 = n22033 ^ n10478 ^ n5270 ;
  assign n28734 = n28733 ^ n24927 ^ n5558 ;
  assign n28735 = ( n20036 & n28732 ) | ( n20036 & n28734 ) | ( n28732 & n28734 ) ;
  assign n28736 = ( ~n6492 & n6861 ) | ( ~n6492 & n28735 ) | ( n6861 & n28735 ) ;
  assign n28738 = n18821 ^ n1740 ^ n1512 ;
  assign n28737 = n19303 ^ n12218 ^ n12067 ;
  assign n28739 = n28738 ^ n28737 ^ n24768 ;
  assign n28740 = n13033 ^ n6863 ^ n680 ;
  assign n28741 = ( n1597 & ~n28351 ) | ( n1597 & n28740 ) | ( ~n28351 & n28740 ) ;
  assign n28742 = ( ~n819 & n2571 ) | ( ~n819 & n24851 ) | ( n2571 & n24851 ) ;
  assign n28743 = ( ~n26600 & n26960 ) | ( ~n26600 & n28742 ) | ( n26960 & n28742 ) ;
  assign n28744 = ( n1347 & n5705 ) | ( n1347 & n15484 ) | ( n5705 & n15484 ) ;
  assign n28745 = ( n1452 & ~n4806 ) | ( n1452 & n6500 ) | ( ~n4806 & n6500 ) ;
  assign n28746 = n9436 ^ n8601 ^ n527 ;
  assign n28747 = n26808 ^ n18523 ^ n3866 ;
  assign n28748 = ( n1139 & ~n5108 ) | ( n1139 & n5677 ) | ( ~n5108 & n5677 ) ;
  assign n28750 = ( ~n1802 & n6588 ) | ( ~n1802 & n17054 ) | ( n6588 & n17054 ) ;
  assign n28749 = n11800 ^ n9747 ^ n8300 ;
  assign n28751 = n28750 ^ n28749 ^ n22397 ;
  assign n28752 = n11714 ^ n11200 ^ n3985 ;
  assign n28753 = ( n8593 & n23466 ) | ( n8593 & n28752 ) | ( n23466 & n28752 ) ;
  assign n28754 = n12649 ^ n9073 ^ n2945 ;
  assign n28755 = ( n2388 & ~n4661 ) | ( n2388 & n13503 ) | ( ~n4661 & n13503 ) ;
  assign n28756 = ( n28753 & n28754 ) | ( n28753 & ~n28755 ) | ( n28754 & ~n28755 ) ;
  assign n28757 = ( ~n11327 & n12981 ) | ( ~n11327 & n22056 ) | ( n12981 & n22056 ) ;
  assign n28758 = n14570 ^ n14041 ^ n10261 ;
  assign n28759 = ( n25290 & ~n26272 ) | ( n25290 & n28758 ) | ( ~n26272 & n28758 ) ;
  assign n28760 = n28759 ^ n14965 ^ n10190 ;
  assign n28761 = ( n9647 & n15435 ) | ( n9647 & ~n23137 ) | ( n15435 & ~n23137 ) ;
  assign n28763 = ( ~n1146 & n2220 ) | ( ~n1146 & n5883 ) | ( n2220 & n5883 ) ;
  assign n28762 = n26814 ^ n15216 ^ n9523 ;
  assign n28764 = n28763 ^ n28762 ^ n17777 ;
  assign n28765 = ( n826 & ~n9826 ) | ( n826 & n14817 ) | ( ~n9826 & n14817 ) ;
  assign n28766 = n28765 ^ n19503 ^ n6159 ;
  assign n28767 = n19450 ^ n9548 ^ n8661 ;
  assign n28768 = ( n5234 & n23541 ) | ( n5234 & n28767 ) | ( n23541 & n28767 ) ;
  assign n28769 = n28768 ^ n9073 ^ n5574 ;
  assign n28770 = n15996 ^ n10714 ^ n9245 ;
  assign n28771 = n28770 ^ n24724 ^ n16055 ;
  assign n28772 = n19020 ^ n11895 ^ n367 ;
  assign n28773 = ( ~n1971 & n5512 ) | ( ~n1971 & n28152 ) | ( n5512 & n28152 ) ;
  assign n28774 = ( ~n11124 & n13478 ) | ( ~n11124 & n28773 ) | ( n13478 & n28773 ) ;
  assign n28775 = n19385 ^ n9780 ^ n5405 ;
  assign n28776 = n28775 ^ n24253 ^ n3817 ;
  assign n28777 = n14246 ^ n8228 ^ n1557 ;
  assign n28778 = ( n3690 & ~n13341 ) | ( n3690 & n15976 ) | ( ~n13341 & n15976 ) ;
  assign n28779 = ( n17373 & n28777 ) | ( n17373 & ~n28778 ) | ( n28777 & ~n28778 ) ;
  assign n28780 = ( n6201 & n8928 ) | ( n6201 & n28779 ) | ( n8928 & n28779 ) ;
  assign n28781 = n28137 ^ n21956 ^ n16099 ;
  assign n28782 = n28781 ^ n24387 ^ n938 ;
  assign n28783 = ( n13169 & n27896 ) | ( n13169 & n28782 ) | ( n27896 & n28782 ) ;
  assign n28784 = ( ~n12692 & n17591 ) | ( ~n12692 & n20310 ) | ( n17591 & n20310 ) ;
  assign n28785 = ( n11072 & ~n11662 ) | ( n11072 & n23409 ) | ( ~n11662 & n23409 ) ;
  assign n28786 = ( ~n174 & n18099 ) | ( ~n174 & n26980 ) | ( n18099 & n26980 ) ;
  assign n28787 = ( n9818 & n15733 ) | ( n9818 & ~n28786 ) | ( n15733 & ~n28786 ) ;
  assign n28788 = n15164 ^ n11081 ^ n10373 ;
  assign n28789 = ( ~n158 & n17799 ) | ( ~n158 & n28788 ) | ( n17799 & n28788 ) ;
  assign n28790 = n3132 ^ n1480 ^ n169 ;
  assign n28791 = ( ~n3090 & n6565 ) | ( ~n3090 & n12148 ) | ( n6565 & n12148 ) ;
  assign n28792 = ( n1933 & ~n3347 ) | ( n1933 & n28791 ) | ( ~n3347 & n28791 ) ;
  assign n28793 = ( ~n3231 & n20519 ) | ( ~n3231 & n28792 ) | ( n20519 & n28792 ) ;
  assign n28794 = ( n24455 & ~n28790 ) | ( n24455 & n28793 ) | ( ~n28790 & n28793 ) ;
  assign n28795 = n19058 ^ n16498 ^ n6120 ;
  assign n28798 = ( n2915 & n11994 ) | ( n2915 & ~n25000 ) | ( n11994 & ~n25000 ) ;
  assign n28796 = n16348 ^ n12070 ^ n9094 ;
  assign n28797 = ( ~n8001 & n20642 ) | ( ~n8001 & n28796 ) | ( n20642 & n28796 ) ;
  assign n28799 = n28798 ^ n28797 ^ n23876 ;
  assign n28800 = ( n1842 & n7332 ) | ( n1842 & ~n22139 ) | ( n7332 & ~n22139 ) ;
  assign n28801 = n28800 ^ n16669 ^ n451 ;
  assign n28802 = ( ~n2108 & n12915 ) | ( ~n2108 & n28801 ) | ( n12915 & n28801 ) ;
  assign n28803 = ( n1289 & n14141 ) | ( n1289 & ~n27561 ) | ( n14141 & ~n27561 ) ;
  assign n28804 = n26931 ^ n19620 ^ n9085 ;
  assign n28805 = ( n14643 & n23590 ) | ( n14643 & ~n23799 ) | ( n23590 & ~n23799 ) ;
  assign n28806 = ( n1252 & ~n2244 ) | ( n1252 & n18596 ) | ( ~n2244 & n18596 ) ;
  assign n28807 = n28806 ^ n4747 ^ n2708 ;
  assign n28808 = ( n2338 & n14350 ) | ( n2338 & ~n18755 ) | ( n14350 & ~n18755 ) ;
  assign n28809 = ( n9414 & n13859 ) | ( n9414 & ~n28808 ) | ( n13859 & ~n28808 ) ;
  assign n28810 = n11572 ^ n917 ^ n681 ;
  assign n28811 = n28810 ^ n24658 ^ n1243 ;
  assign n28812 = n25384 ^ n24199 ^ n14288 ;
  assign n28814 = n16144 ^ n6533 ^ n1071 ;
  assign n28813 = n15203 ^ n1295 ^ n404 ;
  assign n28815 = n28814 ^ n28813 ^ n5850 ;
  assign n28816 = ( n13651 & n14842 ) | ( n13651 & n22050 ) | ( n14842 & n22050 ) ;
  assign n28817 = n28816 ^ n24714 ^ n5278 ;
  assign n28818 = ( ~n1718 & n3486 ) | ( ~n1718 & n28817 ) | ( n3486 & n28817 ) ;
  assign n28819 = ( ~n14425 & n17986 ) | ( ~n14425 & n24090 ) | ( n17986 & n24090 ) ;
  assign n28820 = ( n3935 & n23562 ) | ( n3935 & n28819 ) | ( n23562 & n28819 ) ;
  assign n28821 = n28820 ^ n22200 ^ n9520 ;
  assign n28822 = ( n15952 & n25564 ) | ( n15952 & n27271 ) | ( n25564 & n27271 ) ;
  assign n28823 = ( n3432 & n13204 ) | ( n3432 & ~n28822 ) | ( n13204 & ~n28822 ) ;
  assign n28824 = ( n2459 & n10502 ) | ( n2459 & n15086 ) | ( n10502 & n15086 ) ;
  assign n28826 = n11200 ^ n6791 ^ n3976 ;
  assign n28825 = ( n1998 & n7980 ) | ( n1998 & ~n14049 ) | ( n7980 & ~n14049 ) ;
  assign n28827 = n28826 ^ n28825 ^ n2484 ;
  assign n28828 = ( n17172 & n28824 ) | ( n17172 & ~n28827 ) | ( n28824 & ~n28827 ) ;
  assign n28829 = n28828 ^ n20106 ^ n9271 ;
  assign n28830 = ( n2850 & n6799 ) | ( n2850 & n14098 ) | ( n6799 & n14098 ) ;
  assign n28831 = n13216 ^ n2450 ^ n812 ;
  assign n28832 = ( n19223 & n25783 ) | ( n19223 & ~n28831 ) | ( n25783 & ~n28831 ) ;
  assign n28833 = n28832 ^ n16871 ^ n6379 ;
  assign n28834 = ( n4695 & ~n5125 ) | ( n4695 & n19962 ) | ( ~n5125 & n19962 ) ;
  assign n28835 = ( n17649 & n23076 ) | ( n17649 & ~n28834 ) | ( n23076 & ~n28834 ) ;
  assign n28836 = n28835 ^ n15801 ^ n4279 ;
  assign n28837 = ( n14400 & n27227 ) | ( n14400 & ~n28836 ) | ( n27227 & ~n28836 ) ;
  assign n28838 = n14212 ^ n12110 ^ n10093 ;
  assign n28839 = ( n2666 & ~n23227 ) | ( n2666 & n28838 ) | ( ~n23227 & n28838 ) ;
  assign n28840 = ( n18959 & n21396 ) | ( n18959 & ~n28839 ) | ( n21396 & ~n28839 ) ;
  assign n28841 = ( ~n14740 & n17627 ) | ( ~n14740 & n28003 ) | ( n17627 & n28003 ) ;
  assign n28842 = n23226 ^ n3321 ^ n2950 ;
  assign n28843 = ( n13646 & n28057 ) | ( n13646 & ~n28842 ) | ( n28057 & ~n28842 ) ;
  assign n28844 = ( n13935 & n21368 ) | ( n13935 & ~n28843 ) | ( n21368 & ~n28843 ) ;
  assign n28845 = n12040 ^ n5607 ^ n884 ;
  assign n28846 = ( n6940 & n8020 ) | ( n6940 & ~n18332 ) | ( n8020 & ~n18332 ) ;
  assign n28847 = ( ~n15023 & n28845 ) | ( ~n15023 & n28846 ) | ( n28845 & n28846 ) ;
  assign n28848 = ( ~n5492 & n17126 ) | ( ~n5492 & n27310 ) | ( n17126 & n27310 ) ;
  assign n28850 = ( x50 & n19007 ) | ( x50 & n28429 ) | ( n19007 & n28429 ) ;
  assign n28851 = n28850 ^ n21957 ^ n11434 ;
  assign n28849 = ( n12804 & ~n15978 ) | ( n12804 & n25815 ) | ( ~n15978 & n25815 ) ;
  assign n28852 = n28851 ^ n28849 ^ n26666 ;
  assign n28853 = ( n22872 & ~n23892 ) | ( n22872 & n28852 ) | ( ~n23892 & n28852 ) ;
  assign n28854 = ( n21332 & n26902 ) | ( n21332 & n28853 ) | ( n26902 & n28853 ) ;
  assign n28855 = ( n28294 & n28848 ) | ( n28294 & ~n28854 ) | ( n28848 & ~n28854 ) ;
  assign n28856 = n17664 ^ n14445 ^ n8594 ;
  assign n28857 = ( ~n5189 & n15727 ) | ( ~n5189 & n28856 ) | ( n15727 & n28856 ) ;
  assign n28858 = ( n7982 & n9408 ) | ( n7982 & n12153 ) | ( n9408 & n12153 ) ;
  assign n28859 = n26980 ^ n26215 ^ n17602 ;
  assign n28860 = ( n1572 & n8481 ) | ( n1572 & n28425 ) | ( n8481 & n28425 ) ;
  assign n28861 = ( ~n6064 & n10627 ) | ( ~n6064 & n22657 ) | ( n10627 & n22657 ) ;
  assign n28862 = ( n1371 & n5342 ) | ( n1371 & ~n14927 ) | ( n5342 & ~n14927 ) ;
  assign n28863 = n28862 ^ n18746 ^ n8553 ;
  assign n28864 = ( n16333 & ~n18621 ) | ( n16333 & n27949 ) | ( ~n18621 & n27949 ) ;
  assign n28865 = n26139 ^ n19322 ^ n5558 ;
  assign n28866 = ( n5366 & ~n9424 ) | ( n5366 & n16335 ) | ( ~n9424 & n16335 ) ;
  assign n28867 = ( ~n27831 & n28865 ) | ( ~n27831 & n28866 ) | ( n28865 & n28866 ) ;
  assign n28868 = n28867 ^ n7890 ^ n7242 ;
  assign n28869 = ( n4336 & n11565 ) | ( n4336 & ~n26836 ) | ( n11565 & ~n26836 ) ;
  assign n28870 = ( n13360 & n27548 ) | ( n13360 & n27766 ) | ( n27548 & n27766 ) ;
  assign n28871 = ( n7340 & n11708 ) | ( n7340 & ~n28870 ) | ( n11708 & ~n28870 ) ;
  assign n28872 = ( n2341 & ~n14399 ) | ( n2341 & n27831 ) | ( ~n14399 & n27831 ) ;
  assign n28873 = n14645 ^ n5235 ^ n3089 ;
  assign n28874 = n15495 ^ n10342 ^ n5542 ;
  assign n28875 = n28874 ^ n24234 ^ n16415 ;
  assign n28876 = ( ~n5653 & n28873 ) | ( ~n5653 & n28875 ) | ( n28873 & n28875 ) ;
  assign n28877 = ( n6093 & n6125 ) | ( n6093 & ~n11701 ) | ( n6125 & ~n11701 ) ;
  assign n28878 = ( n5460 & ~n17695 ) | ( n5460 & n28877 ) | ( ~n17695 & n28877 ) ;
  assign n28879 = n17442 ^ n15515 ^ n1148 ;
  assign n28880 = ( n2337 & n11744 ) | ( n2337 & n15999 ) | ( n11744 & n15999 ) ;
  assign n28881 = ( ~n14504 & n28879 ) | ( ~n14504 & n28880 ) | ( n28879 & n28880 ) ;
  assign n28882 = ( ~n19931 & n20521 ) | ( ~n19931 & n28881 ) | ( n20521 & n28881 ) ;
  assign n28883 = n25718 ^ n15218 ^ n3085 ;
  assign n28884 = ( n3988 & n28882 ) | ( n3988 & ~n28883 ) | ( n28882 & ~n28883 ) ;
  assign n28885 = ( n7135 & ~n28878 ) | ( n7135 & n28884 ) | ( ~n28878 & n28884 ) ;
  assign n28886 = ( n3511 & n13757 ) | ( n3511 & ~n19752 ) | ( n13757 & ~n19752 ) ;
  assign n28887 = n28886 ^ n11240 ^ n4467 ;
  assign n28888 = ( ~n8050 & n26062 ) | ( ~n8050 & n27308 ) | ( n26062 & n27308 ) ;
  assign n28889 = ( ~n1079 & n9103 ) | ( ~n1079 & n22259 ) | ( n9103 & n22259 ) ;
  assign n28890 = ( ~n4622 & n6740 ) | ( ~n4622 & n10116 ) | ( n6740 & n10116 ) ;
  assign n28891 = n28890 ^ n21130 ^ n131 ;
  assign n28892 = ( n16349 & ~n28889 ) | ( n16349 & n28891 ) | ( ~n28889 & n28891 ) ;
  assign n28893 = ( ~n3164 & n12675 ) | ( ~n3164 & n28892 ) | ( n12675 & n28892 ) ;
  assign n28894 = ( n4358 & n17507 ) | ( n4358 & n23080 ) | ( n17507 & n23080 ) ;
  assign n28895 = n28894 ^ n22005 ^ n10572 ;
  assign n28896 = ( ~n716 & n1530 ) | ( ~n716 & n19330 ) | ( n1530 & n19330 ) ;
  assign n28897 = n28896 ^ n15139 ^ n10694 ;
  assign n28898 = n18133 ^ n12935 ^ n3682 ;
  assign n28899 = ( n8725 & ~n9976 ) | ( n8725 & n10165 ) | ( ~n9976 & n10165 ) ;
  assign n28900 = n12387 ^ n4669 ^ n3366 ;
  assign n28901 = n28900 ^ n16144 ^ n2569 ;
  assign n28902 = ( ~n28898 & n28899 ) | ( ~n28898 & n28901 ) | ( n28899 & n28901 ) ;
  assign n28903 = n26629 ^ n14113 ^ n5851 ;
  assign n28904 = ( n1419 & n10802 ) | ( n1419 & n28903 ) | ( n10802 & n28903 ) ;
  assign n28905 = n13053 ^ n5419 ^ n3223 ;
  assign n28906 = n14912 ^ n7123 ^ n1734 ;
  assign n28907 = ( ~n1387 & n11853 ) | ( ~n1387 & n14708 ) | ( n11853 & n14708 ) ;
  assign n28908 = ( ~n1665 & n9908 ) | ( ~n1665 & n12126 ) | ( n9908 & n12126 ) ;
  assign n28909 = ( n1168 & n3534 ) | ( n1168 & ~n28908 ) | ( n3534 & ~n28908 ) ;
  assign n28910 = ( ~n4706 & n6475 ) | ( ~n4706 & n28909 ) | ( n6475 & n28909 ) ;
  assign n28911 = ( n15605 & n23124 ) | ( n15605 & n28910 ) | ( n23124 & n28910 ) ;
  assign n28912 = n28911 ^ n13567 ^ n4544 ;
  assign n28913 = ( n3678 & ~n5618 ) | ( n3678 & n17252 ) | ( ~n5618 & n17252 ) ;
  assign n28914 = n7210 ^ n5487 ^ n3628 ;
  assign n28915 = ( n4412 & ~n17564 ) | ( n4412 & n28914 ) | ( ~n17564 & n28914 ) ;
  assign n28916 = ( n11825 & n25703 ) | ( n11825 & ~n28915 ) | ( n25703 & ~n28915 ) ;
  assign n28917 = n20114 ^ n13015 ^ n12547 ;
  assign n28918 = n7277 ^ n3681 ^ n1619 ;
  assign n28919 = n28918 ^ n28911 ^ n7100 ;
  assign n28920 = n28919 ^ n15269 ^ n535 ;
  assign n28921 = ( n1259 & n22548 ) | ( n1259 & ~n27121 ) | ( n22548 & ~n27121 ) ;
  assign n28922 = n9126 ^ n1883 ^ n587 ;
  assign n28923 = ( n15310 & n16637 ) | ( n15310 & ~n28922 ) | ( n16637 & ~n28922 ) ;
  assign n28924 = ( ~n3278 & n16101 ) | ( ~n3278 & n16608 ) | ( n16101 & n16608 ) ;
  assign n28925 = n16889 ^ n11754 ^ n6332 ;
  assign n28926 = n9518 ^ n6422 ^ n5364 ;
  assign n28927 = ( ~n3576 & n6310 ) | ( ~n3576 & n6980 ) | ( n6310 & n6980 ) ;
  assign n28928 = n28927 ^ n259 ^ x63 ;
  assign n28929 = n28928 ^ n1009 ^ n959 ;
  assign n28930 = ( n10599 & n24462 ) | ( n10599 & ~n28929 ) | ( n24462 & ~n28929 ) ;
  assign n28931 = n12503 ^ n9905 ^ n906 ;
  assign n28932 = ( n28926 & n28930 ) | ( n28926 & ~n28931 ) | ( n28930 & ~n28931 ) ;
  assign n28933 = n26920 ^ n15780 ^ n15289 ;
  assign n28934 = n25827 ^ n7966 ^ n2694 ;
  assign n28935 = ( n2955 & n6634 ) | ( n2955 & n18805 ) | ( n6634 & n18805 ) ;
  assign n28936 = n28935 ^ n23945 ^ n16700 ;
  assign n28937 = ( n4590 & ~n4902 ) | ( n4590 & n11823 ) | ( ~n4902 & n11823 ) ;
  assign n28938 = n5072 ^ n3734 ^ n1566 ;
  assign n28939 = n28938 ^ n26001 ^ n8040 ;
  assign n28940 = ( n5564 & ~n28937 ) | ( n5564 & n28939 ) | ( ~n28937 & n28939 ) ;
  assign n28941 = n25371 ^ n5252 ^ n2872 ;
  assign n28942 = ( n2269 & ~n7992 ) | ( n2269 & n11557 ) | ( ~n7992 & n11557 ) ;
  assign n28943 = ( n4864 & n28941 ) | ( n4864 & n28942 ) | ( n28941 & n28942 ) ;
  assign n28944 = n13316 ^ n6231 ^ n4690 ;
  assign n28945 = ( x107 & ~n16885 ) | ( x107 & n28944 ) | ( ~n16885 & n28944 ) ;
  assign n28946 = n9100 ^ n5159 ^ n3284 ;
  assign n28947 = n21444 ^ n14548 ^ n5830 ;
  assign n28948 = ( ~n11454 & n28946 ) | ( ~n11454 & n28947 ) | ( n28946 & n28947 ) ;
  assign n28949 = ( ~n9404 & n10566 ) | ( ~n9404 & n28948 ) | ( n10566 & n28948 ) ;
  assign n28950 = ( n1311 & n3841 ) | ( n1311 & n28949 ) | ( n3841 & n28949 ) ;
  assign n28951 = ( n9838 & ~n22307 ) | ( n9838 & n28950 ) | ( ~n22307 & n28950 ) ;
  assign n28953 = n14673 ^ n1205 ^ n563 ;
  assign n28952 = ( n1014 & ~n18434 ) | ( n1014 & n18688 ) | ( ~n18434 & n18688 ) ;
  assign n28954 = n28953 ^ n28952 ^ n27039 ;
  assign n28955 = n23456 ^ n13704 ^ n10962 ;
  assign n28956 = ( n11883 & n18414 ) | ( n11883 & ~n28955 ) | ( n18414 & ~n28955 ) ;
  assign n28957 = ( n6658 & ~n26357 ) | ( n6658 & n28956 ) | ( ~n26357 & n28956 ) ;
  assign n28959 = n12522 ^ n6904 ^ n6391 ;
  assign n28958 = n12344 ^ n7146 ^ n2824 ;
  assign n28960 = n28959 ^ n28958 ^ n2355 ;
  assign n28961 = n13169 ^ n5506 ^ n3675 ;
  assign n28962 = ( ~n6215 & n15316 ) | ( ~n6215 & n26338 ) | ( n15316 & n26338 ) ;
  assign n28963 = ( n13764 & ~n18600 ) | ( n13764 & n20183 ) | ( ~n18600 & n20183 ) ;
  assign n28964 = n17172 ^ n6189 ^ n507 ;
  assign n28965 = ( n5108 & n20008 ) | ( n5108 & n28964 ) | ( n20008 & n28964 ) ;
  assign n28966 = n20236 ^ n16159 ^ n5054 ;
  assign n28967 = ( n8851 & n13439 ) | ( n8851 & n28966 ) | ( n13439 & n28966 ) ;
  assign n28968 = n27669 ^ n27164 ^ n8391 ;
  assign n28969 = ( ~n4842 & n4942 ) | ( ~n4842 & n28968 ) | ( n4942 & n28968 ) ;
  assign n28970 = ( n16188 & n25463 ) | ( n16188 & ~n28319 ) | ( n25463 & ~n28319 ) ;
  assign n28971 = n15483 ^ n11955 ^ n307 ;
  assign n28972 = ( n11383 & n23312 ) | ( n11383 & ~n28314 ) | ( n23312 & ~n28314 ) ;
  assign n28973 = n28972 ^ n10304 ^ n3668 ;
  assign n28974 = ( n17841 & n23169 ) | ( n17841 & ~n28973 ) | ( n23169 & ~n28973 ) ;
  assign n28975 = ( ~n22388 & n28971 ) | ( ~n22388 & n28974 ) | ( n28971 & n28974 ) ;
  assign n28976 = ( n10988 & n12038 ) | ( n10988 & n12882 ) | ( n12038 & n12882 ) ;
  assign n28977 = n28976 ^ n25848 ^ n16332 ;
  assign n28978 = ( n1409 & n12286 ) | ( n1409 & n24166 ) | ( n12286 & n24166 ) ;
  assign n28979 = n18515 ^ n15419 ^ n7563 ;
  assign n28980 = n28979 ^ n19828 ^ n4718 ;
  assign n28981 = ( n5799 & n14366 ) | ( n5799 & ~n23672 ) | ( n14366 & ~n23672 ) ;
  assign n28982 = ( n13429 & n26038 ) | ( n13429 & n28981 ) | ( n26038 & n28981 ) ;
  assign n28983 = n12910 ^ n1473 ^ n1016 ;
  assign n28984 = n7421 ^ n4187 ^ n2144 ;
  assign n28985 = n23552 ^ n16302 ^ n3226 ;
  assign n28986 = ( ~n7561 & n11346 ) | ( ~n7561 & n13036 ) | ( n11346 & n13036 ) ;
  assign n28987 = ( n3194 & ~n17215 ) | ( n3194 & n19626 ) | ( ~n17215 & n19626 ) ;
  assign n28988 = n28658 ^ n27776 ^ n2519 ;
  assign n28989 = ( ~n1581 & n6980 ) | ( ~n1581 & n11662 ) | ( n6980 & n11662 ) ;
  assign n28990 = ( n4453 & ~n19875 ) | ( n4453 & n28989 ) | ( ~n19875 & n28989 ) ;
  assign n28991 = ( n7455 & n12745 ) | ( n7455 & ~n14501 ) | ( n12745 & ~n14501 ) ;
  assign n28992 = ( ~n25525 & n26850 ) | ( ~n25525 & n28991 ) | ( n26850 & n28991 ) ;
  assign n28993 = n20879 ^ n9536 ^ n4345 ;
  assign n28994 = n11306 ^ n6201 ^ n5051 ;
  assign n28995 = ( n26092 & n28013 ) | ( n26092 & n28994 ) | ( n28013 & n28994 ) ;
  assign n28996 = n28995 ^ n25160 ^ n13945 ;
  assign n28997 = ( ~n25680 & n28993 ) | ( ~n25680 & n28996 ) | ( n28993 & n28996 ) ;
  assign n28998 = ( n27451 & n28992 ) | ( n27451 & n28997 ) | ( n28992 & n28997 ) ;
  assign n28999 = ( n3193 & ~n20250 ) | ( n3193 & n21771 ) | ( ~n20250 & n21771 ) ;
  assign n29000 = ( ~n932 & n21616 ) | ( ~n932 & n28999 ) | ( n21616 & n28999 ) ;
  assign n29001 = ( n16161 & ~n17168 ) | ( n16161 & n20765 ) | ( ~n17168 & n20765 ) ;
  assign n29004 = ( n2480 & n3244 ) | ( n2480 & n5918 ) | ( n3244 & n5918 ) ;
  assign n29002 = n19701 ^ n9713 ^ n943 ;
  assign n29003 = n29002 ^ n24390 ^ n12419 ;
  assign n29005 = n29004 ^ n29003 ^ n2701 ;
  assign n29006 = ( n1729 & ~n2322 ) | ( n1729 & n13127 ) | ( ~n2322 & n13127 ) ;
  assign n29007 = n29006 ^ n5583 ^ n4536 ;
  assign n29010 = n19954 ^ n11459 ^ n6216 ;
  assign n29011 = n29010 ^ n22818 ^ n11335 ;
  assign n29008 = ( n8244 & n19409 ) | ( n8244 & n24829 ) | ( n19409 & n24829 ) ;
  assign n29009 = n29008 ^ n11019 ^ n1527 ;
  assign n29012 = n29011 ^ n29009 ^ n8198 ;
  assign n29013 = ( n11013 & n14495 ) | ( n11013 & n29012 ) | ( n14495 & n29012 ) ;
  assign n29016 = ( n1279 & n3078 ) | ( n1279 & n14599 ) | ( n3078 & n14599 ) ;
  assign n29014 = n23469 ^ n11244 ^ n5749 ;
  assign n29015 = n29014 ^ n24357 ^ n8848 ;
  assign n29017 = n29016 ^ n29015 ^ n7759 ;
  assign n29018 = ( ~n4044 & n4242 ) | ( ~n4044 & n9790 ) | ( n4242 & n9790 ) ;
  assign n29019 = n29018 ^ n4997 ^ n4768 ;
  assign n29020 = n29019 ^ n10714 ^ n3011 ;
  assign n29021 = n21319 ^ n20011 ^ n16537 ;
  assign n29022 = ( ~n5997 & n15675 ) | ( ~n5997 & n28754 ) | ( n15675 & n28754 ) ;
  assign n29023 = n8925 ^ n6446 ^ n2124 ;
  assign n29024 = n29023 ^ n11356 ^ n3034 ;
  assign n29025 = ( n7687 & ~n16266 ) | ( n7687 & n22324 ) | ( ~n16266 & n22324 ) ;
  assign n29026 = ( n5202 & n13104 ) | ( n5202 & n15460 ) | ( n13104 & n15460 ) ;
  assign n29027 = n24318 ^ n19444 ^ n11875 ;
  assign n29028 = ( n1989 & n3906 ) | ( n1989 & ~n16301 ) | ( n3906 & ~n16301 ) ;
  assign n29029 = ( n6158 & n8664 ) | ( n6158 & n11686 ) | ( n8664 & n11686 ) ;
  assign n29030 = n27825 ^ n26123 ^ n10258 ;
  assign n29031 = n24490 ^ n10068 ^ n3438 ;
  assign n29032 = n29031 ^ n23949 ^ n12916 ;
  assign n29033 = ( n1222 & n15954 ) | ( n1222 & n21796 ) | ( n15954 & n21796 ) ;
  assign n29034 = n29033 ^ n12177 ^ n693 ;
  assign n29035 = n21983 ^ n17302 ^ n4550 ;
  assign n29036 = ( n1774 & n1817 ) | ( n1774 & ~n16863 ) | ( n1817 & ~n16863 ) ;
  assign n29037 = n14986 ^ n6238 ^ n2225 ;
  assign n29038 = n29037 ^ n12918 ^ n12012 ;
  assign n29039 = ( n4808 & n13312 ) | ( n4808 & ~n14702 ) | ( n13312 & ~n14702 ) ;
  assign n29040 = n12682 ^ n10259 ^ n1932 ;
  assign n29041 = ( n6790 & n24761 ) | ( n6790 & ~n29040 ) | ( n24761 & ~n29040 ) ;
  assign n29042 = ( n3335 & ~n22111 ) | ( n3335 & n29041 ) | ( ~n22111 & n29041 ) ;
  assign n29043 = ( ~n2112 & n12739 ) | ( ~n2112 & n20480 ) | ( n12739 & n20480 ) ;
  assign n29044 = n29043 ^ n5839 ^ n4813 ;
  assign n29045 = ( n13610 & n25898 ) | ( n13610 & ~n26506 ) | ( n25898 & ~n26506 ) ;
  assign n29046 = ( n10489 & n18034 ) | ( n10489 & n21137 ) | ( n18034 & n21137 ) ;
  assign n29047 = ( n3348 & ~n13391 ) | ( n3348 & n17863 ) | ( ~n13391 & n17863 ) ;
  assign n29048 = ( ~n12834 & n22293 ) | ( ~n12834 & n24428 ) | ( n22293 & n24428 ) ;
  assign n29050 = n22935 ^ n20030 ^ n14510 ;
  assign n29049 = n7578 ^ n7025 ^ n997 ;
  assign n29051 = n29050 ^ n29049 ^ n10021 ;
  assign n29052 = ( ~n991 & n6195 ) | ( ~n991 & n27678 ) | ( n6195 & n27678 ) ;
  assign n29053 = n20281 ^ n18080 ^ n360 ;
  assign n29054 = n29053 ^ n23900 ^ n1260 ;
  assign n29055 = n29054 ^ n24013 ^ n1470 ;
  assign n29056 = ( n22234 & ~n25126 ) | ( n22234 & n27425 ) | ( ~n25126 & n27425 ) ;
  assign n29057 = n24685 ^ n18773 ^ n2863 ;
  assign n29058 = n22871 ^ n12257 ^ n9326 ;
  assign n29059 = n29058 ^ n16280 ^ n14327 ;
  assign n29060 = n18419 ^ n4101 ^ n3714 ;
  assign n29061 = n8253 ^ n2873 ^ n1130 ;
  assign n29062 = ( n434 & n6454 ) | ( n434 & ~n19476 ) | ( n6454 & ~n19476 ) ;
  assign n29063 = ( n18705 & n29061 ) | ( n18705 & ~n29062 ) | ( n29061 & ~n29062 ) ;
  assign n29064 = ( n722 & n9110 ) | ( n722 & ~n13093 ) | ( n9110 & ~n13093 ) ;
  assign n29065 = n26289 ^ n21084 ^ n1700 ;
  assign n29066 = ( n2623 & n9710 ) | ( n2623 & n18446 ) | ( n9710 & n18446 ) ;
  assign n29067 = n6803 ^ n6416 ^ x74 ;
  assign n29068 = ( n9637 & ~n29066 ) | ( n9637 & n29067 ) | ( ~n29066 & n29067 ) ;
  assign n29069 = n29068 ^ n13952 ^ n9747 ;
  assign n29070 = n23396 ^ n13123 ^ n2034 ;
  assign n29071 = n5503 ^ n760 ^ n350 ;
  assign n29072 = n25948 ^ n19425 ^ n6680 ;
  assign n29073 = ( n29070 & ~n29071 ) | ( n29070 & n29072 ) | ( ~n29071 & n29072 ) ;
  assign n29074 = n19901 ^ n2470 ^ n313 ;
  assign n29075 = n14837 ^ n14789 ^ n8622 ;
  assign n29076 = ( ~n6338 & n29074 ) | ( ~n6338 & n29075 ) | ( n29074 & n29075 ) ;
  assign n29077 = n27758 ^ n21182 ^ n20119 ;
  assign n29078 = ( n25944 & n29076 ) | ( n25944 & n29077 ) | ( n29076 & n29077 ) ;
  assign n29079 = ( n7736 & n17581 ) | ( n7736 & n29078 ) | ( n17581 & n29078 ) ;
  assign n29080 = n24763 ^ n15114 ^ n14883 ;
  assign n29081 = ( n4593 & ~n7472 ) | ( n4593 & n29080 ) | ( ~n7472 & n29080 ) ;
  assign n29082 = n19932 ^ n13498 ^ n3684 ;
  assign n29083 = ( n14276 & n24990 ) | ( n14276 & n27387 ) | ( n24990 & n27387 ) ;
  assign n29084 = ( ~n447 & n2732 ) | ( ~n447 & n21600 ) | ( n2732 & n21600 ) ;
  assign n29087 = ( n5662 & ~n9204 ) | ( n5662 & n17848 ) | ( ~n9204 & n17848 ) ;
  assign n29085 = n7361 ^ n527 ^ n490 ;
  assign n29086 = n29085 ^ n25337 ^ n4947 ;
  assign n29088 = n29087 ^ n29086 ^ n9333 ;
  assign n29089 = ( ~n5849 & n11001 ) | ( ~n5849 & n17532 ) | ( n11001 & n17532 ) ;
  assign n29090 = n29089 ^ n26858 ^ n18637 ;
  assign n29091 = n29090 ^ n24854 ^ n305 ;
  assign n29092 = n16627 ^ n11829 ^ n6427 ;
  assign n29093 = n9912 ^ n8593 ^ n8041 ;
  assign n29094 = n29093 ^ n11646 ^ n5080 ;
  assign n29095 = n9230 ^ n5855 ^ n5815 ;
  assign n29096 = ( n11073 & ~n16487 ) | ( n11073 & n29095 ) | ( ~n16487 & n29095 ) ;
  assign n29099 = n11033 ^ n4701 ^ n4690 ;
  assign n29097 = n10433 ^ n7103 ^ n1841 ;
  assign n29098 = n29097 ^ n16539 ^ n7543 ;
  assign n29100 = n29099 ^ n29098 ^ n18084 ;
  assign n29101 = ( ~n17562 & n29096 ) | ( ~n17562 & n29100 ) | ( n29096 & n29100 ) ;
  assign n29102 = ( n1422 & ~n5480 ) | ( n1422 & n10421 ) | ( ~n5480 & n10421 ) ;
  assign n29103 = ( n17410 & n23161 ) | ( n17410 & n29102 ) | ( n23161 & n29102 ) ;
  assign n29104 = n29103 ^ n18079 ^ n12559 ;
  assign n29105 = n29104 ^ n26092 ^ n5823 ;
  assign n29106 = n19353 ^ n16523 ^ n14556 ;
  assign n29107 = ( n24491 & ~n26874 ) | ( n24491 & n29106 ) | ( ~n26874 & n29106 ) ;
  assign n29108 = n9925 ^ n8322 ^ n2611 ;
  assign n29109 = ( n5312 & n5866 ) | ( n5312 & ~n29108 ) | ( n5866 & ~n29108 ) ;
  assign n29111 = ( ~n3396 & n7322 ) | ( ~n3396 & n11955 ) | ( n7322 & n11955 ) ;
  assign n29110 = n21118 ^ n15128 ^ n14413 ;
  assign n29112 = n29111 ^ n29110 ^ n1403 ;
  assign n29113 = ( n7246 & n15435 ) | ( n7246 & n29112 ) | ( n15435 & n29112 ) ;
  assign n29114 = n17365 ^ n8102 ^ x83 ;
  assign n29115 = n14214 ^ n8982 ^ n7720 ;
  assign n29116 = ( n25022 & n28136 ) | ( n25022 & ~n29115 ) | ( n28136 & ~n29115 ) ;
  assign n29117 = ( n787 & n11036 ) | ( n787 & n27037 ) | ( n11036 & n27037 ) ;
  assign n29118 = ( n4149 & n5542 ) | ( n4149 & ~n7348 ) | ( n5542 & ~n7348 ) ;
  assign n29119 = ( n7221 & ~n23381 ) | ( n7221 & n29118 ) | ( ~n23381 & n29118 ) ;
  assign n29120 = ( n813 & n29117 ) | ( n813 & ~n29119 ) | ( n29117 & ~n29119 ) ;
  assign n29121 = n20301 ^ n15353 ^ n1820 ;
  assign n29122 = ( n16564 & n24938 ) | ( n16564 & n29040 ) | ( n24938 & n29040 ) ;
  assign n29123 = ( n7104 & n15040 ) | ( n7104 & ~n17813 ) | ( n15040 & ~n17813 ) ;
  assign n29124 = ( ~n2259 & n11476 ) | ( ~n2259 & n14369 ) | ( n11476 & n14369 ) ;
  assign n29125 = ( ~n11764 & n26640 ) | ( ~n11764 & n29124 ) | ( n26640 & n29124 ) ;
  assign n29126 = ( n1067 & n5108 ) | ( n1067 & n16355 ) | ( n5108 & n16355 ) ;
  assign n29127 = n29126 ^ n19409 ^ n4210 ;
  assign n29128 = n29127 ^ n14713 ^ n3190 ;
  assign n29130 = n17199 ^ n1756 ^ n1320 ;
  assign n29129 = ( n1536 & ~n15301 ) | ( n1536 & n16779 ) | ( ~n15301 & n16779 ) ;
  assign n29131 = n29130 ^ n29129 ^ n21398 ;
  assign n29132 = n14984 ^ n5866 ^ n4097 ;
  assign n29133 = n29132 ^ n25431 ^ n21667 ;
  assign n29134 = ( n25475 & n29131 ) | ( n25475 & ~n29133 ) | ( n29131 & ~n29133 ) ;
  assign n29135 = n19905 ^ n19123 ^ n7763 ;
  assign n29136 = n20755 ^ n12576 ^ n4010 ;
  assign n29137 = ( n13383 & ~n16918 ) | ( n13383 & n29136 ) | ( ~n16918 & n29136 ) ;
  assign n29138 = ( n15540 & n24462 ) | ( n15540 & ~n29137 ) | ( n24462 & ~n29137 ) ;
  assign n29139 = ( n16862 & n29135 ) | ( n16862 & ~n29138 ) | ( n29135 & ~n29138 ) ;
  assign n29140 = n12668 ^ n8801 ^ n8285 ;
  assign n29141 = n28659 ^ n3434 ^ n2492 ;
  assign n29142 = n26477 ^ n13796 ^ n272 ;
  assign n29143 = ( ~n25983 & n29141 ) | ( ~n25983 & n29142 ) | ( n29141 & n29142 ) ;
  assign n29144 = n21737 ^ n19774 ^ n18479 ;
  assign n29145 = n8032 ^ n3430 ^ n1974 ;
  assign n29146 = ( n3416 & n21036 ) | ( n3416 & ~n29145 ) | ( n21036 & ~n29145 ) ;
  assign n29147 = n29146 ^ n9731 ^ n1511 ;
  assign n29148 = n26864 ^ n25409 ^ n13165 ;
  assign n29149 = n22046 ^ n5302 ^ x11 ;
  assign n29150 = n25504 ^ n14710 ^ n355 ;
  assign n29151 = ( n4596 & ~n5509 ) | ( n4596 & n6420 ) | ( ~n5509 & n6420 ) ;
  assign n29152 = ( ~n1100 & n3586 ) | ( ~n1100 & n29151 ) | ( n3586 & n29151 ) ;
  assign n29153 = ( n3695 & n4811 ) | ( n3695 & ~n19766 ) | ( n4811 & ~n19766 ) ;
  assign n29154 = n8510 ^ n6226 ^ n3199 ;
  assign n29155 = ( n2648 & ~n23621 ) | ( n2648 & n29154 ) | ( ~n23621 & n29154 ) ;
  assign n29156 = ( n8627 & ~n8955 ) | ( n8627 & n21207 ) | ( ~n8955 & n21207 ) ;
  assign n29157 = n29156 ^ n19053 ^ n4682 ;
  assign n29158 = n26409 ^ n11707 ^ n2445 ;
  assign n29159 = ( n1637 & n28180 ) | ( n1637 & n29158 ) | ( n28180 & n29158 ) ;
  assign n29160 = n8243 ^ n6917 ^ n2289 ;
  assign n29161 = ( n1627 & n19638 ) | ( n1627 & n29160 ) | ( n19638 & n29160 ) ;
  assign n29162 = n9206 ^ n1430 ^ n191 ;
  assign n29163 = ( n8206 & ~n17566 ) | ( n8206 & n29162 ) | ( ~n17566 & n29162 ) ;
  assign n29164 = ( ~n3385 & n7217 ) | ( ~n3385 & n29163 ) | ( n7217 & n29163 ) ;
  assign n29165 = n29164 ^ n21372 ^ n14365 ;
  assign n29166 = ( n11986 & n17343 ) | ( n11986 & n18382 ) | ( n17343 & n18382 ) ;
  assign n29167 = ( n1866 & n20683 ) | ( n1866 & n29166 ) | ( n20683 & n29166 ) ;
  assign n29168 = ( n5421 & n10788 ) | ( n5421 & n29167 ) | ( n10788 & n29167 ) ;
  assign n29169 = ( n7475 & n13896 ) | ( n7475 & n28653 ) | ( n13896 & n28653 ) ;
  assign n29170 = ( n27983 & ~n29168 ) | ( n27983 & n29169 ) | ( ~n29168 & n29169 ) ;
  assign n29171 = ( n2752 & n7231 ) | ( n2752 & n20194 ) | ( n7231 & n20194 ) ;
  assign n29172 = ( n11056 & n16965 ) | ( n11056 & ~n18142 ) | ( n16965 & ~n18142 ) ;
  assign n29173 = ( n22081 & ~n25184 ) | ( n22081 & n29172 ) | ( ~n25184 & n29172 ) ;
  assign n29174 = n29173 ^ n26547 ^ n3459 ;
  assign n29175 = n19780 ^ n1894 ^ n1736 ;
  assign n29176 = n29175 ^ n22749 ^ n17980 ;
  assign n29177 = n16272 ^ n4386 ^ n2746 ;
  assign n29178 = ( n5770 & n18583 ) | ( n5770 & ~n29177 ) | ( n18583 & ~n29177 ) ;
  assign n29179 = n10673 ^ n4350 ^ n274 ;
  assign n29180 = ( n23900 & n25074 ) | ( n23900 & ~n29179 ) | ( n25074 & ~n29179 ) ;
  assign n29181 = ( n2854 & n19651 ) | ( n2854 & n29180 ) | ( n19651 & n29180 ) ;
  assign n29183 = n25689 ^ n16288 ^ n11758 ;
  assign n29182 = n15201 ^ n6464 ^ n2583 ;
  assign n29184 = n29183 ^ n29182 ^ n16917 ;
  assign n29185 = n19431 ^ n15772 ^ n7675 ;
  assign n29186 = n5858 ^ n4843 ^ n4604 ;
  assign n29187 = ( n5066 & n16671 ) | ( n5066 & n21398 ) | ( n16671 & n21398 ) ;
  assign n29188 = ( ~n1333 & n8189 ) | ( ~n1333 & n21902 ) | ( n8189 & n21902 ) ;
  assign n29189 = ( n12480 & n21652 ) | ( n12480 & n29188 ) | ( n21652 & n29188 ) ;
  assign n29190 = ( n2680 & ~n6748 ) | ( n2680 & n13974 ) | ( ~n6748 & n13974 ) ;
  assign n29191 = n20463 ^ n13801 ^ n11509 ;
  assign n29192 = ( n1710 & n6280 ) | ( n1710 & ~n13233 ) | ( n6280 & ~n13233 ) ;
  assign n29194 = ( n9704 & n16033 ) | ( n9704 & ~n16063 ) | ( n16033 & ~n16063 ) ;
  assign n29193 = ( n1725 & n6593 ) | ( n1725 & ~n9878 ) | ( n6593 & ~n9878 ) ;
  assign n29195 = n29194 ^ n29193 ^ n1323 ;
  assign n29196 = ( ~n10468 & n11779 ) | ( ~n10468 & n18173 ) | ( n11779 & n18173 ) ;
  assign n29197 = n29196 ^ n3489 ^ n141 ;
  assign n29198 = n29197 ^ n14126 ^ n6465 ;
  assign n29199 = ( ~n13811 & n14132 ) | ( ~n13811 & n21888 ) | ( n14132 & n21888 ) ;
  assign n29200 = ( ~n2207 & n11182 ) | ( ~n2207 & n17785 ) | ( n11182 & n17785 ) ;
  assign n29201 = n8791 ^ n6077 ^ n3810 ;
  assign n29202 = ( n5559 & n29200 ) | ( n5559 & n29201 ) | ( n29200 & n29201 ) ;
  assign n29203 = ( n6370 & n26805 ) | ( n6370 & ~n27572 ) | ( n26805 & ~n27572 ) ;
  assign n29204 = ( n2943 & n8898 ) | ( n2943 & ~n9630 ) | ( n8898 & ~n9630 ) ;
  assign n29205 = ( x15 & ~n3641 ) | ( x15 & n5980 ) | ( ~n3641 & n5980 ) ;
  assign n29206 = n9441 ^ n4222 ^ n305 ;
  assign n29207 = ( ~n16511 & n29205 ) | ( ~n16511 & n29206 ) | ( n29205 & n29206 ) ;
  assign n29208 = ( n408 & ~n15675 ) | ( n408 & n17815 ) | ( ~n15675 & n17815 ) ;
  assign n29209 = n12154 ^ n6980 ^ n3020 ;
  assign n29210 = n21560 ^ n4209 ^ n2045 ;
  assign n29211 = n29210 ^ n21851 ^ n4883 ;
  assign n29212 = ( ~x105 & n29209 ) | ( ~x105 & n29211 ) | ( n29209 & n29211 ) ;
  assign n29213 = n29212 ^ n26627 ^ n22045 ;
  assign n29214 = n14257 ^ n12288 ^ n4108 ;
  assign n29215 = ( n7538 & n9793 ) | ( n7538 & ~n29214 ) | ( n9793 & ~n29214 ) ;
  assign n29216 = ( ~n901 & n5327 ) | ( ~n901 & n9315 ) | ( n5327 & n9315 ) ;
  assign n29217 = n29216 ^ n15440 ^ n5354 ;
  assign n29218 = ( n16296 & ~n25920 ) | ( n16296 & n29217 ) | ( ~n25920 & n29217 ) ;
  assign n29219 = n29218 ^ n28594 ^ n548 ;
  assign n29220 = n28937 ^ n14122 ^ n10518 ;
  assign n29221 = n29220 ^ n26453 ^ n15116 ;
  assign n29222 = n15867 ^ n9500 ^ n637 ;
  assign n29223 = ( n493 & n9793 ) | ( n493 & n13027 ) | ( n9793 & n13027 ) ;
  assign n29224 = n29223 ^ n15338 ^ n9517 ;
  assign n29225 = ( n3383 & n6823 ) | ( n3383 & n29224 ) | ( n6823 & n29224 ) ;
  assign n29228 = n24289 ^ n1338 ^ n158 ;
  assign n29226 = ( n2675 & n5155 ) | ( n2675 & n6125 ) | ( n5155 & n6125 ) ;
  assign n29227 = n29226 ^ n16817 ^ n5364 ;
  assign n29229 = n29228 ^ n29227 ^ n28433 ;
  assign n29230 = n16420 ^ n3267 ^ n1205 ;
  assign n29231 = n6213 ^ n6083 ^ n5857 ;
  assign n29232 = n19347 ^ n19048 ^ n3735 ;
  assign n29233 = ( n17372 & ~n29231 ) | ( n17372 & n29232 ) | ( ~n29231 & n29232 ) ;
  assign n29234 = n25942 ^ n17710 ^ n16572 ;
  assign n29235 = ( n1676 & n4686 ) | ( n1676 & n28587 ) | ( n4686 & n28587 ) ;
  assign n29236 = n29235 ^ n2324 ^ n964 ;
  assign n29238 = n12852 ^ n10598 ^ n9785 ;
  assign n29239 = n29238 ^ n24969 ^ n23387 ;
  assign n29237 = ( n3724 & n5437 ) | ( n3724 & ~n24610 ) | ( n5437 & ~n24610 ) ;
  assign n29240 = n29239 ^ n29237 ^ n1672 ;
  assign n29241 = ( n10744 & ~n22215 ) | ( n10744 & n29240 ) | ( ~n22215 & n29240 ) ;
  assign n29242 = n25701 ^ n20435 ^ n7503 ;
  assign n29243 = ( ~n467 & n3830 ) | ( ~n467 & n6754 ) | ( n3830 & n6754 ) ;
  assign n29244 = n13270 ^ n11162 ^ n10477 ;
  assign n29245 = ( n13494 & n29243 ) | ( n13494 & ~n29244 ) | ( n29243 & ~n29244 ) ;
  assign n29246 = ( n11036 & n13322 ) | ( n11036 & ~n29245 ) | ( n13322 & ~n29245 ) ;
  assign n29247 = n29246 ^ n13636 ^ n8883 ;
  assign n29248 = n20160 ^ n13585 ^ n12402 ;
  assign n29249 = ( n5388 & ~n18283 ) | ( n5388 & n25625 ) | ( ~n18283 & n25625 ) ;
  assign n29250 = n15197 ^ n14255 ^ n5541 ;
  assign n29251 = ( n14425 & ~n21475 ) | ( n14425 & n23718 ) | ( ~n21475 & n23718 ) ;
  assign n29252 = ( n28152 & n29250 ) | ( n28152 & n29251 ) | ( n29250 & n29251 ) ;
  assign n29253 = n29252 ^ n20445 ^ n6716 ;
  assign n29256 = ( ~n375 & n2174 ) | ( ~n375 & n3939 ) | ( n2174 & n3939 ) ;
  assign n29254 = n15706 ^ n13016 ^ n9496 ;
  assign n29255 = ( n5506 & ~n5955 ) | ( n5506 & n29254 ) | ( ~n5955 & n29254 ) ;
  assign n29257 = n29256 ^ n29255 ^ n2531 ;
  assign n29258 = n18220 ^ n5695 ^ n1103 ;
  assign n29259 = n28512 ^ n15713 ^ n3475 ;
  assign n29260 = ( n3517 & n11544 ) | ( n3517 & n23345 ) | ( n11544 & n23345 ) ;
  assign n29262 = n6714 ^ n5195 ^ n3257 ;
  assign n29261 = ( n7450 & n21292 ) | ( n7450 & ~n25834 ) | ( n21292 & ~n25834 ) ;
  assign n29263 = n29262 ^ n29261 ^ n20271 ;
  assign n29264 = ( ~n2190 & n17697 ) | ( ~n2190 & n29262 ) | ( n17697 & n29262 ) ;
  assign n29265 = n29264 ^ n11451 ^ n7024 ;
  assign n29266 = ( n4909 & n12725 ) | ( n4909 & n25236 ) | ( n12725 & n25236 ) ;
  assign n29267 = ( n1630 & ~n10878 ) | ( n1630 & n29266 ) | ( ~n10878 & n29266 ) ;
  assign n29268 = ( n769 & n1204 ) | ( n769 & ~n7569 ) | ( n1204 & ~n7569 ) ;
  assign n29269 = n29268 ^ n10525 ^ n5905 ;
  assign n29270 = n10796 ^ n2186 ^ n394 ;
  assign n29271 = ( ~n2358 & n20158 ) | ( ~n2358 & n27812 ) | ( n20158 & n27812 ) ;
  assign n29272 = n29271 ^ n18460 ^ n15301 ;
  assign n29273 = n25642 ^ n15813 ^ n3182 ;
  assign n29274 = ( n3884 & ~n13115 ) | ( n3884 & n14420 ) | ( ~n13115 & n14420 ) ;
  assign n29275 = n17731 ^ n3749 ^ n353 ;
  assign n29276 = n29275 ^ n2029 ^ n787 ;
  assign n29277 = n16596 ^ n4247 ^ n1233 ;
  assign n29278 = n29277 ^ n21755 ^ n5348 ;
  assign n29279 = ( n7501 & n18876 ) | ( n7501 & ~n29278 ) | ( n18876 & ~n29278 ) ;
  assign n29280 = n27708 ^ n26804 ^ n17373 ;
  assign n29281 = ( n4833 & ~n6561 ) | ( n4833 & n14357 ) | ( ~n6561 & n14357 ) ;
  assign n29282 = ( n5422 & n10792 ) | ( n5422 & n29281 ) | ( n10792 & n29281 ) ;
  assign n29283 = ( n3471 & n5975 ) | ( n3471 & n10259 ) | ( n5975 & n10259 ) ;
  assign n29284 = ( ~n240 & n7147 ) | ( ~n240 & n29283 ) | ( n7147 & n29283 ) ;
  assign n29285 = n29284 ^ n19494 ^ n14896 ;
  assign n29286 = ( n2076 & n8039 ) | ( n2076 & ~n14460 ) | ( n8039 & ~n14460 ) ;
  assign n29287 = n29286 ^ n25067 ^ n4342 ;
  assign n29288 = n12750 ^ n6932 ^ n6404 ;
  assign n29289 = n29288 ^ n19364 ^ n1082 ;
  assign n29290 = ( ~n2659 & n22382 ) | ( ~n2659 & n29289 ) | ( n22382 & n29289 ) ;
  assign n29291 = n26639 ^ n17747 ^ n565 ;
  assign n29292 = n29291 ^ n25941 ^ n8931 ;
  assign n29293 = ( ~n2892 & n12095 ) | ( ~n2892 & n29062 ) | ( n12095 & n29062 ) ;
  assign n29294 = ( n28599 & n29292 ) | ( n28599 & n29293 ) | ( n29292 & n29293 ) ;
  assign n29295 = n20478 ^ n13474 ^ n12643 ;
  assign n29296 = ( n705 & ~n7185 ) | ( n705 & n15018 ) | ( ~n7185 & n15018 ) ;
  assign n29297 = ( n12197 & n14411 ) | ( n12197 & n29296 ) | ( n14411 & n29296 ) ;
  assign n29298 = ( ~n16862 & n18281 ) | ( ~n16862 & n20941 ) | ( n18281 & n20941 ) ;
  assign n29299 = n29298 ^ n29054 ^ n26444 ;
  assign n29300 = n18944 ^ n5936 ^ n4541 ;
  assign n29301 = ( n3387 & n20280 ) | ( n3387 & ~n29300 ) | ( n20280 & ~n29300 ) ;
  assign n29302 = n29301 ^ n24292 ^ n2412 ;
  assign n29303 = n18083 ^ n10458 ^ n8694 ;
  assign n29304 = n29303 ^ n25407 ^ n24831 ;
  assign n29305 = ( n12626 & n16325 ) | ( n12626 & ~n27193 ) | ( n16325 & ~n27193 ) ;
  assign n29306 = n12560 ^ n8552 ^ n2683 ;
  assign n29307 = ( n3292 & n4307 ) | ( n3292 & ~n29306 ) | ( n4307 & ~n29306 ) ;
  assign n29308 = n29307 ^ n28354 ^ n10373 ;
  assign n29309 = ( n8045 & n16654 ) | ( n8045 & n29308 ) | ( n16654 & n29308 ) ;
  assign n29310 = n21925 ^ n19566 ^ n19445 ;
  assign n29311 = n29310 ^ n28972 ^ n12424 ;
  assign n29312 = ( n4005 & n16072 ) | ( n4005 & n18852 ) | ( n16072 & n18852 ) ;
  assign n29313 = n18020 ^ n11419 ^ x107 ;
  assign n29314 = n29313 ^ n21060 ^ n20895 ;
  assign n29315 = ( n10298 & ~n16155 ) | ( n10298 & n29314 ) | ( ~n16155 & n29314 ) ;
  assign n29316 = n29315 ^ n18883 ^ n14251 ;
  assign n29317 = ( n8539 & ~n9168 ) | ( n8539 & n15148 ) | ( ~n9168 & n15148 ) ;
  assign n29318 = n29317 ^ n26453 ^ n14198 ;
  assign n29319 = n24536 ^ n12596 ^ n9265 ;
  assign n29320 = n29319 ^ n19720 ^ n18345 ;
  assign n29321 = n17943 ^ n9239 ^ n9100 ;
  assign n29322 = ( ~n19882 & n23849 ) | ( ~n19882 & n29321 ) | ( n23849 & n29321 ) ;
  assign n29323 = n11737 ^ n1384 ^ n546 ;
  assign n29324 = ( n14548 & n18783 ) | ( n14548 & ~n29323 ) | ( n18783 & ~n29323 ) ;
  assign n29325 = ( ~n7368 & n8557 ) | ( ~n7368 & n20639 ) | ( n8557 & n20639 ) ;
  assign n29326 = ( n8551 & n19753 ) | ( n8551 & ~n29325 ) | ( n19753 & ~n29325 ) ;
  assign n29327 = n24795 ^ n18596 ^ n7357 ;
  assign n29328 = ( n456 & n26799 ) | ( n456 & ~n29327 ) | ( n26799 & ~n29327 ) ;
  assign n29329 = ( ~n21206 & n27316 ) | ( ~n21206 & n29328 ) | ( n27316 & n29328 ) ;
  assign n29330 = ( n14124 & n29326 ) | ( n14124 & n29329 ) | ( n29326 & n29329 ) ;
  assign n29331 = n8997 ^ n6904 ^ n2141 ;
  assign n29332 = n18730 ^ n13245 ^ n12992 ;
  assign n29333 = n29332 ^ n16941 ^ n15114 ;
  assign n29334 = n24610 ^ n7858 ^ n1802 ;
  assign n29335 = ( n4609 & ~n26505 ) | ( n4609 & n29334 ) | ( ~n26505 & n29334 ) ;
  assign n29336 = n14025 ^ n8734 ^ n7914 ;
  assign n29337 = n29336 ^ n11079 ^ n5684 ;
  assign n29338 = n21923 ^ n13251 ^ n3683 ;
  assign n29339 = n15893 ^ n9728 ^ n5195 ;
  assign n29340 = n29339 ^ n26006 ^ n17460 ;
  assign n29341 = ( n3975 & n17160 ) | ( n3975 & ~n29340 ) | ( n17160 & ~n29340 ) ;
  assign n29342 = n26704 ^ n20951 ^ n5205 ;
  assign n29343 = n29342 ^ n24608 ^ n8432 ;
  assign n29344 = n20869 ^ n16757 ^ n1828 ;
  assign n29345 = n20530 ^ n9741 ^ n2973 ;
  assign n29346 = ( n17934 & n18191 ) | ( n17934 & n29345 ) | ( n18191 & n29345 ) ;
  assign n29347 = ( n26770 & n29344 ) | ( n26770 & ~n29346 ) | ( n29344 & ~n29346 ) ;
  assign n29348 = n12483 ^ n12100 ^ n1144 ;
  assign n29349 = n29348 ^ n25209 ^ n17540 ;
  assign n29350 = n29349 ^ n3080 ^ n2102 ;
  assign n29351 = ( n5963 & n7531 ) | ( n5963 & n26177 ) | ( n7531 & n26177 ) ;
  assign n29352 = ( x41 & n7895 ) | ( x41 & n13203 ) | ( n7895 & n13203 ) ;
  assign n29353 = n18721 ^ n9454 ^ n3479 ;
  assign n29354 = n26557 ^ n25351 ^ n17879 ;
  assign n29355 = ( n6819 & n9466 ) | ( n6819 & n29354 ) | ( n9466 & n29354 ) ;
  assign n29356 = ( n6122 & ~n29353 ) | ( n6122 & n29355 ) | ( ~n29353 & n29355 ) ;
  assign n29357 = ( ~n20233 & n27482 ) | ( ~n20233 & n29356 ) | ( n27482 & n29356 ) ;
  assign n29358 = ( ~n5552 & n7154 ) | ( ~n5552 & n9180 ) | ( n7154 & n9180 ) ;
  assign n29359 = n15644 ^ n6032 ^ n3964 ;
  assign n29360 = ( ~n1380 & n8992 ) | ( ~n1380 & n11826 ) | ( n8992 & n11826 ) ;
  assign n29361 = n22557 ^ n13311 ^ n2365 ;
  assign n29362 = n26836 ^ n17397 ^ n13493 ;
  assign n29363 = ( n2687 & n13116 ) | ( n2687 & n29362 ) | ( n13116 & n29362 ) ;
  assign n29364 = ( n1189 & n5061 ) | ( n1189 & ~n21912 ) | ( n5061 & ~n21912 ) ;
  assign n29365 = ( n602 & ~n680 ) | ( n602 & n21753 ) | ( ~n680 & n21753 ) ;
  assign n29366 = ( ~n11915 & n29364 ) | ( ~n11915 & n29365 ) | ( n29364 & n29365 ) ;
  assign n29368 = ( ~n5617 & n8553 ) | ( ~n5617 & n20791 ) | ( n8553 & n20791 ) ;
  assign n29367 = n29264 ^ n18260 ^ n1739 ;
  assign n29369 = n29368 ^ n29367 ^ n10368 ;
  assign n29370 = n13614 ^ n6514 ^ n5813 ;
  assign n29371 = n29370 ^ n27693 ^ n18751 ;
  assign n29372 = ( n13261 & ~n23492 ) | ( n13261 & n29371 ) | ( ~n23492 & n29371 ) ;
  assign n29373 = n29372 ^ n9245 ^ n8876 ;
  assign n29374 = ( ~n4475 & n8491 ) | ( ~n4475 & n23141 ) | ( n8491 & n23141 ) ;
  assign n29375 = ( ~x99 & n7219 ) | ( ~x99 & n29374 ) | ( n7219 & n29374 ) ;
  assign n29376 = ( n2498 & ~n11786 ) | ( n2498 & n29375 ) | ( ~n11786 & n29375 ) ;
  assign n29377 = ( n16856 & ~n19674 ) | ( n16856 & n29376 ) | ( ~n19674 & n29376 ) ;
  assign n29378 = n23731 ^ n11838 ^ n10941 ;
  assign n29379 = ( n9565 & n29377 ) | ( n9565 & n29378 ) | ( n29377 & n29378 ) ;
  assign n29380 = n16391 ^ n10353 ^ n4555 ;
  assign n29381 = n18258 ^ n9561 ^ n3160 ;
  assign n29382 = ( n3354 & n6660 ) | ( n3354 & ~n19403 ) | ( n6660 & ~n19403 ) ;
  assign n29385 = n16852 ^ n13522 ^ n2440 ;
  assign n29383 = ( ~n8153 & n10795 ) | ( ~n8153 & n12193 ) | ( n10795 & n12193 ) ;
  assign n29384 = ( n22228 & ~n22944 ) | ( n22228 & n29383 ) | ( ~n22944 & n29383 ) ;
  assign n29386 = n29385 ^ n29384 ^ n13962 ;
  assign n29387 = ( n778 & ~n6714 ) | ( n778 & n25258 ) | ( ~n6714 & n25258 ) ;
  assign n29388 = ( n14788 & ~n16453 ) | ( n14788 & n29387 ) | ( ~n16453 & n29387 ) ;
  assign n29389 = ( ~n258 & n11797 ) | ( ~n258 & n27145 ) | ( n11797 & n27145 ) ;
  assign n29390 = ( n1701 & ~n22086 ) | ( n1701 & n25662 ) | ( ~n22086 & n25662 ) ;
  assign n29391 = ( n8270 & ~n17695 ) | ( n8270 & n23669 ) | ( ~n17695 & n23669 ) ;
  assign n29392 = n16885 ^ n11485 ^ n10764 ;
  assign n29393 = ( ~n6159 & n27888 ) | ( ~n6159 & n29392 ) | ( n27888 & n29392 ) ;
  assign n29394 = n29393 ^ n17730 ^ n2532 ;
  assign n29395 = n18059 ^ n10479 ^ n861 ;
  assign n29396 = n29395 ^ n4325 ^ n418 ;
  assign n29397 = n24225 ^ n11491 ^ n666 ;
  assign n29398 = n29397 ^ n20207 ^ n8761 ;
  assign n29399 = ( n6919 & n14028 ) | ( n6919 & n29398 ) | ( n14028 & n29398 ) ;
  assign n29400 = ( n5291 & ~n5930 ) | ( n5291 & n12533 ) | ( ~n5930 & n12533 ) ;
  assign n29401 = n26631 ^ n16485 ^ n11663 ;
  assign n29402 = n19694 ^ n6009 ^ n5470 ;
  assign n29403 = ( n1228 & n1980 ) | ( n1228 & n10645 ) | ( n1980 & n10645 ) ;
  assign n29404 = ( n2795 & n18106 ) | ( n2795 & n28886 ) | ( n18106 & n28886 ) ;
  assign n29405 = ( n29402 & ~n29403 ) | ( n29402 & n29404 ) | ( ~n29403 & n29404 ) ;
  assign n29406 = ( n20540 & ~n21891 ) | ( n20540 & n23955 ) | ( ~n21891 & n23955 ) ;
  assign n29407 = n20934 ^ n12603 ^ n8704 ;
  assign n29408 = ( ~n26640 & n29406 ) | ( ~n26640 & n29407 ) | ( n29406 & n29407 ) ;
  assign n29409 = ( n3510 & n16218 ) | ( n3510 & ~n27067 ) | ( n16218 & ~n27067 ) ;
  assign n29410 = ( n9846 & n12672 ) | ( n9846 & n16889 ) | ( n12672 & n16889 ) ;
  assign n29411 = n29410 ^ n6636 ^ n6217 ;
  assign n29412 = ( n9069 & n10307 ) | ( n9069 & n13684 ) | ( n10307 & n13684 ) ;
  assign n29413 = n8638 ^ n7678 ^ n3084 ;
  assign n29414 = ( n1024 & n15682 ) | ( n1024 & n17501 ) | ( n15682 & n17501 ) ;
  assign n29415 = n29414 ^ n3902 ^ n2129 ;
  assign n29416 = ( n14413 & n16816 ) | ( n14413 & ~n18973 ) | ( n16816 & ~n18973 ) ;
  assign n29417 = n24784 ^ n17100 ^ n16540 ;
  assign n29418 = ( n11635 & n20478 ) | ( n11635 & ~n24630 ) | ( n20478 & ~n24630 ) ;
  assign n29419 = n16167 ^ n6833 ^ n1464 ;
  assign n29420 = ( n23737 & ~n24285 ) | ( n23737 & n29419 ) | ( ~n24285 & n29419 ) ;
  assign n29421 = n11235 ^ n5025 ^ n1073 ;
  assign n29422 = ( n9786 & n17734 ) | ( n9786 & ~n29421 ) | ( n17734 & ~n29421 ) ;
  assign n29424 = ( ~n268 & n11156 ) | ( ~n268 & n17622 ) | ( n11156 & n17622 ) ;
  assign n29423 = n11522 ^ n3852 ^ n744 ;
  assign n29425 = n29424 ^ n29423 ^ n13843 ;
  assign n29426 = ( ~n14117 & n29422 ) | ( ~n14117 & n29425 ) | ( n29422 & n29425 ) ;
  assign n29427 = n24761 ^ n17130 ^ n11033 ;
  assign n29428 = ( n3388 & ~n11003 ) | ( n3388 & n22363 ) | ( ~n11003 & n22363 ) ;
  assign n29429 = ( n3840 & n7362 ) | ( n3840 & n29428 ) | ( n7362 & n29428 ) ;
  assign n29433 = n21867 ^ n2522 ^ n1268 ;
  assign n29432 = ( n10409 & n12192 ) | ( n10409 & n16472 ) | ( n12192 & n16472 ) ;
  assign n29430 = n12492 ^ n12275 ^ n2030 ;
  assign n29431 = ( n10151 & ~n21576 ) | ( n10151 & n29430 ) | ( ~n21576 & n29430 ) ;
  assign n29434 = n29433 ^ n29432 ^ n29431 ;
  assign n29435 = n27555 ^ n11202 ^ n9637 ;
  assign n29436 = n16403 ^ n13341 ^ n10558 ;
  assign n29437 = ( n1946 & n9066 ) | ( n1946 & ~n17022 ) | ( n9066 & ~n17022 ) ;
  assign n29438 = n29437 ^ n19511 ^ n5314 ;
  assign n29439 = n24769 ^ n17897 ^ n3216 ;
  assign n29440 = ( n1048 & n7020 ) | ( n1048 & n16488 ) | ( n7020 & n16488 ) ;
  assign n29441 = ( n1499 & ~n20701 ) | ( n1499 & n29440 ) | ( ~n20701 & n29440 ) ;
  assign n29442 = n26641 ^ n19471 ^ n13532 ;
  assign n29443 = n29442 ^ n16156 ^ n2301 ;
  assign n29444 = n29443 ^ n16554 ^ n3888 ;
  assign n29445 = ( n279 & n1479 ) | ( n279 & ~n6752 ) | ( n1479 & ~n6752 ) ;
  assign n29446 = ( n3873 & ~n12755 ) | ( n3873 & n29445 ) | ( ~n12755 & n29445 ) ;
  assign n29447 = n28255 ^ n25178 ^ n17724 ;
  assign n29448 = ( n416 & n15087 ) | ( n416 & ~n27906 ) | ( n15087 & ~n27906 ) ;
  assign n29449 = ( n9865 & n12210 ) | ( n9865 & ~n29448 ) | ( n12210 & ~n29448 ) ;
  assign n29450 = ( n5700 & ~n15151 ) | ( n5700 & n18752 ) | ( ~n15151 & n18752 ) ;
  assign n29451 = ( n11767 & n16562 ) | ( n11767 & ~n29450 ) | ( n16562 & ~n29450 ) ;
  assign n29452 = n20422 ^ n15927 ^ n173 ;
  assign n29453 = n29452 ^ n27561 ^ n15895 ;
  assign n29454 = n26081 ^ n15852 ^ x27 ;
  assign n29455 = ( n5836 & ~n21748 ) | ( n5836 & n22592 ) | ( ~n21748 & n22592 ) ;
  assign n29456 = ( n593 & ~n5652 ) | ( n593 & n19086 ) | ( ~n5652 & n19086 ) ;
  assign n29457 = n29328 ^ n19201 ^ n953 ;
  assign n29458 = ( n29455 & n29456 ) | ( n29455 & n29457 ) | ( n29456 & n29457 ) ;
  assign n29459 = n25328 ^ n15876 ^ n2783 ;
  assign n29460 = ( ~n1429 & n2981 ) | ( ~n1429 & n13888 ) | ( n2981 & n13888 ) ;
  assign n29461 = n29460 ^ n13506 ^ n11253 ;
  assign n29462 = n19602 ^ n17226 ^ n12848 ;
  assign n29463 = n14263 ^ n11663 ^ n137 ;
  assign n29464 = n29463 ^ n26059 ^ n21918 ;
  assign n29465 = ( n3126 & n17652 ) | ( n3126 & n29464 ) | ( n17652 & n29464 ) ;
  assign n29466 = ( ~n1945 & n17652 ) | ( ~n1945 & n21006 ) | ( n17652 & n21006 ) ;
  assign n29467 = ( n18960 & ~n19952 ) | ( n18960 & n29466 ) | ( ~n19952 & n29466 ) ;
  assign n29468 = ( ~n8185 & n19969 ) | ( ~n8185 & n23132 ) | ( n19969 & n23132 ) ;
  assign n29469 = ( ~n9198 & n15630 ) | ( ~n9198 & n29468 ) | ( n15630 & n29468 ) ;
  assign n29470 = ( ~n5644 & n11032 ) | ( ~n5644 & n17260 ) | ( n11032 & n17260 ) ;
  assign n29471 = n29470 ^ n14630 ^ n2572 ;
  assign n29472 = n28899 ^ n11720 ^ n1087 ;
  assign n29473 = ( ~n2920 & n3205 ) | ( ~n2920 & n3641 ) | ( n3205 & n3641 ) ;
  assign n29474 = ( ~n6466 & n20870 ) | ( ~n6466 & n29473 ) | ( n20870 & n29473 ) ;
  assign n29475 = n13328 ^ n10591 ^ n2841 ;
  assign n29476 = n7301 ^ n3897 ^ n3163 ;
  assign n29477 = ( ~n4385 & n11564 ) | ( ~n4385 & n29476 ) | ( n11564 & n29476 ) ;
  assign n29478 = n23689 ^ n11481 ^ n10701 ;
  assign n29479 = n20143 ^ n15644 ^ n7748 ;
  assign n29480 = n29479 ^ n22325 ^ n19134 ;
  assign n29481 = ( n623 & n17614 ) | ( n623 & ~n18032 ) | ( n17614 & ~n18032 ) ;
  assign n29482 = ( n197 & ~n6153 ) | ( n197 & n14529 ) | ( ~n6153 & n14529 ) ;
  assign n29483 = n29482 ^ n21534 ^ n15086 ;
  assign n29484 = ( n996 & n8865 ) | ( n996 & n11510 ) | ( n8865 & n11510 ) ;
  assign n29485 = ( n16228 & n18559 ) | ( n16228 & ~n29484 ) | ( n18559 & ~n29484 ) ;
  assign n29486 = n29485 ^ n29154 ^ n27430 ;
  assign n29487 = ( n329 & n7768 ) | ( n329 & ~n10783 ) | ( n7768 & ~n10783 ) ;
  assign n29488 = n14268 ^ n8648 ^ n3725 ;
  assign n29489 = n29488 ^ n12533 ^ n4824 ;
  assign n29490 = ( n16270 & n18535 ) | ( n16270 & n18875 ) | ( n18535 & n18875 ) ;
  assign n29491 = ( n9115 & n25592 ) | ( n9115 & ~n27529 ) | ( n25592 & ~n27529 ) ;
  assign n29492 = n29491 ^ n27246 ^ n920 ;
  assign n29493 = ( n5928 & n6408 ) | ( n5928 & n7220 ) | ( n6408 & n7220 ) ;
  assign n29494 = ( n4951 & n27913 ) | ( n4951 & n29493 ) | ( n27913 & n29493 ) ;
  assign n29495 = n12717 ^ n3256 ^ n1414 ;
  assign n29496 = ( n2582 & n12548 ) | ( n2582 & ~n29495 ) | ( n12548 & ~n29495 ) ;
  assign n29497 = ( ~n14954 & n20862 ) | ( ~n14954 & n29496 ) | ( n20862 & n29496 ) ;
  assign n29498 = n13550 ^ n7817 ^ n7368 ;
  assign n29499 = n22171 ^ n16032 ^ n3816 ;
  assign n29500 = n29499 ^ n22028 ^ n2328 ;
  assign n29501 = n20218 ^ n7319 ^ n5798 ;
  assign n29502 = ( ~n16509 & n18457 ) | ( ~n16509 & n29501 ) | ( n18457 & n29501 ) ;
  assign n29503 = n23018 ^ n8486 ^ n280 ;
  assign n29504 = n27297 ^ n21754 ^ n19245 ;
  assign n29505 = n11480 ^ n6388 ^ n6037 ;
  assign n29506 = n29505 ^ n23726 ^ n8589 ;
  assign n29507 = ( n3021 & n7063 ) | ( n3021 & ~n9050 ) | ( n7063 & ~n9050 ) ;
  assign n29508 = n29507 ^ n715 ^ n656 ;
  assign n29509 = ( n18488 & ~n25726 ) | ( n18488 & n29508 ) | ( ~n25726 & n29508 ) ;
  assign n29510 = ( n4835 & n6576 ) | ( n4835 & ~n7719 ) | ( n6576 & ~n7719 ) ;
  assign n29511 = ( ~n9556 & n27753 ) | ( ~n9556 & n29510 ) | ( n27753 & n29510 ) ;
  assign n29512 = ( n7596 & n9335 ) | ( n7596 & ~n11846 ) | ( n9335 & ~n11846 ) ;
  assign n29513 = n11710 ^ n9232 ^ n1196 ;
  assign n29514 = n29513 ^ n8634 ^ n1103 ;
  assign n29515 = ( n7506 & ~n15308 ) | ( n7506 & n29514 ) | ( ~n15308 & n29514 ) ;
  assign n29516 = n11743 ^ n10891 ^ n6500 ;
  assign n29517 = n29516 ^ n6920 ^ n4412 ;
  assign n29518 = n25772 ^ n13663 ^ n2440 ;
  assign n29519 = ( ~n511 & n23370 ) | ( ~n511 & n29518 ) | ( n23370 & n29518 ) ;
  assign n29521 = ( n1014 & n5056 ) | ( n1014 & n9104 ) | ( n5056 & n9104 ) ;
  assign n29520 = ( ~n4114 & n9510 ) | ( ~n4114 & n20760 ) | ( n9510 & n20760 ) ;
  assign n29522 = n29521 ^ n29520 ^ n17939 ;
  assign n29523 = ( n12112 & n20439 ) | ( n12112 & ~n25262 ) | ( n20439 & ~n25262 ) ;
  assign n29524 = ( n1988 & n22312 ) | ( n1988 & n22455 ) | ( n22312 & n22455 ) ;
  assign n29525 = n29524 ^ n27407 ^ n705 ;
  assign n29526 = n18732 ^ n14498 ^ n2491 ;
  assign n29527 = ( ~n16888 & n23884 ) | ( ~n16888 & n29526 ) | ( n23884 & n29526 ) ;
  assign n29528 = n17780 ^ n10260 ^ n9107 ;
  assign n29529 = n18490 ^ n7960 ^ n4618 ;
  assign n29530 = n27733 ^ n20008 ^ n6325 ;
  assign n29531 = ( n11326 & n22510 ) | ( n11326 & ~n29530 ) | ( n22510 & ~n29530 ) ;
  assign n29532 = ( n835 & n4151 ) | ( n835 & ~n7967 ) | ( n4151 & ~n7967 ) ;
  assign n29533 = n29532 ^ n19468 ^ n3895 ;
  assign n29534 = ( n11658 & n19740 ) | ( n11658 & ~n29533 ) | ( n19740 & ~n29533 ) ;
  assign n29535 = ( n2385 & n12814 ) | ( n2385 & n29534 ) | ( n12814 & n29534 ) ;
  assign n29536 = ( n7335 & ~n16805 ) | ( n7335 & n19601 ) | ( ~n16805 & n19601 ) ;
  assign n29537 = n29536 ^ n13812 ^ n2287 ;
  assign n29538 = n4991 ^ n1375 ^ n1371 ;
  assign n29539 = ( ~n6666 & n10241 ) | ( ~n6666 & n10489 ) | ( n10241 & n10489 ) ;
  assign n29540 = n29539 ^ n9179 ^ n6725 ;
  assign n29541 = ( ~n4741 & n29538 ) | ( ~n4741 & n29540 ) | ( n29538 & n29540 ) ;
  assign n29542 = n26363 ^ n17537 ^ n493 ;
  assign n29543 = n29542 ^ n27994 ^ n2475 ;
  assign n29544 = n29543 ^ n13180 ^ n5870 ;
  assign n29546 = ( n21843 & n23783 ) | ( n21843 & n24509 ) | ( n23783 & n24509 ) ;
  assign n29545 = ( n3881 & n4107 ) | ( n3881 & n19698 ) | ( n4107 & n19698 ) ;
  assign n29547 = n29546 ^ n29545 ^ n26962 ;
  assign n29548 = ( n6723 & ~n20426 ) | ( n6723 & n21590 ) | ( ~n20426 & n21590 ) ;
  assign n29549 = ( n6445 & n8302 ) | ( n6445 & ~n29548 ) | ( n8302 & ~n29548 ) ;
  assign n29550 = n29549 ^ n28979 ^ n13067 ;
  assign n29551 = n10684 ^ n8326 ^ n3417 ;
  assign n29552 = n21717 ^ n8566 ^ n1654 ;
  assign n29553 = ( n373 & n2704 ) | ( n373 & n6402 ) | ( n2704 & n6402 ) ;
  assign n29554 = n29553 ^ n19129 ^ n18679 ;
  assign n29555 = n29554 ^ n2529 ^ n2314 ;
  assign n29556 = n26453 ^ n18920 ^ n15057 ;
  assign n29557 = n29556 ^ n9872 ^ n3081 ;
  assign n29560 = ( n1287 & n4460 ) | ( n1287 & n9064 ) | ( n4460 & n9064 ) ;
  assign n29559 = ( n8782 & n15696 ) | ( n8782 & ~n18893 ) | ( n15696 & ~n18893 ) ;
  assign n29561 = n29560 ^ n29559 ^ n18252 ;
  assign n29558 = n25042 ^ n8917 ^ n3665 ;
  assign n29562 = n29561 ^ n29558 ^ n7823 ;
  assign n29563 = n21801 ^ n6636 ^ n3100 ;
  assign n29564 = ( n1973 & ~n7469 ) | ( n1973 & n14131 ) | ( ~n7469 & n14131 ) ;
  assign n29565 = ( ~n5181 & n19753 ) | ( ~n5181 & n29564 ) | ( n19753 & n29564 ) ;
  assign n29566 = n21029 ^ n9995 ^ n9847 ;
  assign n29567 = ( n23625 & ~n26375 ) | ( n23625 & n29566 ) | ( ~n26375 & n29566 ) ;
  assign n29568 = ( n1724 & n3303 ) | ( n1724 & n11308 ) | ( n3303 & n11308 ) ;
  assign n29569 = n29568 ^ n26781 ^ n14420 ;
  assign n29570 = n21686 ^ n18565 ^ n13823 ;
  assign n29571 = n18447 ^ n9340 ^ n7206 ;
  assign n29572 = n22171 ^ n10281 ^ n8714 ;
  assign n29573 = ( n16601 & n23415 ) | ( n16601 & n29572 ) | ( n23415 & n29572 ) ;
  assign n29574 = n17251 ^ n14111 ^ n3005 ;
  assign n29575 = ( n10011 & n17770 ) | ( n10011 & n29574 ) | ( n17770 & n29574 ) ;
  assign n29578 = n14482 ^ n9102 ^ n654 ;
  assign n29577 = n25146 ^ n24012 ^ n12367 ;
  assign n29576 = n17660 ^ n12823 ^ n11731 ;
  assign n29579 = n29578 ^ n29577 ^ n29576 ;
  assign n29580 = n29579 ^ n18197 ^ n12165 ;
  assign n29581 = ( ~n1304 & n6066 ) | ( ~n1304 & n11157 ) | ( n6066 & n11157 ) ;
  assign n29582 = ( n210 & ~n26238 ) | ( n210 & n29581 ) | ( ~n26238 & n29581 ) ;
  assign n29583 = n29582 ^ n6433 ^ n3192 ;
  assign n29584 = n25403 ^ n9780 ^ n6621 ;
  assign n29585 = n29584 ^ n29464 ^ n7308 ;
  assign n29586 = ( n1979 & ~n4635 ) | ( n1979 & n18376 ) | ( ~n4635 & n18376 ) ;
  assign n29587 = n29586 ^ n24769 ^ n3485 ;
  assign n29589 = n10579 ^ n1326 ^ n896 ;
  assign n29588 = ( ~n1304 & n1471 ) | ( ~n1304 & n3621 ) | ( n1471 & n3621 ) ;
  assign n29590 = n29589 ^ n29588 ^ n26171 ;
  assign n29591 = ( n2424 & ~n2548 ) | ( n2424 & n12008 ) | ( ~n2548 & n12008 ) ;
  assign n29592 = ( n4935 & n13274 ) | ( n4935 & n29591 ) | ( n13274 & n29591 ) ;
  assign n29593 = ( ~n634 & n12869 ) | ( ~n634 & n13229 ) | ( n12869 & n13229 ) ;
  assign n29594 = n29593 ^ n16048 ^ n4249 ;
  assign n29595 = ( n16620 & n29592 ) | ( n16620 & n29594 ) | ( n29592 & n29594 ) ;
  assign n29596 = ( n11389 & n19448 ) | ( n11389 & n19672 ) | ( n19448 & n19672 ) ;
  assign n29597 = ( n18836 & ~n28481 ) | ( n18836 & n29596 ) | ( ~n28481 & n29596 ) ;
  assign n29598 = ( ~n8320 & n22269 ) | ( ~n8320 & n28086 ) | ( n22269 & n28086 ) ;
  assign n29599 = n14666 ^ n11179 ^ n6332 ;
  assign n29600 = ( ~n7518 & n8391 ) | ( ~n7518 & n29599 ) | ( n8391 & n29599 ) ;
  assign n29601 = n29600 ^ n8153 ^ n6186 ;
  assign n29602 = ( n7781 & n10692 ) | ( n7781 & n14660 ) | ( n10692 & n14660 ) ;
  assign n29603 = n29602 ^ n24714 ^ n1924 ;
  assign n29604 = n16014 ^ n12185 ^ n7225 ;
  assign n29605 = n26381 ^ n18937 ^ n14330 ;
  assign n29609 = ( n2694 & n15303 ) | ( n2694 & n23978 ) | ( n15303 & n23978 ) ;
  assign n29606 = ( n7319 & n10989 ) | ( n7319 & n15477 ) | ( n10989 & n15477 ) ;
  assign n29607 = n29606 ^ n23153 ^ n2328 ;
  assign n29608 = ( ~n2743 & n14103 ) | ( ~n2743 & n29607 ) | ( n14103 & n29607 ) ;
  assign n29610 = n29609 ^ n29608 ^ n15921 ;
  assign n29611 = ( n3429 & n7538 ) | ( n3429 & ~n29610 ) | ( n7538 & ~n29610 ) ;
  assign n29612 = n23120 ^ n19493 ^ n5457 ;
  assign n29613 = ( ~n14923 & n17387 ) | ( ~n14923 & n29612 ) | ( n17387 & n29612 ) ;
  assign n29614 = n29613 ^ n16555 ^ n1318 ;
  assign n29615 = ( ~n1100 & n13740 ) | ( ~n1100 & n23381 ) | ( n13740 & n23381 ) ;
  assign n29616 = n5571 ^ n3413 ^ n2203 ;
  assign n29617 = ( x29 & n29329 ) | ( x29 & ~n29616 ) | ( n29329 & ~n29616 ) ;
  assign n29618 = n29617 ^ n11588 ^ n10367 ;
  assign n29619 = n17083 ^ n8780 ^ n4361 ;
  assign n29620 = n23167 ^ n5732 ^ n2502 ;
  assign n29621 = n29620 ^ n28593 ^ n20908 ;
  assign n29622 = ( n8246 & n8396 ) | ( n8246 & ~n15098 ) | ( n8396 & ~n15098 ) ;
  assign n29623 = ( n5861 & n20620 ) | ( n5861 & n29622 ) | ( n20620 & n29622 ) ;
  assign n29624 = n24012 ^ n10548 ^ n7964 ;
  assign n29625 = ( ~n2694 & n8617 ) | ( ~n2694 & n14780 ) | ( n8617 & n14780 ) ;
  assign n29626 = ( ~n11765 & n16480 ) | ( ~n11765 & n19805 ) | ( n16480 & n19805 ) ;
  assign n29627 = ( n14373 & ~n16650 ) | ( n14373 & n29626 ) | ( ~n16650 & n29626 ) ;
  assign n29628 = n25536 ^ n7433 ^ n680 ;
  assign n29629 = ( n736 & ~n14816 ) | ( n736 & n20061 ) | ( ~n14816 & n20061 ) ;
  assign n29631 = ( n1796 & n2725 ) | ( n1796 & n4658 ) | ( n2725 & n4658 ) ;
  assign n29630 = n15012 ^ n2554 ^ n2149 ;
  assign n29632 = n29631 ^ n29630 ^ n13548 ;
  assign n29633 = ( ~n8739 & n29629 ) | ( ~n8739 & n29632 ) | ( n29629 & n29632 ) ;
  assign n29634 = ( ~n2714 & n11975 ) | ( ~n2714 & n14752 ) | ( n11975 & n14752 ) ;
  assign n29635 = n6540 ^ n4853 ^ n1909 ;
  assign n29636 = n29635 ^ n20746 ^ n19539 ;
  assign n29637 = ( n12530 & n13757 ) | ( n12530 & n15550 ) | ( n13757 & n15550 ) ;
  assign n29638 = ( n6414 & n13606 ) | ( n6414 & ~n29637 ) | ( n13606 & ~n29637 ) ;
  assign n29639 = ( n9155 & n17166 ) | ( n9155 & ~n18215 ) | ( n17166 & ~n18215 ) ;
  assign n29640 = ( n267 & n5030 ) | ( n267 & ~n7074 ) | ( n5030 & ~n7074 ) ;
  assign n29641 = ( n1889 & n7614 ) | ( n1889 & n29640 ) | ( n7614 & n29640 ) ;
  assign n29642 = n29641 ^ n24949 ^ n17591 ;
  assign n29643 = n16513 ^ n15106 ^ n6387 ;
  assign n29644 = n29643 ^ n28037 ^ n23421 ;
  assign n29645 = n24903 ^ n18396 ^ n7174 ;
  assign n29646 = ( x66 & ~n1751 ) | ( x66 & n3911 ) | ( ~n1751 & n3911 ) ;
  assign n29647 = ( n8722 & ~n10704 ) | ( n8722 & n29646 ) | ( ~n10704 & n29646 ) ;
  assign n29648 = ( n6741 & n10445 ) | ( n6741 & ~n29647 ) | ( n10445 & ~n29647 ) ;
  assign n29649 = ( n480 & ~n6501 ) | ( n480 & n29648 ) | ( ~n6501 & n29648 ) ;
  assign n29650 = ( n13265 & n13323 ) | ( n13265 & ~n16591 ) | ( n13323 & ~n16591 ) ;
  assign n29651 = n16330 ^ n15266 ^ n10365 ;
  assign n29652 = n14687 ^ n9358 ^ n3320 ;
  assign n29653 = ( n978 & n5052 ) | ( n978 & n5869 ) | ( n5052 & n5869 ) ;
  assign n29654 = n12879 ^ n5731 ^ n1216 ;
  assign n29655 = ( n16938 & n29653 ) | ( n16938 & ~n29654 ) | ( n29653 & ~n29654 ) ;
  assign n29656 = ( ~n3172 & n6079 ) | ( ~n3172 & n29655 ) | ( n6079 & n29655 ) ;
  assign n29657 = n28234 ^ n18416 ^ n8664 ;
  assign n29658 = n26064 ^ n4732 ^ n3432 ;
  assign n29659 = n21396 ^ n18565 ^ n4461 ;
  assign n29660 = ( n5016 & n5557 ) | ( n5016 & ~n9573 ) | ( n5557 & ~n9573 ) ;
  assign n29661 = n17785 ^ n5074 ^ n4615 ;
  assign n29664 = n26822 ^ n18024 ^ n12331 ;
  assign n29665 = ( n8217 & ~n10696 ) | ( n8217 & n12013 ) | ( ~n10696 & n12013 ) ;
  assign n29666 = ( ~n12184 & n29664 ) | ( ~n12184 & n29665 ) | ( n29664 & n29665 ) ;
  assign n29662 = ( n4133 & ~n6561 ) | ( n4133 & n11414 ) | ( ~n6561 & n11414 ) ;
  assign n29663 = ( n17866 & ~n24597 ) | ( n17866 & n29662 ) | ( ~n24597 & n29662 ) ;
  assign n29667 = n29666 ^ n29663 ^ n17432 ;
  assign n29668 = n13091 ^ n5862 ^ n2225 ;
  assign n29669 = n20886 ^ n5419 ^ x101 ;
  assign n29670 = n22732 ^ n13139 ^ n12810 ;
  assign n29671 = ( n12903 & n19467 ) | ( n12903 & ~n29670 ) | ( n19467 & ~n29670 ) ;
  assign n29672 = ( n9172 & n23957 ) | ( n9172 & n29671 ) | ( n23957 & n29671 ) ;
  assign n29673 = ( ~x28 & n5330 ) | ( ~x28 & n12281 ) | ( n5330 & n12281 ) ;
  assign n29674 = n1764 ^ n447 ^ x39 ;
  assign n29675 = ( ~n21148 & n29484 ) | ( ~n21148 & n29674 ) | ( n29484 & n29674 ) ;
  assign n29679 = n13445 ^ n7172 ^ n2926 ;
  assign n29676 = n20328 ^ n16577 ^ n11650 ;
  assign n29677 = ( n5935 & n18498 ) | ( n5935 & n23323 ) | ( n18498 & n23323 ) ;
  assign n29678 = ( n6399 & n29676 ) | ( n6399 & ~n29677 ) | ( n29676 & ~n29677 ) ;
  assign n29680 = n29679 ^ n29678 ^ n19041 ;
  assign n29681 = n11482 ^ n2418 ^ n2030 ;
  assign n29682 = ( n13537 & n23557 ) | ( n13537 & ~n24613 ) | ( n23557 & ~n24613 ) ;
  assign n29683 = n26950 ^ n4737 ^ n4266 ;
  assign n29684 = ( n10128 & ~n15416 ) | ( n10128 & n29683 ) | ( ~n15416 & n29683 ) ;
  assign n29685 = ( n2440 & ~n5484 ) | ( n2440 & n29684 ) | ( ~n5484 & n29684 ) ;
  assign n29686 = ( n222 & n3596 ) | ( n222 & n25888 ) | ( n3596 & n25888 ) ;
  assign n29687 = n22968 ^ n2742 ^ n910 ;
  assign n29688 = n29687 ^ n26952 ^ n25045 ;
  assign n29689 = n26995 ^ n22599 ^ n7307 ;
  assign n29690 = ( ~n10151 & n11937 ) | ( ~n10151 & n27566 ) | ( n11937 & n27566 ) ;
  assign n29691 = ( n1667 & ~n19825 ) | ( n1667 & n29690 ) | ( ~n19825 & n29690 ) ;
  assign n29692 = n29691 ^ n22299 ^ n8318 ;
  assign n29693 = n7449 ^ n661 ^ n352 ;
  assign n29694 = n29693 ^ n18196 ^ n16669 ;
  assign n29695 = ( n13501 & n22926 ) | ( n13501 & ~n29694 ) | ( n22926 & ~n29694 ) ;
  assign n29696 = ( n13862 & ~n29692 ) | ( n13862 & n29695 ) | ( ~n29692 & n29695 ) ;
  assign n29697 = n7375 ^ n2448 ^ n932 ;
  assign n29698 = ( n2943 & n7280 ) | ( n2943 & n23949 ) | ( n7280 & n23949 ) ;
  assign n29699 = ( ~n20338 & n29697 ) | ( ~n20338 & n29698 ) | ( n29697 & n29698 ) ;
  assign n29700 = n9094 ^ n4652 ^ n3363 ;
  assign n29701 = ( n865 & ~n6664 ) | ( n865 & n29700 ) | ( ~n6664 & n29700 ) ;
  assign n29702 = ( n11447 & n29699 ) | ( n11447 & n29701 ) | ( n29699 & n29701 ) ;
  assign n29703 = n29702 ^ n16705 ^ n11519 ;
  assign n29704 = ( x34 & ~n6871 ) | ( x34 & n22154 ) | ( ~n6871 & n22154 ) ;
  assign n29705 = n29704 ^ n28104 ^ n2582 ;
  assign n29706 = n29705 ^ n20872 ^ n15387 ;
  assign n29707 = ( ~n453 & n487 ) | ( ~n453 & n1458 ) | ( n487 & n1458 ) ;
  assign n29708 = n29707 ^ n18087 ^ n15206 ;
  assign n29709 = ( ~n12300 & n27198 ) | ( ~n12300 & n29708 ) | ( n27198 & n29708 ) ;
  assign n29710 = n26899 ^ n5742 ^ n5090 ;
  assign n29711 = n12882 ^ n3351 ^ n1720 ;
  assign n29712 = n19863 ^ n16880 ^ n9905 ;
  assign n29713 = ( n2091 & n5514 ) | ( n2091 & ~n25158 ) | ( n5514 & ~n25158 ) ;
  assign n29714 = n11621 ^ n4039 ^ x127 ;
  assign n29715 = n29714 ^ n28230 ^ n1506 ;
  assign n29716 = n29715 ^ n17839 ^ n4635 ;
  assign n29717 = ( n1664 & n10557 ) | ( n1664 & ~n20191 ) | ( n10557 & ~n20191 ) ;
  assign n29720 = n19608 ^ n8225 ^ n5548 ;
  assign n29721 = n29720 ^ n14821 ^ n13801 ;
  assign n29719 = ( n10462 & ~n17004 ) | ( n10462 & n21336 ) | ( ~n17004 & n21336 ) ;
  assign n29722 = n29721 ^ n29719 ^ n13383 ;
  assign n29723 = ( n11447 & n17327 ) | ( n11447 & ~n29722 ) | ( n17327 & ~n29722 ) ;
  assign n29718 = ( ~n10735 & n17552 ) | ( ~n10735 & n20524 ) | ( n17552 & n20524 ) ;
  assign n29724 = n29723 ^ n29718 ^ n28625 ;
  assign n29725 = n29724 ^ n12771 ^ n7856 ;
  assign n29726 = ( n3655 & n6874 ) | ( n3655 & n29725 ) | ( n6874 & n29725 ) ;
  assign n29727 = ( ~n632 & n987 ) | ( ~n632 & n23884 ) | ( n987 & n23884 ) ;
  assign n29728 = ( n3264 & n6193 ) | ( n3264 & ~n15957 ) | ( n6193 & ~n15957 ) ;
  assign n29729 = n21283 ^ n11552 ^ n434 ;
  assign n29730 = n16759 ^ n7990 ^ n667 ;
  assign n29731 = ( n9133 & n18937 ) | ( n9133 & ~n29730 ) | ( n18937 & ~n29730 ) ;
  assign n29733 = ( n1223 & n8773 ) | ( n1223 & n21892 ) | ( n8773 & n21892 ) ;
  assign n29732 = n24458 ^ n15513 ^ n12494 ;
  assign n29734 = n29733 ^ n29732 ^ n19355 ;
  assign n29735 = ( ~n7987 & n14543 ) | ( ~n7987 & n14547 ) | ( n14543 & n14547 ) ;
  assign n29736 = ( n2942 & ~n21728 ) | ( n2942 & n29735 ) | ( ~n21728 & n29735 ) ;
  assign n29737 = n29736 ^ n17133 ^ n2260 ;
  assign n29738 = n27505 ^ n19570 ^ n13596 ;
  assign n29739 = n13975 ^ n13037 ^ n5754 ;
  assign n29740 = ( n9754 & n14024 ) | ( n9754 & ~n16979 ) | ( n14024 & ~n16979 ) ;
  assign n29741 = n26866 ^ n26212 ^ n6296 ;
  assign n29742 = ( n5889 & n9579 ) | ( n5889 & ~n29741 ) | ( n9579 & ~n29741 ) ;
  assign n29743 = ( n6472 & ~n8730 ) | ( n6472 & n9516 ) | ( ~n8730 & n9516 ) ;
  assign n29744 = n29684 ^ n15435 ^ n6914 ;
  assign n29745 = ( n29255 & n29743 ) | ( n29255 & ~n29744 ) | ( n29743 & ~n29744 ) ;
  assign n29746 = n9186 ^ n5862 ^ n5849 ;
  assign n29747 = n26261 ^ n19975 ^ n4009 ;
  assign n29748 = n25780 ^ n12345 ^ n7453 ;
  assign n29749 = n29748 ^ n17700 ^ n10562 ;
  assign n29750 = ( n9115 & n21845 ) | ( n9115 & ~n23468 ) | ( n21845 & ~n23468 ) ;
  assign n29751 = n29750 ^ n14163 ^ n4369 ;
  assign n29752 = ( ~n5758 & n7717 ) | ( ~n5758 & n13092 ) | ( n7717 & n13092 ) ;
  assign n29753 = ( n9330 & ~n17494 ) | ( n9330 & n25066 ) | ( ~n17494 & n25066 ) ;
  assign n29754 = n20705 ^ n20539 ^ n9212 ;
  assign n29755 = n26134 ^ n22030 ^ n1235 ;
  assign n29756 = ( ~n3335 & n15174 ) | ( ~n3335 & n29755 ) | ( n15174 & n29755 ) ;
  assign n29757 = ( n14644 & ~n24605 ) | ( n14644 & n29756 ) | ( ~n24605 & n29756 ) ;
  assign n29758 = n12766 ^ n7711 ^ n6409 ;
  assign n29759 = n12732 ^ n3028 ^ n2295 ;
  assign n29760 = n27713 ^ n5701 ^ n2467 ;
  assign n29761 = n7083 ^ n3123 ^ n2037 ;
  assign n29762 = ( n9406 & n17901 ) | ( n9406 & ~n29761 ) | ( n17901 & ~n29761 ) ;
  assign n29763 = ( ~n4237 & n6416 ) | ( ~n4237 & n14018 ) | ( n6416 & n14018 ) ;
  assign n29766 = n20255 ^ n12744 ^ n7673 ;
  assign n29765 = ( n8328 & ~n11780 ) | ( n8328 & n22200 ) | ( ~n11780 & n22200 ) ;
  assign n29764 = n6548 ^ n3341 ^ n796 ;
  assign n29767 = n29766 ^ n29765 ^ n29764 ;
  assign n29768 = ( n12909 & ~n13893 ) | ( n12909 & n24899 ) | ( ~n13893 & n24899 ) ;
  assign n29769 = n29768 ^ n4821 ^ n3019 ;
  assign n29770 = n13591 ^ n8914 ^ n5080 ;
  assign n29771 = ( n9819 & ~n29769 ) | ( n9819 & n29770 ) | ( ~n29769 & n29770 ) ;
  assign n29772 = n29771 ^ n14739 ^ n2092 ;
  assign n29773 = ( n13961 & ~n21745 ) | ( n13961 & n29772 ) | ( ~n21745 & n29772 ) ;
  assign n29774 = n28169 ^ n12874 ^ n5451 ;
  assign n29775 = n29774 ^ n15473 ^ n2118 ;
  assign n29776 = n21361 ^ n8335 ^ n1637 ;
  assign n29777 = ( ~n10330 & n13439 ) | ( ~n10330 & n25981 ) | ( n13439 & n25981 ) ;
  assign n29778 = ( n27130 & ~n29776 ) | ( n27130 & n29777 ) | ( ~n29776 & n29777 ) ;
  assign n29779 = ( ~n8836 & n11129 ) | ( ~n8836 & n12548 ) | ( n11129 & n12548 ) ;
  assign n29780 = n14001 ^ n9000 ^ n5587 ;
  assign n29781 = n29780 ^ n19457 ^ n13241 ;
  assign n29784 = n13454 ^ n12131 ^ n8018 ;
  assign n29782 = ( n10072 & ~n13512 ) | ( n10072 & n20573 ) | ( ~n13512 & n20573 ) ;
  assign n29783 = n29782 ^ n5783 ^ n1140 ;
  assign n29785 = n29784 ^ n29783 ^ n12498 ;
  assign n29786 = n14507 ^ n5102 ^ n2080 ;
  assign n29787 = n29786 ^ n25577 ^ n21488 ;
  assign n29788 = ( n3906 & ~n14992 ) | ( n3906 & n20659 ) | ( ~n14992 & n20659 ) ;
  assign n29789 = n24706 ^ n4612 ^ n1366 ;
  assign n29790 = ( ~n27907 & n29788 ) | ( ~n27907 & n29789 ) | ( n29788 & n29789 ) ;
  assign n29793 = ( n3723 & ~n7798 ) | ( n3723 & n13998 ) | ( ~n7798 & n13998 ) ;
  assign n29792 = ( ~n17216 & n19807 ) | ( ~n17216 & n25039 ) | ( n19807 & n25039 ) ;
  assign n29794 = n29793 ^ n29792 ^ n22488 ;
  assign n29791 = ( n9443 & n12698 ) | ( n9443 & n21739 ) | ( n12698 & n21739 ) ;
  assign n29795 = n29794 ^ n29791 ^ n13729 ;
  assign n29796 = ( n9112 & ~n9127 ) | ( n9112 & n12799 ) | ( ~n9127 & n12799 ) ;
  assign n29797 = ( n818 & n1064 ) | ( n818 & n3208 ) | ( n1064 & n3208 ) ;
  assign n29798 = n29797 ^ n17855 ^ n4221 ;
  assign n29799 = ( n3505 & n16613 ) | ( n3505 & n23907 ) | ( n16613 & n23907 ) ;
  assign n29800 = n29799 ^ n24388 ^ n20426 ;
  assign n29801 = n29800 ^ n19087 ^ n2179 ;
  assign n29802 = ( n11916 & n21688 ) | ( n11916 & ~n24946 ) | ( n21688 & ~n24946 ) ;
  assign n29803 = ( ~n4741 & n5682 ) | ( ~n4741 & n14349 ) | ( n5682 & n14349 ) ;
  assign n29804 = ( ~n5155 & n20391 ) | ( ~n5155 & n29803 ) | ( n20391 & n29803 ) ;
  assign n29805 = n28862 ^ n22710 ^ n10159 ;
  assign n29806 = n18524 ^ n11523 ^ n3614 ;
  assign n29807 = ( n15234 & n22939 ) | ( n15234 & n29806 ) | ( n22939 & n29806 ) ;
  assign n29808 = n19695 ^ n15015 ^ n9955 ;
  assign n29809 = n17098 ^ n1066 ^ n974 ;
  assign n29810 = ( n14718 & n29808 ) | ( n14718 & ~n29809 ) | ( n29808 & ~n29809 ) ;
  assign n29811 = ( n2012 & n2955 ) | ( n2012 & n23940 ) | ( n2955 & n23940 ) ;
  assign n29812 = ( ~n2692 & n26641 ) | ( ~n2692 & n29811 ) | ( n26641 & n29811 ) ;
  assign n29815 = ( n10663 & ~n16873 ) | ( n10663 & n22813 ) | ( ~n16873 & n22813 ) ;
  assign n29816 = ( ~n1607 & n15396 ) | ( ~n1607 & n29815 ) | ( n15396 & n29815 ) ;
  assign n29813 = ( n1036 & n8604 ) | ( n1036 & ~n16024 ) | ( n8604 & ~n16024 ) ;
  assign n29814 = n29813 ^ n19531 ^ n5162 ;
  assign n29817 = n29816 ^ n29814 ^ n19495 ;
  assign n29818 = ( n17533 & ~n18270 ) | ( n17533 & n18518 ) | ( ~n18270 & n18518 ) ;
  assign n29819 = ( n2732 & ~n3875 ) | ( n2732 & n29818 ) | ( ~n3875 & n29818 ) ;
  assign n29820 = n29819 ^ n12937 ^ n12580 ;
  assign n29822 = ( n3543 & n29238 ) | ( n3543 & n29578 ) | ( n29238 & n29578 ) ;
  assign n29823 = n29822 ^ n22111 ^ n12704 ;
  assign n29821 = n20185 ^ n18834 ^ n11603 ;
  assign n29824 = n29823 ^ n29821 ^ n2195 ;
  assign n29825 = n10359 ^ n2660 ^ n154 ;
  assign n29826 = n29825 ^ n27090 ^ n9490 ;
  assign n29827 = ( ~n4271 & n19882 ) | ( ~n4271 & n26846 ) | ( n19882 & n26846 ) ;
  assign n29828 = ( n3316 & n7217 ) | ( n3316 & n25580 ) | ( n7217 & n25580 ) ;
  assign n29829 = n27749 ^ n20309 ^ n13645 ;
  assign n29830 = ( ~x65 & n8403 ) | ( ~x65 & n15034 ) | ( n8403 & n15034 ) ;
  assign n29831 = n15714 ^ n7391 ^ n978 ;
  assign n29832 = ( n3149 & ~n3614 ) | ( n3149 & n3802 ) | ( ~n3614 & n3802 ) ;
  assign n29833 = ( n9371 & ~n29831 ) | ( n9371 & n29832 ) | ( ~n29831 & n29832 ) ;
  assign n29834 = ( n12944 & ~n17461 ) | ( n12944 & n24723 ) | ( ~n17461 & n24723 ) ;
  assign n29835 = ( n26077 & ~n29833 ) | ( n26077 & n29834 ) | ( ~n29833 & n29834 ) ;
  assign n29836 = n12190 ^ n729 ^ n506 ;
  assign n29837 = n29836 ^ n25622 ^ n5113 ;
  assign n29839 = n11563 ^ n8127 ^ n4025 ;
  assign n29838 = ( ~n2949 & n3597 ) | ( ~n2949 & n11428 ) | ( n3597 & n11428 ) ;
  assign n29840 = n29839 ^ n29838 ^ n19048 ;
  assign n29841 = n28836 ^ n26212 ^ n15657 ;
  assign n29842 = n29841 ^ n2920 ^ n2096 ;
  assign n29843 = ( x1 & n828 ) | ( x1 & n28670 ) | ( n828 & n28670 ) ;
  assign n29844 = n22707 ^ n11183 ^ n4324 ;
  assign n29845 = ( n796 & n4629 ) | ( n796 & n11038 ) | ( n4629 & n11038 ) ;
  assign n29846 = ( n2123 & n24770 ) | ( n2123 & n29845 ) | ( n24770 & n29845 ) ;
  assign n29847 = n25342 ^ n15687 ^ n4123 ;
  assign n29848 = n20024 ^ n15873 ^ n8101 ;
  assign n29849 = ( n28539 & n29847 ) | ( n28539 & ~n29848 ) | ( n29847 & ~n29848 ) ;
  assign n29850 = ( ~n7107 & n7678 ) | ( ~n7107 & n21901 ) | ( n7678 & n21901 ) ;
  assign n29851 = n29850 ^ n27756 ^ n15678 ;
  assign n29852 = n20334 ^ n11546 ^ n1150 ;
  assign n29853 = n29852 ^ n23731 ^ n16077 ;
  assign n29854 = ( ~n2996 & n14966 ) | ( ~n2996 & n29066 ) | ( n14966 & n29066 ) ;
  assign n29855 = ( n2344 & n18721 ) | ( n2344 & n29854 ) | ( n18721 & n29854 ) ;
  assign n29856 = n22306 ^ n10353 ^ n2279 ;
  assign n29857 = ( n765 & n2423 ) | ( n765 & ~n18999 ) | ( n2423 & ~n18999 ) ;
  assign n29858 = ( n12155 & n19299 ) | ( n12155 & n29857 ) | ( n19299 & n29857 ) ;
  assign n29859 = ( n5260 & n21207 ) | ( n5260 & ~n26849 ) | ( n21207 & ~n26849 ) ;
  assign n29860 = n26380 ^ n14617 ^ n2092 ;
  assign n29861 = n25589 ^ n19385 ^ n5296 ;
  assign n29862 = n29861 ^ n13611 ^ n7813 ;
  assign n29864 = ( ~n3203 & n14436 ) | ( ~n3203 & n20460 ) | ( n14436 & n20460 ) ;
  assign n29865 = ( n5836 & n7219 ) | ( n5836 & ~n29864 ) | ( n7219 & ~n29864 ) ;
  assign n29863 = ( n1835 & n2911 ) | ( n1835 & ~n22101 ) | ( n2911 & ~n22101 ) ;
  assign n29866 = n29865 ^ n29863 ^ n10269 ;
  assign n29867 = ( n940 & ~n29862 ) | ( n940 & n29866 ) | ( ~n29862 & n29866 ) ;
  assign n29868 = ( ~n2728 & n5873 ) | ( ~n2728 & n6468 ) | ( n5873 & n6468 ) ;
  assign n29869 = ( n2675 & n9380 ) | ( n2675 & n29868 ) | ( n9380 & n29868 ) ;
  assign n29870 = n29869 ^ n10298 ^ n2137 ;
  assign n29871 = ( n1445 & ~n1497 ) | ( n1445 & n29870 ) | ( ~n1497 & n29870 ) ;
  assign n29872 = n20566 ^ n12210 ^ n4272 ;
  assign n29873 = ( n25111 & ~n29871 ) | ( n25111 & n29872 ) | ( ~n29871 & n29872 ) ;
  assign n29874 = n18999 ^ n15571 ^ n9990 ;
  assign n29875 = ( n20709 & n29854 ) | ( n20709 & ~n29874 ) | ( n29854 & ~n29874 ) ;
  assign n29876 = ( n3115 & n3374 ) | ( n3115 & n20304 ) | ( n3374 & n20304 ) ;
  assign n29877 = ( ~n3919 & n20609 ) | ( ~n3919 & n28926 ) | ( n20609 & n28926 ) ;
  assign n29878 = n29877 ^ n12249 ^ n7091 ;
  assign n29879 = ( n324 & n1696 ) | ( n324 & ~n3576 ) | ( n1696 & ~n3576 ) ;
  assign n29880 = n29879 ^ n13494 ^ n6176 ;
  assign n29881 = n29880 ^ n25717 ^ n14688 ;
  assign n29882 = ( n730 & ~n3742 ) | ( n730 & n15800 ) | ( ~n3742 & n15800 ) ;
  assign n29883 = ( n2840 & ~n12096 ) | ( n2840 & n29882 ) | ( ~n12096 & n29882 ) ;
  assign n29884 = ( n7352 & n9484 ) | ( n7352 & n13102 ) | ( n9484 & n13102 ) ;
  assign n29885 = ( ~n1366 & n2028 ) | ( ~n1366 & n8762 ) | ( n2028 & n8762 ) ;
  assign n29886 = n13366 ^ n9057 ^ n1999 ;
  assign n29887 = ( n15071 & ~n29885 ) | ( n15071 & n29886 ) | ( ~n29885 & n29886 ) ;
  assign n29888 = ( ~n28283 & n28686 ) | ( ~n28283 & n29887 ) | ( n28686 & n29887 ) ;
  assign n29889 = n20660 ^ n20454 ^ n19885 ;
  assign n29890 = ( n12062 & n29888 ) | ( n12062 & ~n29889 ) | ( n29888 & ~n29889 ) ;
  assign n29891 = n20099 ^ n13203 ^ n1134 ;
  assign n29892 = ( n499 & ~n11276 ) | ( n499 & n27716 ) | ( ~n11276 & n27716 ) ;
  assign n29893 = ( n7899 & n18970 ) | ( n7899 & ~n20029 ) | ( n18970 & ~n20029 ) ;
  assign n29894 = n6689 ^ n5626 ^ n3198 ;
  assign n29895 = n29894 ^ n13647 ^ n12901 ;
  assign n29896 = ( n787 & ~n3112 ) | ( n787 & n29895 ) | ( ~n3112 & n29895 ) ;
  assign n29897 = n22990 ^ n20154 ^ n19875 ;
  assign n29898 = n29897 ^ n26759 ^ n13779 ;
  assign n29899 = n27005 ^ n7896 ^ n5627 ;
  assign n29901 = n20305 ^ n15147 ^ n2930 ;
  assign n29900 = ( n7362 & n18756 ) | ( n7362 & n28838 ) | ( n18756 & n28838 ) ;
  assign n29902 = n29901 ^ n29900 ^ n16152 ;
  assign n29903 = n26401 ^ n6028 ^ n3019 ;
  assign n29904 = n27709 ^ n12432 ^ n1414 ;
  assign n29905 = ( n15244 & n27165 ) | ( n15244 & n29904 ) | ( n27165 & n29904 ) ;
  assign n29906 = ( n5405 & ~n17759 ) | ( n5405 & n22325 ) | ( ~n17759 & n22325 ) ;
  assign n29907 = n12535 ^ n12083 ^ n8167 ;
  assign n29908 = n29907 ^ n15510 ^ n14581 ;
  assign n29909 = ( n3466 & n6004 ) | ( n3466 & ~n16706 ) | ( n6004 & ~n16706 ) ;
  assign n29910 = ( n5765 & ~n7978 ) | ( n5765 & n21127 ) | ( ~n7978 & n21127 ) ;
  assign n29911 = ( n5801 & ~n28142 ) | ( n5801 & n29910 ) | ( ~n28142 & n29910 ) ;
  assign n29912 = ( n17759 & ~n19599 ) | ( n17759 & n23878 ) | ( ~n19599 & n23878 ) ;
  assign n29913 = ( n19037 & ~n24744 ) | ( n19037 & n25932 ) | ( ~n24744 & n25932 ) ;
  assign n29914 = n29321 ^ n10791 ^ n7469 ;
  assign n29915 = n18416 ^ n9872 ^ n2607 ;
  assign n29916 = n19012 ^ n15390 ^ n4723 ;
  assign n29917 = ( n2323 & n21269 ) | ( n2323 & ~n29916 ) | ( n21269 & ~n29916 ) ;
  assign n29918 = ( ~n10260 & n29915 ) | ( ~n10260 & n29917 ) | ( n29915 & n29917 ) ;
  assign n29919 = ( n17305 & n24482 ) | ( n17305 & ~n29918 ) | ( n24482 & ~n29918 ) ;
  assign n29920 = ( n25258 & ~n28390 ) | ( n25258 & n29720 ) | ( ~n28390 & n29720 ) ;
  assign n29921 = n9839 ^ n1221 ^ x103 ;
  assign n29922 = ( n3110 & n10811 ) | ( n3110 & ~n20699 ) | ( n10811 & ~n20699 ) ;
  assign n29923 = ( n18781 & n26789 ) | ( n18781 & n29922 ) | ( n26789 & n29922 ) ;
  assign n29924 = ( n29920 & n29921 ) | ( n29920 & ~n29923 ) | ( n29921 & ~n29923 ) ;
  assign n29927 = n19364 ^ n12279 ^ n7123 ;
  assign n29925 = n19877 ^ n16738 ^ n11844 ;
  assign n29926 = ( n10851 & n16472 ) | ( n10851 & n29925 ) | ( n16472 & n29925 ) ;
  assign n29928 = n29927 ^ n29926 ^ n8890 ;
  assign n29929 = ( ~n2390 & n14103 ) | ( ~n2390 & n21865 ) | ( n14103 & n21865 ) ;
  assign n29930 = ( n10908 & n14659 ) | ( n10908 & n23843 ) | ( n14659 & n23843 ) ;
  assign n29931 = n14036 ^ n9746 ^ n3331 ;
  assign n29932 = n18356 ^ n16864 ^ n11636 ;
  assign n29933 = n29932 ^ n12965 ^ n8175 ;
  assign n29934 = ( n3298 & n12913 ) | ( n3298 & n28597 ) | ( n12913 & n28597 ) ;
  assign n29935 = n28658 ^ n7889 ^ n3225 ;
  assign n29936 = ( ~n3287 & n4819 ) | ( ~n3287 & n6516 ) | ( n4819 & n6516 ) ;
  assign n29937 = n20729 ^ n13715 ^ n5909 ;
  assign n29938 = ( n5293 & ~n9868 ) | ( n5293 & n29937 ) | ( ~n9868 & n29937 ) ;
  assign n29939 = n16093 ^ n13757 ^ n6540 ;
  assign n29940 = n29939 ^ n13061 ^ n7068 ;
  assign n29941 = n14686 ^ n5055 ^ n2703 ;
  assign n29943 = n8739 ^ n7266 ^ n2410 ;
  assign n29942 = n22270 ^ n20539 ^ n8650 ;
  assign n29944 = n29943 ^ n29942 ^ n19287 ;
  assign n29945 = ( n25066 & ~n29941 ) | ( n25066 & n29944 ) | ( ~n29941 & n29944 ) ;
  assign n29946 = ( n4048 & ~n16323 ) | ( n4048 & n26282 ) | ( ~n16323 & n26282 ) ;
  assign n29947 = n29946 ^ n28946 ^ n19508 ;
  assign n29948 = ( n8522 & n10106 ) | ( n8522 & n21039 ) | ( n10106 & n21039 ) ;
  assign n29949 = n29948 ^ n2504 ^ n1350 ;
  assign n29950 = n22173 ^ n9113 ^ n2302 ;
  assign n29951 = ( n15268 & ~n26929 ) | ( n15268 & n29950 ) | ( ~n26929 & n29950 ) ;
  assign n29952 = n10478 ^ n10312 ^ n6146 ;
  assign n29953 = n29952 ^ n10480 ^ n581 ;
  assign n29954 = n28484 ^ n27662 ^ n18854 ;
  assign n29955 = n17551 ^ n13484 ^ n5032 ;
  assign n29956 = ( n14343 & n28522 ) | ( n14343 & n29955 ) | ( n28522 & n29955 ) ;
  assign n29959 = ( n1195 & n2360 ) | ( n1195 & ~n4636 ) | ( n2360 & ~n4636 ) ;
  assign n29960 = ( n11357 & n12752 ) | ( n11357 & ~n29959 ) | ( n12752 & ~n29959 ) ;
  assign n29957 = n22107 ^ n5596 ^ n2433 ;
  assign n29958 = n29957 ^ n24731 ^ n15348 ;
  assign n29961 = n29960 ^ n29958 ^ n3149 ;
  assign n29962 = n21427 ^ n7818 ^ n213 ;
  assign n29963 = n24159 ^ n11735 ^ n2317 ;
  assign n29964 = ( n3222 & n5066 ) | ( n3222 & ~n29963 ) | ( n5066 & ~n29963 ) ;
  assign n29965 = n7824 ^ n2414 ^ n2007 ;
  assign n29966 = n29965 ^ n27689 ^ n24726 ;
  assign n29967 = n10358 ^ n8189 ^ n1819 ;
  assign n29968 = ( n14880 & n19637 ) | ( n14880 & ~n29967 ) | ( n19637 & ~n29967 ) ;
  assign n29970 = ( n8338 & n17529 ) | ( n8338 & n21018 ) | ( n17529 & n21018 ) ;
  assign n29969 = n20503 ^ n16155 ^ n12927 ;
  assign n29971 = n29970 ^ n29969 ^ n3462 ;
  assign n29972 = ( n5974 & n15322 ) | ( n5974 & ~n24564 ) | ( n15322 & ~n24564 ) ;
  assign n29973 = n27588 ^ n7413 ^ n4873 ;
  assign n29974 = n29973 ^ n26809 ^ n16454 ;
  assign n29975 = ( n1132 & ~n12221 ) | ( n1132 & n17318 ) | ( ~n12221 & n17318 ) ;
  assign n29976 = ( ~n10452 & n16222 ) | ( ~n10452 & n29975 ) | ( n16222 & n29975 ) ;
  assign n29977 = n19029 ^ n15123 ^ n13667 ;
  assign n29978 = ( n5895 & n12683 ) | ( n5895 & ~n24765 ) | ( n12683 & ~n24765 ) ;
  assign n29979 = ( ~n1492 & n3009 ) | ( ~n1492 & n9187 ) | ( n3009 & n9187 ) ;
  assign n29980 = ( ~n21582 & n22297 ) | ( ~n21582 & n29979 ) | ( n22297 & n29979 ) ;
  assign n29981 = n23839 ^ n11919 ^ n3293 ;
  assign n29982 = ( ~n9419 & n15836 ) | ( ~n9419 & n17462 ) | ( n15836 & n17462 ) ;
  assign n29983 = ( ~n3296 & n11472 ) | ( ~n3296 & n17444 ) | ( n11472 & n17444 ) ;
  assign n29984 = ( ~n1436 & n29982 ) | ( ~n1436 & n29983 ) | ( n29982 & n29983 ) ;
  assign n29985 = n10808 ^ n10001 ^ x72 ;
  assign n29986 = n14553 ^ n8381 ^ n7508 ;
  assign n29987 = n29986 ^ n5231 ^ n792 ;
  assign n29988 = n26794 ^ n19321 ^ n8576 ;
  assign n29989 = ( n3802 & n4015 ) | ( n3802 & ~n4734 ) | ( n4015 & ~n4734 ) ;
  assign n29990 = n29989 ^ n14923 ^ n4140 ;
  assign n29991 = n21577 ^ n7418 ^ n2495 ;
  assign n29992 = n29991 ^ n14972 ^ n13376 ;
  assign n29993 = n29992 ^ n6850 ^ n169 ;
  assign n29994 = n23965 ^ n5044 ^ n2104 ;
  assign n29995 = ( n8006 & ~n22656 ) | ( n8006 & n29994 ) | ( ~n22656 & n29994 ) ;
  assign n29996 = n29995 ^ n1347 ^ n262 ;
  assign n29997 = ( ~n13661 & n20871 ) | ( ~n13661 & n29704 ) | ( n20871 & n29704 ) ;
  assign n29998 = n29997 ^ n16736 ^ n5137 ;
  assign n29999 = ( n14584 & ~n19788 ) | ( n14584 & n20885 ) | ( ~n19788 & n20885 ) ;
  assign n30000 = n25312 ^ n9404 ^ n5151 ;
  assign n30001 = n30000 ^ n23227 ^ n6365 ;
  assign n30002 = ( ~n1406 & n13475 ) | ( ~n1406 & n13762 ) | ( n13475 & n13762 ) ;
  assign n30003 = ( n2948 & n4104 ) | ( n2948 & ~n14976 ) | ( n4104 & ~n14976 ) ;
  assign n30004 = ( n5065 & n11205 ) | ( n5065 & ~n30003 ) | ( n11205 & ~n30003 ) ;
  assign n30005 = n20569 ^ n19611 ^ n13692 ;
  assign n30007 = ( n978 & ~n4577 ) | ( n978 & n17632 ) | ( ~n4577 & n17632 ) ;
  assign n30006 = ( n623 & n10049 ) | ( n623 & n14494 ) | ( n10049 & n14494 ) ;
  assign n30008 = n30007 ^ n30006 ^ n14284 ;
  assign n30009 = n14806 ^ n3290 ^ n2512 ;
  assign n30010 = ( ~n1201 & n27639 ) | ( ~n1201 & n30009 ) | ( n27639 & n30009 ) ;
  assign n30011 = n22056 ^ n20498 ^ n17331 ;
  assign n30012 = ( n6795 & n8881 ) | ( n6795 & n22751 ) | ( n8881 & n22751 ) ;
  assign n30013 = ( n4952 & n5229 ) | ( n4952 & n17835 ) | ( n5229 & n17835 ) ;
  assign n30014 = ( ~n1307 & n5950 ) | ( ~n1307 & n16213 ) | ( n5950 & n16213 ) ;
  assign n30015 = ( n1482 & ~n30013 ) | ( n1482 & n30014 ) | ( ~n30013 & n30014 ) ;
  assign n30016 = ( ~n806 & n17771 ) | ( ~n806 & n30015 ) | ( n17771 & n30015 ) ;
  assign n30017 = n18524 ^ n8475 ^ n5174 ;
  assign n30018 = n30017 ^ n23469 ^ n9090 ;
  assign n30019 = ( n8753 & n17538 ) | ( n8753 & n30018 ) | ( n17538 & n30018 ) ;
  assign n30020 = ( n320 & ~n14968 ) | ( n320 & n24002 ) | ( ~n14968 & n24002 ) ;
  assign n30021 = ( ~n1489 & n2286 ) | ( ~n1489 & n30020 ) | ( n2286 & n30020 ) ;
  assign n30022 = n27120 ^ n16495 ^ n6111 ;
  assign n30023 = ( n2066 & n20520 ) | ( n2066 & ~n30022 ) | ( n20520 & ~n30022 ) ;
  assign n30024 = n30023 ^ n13564 ^ n6051 ;
  assign n30025 = n10206 ^ n9040 ^ n7570 ;
  assign n30026 = ( n16779 & ~n28966 ) | ( n16779 & n30025 ) | ( ~n28966 & n30025 ) ;
  assign n30027 = n29813 ^ n3946 ^ n1745 ;
  assign n30028 = n19514 ^ n18319 ^ n3314 ;
  assign n30029 = ( n2081 & n14761 ) | ( n2081 & ~n30028 ) | ( n14761 & ~n30028 ) ;
  assign n30031 = ( n5526 & n6564 ) | ( n5526 & n17747 ) | ( n6564 & n17747 ) ;
  assign n30030 = n8596 ^ n8351 ^ n6589 ;
  assign n30032 = n30031 ^ n30030 ^ n6579 ;
  assign n30033 = ( n3796 & n16188 ) | ( n3796 & n30032 ) | ( n16188 & n30032 ) ;
  assign n30034 = n30033 ^ n17872 ^ n2008 ;
  assign n30035 = n15614 ^ n6981 ^ n4997 ;
  assign n30037 = ( n11159 & n20731 ) | ( n11159 & ~n21717 ) | ( n20731 & ~n21717 ) ;
  assign n30036 = n23852 ^ n19977 ^ n6247 ;
  assign n30038 = n30037 ^ n30036 ^ n26985 ;
  assign n30039 = ( n16328 & n16378 ) | ( n16328 & n25361 ) | ( n16378 & n25361 ) ;
  assign n30040 = ( ~n11354 & n22081 ) | ( ~n11354 & n30039 ) | ( n22081 & n30039 ) ;
  assign n30041 = n28735 ^ n21049 ^ n11022 ;
  assign n30044 = ( ~n1147 & n9039 ) | ( ~n1147 & n10196 ) | ( n9039 & n10196 ) ;
  assign n30042 = ( n6058 & n18251 ) | ( n6058 & ~n26834 ) | ( n18251 & ~n26834 ) ;
  assign n30043 = ( ~n831 & n7629 ) | ( ~n831 & n30042 ) | ( n7629 & n30042 ) ;
  assign n30045 = n30044 ^ n30043 ^ n244 ;
  assign n30046 = n30045 ^ n14288 ^ n11012 ;
  assign n30047 = ( n5742 & n8483 ) | ( n5742 & n30046 ) | ( n8483 & n30046 ) ;
  assign n30048 = ( n3584 & ~n4628 ) | ( n3584 & n10148 ) | ( ~n4628 & n10148 ) ;
  assign n30049 = n30048 ^ n27305 ^ n26236 ;
  assign n30050 = n19272 ^ n3244 ^ n2127 ;
  assign n30051 = n13187 ^ n8890 ^ n335 ;
  assign n30052 = n30051 ^ n14651 ^ n5041 ;
  assign n30053 = ( ~n15182 & n15759 ) | ( ~n15182 & n21473 ) | ( n15759 & n21473 ) ;
  assign n30054 = ( ~n4548 & n15261 ) | ( ~n4548 & n25842 ) | ( n15261 & n25842 ) ;
  assign n30055 = ( n11720 & n16228 ) | ( n11720 & ~n30054 ) | ( n16228 & ~n30054 ) ;
  assign n30056 = n30055 ^ n16598 ^ n3653 ;
  assign n30057 = n11021 ^ n9576 ^ n5703 ;
  assign n30058 = ( ~n5076 & n24484 ) | ( ~n5076 & n29635 ) | ( n24484 & n29635 ) ;
  assign n30059 = n29246 ^ n26343 ^ n2739 ;
  assign n30060 = n25856 ^ n14109 ^ n11527 ;
  assign n30061 = n30060 ^ n27077 ^ n15123 ;
  assign n30062 = n30061 ^ n19845 ^ n1507 ;
  assign n30064 = ( n5030 & ~n6370 ) | ( n5030 & n11061 ) | ( ~n6370 & n11061 ) ;
  assign n30063 = n28302 ^ n25321 ^ n9776 ;
  assign n30065 = n30064 ^ n30063 ^ n25582 ;
  assign n30066 = n23709 ^ n14332 ^ n5548 ;
  assign n30067 = n30066 ^ n13296 ^ n6820 ;
  assign n30068 = n30067 ^ n20506 ^ n3734 ;
  assign n30069 = n4261 ^ n3052 ^ n266 ;
  assign n30070 = n30069 ^ n19318 ^ n3274 ;
  assign n30071 = n8817 ^ n4371 ^ n2169 ;
  assign n30072 = n30071 ^ n5841 ^ n4247 ;
  assign n30073 = n11205 ^ n5022 ^ n131 ;
  assign n30074 = n30073 ^ n29087 ^ n11586 ;
  assign n30075 = ( n5491 & n5617 ) | ( n5491 & n25692 ) | ( n5617 & n25692 ) ;
  assign n30076 = n22594 ^ n13123 ^ n2238 ;
  assign n30077 = n30076 ^ n29838 ^ n23776 ;
  assign n30079 = n10324 ^ n2751 ^ n1484 ;
  assign n30078 = n20582 ^ n6522 ^ n3023 ;
  assign n30080 = n30079 ^ n30078 ^ n3443 ;
  assign n30081 = ( n6358 & n8506 ) | ( n6358 & n18884 ) | ( n8506 & n18884 ) ;
  assign n30082 = n10193 ^ n3425 ^ n2824 ;
  assign n30083 = ( n14278 & n15431 ) | ( n14278 & n16460 ) | ( n15431 & n16460 ) ;
  assign n30084 = n13555 ^ n6169 ^ n5011 ;
  assign n30085 = ( n246 & ~n13018 ) | ( n246 & n30084 ) | ( ~n13018 & n30084 ) ;
  assign n30086 = ( n20558 & ~n30083 ) | ( n20558 & n30085 ) | ( ~n30083 & n30085 ) ;
  assign n30087 = ( n4391 & ~n6937 ) | ( n4391 & n9627 ) | ( ~n6937 & n9627 ) ;
  assign n30088 = n23607 ^ n15152 ^ n6142 ;
  assign n30089 = n30088 ^ n6731 ^ n823 ;
  assign n30090 = ( n1316 & n1338 ) | ( n1316 & ~n1926 ) | ( n1338 & ~n1926 ) ;
  assign n30091 = n30090 ^ n25661 ^ n16905 ;
  assign n30092 = n30091 ^ n24766 ^ n7884 ;
  assign n30093 = ( n3153 & ~n5351 ) | ( n3153 & n6867 ) | ( ~n5351 & n6867 ) ;
  assign n30094 = n30093 ^ n25244 ^ n18677 ;
  assign n30095 = ( n24883 & n26380 ) | ( n24883 & ~n30094 ) | ( n26380 & ~n30094 ) ;
  assign n30096 = n30095 ^ n27200 ^ n26772 ;
  assign n30097 = ( n8681 & n23169 ) | ( n8681 & n24766 ) | ( n23169 & n24766 ) ;
  assign n30098 = n30097 ^ n18625 ^ n2548 ;
  assign n30099 = ( n10485 & n20683 ) | ( n10485 & n30098 ) | ( n20683 & n30098 ) ;
  assign n30100 = n14547 ^ n10451 ^ n5455 ;
  assign n30101 = n30100 ^ n9339 ^ n8595 ;
  assign n30102 = ( n4367 & n5220 ) | ( n4367 & ~n7744 ) | ( n5220 & ~n7744 ) ;
  assign n30103 = ( n3208 & ~n8822 ) | ( n3208 & n30102 ) | ( ~n8822 & n30102 ) ;
  assign n30104 = ( n18226 & n28773 ) | ( n18226 & n30103 ) | ( n28773 & n30103 ) ;
  assign n30105 = ( n1325 & n14639 ) | ( n1325 & n17548 ) | ( n14639 & n17548 ) ;
  assign n30106 = n17115 ^ n13041 ^ n12163 ;
  assign n30107 = ( ~n25584 & n30105 ) | ( ~n25584 & n30106 ) | ( n30105 & n30106 ) ;
  assign n30108 = ( n1648 & n2373 ) | ( n1648 & ~n9797 ) | ( n2373 & ~n9797 ) ;
  assign n30109 = ( n6256 & n12183 ) | ( n6256 & n23172 ) | ( n12183 & n23172 ) ;
  assign n30110 = n30109 ^ n21824 ^ n13813 ;
  assign n30111 = ( n10220 & n26380 ) | ( n10220 & n30110 ) | ( n26380 & n30110 ) ;
  assign n30112 = n30111 ^ n24598 ^ n6920 ;
  assign n30117 = n24564 ^ n14590 ^ n1921 ;
  assign n30118 = n30117 ^ n19904 ^ n4517 ;
  assign n30115 = n11078 ^ n8005 ^ n7121 ;
  assign n30114 = ( n4682 & ~n7034 ) | ( n4682 & n15969 ) | ( ~n7034 & n15969 ) ;
  assign n30116 = n30115 ^ n30114 ^ n21856 ;
  assign n30113 = ( n2440 & ~n11154 ) | ( n2440 & n21487 ) | ( ~n11154 & n21487 ) ;
  assign n30119 = n30118 ^ n30116 ^ n30113 ;
  assign n30120 = n2386 ^ n1994 ^ n762 ;
  assign n30121 = n25379 ^ n18507 ^ n4765 ;
  assign n30122 = ( n11963 & n18799 ) | ( n11963 & ~n30121 ) | ( n18799 & ~n30121 ) ;
  assign n30123 = ( n5047 & n11445 ) | ( n5047 & n23746 ) | ( n11445 & n23746 ) ;
  assign n30124 = ( n3001 & n5009 ) | ( n3001 & n16107 ) | ( n5009 & n16107 ) ;
  assign n30125 = ( ~n2643 & n20031 ) | ( ~n2643 & n30124 ) | ( n20031 & n30124 ) ;
  assign n30126 = ( ~n3236 & n16187 ) | ( ~n3236 & n30125 ) | ( n16187 & n30125 ) ;
  assign n30127 = n28483 ^ n23978 ^ n392 ;
  assign n30128 = n30127 ^ n13314 ^ n8453 ;
  assign n30129 = n13183 ^ n4744 ^ n3544 ;
  assign n30130 = n6824 ^ n3368 ^ n2923 ;
  assign n30131 = ( n19820 & n28169 ) | ( n19820 & n30130 ) | ( n28169 & n30130 ) ;
  assign n30132 = ( n20231 & n30129 ) | ( n20231 & ~n30131 ) | ( n30129 & ~n30131 ) ;
  assign n30133 = n12583 ^ n6336 ^ n4598 ;
  assign n30134 = n11895 ^ n11158 ^ n1494 ;
  assign n30135 = n30134 ^ n17102 ^ n7024 ;
  assign n30136 = n30135 ^ n14676 ^ n10060 ;
  assign n30137 = ( n9370 & n23935 ) | ( n9370 & n30136 ) | ( n23935 & n30136 ) ;
  assign n30138 = ( ~n8652 & n10754 ) | ( ~n8652 & n12165 ) | ( n10754 & n12165 ) ;
  assign n30139 = n30138 ^ n7597 ^ n903 ;
  assign n30140 = ( ~n30133 & n30137 ) | ( ~n30133 & n30139 ) | ( n30137 & n30139 ) ;
  assign n30141 = n22960 ^ n9203 ^ n710 ;
  assign n30142 = n28167 ^ n21663 ^ n9043 ;
  assign n30143 = ( n7781 & n30141 ) | ( n7781 & n30142 ) | ( n30141 & n30142 ) ;
  assign n30144 = ( n1831 & n19002 ) | ( n1831 & n22249 ) | ( n19002 & n22249 ) ;
  assign n30145 = n17800 ^ n4914 ^ n1429 ;
  assign n30146 = n30145 ^ n7756 ^ n5703 ;
  assign n30147 = ( n1097 & n25625 ) | ( n1097 & n26660 ) | ( n25625 & n26660 ) ;
  assign n30148 = ( n22444 & ~n30146 ) | ( n22444 & n30147 ) | ( ~n30146 & n30147 ) ;
  assign n30149 = ( n3006 & n13685 ) | ( n3006 & n19149 ) | ( n13685 & n19149 ) ;
  assign n30150 = ( n9582 & ~n16326 ) | ( n9582 & n30149 ) | ( ~n16326 & n30149 ) ;
  assign n30151 = ( n751 & n997 ) | ( n751 & n25474 ) | ( n997 & n25474 ) ;
  assign n30152 = ( ~n1088 & n4568 ) | ( ~n1088 & n9707 ) | ( n4568 & n9707 ) ;
  assign n30153 = ( ~n19330 & n26907 ) | ( ~n19330 & n30152 ) | ( n26907 & n30152 ) ;
  assign n30154 = ( n1491 & n6949 ) | ( n1491 & ~n13780 ) | ( n6949 & ~n13780 ) ;
  assign n30155 = n12620 ^ n9473 ^ n1071 ;
  assign n30156 = ( n7095 & ~n7895 ) | ( n7095 & n15086 ) | ( ~n7895 & n15086 ) ;
  assign n30157 = n30156 ^ n18658 ^ n152 ;
  assign n30158 = n24482 ^ n19025 ^ n1894 ;
  assign n30159 = n30158 ^ n25210 ^ n16014 ;
  assign n30160 = ( n5309 & n10739 ) | ( n5309 & ~n16284 ) | ( n10739 & ~n16284 ) ;
  assign n30161 = n12836 ^ n10876 ^ n5542 ;
  assign n30163 = n21869 ^ n17791 ^ n17288 ;
  assign n30162 = n16815 ^ n16303 ^ n13467 ;
  assign n30164 = n30163 ^ n30162 ^ n24913 ;
  assign n30165 = n20361 ^ n14425 ^ n4665 ;
  assign n30166 = ( n7715 & ~n10827 ) | ( n7715 & n29145 ) | ( ~n10827 & n29145 ) ;
  assign n30167 = n30166 ^ n16884 ^ n3919 ;
  assign n30168 = ( n755 & n30165 ) | ( n755 & n30167 ) | ( n30165 & n30167 ) ;
  assign n30169 = ( ~n3761 & n8548 ) | ( ~n3761 & n22168 ) | ( n8548 & n22168 ) ;
  assign n30170 = ( n7022 & ~n15749 ) | ( n7022 & n17419 ) | ( ~n15749 & n17419 ) ;
  assign n30171 = n15733 ^ n13150 ^ n2064 ;
  assign n30172 = n30171 ^ n19735 ^ n8931 ;
  assign n30173 = ( n2892 & n8128 ) | ( n2892 & ~n30172 ) | ( n8128 & ~n30172 ) ;
  assign n30174 = n13383 ^ n10771 ^ n2182 ;
  assign n30175 = n30174 ^ n21267 ^ n7216 ;
  assign n30176 = ( ~n8289 & n15437 ) | ( ~n8289 & n30175 ) | ( n15437 & n30175 ) ;
  assign n30180 = ( n2877 & n9047 ) | ( n2877 & n14535 ) | ( n9047 & n14535 ) ;
  assign n30178 = n21523 ^ n12476 ^ n5382 ;
  assign n30177 = ( n9348 & n14437 ) | ( n9348 & n17100 ) | ( n14437 & n17100 ) ;
  assign n30179 = n30178 ^ n30177 ^ n2022 ;
  assign n30181 = n30180 ^ n30179 ^ n711 ;
  assign n30182 = n23196 ^ n12564 ^ n2733 ;
  assign n30183 = ( n8473 & ~n15089 ) | ( n8473 & n24617 ) | ( ~n15089 & n24617 ) ;
  assign n30184 = ( n326 & n4067 ) | ( n326 & ~n10393 ) | ( n4067 & ~n10393 ) ;
  assign n30185 = n10392 ^ n8574 ^ n1803 ;
  assign n30186 = n30185 ^ n29566 ^ n19843 ;
  assign n30187 = n30186 ^ n16959 ^ n13482 ;
  assign n30188 = n29609 ^ n18488 ^ n6972 ;
  assign n30190 = ( n896 & ~n3371 ) | ( n896 & n3902 ) | ( ~n3371 & n3902 ) ;
  assign n30189 = ( n2606 & ~n4251 ) | ( n2606 & n8198 ) | ( ~n4251 & n8198 ) ;
  assign n30191 = n30190 ^ n30189 ^ n865 ;
  assign n30192 = n30191 ^ n25849 ^ n23252 ;
  assign n30193 = n22602 ^ n4018 ^ n2278 ;
  assign n30194 = ( ~n5287 & n14305 ) | ( ~n5287 & n30193 ) | ( n14305 & n30193 ) ;
  assign n30195 = ( ~n6593 & n18354 ) | ( ~n6593 & n21117 ) | ( n18354 & n21117 ) ;
  assign n30196 = ( n3015 & ~n6117 ) | ( n3015 & n7730 ) | ( ~n6117 & n7730 ) ;
  assign n30197 = n16772 ^ n16759 ^ n3888 ;
  assign n30198 = ( n22451 & n24203 ) | ( n22451 & ~n30197 ) | ( n24203 & ~n30197 ) ;
  assign n30199 = ( n5210 & n17031 ) | ( n5210 & n30198 ) | ( n17031 & n30198 ) ;
  assign n30200 = n30199 ^ n25634 ^ n16066 ;
  assign n30201 = n9096 ^ n3842 ^ n161 ;
  assign n30202 = ( n4721 & n9223 ) | ( n4721 & ~n30201 ) | ( n9223 & ~n30201 ) ;
  assign n30203 = ( n14837 & ~n20699 ) | ( n14837 & n26632 ) | ( ~n20699 & n26632 ) ;
  assign n30204 = ( n6786 & ~n26061 ) | ( n6786 & n30203 ) | ( ~n26061 & n30203 ) ;
  assign n30205 = ( n4197 & n17409 ) | ( n4197 & ~n28831 ) | ( n17409 & ~n28831 ) ;
  assign n30206 = n30205 ^ n8397 ^ n8047 ;
  assign n30207 = n30206 ^ n26177 ^ n15560 ;
  assign n30208 = n19373 ^ n4773 ^ n575 ;
  assign n30209 = ( n144 & n11530 ) | ( n144 & n13388 ) | ( n11530 & n13388 ) ;
  assign n30210 = n30209 ^ n26379 ^ n22422 ;
  assign n30211 = ( ~n6147 & n10855 ) | ( ~n6147 & n30210 ) | ( n10855 & n30210 ) ;
  assign n30212 = ( n3105 & ~n6794 ) | ( n3105 & n15431 ) | ( ~n6794 & n15431 ) ;
  assign n30213 = ( n9455 & n14605 ) | ( n9455 & n30212 ) | ( n14605 & n30212 ) ;
  assign n30214 = n22343 ^ n1645 ^ x79 ;
  assign n30215 = n28540 ^ n16897 ^ n1044 ;
  assign n30216 = n30215 ^ n23213 ^ n17557 ;
  assign n30217 = n16479 ^ n1588 ^ n978 ;
  assign n30218 = n30217 ^ n11726 ^ n7466 ;
  assign n30219 = ( ~n2219 & n5944 ) | ( ~n2219 & n30218 ) | ( n5944 & n30218 ) ;
  assign n30220 = ( n957 & ~n16989 ) | ( n957 & n23690 ) | ( ~n16989 & n23690 ) ;
  assign n30221 = ( n15839 & n16486 ) | ( n15839 & n30220 ) | ( n16486 & n30220 ) ;
  assign n30222 = n30221 ^ n23521 ^ n11129 ;
  assign n30223 = n28159 ^ n25429 ^ n14101 ;
  assign n30224 = ( ~n8565 & n17957 ) | ( ~n8565 & n30223 ) | ( n17957 & n30223 ) ;
  assign n30225 = ( x83 & ~n3746 ) | ( x83 & n10004 ) | ( ~n3746 & n10004 ) ;
  assign n30226 = n20322 ^ n18319 ^ n7993 ;
  assign n30227 = ( n545 & n9428 ) | ( n545 & n14684 ) | ( n9428 & n14684 ) ;
  assign n30228 = n21757 ^ n14379 ^ n10186 ;
  assign n30229 = n14839 ^ n11931 ^ n9149 ;
  assign n30230 = ( n14643 & ~n18100 ) | ( n14643 & n18797 ) | ( ~n18100 & n18797 ) ;
  assign n30231 = ( n7709 & n15068 ) | ( n7709 & ~n21054 ) | ( n15068 & ~n21054 ) ;
  assign n30232 = ( n4357 & n13947 ) | ( n4357 & n14878 ) | ( n13947 & n14878 ) ;
  assign n30233 = ( n20626 & ~n25116 ) | ( n20626 & n30232 ) | ( ~n25116 & n30232 ) ;
  assign n30234 = ( ~n1688 & n9517 ) | ( ~n1688 & n30233 ) | ( n9517 & n30233 ) ;
  assign n30235 = n26799 ^ n13646 ^ n12165 ;
  assign n30236 = ( n9459 & n21331 ) | ( n9459 & ~n30235 ) | ( n21331 & ~n30235 ) ;
  assign n30237 = n30236 ^ n4207 ^ n174 ;
  assign n30238 = n30237 ^ n25026 ^ n12947 ;
  assign n30242 = n9089 ^ n6366 ^ n3062 ;
  assign n30239 = ( n3095 & ~n11032 ) | ( n3095 & n17944 ) | ( ~n11032 & n17944 ) ;
  assign n30240 = ( n10701 & n15476 ) | ( n10701 & n17564 ) | ( n15476 & n17564 ) ;
  assign n30241 = ( n6624 & n30239 ) | ( n6624 & n30240 ) | ( n30239 & n30240 ) ;
  assign n30243 = n30242 ^ n30241 ^ n25989 ;
  assign n30244 = n19838 ^ n10809 ^ n8758 ;
  assign n30245 = n30244 ^ n20447 ^ n12818 ;
  assign n30247 = ( n4099 & n5671 ) | ( n4099 & ~n12752 ) | ( n5671 & ~n12752 ) ;
  assign n30246 = ( n2336 & ~n5869 ) | ( n2336 & n15729 ) | ( ~n5869 & n15729 ) ;
  assign n30248 = n30247 ^ n30246 ^ n27803 ;
  assign n30249 = ( n12153 & n27735 ) | ( n12153 & n28612 ) | ( n27735 & n28612 ) ;
  assign n30250 = n10319 ^ n5701 ^ n3164 ;
  assign n30251 = n30250 ^ n24740 ^ n2698 ;
  assign n30252 = n27234 ^ n10547 ^ n5383 ;
  assign n30253 = ( n19186 & n24478 ) | ( n19186 & n27427 ) | ( n24478 & n27427 ) ;
  assign n30254 = ( n12017 & n19681 ) | ( n12017 & n20280 ) | ( n19681 & n20280 ) ;
  assign n30255 = n30254 ^ n24783 ^ n17023 ;
  assign n30256 = ( n5554 & ~n9485 ) | ( n5554 & n15421 ) | ( ~n9485 & n15421 ) ;
  assign n30257 = n16148 ^ n15636 ^ n12715 ;
  assign n30258 = ( n9196 & n24515 ) | ( n9196 & n30257 ) | ( n24515 & n30257 ) ;
  assign y0 = ~n432 ;
  assign y1 = n498 ;
  assign y2 = ~n606 ;
  assign y3 = ~n659 ;
  assign y4 = n689 ;
  assign y5 = ~n843 ;
  assign y6 = n930 ;
  assign y7 = ~n1038 ;
  assign y8 = n1086 ;
  assign y9 = n1160 ;
  assign y10 = ~n1194 ;
  assign y11 = ~n1217 ;
  assign y12 = n1250 ;
  assign y13 = n1255 ;
  assign y14 = n1282 ;
  assign y15 = n1340 ;
  assign y16 = n1398 ;
  assign y17 = ~n1518 ;
  assign y18 = ~n1519 ;
  assign y19 = n1538 ;
  assign y20 = n1548 ;
  assign y21 = ~n1574 ;
  assign y22 = ~n1618 ;
  assign y23 = n1658 ;
  assign y24 = n1687 ;
  assign y25 = ~n1711 ;
  assign y26 = ~n1726 ;
  assign y27 = n1746 ;
  assign y28 = ~n1797 ;
  assign y29 = ~n1826 ;
  assign y30 = n1849 ;
  assign y31 = ~n1856 ;
  assign y32 = ~n1890 ;
  assign y33 = ~n1918 ;
  assign y34 = ~n1963 ;
  assign y35 = ~n1970 ;
  assign y36 = n1976 ;
  assign y37 = n2004 ;
  assign y38 = n2031 ;
  assign y39 = ~n2063 ;
  assign y40 = ~n2078 ;
  assign y41 = n2086 ;
  assign y42 = ~n2100 ;
  assign y43 = ~n2135 ;
  assign y44 = n2172 ;
  assign y45 = ~n2192 ;
  assign y46 = n2251 ;
  assign y47 = n2267 ;
  assign y48 = n2272 ;
  assign y49 = ~n2312 ;
  assign y50 = n2350 ;
  assign y51 = ~n2382 ;
  assign y52 = ~n2392 ;
  assign y53 = ~n2426 ;
  assign y54 = ~n2443 ;
  assign y55 = ~n2471 ;
  assign y56 = n2500 ;
  assign y57 = ~n2510 ;
  assign y58 = ~n2544 ;
  assign y59 = ~n2551 ;
  assign y60 = ~n2613 ;
  assign y61 = ~n2618 ;
  assign y62 = n2625 ;
  assign y63 = ~n2640 ;
  assign y64 = n2653 ;
  assign y65 = n2655 ;
  assign y66 = n2700 ;
  assign y67 = ~n2709 ;
  assign y68 = n2716 ;
  assign y69 = ~n2729 ;
  assign y70 = ~n2740 ;
  assign y71 = n2756 ;
  assign y72 = ~n2775 ;
  assign y73 = ~n2823 ;
  assign y74 = n2825 ;
  assign y75 = ~n2833 ;
  assign y76 = n2847 ;
  assign y77 = ~n2851 ;
  assign y78 = n2895 ;
  assign y79 = n2909 ;
  assign y80 = ~n2922 ;
  assign y81 = n2936 ;
  assign y82 = n2940 ;
  assign y83 = n2963 ;
  assign y84 = n2979 ;
  assign y85 = ~n2980 ;
  assign y86 = n2992 ;
  assign y87 = n3012 ;
  assign y88 = ~n3032 ;
  assign y89 = n3040 ;
  assign y90 = ~n3075 ;
  assign y91 = n3099 ;
  assign y92 = n3121 ;
  assign y93 = ~n3146 ;
  assign y94 = ~n3158 ;
  assign y95 = ~n3171 ;
  assign y96 = n3173 ;
  assign y97 = n3176 ;
  assign y98 = ~n3195 ;
  assign y99 = n3197 ;
  assign y100 = n3224 ;
  assign y101 = n3251 ;
  assign y102 = n3266 ;
  assign y103 = ~n3279 ;
  assign y104 = ~n3302 ;
  assign y105 = ~n3330 ;
  assign y106 = n3337 ;
  assign y107 = ~n3390 ;
  assign y108 = n3402 ;
  assign y109 = n3410 ;
  assign y110 = n3411 ;
  assign y111 = ~n3415 ;
  assign y112 = n3465 ;
  assign y113 = ~n3474 ;
  assign y114 = n3500 ;
  assign y115 = ~n3538 ;
  assign y116 = n3558 ;
  assign y117 = n3573 ;
  assign y118 = n3580 ;
  assign y119 = n3583 ;
  assign y120 = ~n3599 ;
  assign y121 = ~n3604 ;
  assign y122 = n3615 ;
  assign y123 = ~n3623 ;
  assign y124 = ~n3646 ;
  assign y125 = n3662 ;
  assign y126 = n3680 ;
  assign y127 = ~n3685 ;
  assign y128 = ~n3709 ;
  assign y129 = n3727 ;
  assign y130 = ~n3751 ;
  assign y131 = ~n3759 ;
  assign y132 = ~n3769 ;
  assign y133 = n3815 ;
  assign y134 = ~n3823 ;
  assign y135 = n3872 ;
  assign y136 = ~n3899 ;
  assign y137 = n3915 ;
  assign y138 = ~n3916 ;
  assign y139 = n3920 ;
  assign y140 = ~n3955 ;
  assign y141 = n3958 ;
  assign y142 = n3983 ;
  assign y143 = n3994 ;
  assign y144 = ~n3998 ;
  assign y145 = ~n4017 ;
  assign y146 = ~n4022 ;
  assign y147 = n4033 ;
  assign y148 = ~n4057 ;
  assign y149 = n4075 ;
  assign y150 = ~n4106 ;
  assign y151 = n4118 ;
  assign y152 = n4138 ;
  assign y153 = n4139 ;
  assign y154 = ~n4164 ;
  assign y155 = ~n4178 ;
  assign y156 = ~n4196 ;
  assign y157 = n4201 ;
  assign y158 = ~n4203 ;
  assign y159 = n4208 ;
  assign y160 = ~n4231 ;
  assign y161 = ~n4246 ;
  assign y162 = n4262 ;
  assign y163 = n4268 ;
  assign y164 = ~n4277 ;
  assign y165 = n4304 ;
  assign y166 = n4317 ;
  assign y167 = ~n4320 ;
  assign y168 = ~n4333 ;
  assign y169 = n4337 ;
  assign y170 = n4356 ;
  assign y171 = n4390 ;
  assign y172 = n4395 ;
  assign y173 = ~n4400 ;
  assign y174 = n4404 ;
  assign y175 = n4427 ;
  assign y176 = n4505 ;
  assign y177 = n4523 ;
  assign y178 = n4528 ;
  assign y179 = ~n4532 ;
  assign y180 = ~n4534 ;
  assign y181 = n4535 ;
  assign y182 = n4547 ;
  assign y183 = n4560 ;
  assign y184 = ~n4575 ;
  assign y185 = ~n4581 ;
  assign y186 = ~n4601 ;
  assign y187 = n4632 ;
  assign y188 = ~n4643 ;
  assign y189 = ~n4655 ;
  assign y190 = ~n4657 ;
  assign y191 = n4668 ;
  assign y192 = n4685 ;
  assign y193 = n4688 ;
  assign y194 = ~n4698 ;
  assign y195 = ~n4719 ;
  assign y196 = ~n4728 ;
  assign y197 = ~n4730 ;
  assign y198 = n4735 ;
  assign y199 = n4754 ;
  assign y200 = n4776 ;
  assign y201 = ~n4788 ;
  assign y202 = ~n4792 ;
  assign y203 = n4802 ;
  assign y204 = ~n4807 ;
  assign y205 = n4815 ;
  assign y206 = n4826 ;
  assign y207 = n4830 ;
  assign y208 = n4836 ;
  assign y209 = ~n4844 ;
  assign y210 = ~n4854 ;
  assign y211 = ~n4877 ;
  assign y212 = ~n4880 ;
  assign y213 = n4889 ;
  assign y214 = n4896 ;
  assign y215 = n4906 ;
  assign y216 = ~n4912 ;
  assign y217 = n4923 ;
  assign y218 = ~n4934 ;
  assign y219 = n4946 ;
  assign y220 = n4964 ;
  assign y221 = n4969 ;
  assign y222 = n4972 ;
  assign y223 = ~n4975 ;
  assign y224 = n4978 ;
  assign y225 = n4987 ;
  assign y226 = ~n5000 ;
  assign y227 = n5012 ;
  assign y228 = n5014 ;
  assign y229 = n5033 ;
  assign y230 = n5036 ;
  assign y231 = n5063 ;
  assign y232 = n5083 ;
  assign y233 = n5085 ;
  assign y234 = ~n5088 ;
  assign y235 = n5094 ;
  assign y236 = ~n5096 ;
  assign y237 = n5098 ;
  assign y238 = n5115 ;
  assign y239 = ~n5145 ;
  assign y240 = n5148 ;
  assign y241 = n5156 ;
  assign y242 = n5158 ;
  assign y243 = n5188 ;
  assign y244 = ~n5192 ;
  assign y245 = n5201 ;
  assign y246 = n5242 ;
  assign y247 = n5250 ;
  assign y248 = n5268 ;
  assign y249 = n5277 ;
  assign y250 = n5290 ;
  assign y251 = n5300 ;
  assign y252 = n5338 ;
  assign y253 = n5355 ;
  assign y254 = ~n5365 ;
  assign y255 = n5389 ;
  assign y256 = n5413 ;
  assign y257 = n5423 ;
  assign y258 = ~n5430 ;
  assign y259 = n5431 ;
  assign y260 = ~n5443 ;
  assign y261 = ~n5453 ;
  assign y262 = ~n5458 ;
  assign y263 = n5481 ;
  assign y264 = n5490 ;
  assign y265 = ~n5499 ;
  assign y266 = n5507 ;
  assign y267 = ~n5517 ;
  assign y268 = ~n5523 ;
  assign y269 = n5532 ;
  assign y270 = ~n5534 ;
  assign y271 = n5535 ;
  assign y272 = n5537 ;
  assign y273 = ~n5543 ;
  assign y274 = ~n5562 ;
  assign y275 = ~n5568 ;
  assign y276 = n5576 ;
  assign y277 = n5591 ;
  assign y278 = n5599 ;
  assign y279 = ~n5602 ;
  assign y280 = n5606 ;
  assign y281 = ~n5611 ;
  assign y282 = n5619 ;
  assign y283 = ~n5629 ;
  assign y284 = n5637 ;
  assign y285 = n5641 ;
  assign y286 = ~n5656 ;
  assign y287 = n5658 ;
  assign y288 = ~n5667 ;
  assign y289 = n5672 ;
  assign y290 = ~n5673 ;
  assign y291 = ~n5688 ;
  assign y292 = n5693 ;
  assign y293 = n5697 ;
  assign y294 = n5707 ;
  assign y295 = n5711 ;
  assign y296 = ~n5717 ;
  assign y297 = ~n5738 ;
  assign y298 = ~n5752 ;
  assign y299 = n5756 ;
  assign y300 = n5760 ;
  assign y301 = ~n5764 ;
  assign y302 = n5778 ;
  assign y303 = n5790 ;
  assign y304 = n5812 ;
  assign y305 = n5821 ;
  assign y306 = ~n5828 ;
  assign y307 = n5852 ;
  assign y308 = ~n5875 ;
  assign y309 = ~n5877 ;
  assign y310 = n5878 ;
  assign y311 = ~n5888 ;
  assign y312 = n5894 ;
  assign y313 = ~n5907 ;
  assign y314 = ~n5910 ;
  assign y315 = ~n5917 ;
  assign y316 = ~n5925 ;
  assign y317 = ~n5929 ;
  assign y318 = n5960 ;
  assign y319 = n5964 ;
  assign y320 = ~n5977 ;
  assign y321 = ~n5986 ;
  assign y322 = n5992 ;
  assign y323 = ~n5995 ;
  assign y324 = ~n6000 ;
  assign y325 = n6006 ;
  assign y326 = ~n6007 ;
  assign y327 = ~n6010 ;
  assign y328 = ~n6027 ;
  assign y329 = ~n6052 ;
  assign y330 = n6061 ;
  assign y331 = ~n6073 ;
  assign y332 = ~n6078 ;
  assign y333 = ~n6091 ;
  assign y334 = ~n6112 ;
  assign y335 = ~n6139 ;
  assign y336 = n6144 ;
  assign y337 = n6151 ;
  assign y338 = n6152 ;
  assign y339 = n6180 ;
  assign y340 = n6182 ;
  assign y341 = n6192 ;
  assign y342 = ~n6198 ;
  assign y343 = ~n6205 ;
  assign y344 = n6233 ;
  assign y345 = n6242 ;
  assign y346 = n6249 ;
  assign y347 = ~n6255 ;
  assign y348 = n6261 ;
  assign y349 = ~n6286 ;
  assign y350 = n6290 ;
  assign y351 = n6307 ;
  assign y352 = n6349 ;
  assign y353 = ~n6354 ;
  assign y354 = ~n6364 ;
  assign y355 = ~n6374 ;
  assign y356 = ~n6378 ;
  assign y357 = ~n6385 ;
  assign y358 = ~n6389 ;
  assign y359 = n6398 ;
  assign y360 = n6407 ;
  assign y361 = ~n6413 ;
  assign y362 = n6418 ;
  assign y363 = ~n6438 ;
  assign y364 = n6449 ;
  assign y365 = n6455 ;
  assign y366 = n6459 ;
  assign y367 = n6476 ;
  assign y368 = n6477 ;
  assign y369 = n6478 ;
  assign y370 = ~n6479 ;
  assign y371 = n6481 ;
  assign y372 = ~n6493 ;
  assign y373 = n6494 ;
  assign y374 = n6503 ;
  assign y375 = n6504 ;
  assign y376 = ~n6508 ;
  assign y377 = n6510 ;
  assign y378 = ~n6523 ;
  assign y379 = ~n6528 ;
  assign y380 = ~n6535 ;
  assign y381 = ~n6536 ;
  assign y382 = ~n6538 ;
  assign y383 = n6551 ;
  assign y384 = n6560 ;
  assign y385 = ~n6587 ;
  assign y386 = ~n6596 ;
  assign y387 = ~n6597 ;
  assign y388 = ~n6599 ;
  assign y389 = ~n6606 ;
  assign y390 = n6608 ;
  assign y391 = n6613 ;
  assign y392 = ~n6626 ;
  assign y393 = ~n6628 ;
  assign y394 = ~n6637 ;
  assign y395 = n6644 ;
  assign y396 = n6647 ;
  assign y397 = n6662 ;
  assign y398 = n6663 ;
  assign y399 = ~n6675 ;
  assign y400 = ~n6677 ;
  assign y401 = ~n6679 ;
  assign y402 = n6683 ;
  assign y403 = ~n6707 ;
  assign y404 = n6718 ;
  assign y405 = n6721 ;
  assign y406 = n6729 ;
  assign y407 = n6730 ;
  assign y408 = n6750 ;
  assign y409 = n6763 ;
  assign y410 = n6764 ;
  assign y411 = n6774 ;
  assign y412 = n6778 ;
  assign y413 = n6779 ;
  assign y414 = n6781 ;
  assign y415 = ~n6782 ;
  assign y416 = n6797 ;
  assign y417 = n6800 ;
  assign y418 = n6813 ;
  assign y419 = ~n6821 ;
  assign y420 = n6827 ;
  assign y421 = ~n6840 ;
  assign y422 = n6841 ;
  assign y423 = n6847 ;
  assign y424 = n6851 ;
  assign y425 = n6858 ;
  assign y426 = ~n6888 ;
  assign y427 = n6900 ;
  assign y428 = n6903 ;
  assign y429 = ~n6908 ;
  assign y430 = n6909 ;
  assign y431 = ~n6916 ;
  assign y432 = n6921 ;
  assign y433 = ~n6931 ;
  assign y434 = ~n6934 ;
  assign y435 = n6938 ;
  assign y436 = n6939 ;
  assign y437 = ~n6951 ;
  assign y438 = ~n6962 ;
  assign y439 = ~n6969 ;
  assign y440 = ~n6985 ;
  assign y441 = n6993 ;
  assign y442 = ~n6998 ;
  assign y443 = ~n7013 ;
  assign y444 = ~n7021 ;
  assign y445 = n7029 ;
  assign y446 = n7047 ;
  assign y447 = ~n7062 ;
  assign y448 = ~n7064 ;
  assign y449 = n7069 ;
  assign y450 = n7073 ;
  assign y451 = ~n7075 ;
  assign y452 = ~n7079 ;
  assign y453 = n7080 ;
  assign y454 = ~n7081 ;
  assign y455 = n7082 ;
  assign y456 = n7101 ;
  assign y457 = ~n7111 ;
  assign y458 = n7122 ;
  assign y459 = ~n7127 ;
  assign y460 = n7128 ;
  assign y461 = ~n7138 ;
  assign y462 = ~n7139 ;
  assign y463 = n7141 ;
  assign y464 = ~n7157 ;
  assign y465 = ~n7167 ;
  assign y466 = n7179 ;
  assign y467 = ~n7193 ;
  assign y468 = ~n7203 ;
  assign y469 = n7208 ;
  assign y470 = n7213 ;
  assign y471 = n7227 ;
  assign y472 = n7233 ;
  assign y473 = n7234 ;
  assign y474 = n7236 ;
  assign y475 = n7237 ;
  assign y476 = n7244 ;
  assign y477 = ~n7249 ;
  assign y478 = ~n7258 ;
  assign y479 = ~n7259 ;
  assign y480 = n7268 ;
  assign y481 = ~n7279 ;
  assign y482 = ~n7284 ;
  assign y483 = n7286 ;
  assign y484 = n7290 ;
  assign y485 = n7291 ;
  assign y486 = n7293 ;
  assign y487 = ~n7305 ;
  assign y488 = ~n7309 ;
  assign y489 = n7341 ;
  assign y490 = ~n7351 ;
  assign y491 = n7366 ;
  assign y492 = n7372 ;
  assign y493 = ~n7373 ;
  assign y494 = n7387 ;
  assign y495 = ~n7400 ;
  assign y496 = n7404 ;
  assign y497 = n7415 ;
  assign y498 = n7417 ;
  assign y499 = ~n7430 ;
  assign y500 = n7439 ;
  assign y501 = ~n7440 ;
  assign y502 = n7442 ;
  assign y503 = n7446 ;
  assign y504 = ~n7448 ;
  assign y505 = n7451 ;
  assign y506 = ~n7462 ;
  assign y507 = ~n7467 ;
  assign y508 = ~n7477 ;
  assign y509 = ~n7478 ;
  assign y510 = n7487 ;
  assign y511 = n7492 ;
  assign y512 = ~n7496 ;
  assign y513 = ~n7504 ;
  assign y514 = ~n7514 ;
  assign y515 = ~n7519 ;
  assign y516 = ~n7521 ;
  assign y517 = n7524 ;
  assign y518 = ~n7527 ;
  assign y519 = n7535 ;
  assign y520 = ~n7540 ;
  assign y521 = ~n7546 ;
  assign y522 = n7553 ;
  assign y523 = n7568 ;
  assign y524 = ~n7580 ;
  assign y525 = n7584 ;
  assign y526 = n7587 ;
  assign y527 = ~n7605 ;
  assign y528 = ~n7617 ;
  assign y529 = ~n7626 ;
  assign y530 = n7637 ;
  assign y531 = n7639 ;
  assign y532 = n7644 ;
  assign y533 = n7645 ;
  assign y534 = n7652 ;
  assign y535 = n7653 ;
  assign y536 = ~n7656 ;
  assign y537 = ~n7661 ;
  assign y538 = n7662 ;
  assign y539 = n7676 ;
  assign y540 = ~n7682 ;
  assign y541 = ~n7690 ;
  assign y542 = ~n7691 ;
  assign y543 = ~n7706 ;
  assign y544 = ~n7708 ;
  assign y545 = n7710 ;
  assign y546 = ~n7718 ;
  assign y547 = n7721 ;
  assign y548 = ~n7733 ;
  assign y549 = n7735 ;
  assign y550 = ~n7739 ;
  assign y551 = ~n7740 ;
  assign y552 = n7742 ;
  assign y553 = ~n7749 ;
  assign y554 = n7757 ;
  assign y555 = n7765 ;
  assign y556 = ~n7771 ;
  assign y557 = n7785 ;
  assign y558 = ~n7786 ;
  assign y559 = n7800 ;
  assign y560 = ~n7806 ;
  assign y561 = ~n7828 ;
  assign y562 = n7837 ;
  assign y563 = ~n7844 ;
  assign y564 = n7860 ;
  assign y565 = n7872 ;
  assign y566 = ~n7876 ;
  assign y567 = ~n7883 ;
  assign y568 = n7888 ;
  assign y569 = n7894 ;
  assign y570 = n7906 ;
  assign y571 = n7916 ;
  assign y572 = n7921 ;
  assign y573 = n7948 ;
  assign y574 = n7963 ;
  assign y575 = ~n7973 ;
  assign y576 = n7977 ;
  assign y577 = ~n7984 ;
  assign y578 = n8002 ;
  assign y579 = n8015 ;
  assign y580 = ~n8021 ;
  assign y581 = ~n8023 ;
  assign y582 = ~n8024 ;
  assign y583 = ~n8034 ;
  assign y584 = ~n8035 ;
  assign y585 = ~n8057 ;
  assign y586 = ~n8071 ;
  assign y587 = ~n8076 ;
  assign y588 = n8078 ;
  assign y589 = ~n8081 ;
  assign y590 = n8085 ;
  assign y591 = n8086 ;
  assign y592 = ~n8096 ;
  assign y593 = n8104 ;
  assign y594 = ~n8111 ;
  assign y595 = n8120 ;
  assign y596 = ~n8124 ;
  assign y597 = ~n8134 ;
  assign y598 = ~n8151 ;
  assign y599 = n8158 ;
  assign y600 = ~n8174 ;
  assign y601 = n8184 ;
  assign y602 = n8188 ;
  assign y603 = ~n8190 ;
  assign y604 = ~n8193 ;
  assign y605 = n8197 ;
  assign y606 = ~n8213 ;
  assign y607 = n8219 ;
  assign y608 = n8223 ;
  assign y609 = n8224 ;
  assign y610 = n8232 ;
  assign y611 = ~n8235 ;
  assign y612 = ~n8241 ;
  assign y613 = n8256 ;
  assign y614 = n8261 ;
  assign y615 = ~n8265 ;
  assign y616 = n8273 ;
  assign y617 = n8279 ;
  assign y618 = n8284 ;
  assign y619 = n8291 ;
  assign y620 = n8297 ;
  assign y621 = ~n8305 ;
  assign y622 = n8307 ;
  assign y623 = ~n8311 ;
  assign y624 = ~n8313 ;
  assign y625 = n8319 ;
  assign y626 = n8321 ;
  assign y627 = ~n8323 ;
  assign y628 = n8343 ;
  assign y629 = n8346 ;
  assign y630 = n8357 ;
  assign y631 = ~n8359 ;
  assign y632 = ~n8373 ;
  assign y633 = n8388 ;
  assign y634 = n8394 ;
  assign y635 = ~n8400 ;
  assign y636 = n8416 ;
  assign y637 = ~n8424 ;
  assign y638 = n8426 ;
  assign y639 = n8440 ;
  assign y640 = ~n8455 ;
  assign y641 = n8469 ;
  assign y642 = n8478 ;
  assign y643 = ~n8482 ;
  assign y644 = n8485 ;
  assign y645 = ~n8492 ;
  assign y646 = n8495 ;
  assign y647 = n8505 ;
  assign y648 = n8519 ;
  assign y649 = ~n8528 ;
  assign y650 = n8531 ;
  assign y651 = ~n8541 ;
  assign y652 = ~n8547 ;
  assign y653 = ~n8550 ;
  assign y654 = n8578 ;
  assign y655 = n8579 ;
  assign y656 = ~n8581 ;
  assign y657 = ~n8592 ;
  assign y658 = n8599 ;
  assign y659 = ~n8602 ;
  assign y660 = ~n8607 ;
  assign y661 = ~n8611 ;
  assign y662 = n8613 ;
  assign y663 = n8623 ;
  assign y664 = ~n8628 ;
  assign y665 = n8640 ;
  assign y666 = ~n8644 ;
  assign y667 = n8646 ;
  assign y668 = n8656 ;
  assign y669 = n8659 ;
  assign y670 = n8663 ;
  assign y671 = n8672 ;
  assign y672 = ~n8676 ;
  assign y673 = ~n8679 ;
  assign y674 = n8683 ;
  assign y675 = ~n8693 ;
  assign y676 = n8699 ;
  assign y677 = n8700 ;
  assign y678 = n8701 ;
  assign y679 = n8706 ;
  assign y680 = ~n8707 ;
  assign y681 = ~n8709 ;
  assign y682 = ~n8710 ;
  assign y683 = n8715 ;
  assign y684 = ~n8720 ;
  assign y685 = ~n8721 ;
  assign y686 = n8726 ;
  assign y687 = ~n8731 ;
  assign y688 = n8744 ;
  assign y689 = ~n8751 ;
  assign y690 = ~n8752 ;
  assign y691 = ~n8764 ;
  assign y692 = n8776 ;
  assign y693 = ~n8784 ;
  assign y694 = ~n8787 ;
  assign y695 = n8793 ;
  assign y696 = ~n8809 ;
  assign y697 = n8812 ;
  assign y698 = ~n8816 ;
  assign y699 = ~n8819 ;
  assign y700 = n8826 ;
  assign y701 = n8832 ;
  assign y702 = n8841 ;
  assign y703 = n8847 ;
  assign y704 = ~n8850 ;
  assign y705 = ~n8862 ;
  assign y706 = n8872 ;
  assign y707 = n8874 ;
  assign y708 = n8887 ;
  assign y709 = ~n8888 ;
  assign y710 = ~n8893 ;
  assign y711 = ~n8894 ;
  assign y712 = n8897 ;
  assign y713 = ~n8909 ;
  assign y714 = n8916 ;
  assign y715 = n8927 ;
  assign y716 = ~n8937 ;
  assign y717 = n8961 ;
  assign y718 = n8964 ;
  assign y719 = n8971 ;
  assign y720 = n8973 ;
  assign y721 = n8976 ;
  assign y722 = n8978 ;
  assign y723 = n8979 ;
  assign y724 = ~n8991 ;
  assign y725 = n8993 ;
  assign y726 = ~n8995 ;
  assign y727 = n8999 ;
  assign y728 = ~n9002 ;
  assign y729 = n9018 ;
  assign y730 = n9023 ;
  assign y731 = n9027 ;
  assign y732 = ~n9030 ;
  assign y733 = n9036 ;
  assign y734 = n9037 ;
  assign y735 = ~n9042 ;
  assign y736 = n9049 ;
  assign y737 = ~n9061 ;
  assign y738 = ~n9071 ;
  assign y739 = n9083 ;
  assign y740 = ~n9084 ;
  assign y741 = n9086 ;
  assign y742 = ~n9088 ;
  assign y743 = n9111 ;
  assign y744 = ~n9118 ;
  assign y745 = ~n9123 ;
  assign y746 = n9140 ;
  assign y747 = ~n9142 ;
  assign y748 = ~n9147 ;
  assign y749 = n9154 ;
  assign y750 = n9159 ;
  assign y751 = ~n9167 ;
  assign y752 = n9171 ;
  assign y753 = n9197 ;
  assign y754 = ~n9202 ;
  assign y755 = ~n9210 ;
  assign y756 = n9214 ;
  assign y757 = n9231 ;
  assign y758 = n9233 ;
  assign y759 = n9240 ;
  assign y760 = n9246 ;
  assign y761 = n9247 ;
  assign y762 = ~n9250 ;
  assign y763 = ~n9254 ;
  assign y764 = n9258 ;
  assign y765 = ~n9260 ;
  assign y766 = ~n9272 ;
  assign y767 = n9276 ;
  assign y768 = n9279 ;
  assign y769 = n9284 ;
  assign y770 = n9286 ;
  assign y771 = ~n9290 ;
  assign y772 = n9296 ;
  assign y773 = n9305 ;
  assign y774 = n9309 ;
  assign y775 = n9311 ;
  assign y776 = ~n9313 ;
  assign y777 = n9317 ;
  assign y778 = n9320 ;
  assign y779 = n9327 ;
  assign y780 = n9331 ;
  assign y781 = n9337 ;
  assign y782 = n9338 ;
  assign y783 = n9342 ;
  assign y784 = n9350 ;
  assign y785 = ~n9361 ;
  assign y786 = n9372 ;
  assign y787 = n9375 ;
  assign y788 = ~n9378 ;
  assign y789 = ~n9379 ;
  assign y790 = ~n9382 ;
  assign y791 = n9385 ;
  assign y792 = n9390 ;
  assign y793 = n9395 ;
  assign y794 = ~n9409 ;
  assign y795 = n9417 ;
  assign y796 = ~n9427 ;
  assign y797 = n9429 ;
  assign y798 = ~n9448 ;
  assign y799 = n9450 ;
  assign y800 = n9457 ;
  assign y801 = ~n9468 ;
  assign y802 = n9481 ;
  assign y803 = n9486 ;
  assign y804 = n9495 ;
  assign y805 = ~n9505 ;
  assign y806 = ~n9515 ;
  assign y807 = ~n9529 ;
  assign y808 = n9533 ;
  assign y809 = ~n9534 ;
  assign y810 = n9535 ;
  assign y811 = ~n9537 ;
  assign y812 = ~n9547 ;
  assign y813 = n9560 ;
  assign y814 = n9566 ;
  assign y815 = n9571 ;
  assign y816 = n9577 ;
  assign y817 = ~n9580 ;
  assign y818 = ~n9585 ;
  assign y819 = ~n9590 ;
  assign y820 = n9603 ;
  assign y821 = n9604 ;
  assign y822 = ~n9608 ;
  assign y823 = n9609 ;
  assign y824 = n9613 ;
  assign y825 = ~n9614 ;
  assign y826 = ~n9616 ;
  assign y827 = ~n9625 ;
  assign y828 = n9632 ;
  assign y829 = n9635 ;
  assign y830 = ~n9641 ;
  assign y831 = n9648 ;
  assign y832 = n9653 ;
  assign y833 = ~n9657 ;
  assign y834 = ~n9661 ;
  assign y835 = ~n9663 ;
  assign y836 = ~n9664 ;
  assign y837 = n9671 ;
  assign y838 = n9672 ;
  assign y839 = ~n9682 ;
  assign y840 = n9694 ;
  assign y841 = ~n9695 ;
  assign y842 = ~n9697 ;
  assign y843 = n9703 ;
  assign y844 = n9705 ;
  assign y845 = n9706 ;
  assign y846 = n9708 ;
  assign y847 = ~n9719 ;
  assign y848 = ~n9721 ;
  assign y849 = ~n9722 ;
  assign y850 = n9732 ;
  assign y851 = ~n9736 ;
  assign y852 = n9743 ;
  assign y853 = n9749 ;
  assign y854 = n9753 ;
  assign y855 = ~n9759 ;
  assign y856 = n9760 ;
  assign y857 = n9763 ;
  assign y858 = ~n9767 ;
  assign y859 = ~n9769 ;
  assign y860 = ~n9784 ;
  assign y861 = n9799 ;
  assign y862 = ~n9809 ;
  assign y863 = n9812 ;
  assign y864 = n9814 ;
  assign y865 = ~n9817 ;
  assign y866 = ~n9821 ;
  assign y867 = ~n9822 ;
  assign y868 = ~n9823 ;
  assign y869 = ~n9825 ;
  assign y870 = ~n9832 ;
  assign y871 = ~n9835 ;
  assign y872 = ~n9837 ;
  assign y873 = ~n9842 ;
  assign y874 = ~n9844 ;
  assign y875 = n9845 ;
  assign y876 = ~n9848 ;
  assign y877 = n9859 ;
  assign y878 = n9864 ;
  assign y879 = ~n9866 ;
  assign y880 = n9870 ;
  assign y881 = ~n9874 ;
  assign y882 = n9899 ;
  assign y883 = n9901 ;
  assign y884 = ~n9902 ;
  assign y885 = ~n9904 ;
  assign y886 = n9906 ;
  assign y887 = ~n9913 ;
  assign y888 = ~n9916 ;
  assign y889 = n9927 ;
  assign y890 = n9934 ;
  assign y891 = ~n9935 ;
  assign y892 = n9939 ;
  assign y893 = n9941 ;
  assign y894 = n9949 ;
  assign y895 = n9951 ;
  assign y896 = n9953 ;
  assign y897 = ~n9964 ;
  assign y898 = ~n9969 ;
  assign y899 = ~n9971 ;
  assign y900 = ~n9973 ;
  assign y901 = ~n9977 ;
  assign y902 = ~n9979 ;
  assign y903 = n9981 ;
  assign y904 = ~n9994 ;
  assign y905 = ~n9998 ;
  assign y906 = n10005 ;
  assign y907 = ~n10008 ;
  assign y908 = n10016 ;
  assign y909 = n10024 ;
  assign y910 = ~n10030 ;
  assign y911 = ~n10034 ;
  assign y912 = n10037 ;
  assign y913 = n10041 ;
  assign y914 = n10046 ;
  assign y915 = n10052 ;
  assign y916 = ~n10055 ;
  assign y917 = n10064 ;
  assign y918 = ~n10069 ;
  assign y919 = ~n10070 ;
  assign y920 = n10076 ;
  assign y921 = n10079 ;
  assign y922 = ~n10081 ;
  assign y923 = ~n10086 ;
  assign y924 = n10097 ;
  assign y925 = n10101 ;
  assign y926 = n10102 ;
  assign y927 = n10104 ;
  assign y928 = n10105 ;
  assign y929 = ~n10113 ;
  assign y930 = n10123 ;
  assign y931 = n10143 ;
  assign y932 = ~n10147 ;
  assign y933 = n10150 ;
  assign y934 = n10155 ;
  assign y935 = n10156 ;
  assign y936 = ~n10158 ;
  assign y937 = ~n10162 ;
  assign y938 = ~n10163 ;
  assign y939 = ~n10179 ;
  assign y940 = n10184 ;
  assign y941 = ~n10187 ;
  assign y942 = n10192 ;
  assign y943 = ~n10195 ;
  assign y944 = n10205 ;
  assign y945 = ~n10209 ;
  assign y946 = ~n10210 ;
  assign y947 = n10214 ;
  assign y948 = ~n10225 ;
  assign y949 = ~n10227 ;
  assign y950 = n10229 ;
  assign y951 = ~n10234 ;
  assign y952 = n10235 ;
  assign y953 = n10246 ;
  assign y954 = n10263 ;
  assign y955 = ~n10270 ;
  assign y956 = n10272 ;
  assign y957 = n10273 ;
  assign y958 = ~n10277 ;
  assign y959 = ~n10279 ;
  assign y960 = ~n10284 ;
  assign y961 = n10285 ;
  assign y962 = n10292 ;
  assign y963 = n10295 ;
  assign y964 = ~n10296 ;
  assign y965 = n10299 ;
  assign y966 = ~n10303 ;
  assign y967 = ~n10317 ;
  assign y968 = ~n10322 ;
  assign y969 = n10323 ;
  assign y970 = ~n10325 ;
  assign y971 = n10333 ;
  assign y972 = ~n10335 ;
  assign y973 = ~n10343 ;
  assign y974 = ~n10344 ;
  assign y975 = n10356 ;
  assign y976 = n10357 ;
  assign y977 = n10361 ;
  assign y978 = ~n10364 ;
  assign y979 = ~n10372 ;
  assign y980 = n10378 ;
  assign y981 = ~n10379 ;
  assign y982 = ~n10381 ;
  assign y983 = ~n10382 ;
  assign y984 = ~n10385 ;
  assign y985 = n10386 ;
  assign y986 = ~n10394 ;
  assign y987 = ~n10399 ;
  assign y988 = ~n10400 ;
  assign y989 = n10402 ;
  assign y990 = ~n10407 ;
  assign y991 = n10413 ;
  assign y992 = ~n10414 ;
  assign y993 = n10420 ;
  assign y994 = n10428 ;
  assign y995 = n10437 ;
  assign y996 = n10443 ;
  assign y997 = ~n10448 ;
  assign y998 = ~n10456 ;
  assign y999 = n10460 ;
  assign y1000 = n10481 ;
  assign y1001 = ~n10487 ;
  assign y1002 = ~n10490 ;
  assign y1003 = n10493 ;
  assign y1004 = n10494 ;
  assign y1005 = ~n10503 ;
  assign y1006 = n10509 ;
  assign y1007 = n10510 ;
  assign y1008 = n10514 ;
  assign y1009 = ~n10520 ;
  assign y1010 = ~n10524 ;
  assign y1011 = ~n10527 ;
  assign y1012 = n10530 ;
  assign y1013 = n10535 ;
  assign y1014 = n10536 ;
  assign y1015 = ~n10538 ;
  assign y1016 = ~n10540 ;
  assign y1017 = ~n10542 ;
  assign y1018 = n10544 ;
  assign y1019 = n10564 ;
  assign y1020 = n10565 ;
  assign y1021 = n10568 ;
  assign y1022 = ~n10576 ;
  assign y1023 = n10577 ;
  assign y1024 = n10585 ;
  assign y1025 = n10592 ;
  assign y1026 = ~n10593 ;
  assign y1027 = ~n10595 ;
  assign y1028 = ~n10600 ;
  assign y1029 = n10604 ;
  assign y1030 = ~n10610 ;
  assign y1031 = ~n10612 ;
  assign y1032 = n10616 ;
  assign y1033 = n10625 ;
  assign y1034 = n10637 ;
  assign y1035 = n10642 ;
  assign y1036 = ~n10646 ;
  assign y1037 = n10656 ;
  assign y1038 = n10672 ;
  assign y1039 = ~n10675 ;
  assign y1040 = n10681 ;
  assign y1041 = ~n10686 ;
  assign y1042 = ~n10689 ;
  assign y1043 = ~n10702 ;
  assign y1044 = ~n10703 ;
  assign y1045 = ~n10705 ;
  assign y1046 = ~n10711 ;
  assign y1047 = n10718 ;
  assign y1048 = n10722 ;
  assign y1049 = ~n10729 ;
  assign y1050 = ~n10730 ;
  assign y1051 = ~n10733 ;
  assign y1052 = ~n10746 ;
  assign y1053 = n10748 ;
  assign y1054 = ~n10751 ;
  assign y1055 = ~n10752 ;
  assign y1056 = n10757 ;
  assign y1057 = n10761 ;
  assign y1058 = ~n10766 ;
  assign y1059 = n10767 ;
  assign y1060 = ~n10770 ;
  assign y1061 = n10776 ;
  assign y1062 = ~n10784 ;
  assign y1063 = n10785 ;
  assign y1064 = ~n10798 ;
  assign y1065 = n10799 ;
  assign y1066 = ~n10805 ;
  assign y1067 = n10812 ;
  assign y1068 = n10815 ;
  assign y1069 = ~n10817 ;
  assign y1070 = ~n10820 ;
  assign y1071 = n10822 ;
  assign y1072 = ~n10824 ;
  assign y1073 = n10826 ;
  assign y1074 = n10833 ;
  assign y1075 = ~n10834 ;
  assign y1076 = n10835 ;
  assign y1077 = ~n10854 ;
  assign y1078 = n10860 ;
  assign y1079 = n10865 ;
  assign y1080 = n10871 ;
  assign y1081 = n10873 ;
  assign y1082 = ~n10883 ;
  assign y1083 = n10888 ;
  assign y1084 = ~n10894 ;
  assign y1085 = n10896 ;
  assign y1086 = n10898 ;
  assign y1087 = ~n10899 ;
  assign y1088 = n10907 ;
  assign y1089 = n10918 ;
  assign y1090 = ~n10919 ;
  assign y1091 = n10921 ;
  assign y1092 = n10924 ;
  assign y1093 = n10928 ;
  assign y1094 = n10929 ;
  assign y1095 = ~n10930 ;
  assign y1096 = n10932 ;
  assign y1097 = n10935 ;
  assign y1098 = n10939 ;
  assign y1099 = ~n10942 ;
  assign y1100 = ~n10947 ;
  assign y1101 = ~n10951 ;
  assign y1102 = n10953 ;
  assign y1103 = ~n10955 ;
  assign y1104 = ~n10968 ;
  assign y1105 = n10975 ;
  assign y1106 = ~n10981 ;
  assign y1107 = ~n10982 ;
  assign y1108 = ~n10987 ;
  assign y1109 = ~n10990 ;
  assign y1110 = ~n11009 ;
  assign y1111 = ~n11014 ;
  assign y1112 = ~n11018 ;
  assign y1113 = ~n11024 ;
  assign y1114 = ~n11028 ;
  assign y1115 = ~n11030 ;
  assign y1116 = ~n11039 ;
  assign y1117 = ~n11048 ;
  assign y1118 = ~n11058 ;
  assign y1119 = n11063 ;
  assign y1120 = n11065 ;
  assign y1121 = ~n11076 ;
  assign y1122 = n11083 ;
  assign y1123 = ~n11086 ;
  assign y1124 = n11090 ;
  assign y1125 = ~n11095 ;
  assign y1126 = n11100 ;
  assign y1127 = n11102 ;
  assign y1128 = n11105 ;
  assign y1129 = ~n11108 ;
  assign y1130 = n11116 ;
  assign y1131 = n11121 ;
  assign y1132 = n11128 ;
  assign y1133 = n11132 ;
  assign y1134 = ~n11133 ;
  assign y1135 = ~n11138 ;
  assign y1136 = n11140 ;
  assign y1137 = n11144 ;
  assign y1138 = ~n11147 ;
  assign y1139 = n11149 ;
  assign y1140 = ~n11160 ;
  assign y1141 = n11163 ;
  assign y1142 = ~n11165 ;
  assign y1143 = n11180 ;
  assign y1144 = n11184 ;
  assign y1145 = n11190 ;
  assign y1146 = ~n11194 ;
  assign y1147 = n11198 ;
  assign y1148 = n11199 ;
  assign y1149 = n11203 ;
  assign y1150 = ~n11206 ;
  assign y1151 = ~n11219 ;
  assign y1152 = n11221 ;
  assign y1153 = n11226 ;
  assign y1154 = n11227 ;
  assign y1155 = n11229 ;
  assign y1156 = ~n11233 ;
  assign y1157 = n11236 ;
  assign y1158 = ~n11249 ;
  assign y1159 = n11254 ;
  assign y1160 = n11261 ;
  assign y1161 = ~n11265 ;
  assign y1162 = ~n11269 ;
  assign y1163 = ~n11274 ;
  assign y1164 = n11277 ;
  assign y1165 = ~n11289 ;
  assign y1166 = n11295 ;
  assign y1167 = ~n11296 ;
  assign y1168 = ~n11305 ;
  assign y1169 = n11312 ;
  assign y1170 = ~n11316 ;
  assign y1171 = n11322 ;
  assign y1172 = ~n11324 ;
  assign y1173 = n11325 ;
  assign y1174 = ~n11332 ;
  assign y1175 = ~n11333 ;
  assign y1176 = n11337 ;
  assign y1177 = ~n11341 ;
  assign y1178 = ~n11345 ;
  assign y1179 = ~n11349 ;
  assign y1180 = n11360 ;
  assign y1181 = ~n11361 ;
  assign y1182 = ~n11368 ;
  assign y1183 = ~n11375 ;
  assign y1184 = n11379 ;
  assign y1185 = n11385 ;
  assign y1186 = ~n11386 ;
  assign y1187 = ~n11388 ;
  assign y1188 = ~n11397 ;
  assign y1189 = ~n11399 ;
  assign y1190 = n11403 ;
  assign y1191 = n11405 ;
  assign y1192 = n11417 ;
  assign y1193 = ~n11421 ;
  assign y1194 = n11435 ;
  assign y1195 = n11436 ;
  assign y1196 = n11440 ;
  assign y1197 = ~n11446 ;
  assign y1198 = n11453 ;
  assign y1199 = n11458 ;
  assign y1200 = ~n11460 ;
  assign y1201 = n11463 ;
  assign y1202 = ~n11471 ;
  assign y1203 = n11474 ;
  assign y1204 = n11483 ;
  assign y1205 = ~n11492 ;
  assign y1206 = n11497 ;
  assign y1207 = n11500 ;
  assign y1208 = n11502 ;
  assign y1209 = ~n11508 ;
  assign y1210 = ~n11512 ;
  assign y1211 = ~n11517 ;
  assign y1212 = n11518 ;
  assign y1213 = ~n11521 ;
  assign y1214 = ~n11526 ;
  assign y1215 = ~n11532 ;
  assign y1216 = ~n11537 ;
  assign y1217 = n11539 ;
  assign y1218 = n11540 ;
  assign y1219 = n11543 ;
  assign y1220 = n11550 ;
  assign y1221 = n11553 ;
  assign y1222 = n11555 ;
  assign y1223 = ~n11558 ;
  assign y1224 = ~n11559 ;
  assign y1225 = n11561 ;
  assign y1226 = ~n11566 ;
  assign y1227 = ~n11573 ;
  assign y1228 = ~n11576 ;
  assign y1229 = n11579 ;
  assign y1230 = n11585 ;
  assign y1231 = n11590 ;
  assign y1232 = n11592 ;
  assign y1233 = ~n11593 ;
  assign y1234 = ~n11595 ;
  assign y1235 = n11601 ;
  assign y1236 = ~n11606 ;
  assign y1237 = n11609 ;
  assign y1238 = n11611 ;
  assign y1239 = n11614 ;
  assign y1240 = n11617 ;
  assign y1241 = n11620 ;
  assign y1242 = n11625 ;
  assign y1243 = ~n11627 ;
  assign y1244 = ~n11628 ;
  assign y1245 = n11631 ;
  assign y1246 = n11633 ;
  assign y1247 = n11643 ;
  assign y1248 = ~n11647 ;
  assign y1249 = n11651 ;
  assign y1250 = ~n11656 ;
  assign y1251 = ~n11659 ;
  assign y1252 = n11671 ;
  assign y1253 = ~n11674 ;
  assign y1254 = ~n11682 ;
  assign y1255 = ~n11683 ;
  assign y1256 = n11685 ;
  assign y1257 = ~n11687 ;
  assign y1258 = n11688 ;
  assign y1259 = ~n11690 ;
  assign y1260 = n11709 ;
  assign y1261 = ~n11713 ;
  assign y1262 = n11724 ;
  assign y1263 = ~n11730 ;
  assign y1264 = ~n11734 ;
  assign y1265 = n11739 ;
  assign y1266 = n11748 ;
  assign y1267 = ~n11751 ;
  assign y1268 = ~n11752 ;
  assign y1269 = n11755 ;
  assign y1270 = n11756 ;
  assign y1271 = ~n11757 ;
  assign y1272 = ~n11759 ;
  assign y1273 = ~n11766 ;
  assign y1274 = ~n11775 ;
  assign y1275 = n11781 ;
  assign y1276 = n11788 ;
  assign y1277 = ~n11792 ;
  assign y1278 = ~n11801 ;
  assign y1279 = n11803 ;
  assign y1280 = n11804 ;
  assign y1281 = n11807 ;
  assign y1282 = ~n11810 ;
  assign y1283 = n11812 ;
  assign y1284 = n11814 ;
  assign y1285 = n11816 ;
  assign y1286 = ~n11818 ;
  assign y1287 = ~n11827 ;
  assign y1288 = ~n11832 ;
  assign y1289 = n11833 ;
  assign y1290 = n11839 ;
  assign y1291 = ~n11841 ;
  assign y1292 = n11850 ;
  assign y1293 = ~n11857 ;
  assign y1294 = ~n11861 ;
  assign y1295 = n11863 ;
  assign y1296 = n11865 ;
  assign y1297 = ~n11868 ;
  assign y1298 = ~n11874 ;
  assign y1299 = ~n11877 ;
  assign y1300 = ~n11880 ;
  assign y1301 = ~n11892 ;
  assign y1302 = ~n11900 ;
  assign y1303 = n11902 ;
  assign y1304 = ~n11905 ;
  assign y1305 = n11912 ;
  assign y1306 = ~n11918 ;
  assign y1307 = n11929 ;
  assign y1308 = n11930 ;
  assign y1309 = n11938 ;
  assign y1310 = ~n11943 ;
  assign y1311 = n11951 ;
  assign y1312 = ~n11954 ;
  assign y1313 = n11959 ;
  assign y1314 = n11962 ;
  assign y1315 = n11966 ;
  assign y1316 = n11968 ;
  assign y1317 = ~n11971 ;
  assign y1318 = n11977 ;
  assign y1319 = n11979 ;
  assign y1320 = ~n11989 ;
  assign y1321 = ~n11991 ;
  assign y1322 = ~n11992 ;
  assign y1323 = n12003 ;
  assign y1324 = ~n12006 ;
  assign y1325 = ~n12007 ;
  assign y1326 = n12009 ;
  assign y1327 = n12014 ;
  assign y1328 = n12021 ;
  assign y1329 = n12023 ;
  assign y1330 = ~n12027 ;
  assign y1331 = n12031 ;
  assign y1332 = ~n12032 ;
  assign y1333 = n12035 ;
  assign y1334 = ~n12041 ;
  assign y1335 = ~n12043 ;
  assign y1336 = n12048 ;
  assign y1337 = n12049 ;
  assign y1338 = n12057 ;
  assign y1339 = ~n12060 ;
  assign y1340 = n12069 ;
  assign y1341 = ~n12073 ;
  assign y1342 = ~n12075 ;
  assign y1343 = n12080 ;
  assign y1344 = ~n12081 ;
  assign y1345 = ~n12085 ;
  assign y1346 = ~n12086 ;
  assign y1347 = ~n12092 ;
  assign y1348 = n12093 ;
  assign y1349 = ~n12111 ;
  assign y1350 = n12113 ;
  assign y1351 = n12117 ;
  assign y1352 = n12120 ;
  assign y1353 = ~n12124 ;
  assign y1354 = n12127 ;
  assign y1355 = ~n12128 ;
  assign y1356 = n12129 ;
  assign y1357 = n12141 ;
  assign y1358 = ~n12144 ;
  assign y1359 = ~n12152 ;
  assign y1360 = ~n12157 ;
  assign y1361 = n12161 ;
  assign y1362 = ~n12166 ;
  assign y1363 = n12169 ;
  assign y1364 = n12175 ;
  assign y1365 = ~n12176 ;
  assign y1366 = n12188 ;
  assign y1367 = n12189 ;
  assign y1368 = n12191 ;
  assign y1369 = ~n12198 ;
  assign y1370 = ~n12199 ;
  assign y1371 = ~n12200 ;
  assign y1372 = n12201 ;
  assign y1373 = ~n12202 ;
  assign y1374 = ~n12207 ;
  assign y1375 = ~n12208 ;
  assign y1376 = n12209 ;
  assign y1377 = n12212 ;
  assign y1378 = ~n12220 ;
  assign y1379 = ~n12223 ;
  assign y1380 = n12227 ;
  assign y1381 = n12230 ;
  assign y1382 = ~n12237 ;
  assign y1383 = n12246 ;
  assign y1384 = n12252 ;
  assign y1385 = ~n12255 ;
  assign y1386 = n12259 ;
  assign y1387 = n12262 ;
  assign y1388 = n12266 ;
  assign y1389 = ~n12268 ;
  assign y1390 = n12272 ;
  assign y1391 = ~n12273 ;
  assign y1392 = ~n12280 ;
  assign y1393 = n12283 ;
  assign y1394 = ~n12290 ;
  assign y1395 = n12298 ;
  assign y1396 = ~n12299 ;
  assign y1397 = ~n12304 ;
  assign y1398 = n12313 ;
  assign y1399 = n12315 ;
  assign y1400 = n12319 ;
  assign y1401 = ~n12322 ;
  assign y1402 = ~n12327 ;
  assign y1403 = n12328 ;
  assign y1404 = n12336 ;
  assign y1405 = ~n12359 ;
  assign y1406 = n12361 ;
  assign y1407 = ~n12362 ;
  assign y1408 = n12363 ;
  assign y1409 = n12369 ;
  assign y1410 = n12375 ;
  assign y1411 = ~n12378 ;
  assign y1412 = ~n12380 ;
  assign y1413 = ~n12381 ;
  assign y1414 = n12382 ;
  assign y1415 = ~n12389 ;
  assign y1416 = ~n12393 ;
  assign y1417 = n12395 ;
  assign y1418 = n12398 ;
  assign y1419 = ~n12403 ;
  assign y1420 = ~n12409 ;
  assign y1421 = n12411 ;
  assign y1422 = n12412 ;
  assign y1423 = n12413 ;
  assign y1424 = n12417 ;
  assign y1425 = ~n12418 ;
  assign y1426 = ~n12423 ;
  assign y1427 = ~n12425 ;
  assign y1428 = n12434 ;
  assign y1429 = ~n12437 ;
  assign y1430 = ~n12445 ;
  assign y1431 = n12451 ;
  assign y1432 = ~n12452 ;
  assign y1433 = ~n12455 ;
  assign y1434 = ~n12459 ;
  assign y1435 = n12460 ;
  assign y1436 = ~n12462 ;
  assign y1437 = ~n12467 ;
  assign y1438 = n12472 ;
  assign y1439 = ~n12484 ;
  assign y1440 = ~n12486 ;
  assign y1441 = ~n12489 ;
  assign y1442 = ~n12500 ;
  assign y1443 = ~n12501 ;
  assign y1444 = ~n12502 ;
  assign y1445 = n12505 ;
  assign y1446 = ~n12510 ;
  assign y1447 = n12512 ;
  assign y1448 = ~n12515 ;
  assign y1449 = ~n12519 ;
  assign y1450 = ~n12520 ;
  assign y1451 = n12521 ;
  assign y1452 = ~n12525 ;
  assign y1453 = n12539 ;
  assign y1454 = n12543 ;
  assign y1455 = n12550 ;
  assign y1456 = ~n12551 ;
  assign y1457 = ~n12554 ;
  assign y1458 = n12561 ;
  assign y1459 = n12567 ;
  assign y1460 = ~n12579 ;
  assign y1461 = n12584 ;
  assign y1462 = ~n12592 ;
  assign y1463 = n12593 ;
  assign y1464 = ~n12594 ;
  assign y1465 = n12598 ;
  assign y1466 = ~n12599 ;
  assign y1467 = ~n12607 ;
  assign y1468 = n12611 ;
  assign y1469 = n12614 ;
  assign y1470 = ~n12618 ;
  assign y1471 = n12619 ;
  assign y1472 = ~n12622 ;
  assign y1473 = ~n12633 ;
  assign y1474 = n12641 ;
  assign y1475 = ~n12646 ;
  assign y1476 = ~n12650 ;
  assign y1477 = ~n12653 ;
  assign y1478 = n12655 ;
  assign y1479 = ~n12669 ;
  assign y1480 = ~n12673 ;
  assign y1481 = n12674 ;
  assign y1482 = n12679 ;
  assign y1483 = n12681 ;
  assign y1484 = ~n12685 ;
  assign y1485 = n12687 ;
  assign y1486 = ~n12689 ;
  assign y1487 = ~n12695 ;
  assign y1488 = ~n12696 ;
  assign y1489 = ~n12697 ;
  assign y1490 = ~n12700 ;
  assign y1491 = n12702 ;
  assign y1492 = n12703 ;
  assign y1493 = n12706 ;
  assign y1494 = n12707 ;
  assign y1495 = n12711 ;
  assign y1496 = n12722 ;
  assign y1497 = n12724 ;
  assign y1498 = n12727 ;
  assign y1499 = n12729 ;
  assign y1500 = ~n12731 ;
  assign y1501 = ~n12735 ;
  assign y1502 = n12737 ;
  assign y1503 = n12741 ;
  assign y1504 = ~n12747 ;
  assign y1505 = n12753 ;
  assign y1506 = n12757 ;
  assign y1507 = ~n12758 ;
  assign y1508 = n12761 ;
  assign y1509 = n12762 ;
  assign y1510 = n12770 ;
  assign y1511 = ~n12772 ;
  assign y1512 = ~n12775 ;
  assign y1513 = n12776 ;
  assign y1514 = n12778 ;
  assign y1515 = ~n12782 ;
  assign y1516 = ~n12786 ;
  assign y1517 = ~n12791 ;
  assign y1518 = ~n12793 ;
  assign y1519 = n12803 ;
  assign y1520 = ~n12809 ;
  assign y1521 = n12812 ;
  assign y1522 = ~n12822 ;
  assign y1523 = n12827 ;
  assign y1524 = n12842 ;
  assign y1525 = n12851 ;
  assign y1526 = n12855 ;
  assign y1527 = n12857 ;
  assign y1528 = n12858 ;
  assign y1529 = n12861 ;
  assign y1530 = ~n12865 ;
  assign y1531 = ~n12871 ;
  assign y1532 = ~n12872 ;
  assign y1533 = n12884 ;
  assign y1534 = ~n12886 ;
  assign y1535 = ~n12891 ;
  assign y1536 = n12893 ;
  assign y1537 = ~n12898 ;
  assign y1538 = n12912 ;
  assign y1539 = ~n12914 ;
  assign y1540 = ~n12917 ;
  assign y1541 = n12923 ;
  assign y1542 = n12928 ;
  assign y1543 = n12931 ;
  assign y1544 = ~n12938 ;
  assign y1545 = n12940 ;
  assign y1546 = ~n12946 ;
  assign y1547 = n12948 ;
  assign y1548 = ~n12952 ;
  assign y1549 = n12956 ;
  assign y1550 = ~n12957 ;
  assign y1551 = n12960 ;
  assign y1552 = ~n12969 ;
  assign y1553 = ~n12980 ;
  assign y1554 = n12983 ;
  assign y1555 = ~n12985 ;
  assign y1556 = ~n12990 ;
  assign y1557 = n12991 ;
  assign y1558 = n12993 ;
  assign y1559 = ~n12996 ;
  assign y1560 = ~n12997 ;
  assign y1561 = n13002 ;
  assign y1562 = n13003 ;
  assign y1563 = n13011 ;
  assign y1564 = n13014 ;
  assign y1565 = n13028 ;
  assign y1566 = ~n13034 ;
  assign y1567 = n13038 ;
  assign y1568 = n13040 ;
  assign y1569 = ~n13047 ;
  assign y1570 = n13050 ;
  assign y1571 = n13052 ;
  assign y1572 = n13056 ;
  assign y1573 = n13060 ;
  assign y1574 = n13071 ;
  assign y1575 = n13076 ;
  assign y1576 = n13079 ;
  assign y1577 = n13084 ;
  assign y1578 = ~n13086 ;
  assign y1579 = ~n13090 ;
  assign y1580 = n13097 ;
  assign y1581 = ~n13108 ;
  assign y1582 = n13110 ;
  assign y1583 = ~n13112 ;
  assign y1584 = ~n13117 ;
  assign y1585 = n13121 ;
  assign y1586 = n13122 ;
  assign y1587 = ~n13126 ;
  assign y1588 = n13128 ;
  assign y1589 = n13131 ;
  assign y1590 = n13144 ;
  assign y1591 = n13147 ;
  assign y1592 = n13148 ;
  assign y1593 = n13157 ;
  assign y1594 = n13158 ;
  assign y1595 = n13162 ;
  assign y1596 = n13164 ;
  assign y1597 = n13166 ;
  assign y1598 = n13167 ;
  assign y1599 = ~n13176 ;
  assign y1600 = ~n13179 ;
  assign y1601 = ~n13181 ;
  assign y1602 = ~n13182 ;
  assign y1603 = n13186 ;
  assign y1604 = ~n13192 ;
  assign y1605 = n13193 ;
  assign y1606 = ~n13196 ;
  assign y1607 = n13199 ;
  assign y1608 = ~n13200 ;
  assign y1609 = n13202 ;
  assign y1610 = ~n13210 ;
  assign y1611 = n13213 ;
  assign y1612 = n13217 ;
  assign y1613 = ~n13222 ;
  assign y1614 = n13230 ;
  assign y1615 = ~n13231 ;
  assign y1616 = ~n13235 ;
  assign y1617 = n13240 ;
  assign y1618 = ~n13242 ;
  assign y1619 = n13247 ;
  assign y1620 = ~n13248 ;
  assign y1621 = n13252 ;
  assign y1622 = ~n13254 ;
  assign y1623 = n13257 ;
  assign y1624 = n13260 ;
  assign y1625 = ~n13263 ;
  assign y1626 = n13266 ;
  assign y1627 = ~n13267 ;
  assign y1628 = ~n13275 ;
  assign y1629 = ~n13278 ;
  assign y1630 = n13281 ;
  assign y1631 = n13290 ;
  assign y1632 = ~n13294 ;
  assign y1633 = ~n13295 ;
  assign y1634 = n13297 ;
  assign y1635 = ~n13299 ;
  assign y1636 = n13300 ;
  assign y1637 = n13303 ;
  assign y1638 = ~n13308 ;
  assign y1639 = ~n13309 ;
  assign y1640 = n13313 ;
  assign y1641 = ~n13317 ;
  assign y1642 = ~n13319 ;
  assign y1643 = ~n13320 ;
  assign y1644 = ~n13321 ;
  assign y1645 = n13326 ;
  assign y1646 = n13331 ;
  assign y1647 = ~n13335 ;
  assign y1648 = n13337 ;
  assign y1649 = ~n13342 ;
  assign y1650 = ~n13343 ;
  assign y1651 = ~n13345 ;
  assign y1652 = ~n13349 ;
  assign y1653 = n13351 ;
  assign y1654 = n13354 ;
  assign y1655 = n13359 ;
  assign y1656 = ~n13362 ;
  assign y1657 = n13364 ;
  assign y1658 = n13374 ;
  assign y1659 = ~n13377 ;
  assign y1660 = ~n13385 ;
  assign y1661 = ~n13393 ;
  assign y1662 = n13395 ;
  assign y1663 = n13397 ;
  assign y1664 = ~n13399 ;
  assign y1665 = n13407 ;
  assign y1666 = n13415 ;
  assign y1667 = ~n13427 ;
  assign y1668 = n13428 ;
  assign y1669 = n13431 ;
  assign y1670 = n13435 ;
  assign y1671 = ~n13438 ;
  assign y1672 = n13441 ;
  assign y1673 = ~n13442 ;
  assign y1674 = n13443 ;
  assign y1675 = n13452 ;
  assign y1676 = ~n13453 ;
  assign y1677 = n13458 ;
  assign y1678 = n13460 ;
  assign y1679 = ~n13462 ;
  assign y1680 = n13464 ;
  assign y1681 = n13471 ;
  assign y1682 = n13473 ;
  assign y1683 = ~n13487 ;
  assign y1684 = ~n13489 ;
  assign y1685 = n13497 ;
  assign y1686 = n13500 ;
  assign y1687 = ~n13502 ;
  assign y1688 = ~n13509 ;
  assign y1689 = n13513 ;
  assign y1690 = ~n13517 ;
  assign y1691 = ~n13520 ;
  assign y1692 = n13526 ;
  assign y1693 = ~n13528 ;
  assign y1694 = n13530 ;
  assign y1695 = n13535 ;
  assign y1696 = ~n13539 ;
  assign y1697 = n13542 ;
  assign y1698 = ~n13545 ;
  assign y1699 = ~n13547 ;
  assign y1700 = ~n13549 ;
  assign y1701 = n13551 ;
  assign y1702 = ~n13557 ;
  assign y1703 = ~n13562 ;
  assign y1704 = ~n13570 ;
  assign y1705 = n13573 ;
  assign y1706 = n13574 ;
  assign y1707 = n13581 ;
  assign y1708 = n13582 ;
  assign y1709 = n13584 ;
  assign y1710 = n13594 ;
  assign y1711 = ~n13597 ;
  assign y1712 = n13600 ;
  assign y1713 = n13602 ;
  assign y1714 = ~n13603 ;
  assign y1715 = ~n13604 ;
  assign y1716 = ~n13613 ;
  assign y1717 = ~n13616 ;
  assign y1718 = n13622 ;
  assign y1719 = n13623 ;
  assign y1720 = ~n13624 ;
  assign y1721 = ~n13625 ;
  assign y1722 = n13628 ;
  assign y1723 = ~n13637 ;
  assign y1724 = ~n13639 ;
  assign y1725 = n13643 ;
  assign y1726 = ~n13650 ;
  assign y1727 = n13652 ;
  assign y1728 = ~n13657 ;
  assign y1729 = ~n13664 ;
  assign y1730 = n13665 ;
  assign y1731 = ~n13672 ;
  assign y1732 = ~n13673 ;
  assign y1733 = n13676 ;
  assign y1734 = n13679 ;
  assign y1735 = n13693 ;
  assign y1736 = n13696 ;
  assign y1737 = n13699 ;
  assign y1738 = ~n13702 ;
  assign y1739 = n13709 ;
  assign y1740 = ~n13712 ;
  assign y1741 = n13716 ;
  assign y1742 = ~n13718 ;
  assign y1743 = n13721 ;
  assign y1744 = ~n13725 ;
  assign y1745 = n13727 ;
  assign y1746 = ~n13733 ;
  assign y1747 = n13736 ;
  assign y1748 = ~n13738 ;
  assign y1749 = n13746 ;
  assign y1750 = n13747 ;
  assign y1751 = ~n13752 ;
  assign y1752 = n13753 ;
  assign y1753 = n13754 ;
  assign y1754 = n13760 ;
  assign y1755 = n13763 ;
  assign y1756 = ~n13767 ;
  assign y1757 = n13768 ;
  assign y1758 = ~n13772 ;
  assign y1759 = ~n13783 ;
  assign y1760 = ~n13788 ;
  assign y1761 = n13792 ;
  assign y1762 = n13794 ;
  assign y1763 = n13800 ;
  assign y1764 = n13802 ;
  assign y1765 = n13805 ;
  assign y1766 = n13810 ;
  assign y1767 = n13824 ;
  assign y1768 = ~n13830 ;
  assign y1769 = n13837 ;
  assign y1770 = n13840 ;
  assign y1771 = ~n13845 ;
  assign y1772 = n13847 ;
  assign y1773 = n13849 ;
  assign y1774 = ~n13854 ;
  assign y1775 = ~n13856 ;
  assign y1776 = n13858 ;
  assign y1777 = n13860 ;
  assign y1778 = n13865 ;
  assign y1779 = n13877 ;
  assign y1780 = n13878 ;
  assign y1781 = n13879 ;
  assign y1782 = ~n13883 ;
  assign y1783 = n13890 ;
  assign y1784 = ~n13892 ;
  assign y1785 = n13895 ;
  assign y1786 = ~n13899 ;
  assign y1787 = n13905 ;
  assign y1788 = n13906 ;
  assign y1789 = ~n13907 ;
  assign y1790 = ~n13911 ;
  assign y1791 = n13919 ;
  assign y1792 = n13921 ;
  assign y1793 = n13924 ;
  assign y1794 = ~n13929 ;
  assign y1795 = n13936 ;
  assign y1796 = ~n13949 ;
  assign y1797 = ~n13950 ;
  assign y1798 = n13954 ;
  assign y1799 = n13957 ;
  assign y1800 = n13958 ;
  assign y1801 = ~n13963 ;
  assign y1802 = ~n13964 ;
  assign y1803 = n13967 ;
  assign y1804 = n13968 ;
  assign y1805 = n13970 ;
  assign y1806 = n13971 ;
  assign y1807 = ~n13979 ;
  assign y1808 = ~n13981 ;
  assign y1809 = n13988 ;
  assign y1810 = n13992 ;
  assign y1811 = ~n13995 ;
  assign y1812 = n14010 ;
  assign y1813 = n14013 ;
  assign y1814 = n14014 ;
  assign y1815 = n14017 ;
  assign y1816 = ~n14030 ;
  assign y1817 = ~n14032 ;
  assign y1818 = n14038 ;
  assign y1819 = n14040 ;
  assign y1820 = ~n14046 ;
  assign y1821 = n14048 ;
  assign y1822 = n14056 ;
  assign y1823 = ~n14057 ;
  assign y1824 = ~n14060 ;
  assign y1825 = ~n14065 ;
  assign y1826 = n14072 ;
  assign y1827 = n14076 ;
  assign y1828 = n14078 ;
  assign y1829 = n14080 ;
  assign y1830 = n14082 ;
  assign y1831 = n14083 ;
  assign y1832 = n14084 ;
  assign y1833 = n14088 ;
  assign y1834 = ~n14093 ;
  assign y1835 = n14100 ;
  assign y1836 = ~n14112 ;
  assign y1837 = ~n14115 ;
  assign y1838 = ~n14120 ;
  assign y1839 = ~n14123 ;
  assign y1840 = ~n14125 ;
  assign y1841 = ~n14130 ;
  assign y1842 = n14135 ;
  assign y1843 = n14145 ;
  assign y1844 = ~n14155 ;
  assign y1845 = ~n14157 ;
  assign y1846 = ~n14158 ;
  assign y1847 = ~n14162 ;
  assign y1848 = ~n14170 ;
  assign y1849 = ~n14172 ;
  assign y1850 = n14176 ;
  assign y1851 = n14178 ;
  assign y1852 = n14182 ;
  assign y1853 = ~n14185 ;
  assign y1854 = n14192 ;
  assign y1855 = ~n14193 ;
  assign y1856 = ~n14194 ;
  assign y1857 = ~n14207 ;
  assign y1858 = ~n14208 ;
  assign y1859 = n14213 ;
  assign y1860 = ~n14219 ;
  assign y1861 = n14221 ;
  assign y1862 = n14222 ;
  assign y1863 = n14223 ;
  assign y1864 = ~n14225 ;
  assign y1865 = ~n14228 ;
  assign y1866 = n14229 ;
  assign y1867 = ~n14231 ;
  assign y1868 = ~n14233 ;
  assign y1869 = ~n14236 ;
  assign y1870 = ~n14238 ;
  assign y1871 = n14241 ;
  assign y1872 = n14245 ;
  assign y1873 = n14247 ;
  assign y1874 = n14249 ;
  assign y1875 = n14253 ;
  assign y1876 = n14256 ;
  assign y1877 = ~n14258 ;
  assign y1878 = n14259 ;
  assign y1879 = ~n14260 ;
  assign y1880 = ~n14261 ;
  assign y1881 = ~n14270 ;
  assign y1882 = n14272 ;
  assign y1883 = n14275 ;
  assign y1884 = ~n14281 ;
  assign y1885 = n14287 ;
  assign y1886 = n14291 ;
  assign y1887 = n14295 ;
  assign y1888 = n14299 ;
  assign y1889 = n14302 ;
  assign y1890 = n14303 ;
  assign y1891 = n14309 ;
  assign y1892 = n14315 ;
  assign y1893 = n14316 ;
  assign y1894 = n14317 ;
  assign y1895 = ~n14318 ;
  assign y1896 = ~n14321 ;
  assign y1897 = ~n14341 ;
  assign y1898 = ~n14342 ;
  assign y1899 = n14345 ;
  assign y1900 = n14346 ;
  assign y1901 = ~n14347 ;
  assign y1902 = n14348 ;
  assign y1903 = n14352 ;
  assign y1904 = n14355 ;
  assign y1905 = ~n14361 ;
  assign y1906 = ~n14372 ;
  assign y1907 = n14375 ;
  assign y1908 = n14376 ;
  assign y1909 = ~n14383 ;
  assign y1910 = n14385 ;
  assign y1911 = ~n14388 ;
  assign y1912 = n14393 ;
  assign y1913 = n14394 ;
  assign y1914 = ~n14395 ;
  assign y1915 = n14402 ;
  assign y1916 = n14403 ;
  assign y1917 = n14406 ;
  assign y1918 = n14409 ;
  assign y1919 = n14410 ;
  assign y1920 = n14415 ;
  assign y1921 = ~n14417 ;
  assign y1922 = ~n14418 ;
  assign y1923 = n14421 ;
  assign y1924 = ~n14427 ;
  assign y1925 = n14428 ;
  assign y1926 = ~n14430 ;
  assign y1927 = ~n14434 ;
  assign y1928 = ~n14442 ;
  assign y1929 = ~n14444 ;
  assign y1930 = n14447 ;
  assign y1931 = n14450 ;
  assign y1932 = n14453 ;
  assign y1933 = ~n14457 ;
  assign y1934 = ~n14458 ;
  assign y1935 = ~n14461 ;
  assign y1936 = ~n14462 ;
  assign y1937 = n14465 ;
  assign y1938 = ~n14466 ;
  assign y1939 = ~n14468 ;
  assign y1940 = ~n14470 ;
  assign y1941 = n14473 ;
  assign y1942 = n14479 ;
  assign y1943 = n14481 ;
  assign y1944 = ~n14483 ;
  assign y1945 = n14486 ;
  assign y1946 = n14490 ;
  assign y1947 = ~n14493 ;
  assign y1948 = n14497 ;
  assign y1949 = ~n14500 ;
  assign y1950 = ~n14512 ;
  assign y1951 = ~n14515 ;
  assign y1952 = ~n14521 ;
  assign y1953 = ~n14525 ;
  assign y1954 = ~n14531 ;
  assign y1955 = ~n14533 ;
  assign y1956 = n14540 ;
  assign y1957 = ~n14546 ;
  assign y1958 = n14551 ;
  assign y1959 = n14557 ;
  assign y1960 = n14560 ;
  assign y1961 = ~n14564 ;
  assign y1962 = ~n14569 ;
  assign y1963 = ~n14572 ;
  assign y1964 = ~n14574 ;
  assign y1965 = ~n14576 ;
  assign y1966 = n14582 ;
  assign y1967 = n14586 ;
  assign y1968 = n14588 ;
  assign y1969 = n14592 ;
  assign y1970 = n14598 ;
  assign y1971 = ~n14601 ;
  assign y1972 = n14603 ;
  assign y1973 = ~n14608 ;
  assign y1974 = ~n14609 ;
  assign y1975 = ~n14611 ;
  assign y1976 = ~n14615 ;
  assign y1977 = n14622 ;
  assign y1978 = n14625 ;
  assign y1979 = n14626 ;
  assign y1980 = ~n14629 ;
  assign y1981 = ~n14642 ;
  assign y1982 = n14647 ;
  assign y1983 = ~n14652 ;
  assign y1984 = ~n14665 ;
  assign y1985 = n14678 ;
  assign y1986 = n14679 ;
  assign y1987 = ~n14690 ;
  assign y1988 = ~n14691 ;
  assign y1989 = ~n14697 ;
  assign y1990 = ~n14700 ;
  assign y1991 = n14704 ;
  assign y1992 = ~n14706 ;
  assign y1993 = n14709 ;
  assign y1994 = ~n14711 ;
  assign y1995 = n14715 ;
  assign y1996 = ~n14723 ;
  assign y1997 = n14726 ;
  assign y1998 = ~n14728 ;
  assign y1999 = ~n14736 ;
  assign y2000 = n14738 ;
  assign y2001 = ~n14741 ;
  assign y2002 = ~n14745 ;
  assign y2003 = n14747 ;
  assign y2004 = n14751 ;
  assign y2005 = n14756 ;
  assign y2006 = n14764 ;
  assign y2007 = n14765 ;
  assign y2008 = n14770 ;
  assign y2009 = ~n14776 ;
  assign y2010 = n14778 ;
  assign y2011 = ~n14783 ;
  assign y2012 = n14786 ;
  assign y2013 = n14797 ;
  assign y2014 = n14798 ;
  assign y2015 = ~n14802 ;
  assign y2016 = ~n14805 ;
  assign y2017 = n14818 ;
  assign y2018 = n14822 ;
  assign y2019 = ~n14824 ;
  assign y2020 = ~n14828 ;
  assign y2021 = ~n14832 ;
  assign y2022 = n14844 ;
  assign y2023 = n14853 ;
  assign y2024 = n14859 ;
  assign y2025 = n14863 ;
  assign y2026 = n14868 ;
  assign y2027 = ~n14877 ;
  assign y2028 = ~n14885 ;
  assign y2029 = n14892 ;
  assign y2030 = ~n14894 ;
  assign y2031 = n14895 ;
  assign y2032 = ~n14900 ;
  assign y2033 = ~n14903 ;
  assign y2034 = n14907 ;
  assign y2035 = n14908 ;
  assign y2036 = n14910 ;
  assign y2037 = n14918 ;
  assign y2038 = ~n14919 ;
  assign y2039 = ~n14925 ;
  assign y2040 = n14929 ;
  assign y2041 = ~n14937 ;
  assign y2042 = ~n14944 ;
  assign y2043 = ~n14946 ;
  assign y2044 = n14947 ;
  assign y2045 = n14951 ;
  assign y2046 = ~n14957 ;
  assign y2047 = ~n14958 ;
  assign y2048 = ~n14961 ;
  assign y2049 = n14963 ;
  assign y2050 = n14964 ;
  assign y2051 = ~n14970 ;
  assign y2052 = ~n14980 ;
  assign y2053 = ~n14987 ;
  assign y2054 = n14988 ;
  assign y2055 = n14998 ;
  assign y2056 = ~n14999 ;
  assign y2057 = ~n15001 ;
  assign y2058 = ~n15005 ;
  assign y2059 = n15010 ;
  assign y2060 = ~n15022 ;
  assign y2061 = ~n15029 ;
  assign y2062 = n15030 ;
  assign y2063 = ~n15032 ;
  assign y2064 = n15036 ;
  assign y2065 = ~n15038 ;
  assign y2066 = n15041 ;
  assign y2067 = n15043 ;
  assign y2068 = ~n15047 ;
  assign y2069 = n15049 ;
  assign y2070 = n15050 ;
  assign y2071 = ~n15053 ;
  assign y2072 = n15056 ;
  assign y2073 = n15059 ;
  assign y2074 = n15060 ;
  assign y2075 = ~n15070 ;
  assign y2076 = n15072 ;
  assign y2077 = n15085 ;
  assign y2078 = n15088 ;
  assign y2079 = n15091 ;
  assign y2080 = n15092 ;
  assign y2081 = n15093 ;
  assign y2082 = ~n15099 ;
  assign y2083 = ~n15101 ;
  assign y2084 = n15105 ;
  assign y2085 = n15108 ;
  assign y2086 = n15109 ;
  assign y2087 = n15111 ;
  assign y2088 = ~n15122 ;
  assign y2089 = ~n15124 ;
  assign y2090 = ~n15127 ;
  assign y2091 = ~n15129 ;
  assign y2092 = n15136 ;
  assign y2093 = n15138 ;
  assign y2094 = n15140 ;
  assign y2095 = n15145 ;
  assign y2096 = ~n15146 ;
  assign y2097 = n15150 ;
  assign y2098 = n15158 ;
  assign y2099 = ~n15160 ;
  assign y2100 = ~n15163 ;
  assign y2101 = ~n15165 ;
  assign y2102 = n15170 ;
  assign y2103 = ~n15171 ;
  assign y2104 = ~n15176 ;
  assign y2105 = n15178 ;
  assign y2106 = ~n15181 ;
  assign y2107 = n15185 ;
  assign y2108 = ~n15196 ;
  assign y2109 = n15210 ;
  assign y2110 = ~n15217 ;
  assign y2111 = n15221 ;
  assign y2112 = ~n15224 ;
  assign y2113 = ~n15225 ;
  assign y2114 = n15227 ;
  assign y2115 = ~n15231 ;
  assign y2116 = n15235 ;
  assign y2117 = ~n15237 ;
  assign y2118 = n15243 ;
  assign y2119 = ~n15247 ;
  assign y2120 = ~n15252 ;
  assign y2121 = n15257 ;
  assign y2122 = ~n15258 ;
  assign y2123 = n15262 ;
  assign y2124 = n15267 ;
  assign y2125 = n15270 ;
  assign y2126 = n15276 ;
  assign y2127 = ~n15280 ;
  assign y2128 = n15286 ;
  assign y2129 = ~n15290 ;
  assign y2130 = ~n15299 ;
  assign y2131 = ~n15302 ;
  assign y2132 = n15309 ;
  assign y2133 = ~n15311 ;
  assign y2134 = ~n15314 ;
  assign y2135 = n15315 ;
  assign y2136 = n15319 ;
  assign y2137 = n15324 ;
  assign y2138 = ~n15325 ;
  assign y2139 = n15327 ;
  assign y2140 = ~n15329 ;
  assign y2141 = ~n15330 ;
  assign y2142 = ~n15331 ;
  assign y2143 = n15332 ;
  assign y2144 = ~n15335 ;
  assign y2145 = ~n15340 ;
  assign y2146 = n15344 ;
  assign y2147 = ~n15349 ;
  assign y2148 = ~n15352 ;
  assign y2149 = ~n15354 ;
  assign y2150 = ~n15357 ;
  assign y2151 = n15363 ;
  assign y2152 = n15366 ;
  assign y2153 = n15369 ;
  assign y2154 = ~n15370 ;
  assign y2155 = ~n15374 ;
  assign y2156 = n15380 ;
  assign y2157 = ~n15386 ;
  assign y2158 = ~n15389 ;
  assign y2159 = ~n15394 ;
  assign y2160 = n15400 ;
  assign y2161 = ~n15403 ;
  assign y2162 = ~n15404 ;
  assign y2163 = n15408 ;
  assign y2164 = ~n15409 ;
  assign y2165 = n15410 ;
  assign y2166 = n15414 ;
  assign y2167 = ~n15425 ;
  assign y2168 = ~n15426 ;
  assign y2169 = n15427 ;
  assign y2170 = n15428 ;
  assign y2171 = n15430 ;
  assign y2172 = ~n15434 ;
  assign y2173 = n15446 ;
  assign y2174 = n15448 ;
  assign y2175 = ~n15454 ;
  assign y2176 = n15455 ;
  assign y2177 = ~n15457 ;
  assign y2178 = n15458 ;
  assign y2179 = n15462 ;
  assign y2180 = ~n15463 ;
  assign y2181 = ~n15464 ;
  assign y2182 = n15466 ;
  assign y2183 = ~n15467 ;
  assign y2184 = ~n15469 ;
  assign y2185 = n15471 ;
  assign y2186 = n15475 ;
  assign y2187 = ~n15479 ;
  assign y2188 = ~n15482 ;
  assign y2189 = ~n15485 ;
  assign y2190 = n15493 ;
  assign y2191 = ~n15497 ;
  assign y2192 = ~n15507 ;
  assign y2193 = n15512 ;
  assign y2194 = n15517 ;
  assign y2195 = ~n15522 ;
  assign y2196 = n15523 ;
  assign y2197 = ~n15527 ;
  assign y2198 = n15532 ;
  assign y2199 = n15536 ;
  assign y2200 = ~n15538 ;
  assign y2201 = ~n15543 ;
  assign y2202 = n15545 ;
  assign y2203 = n15547 ;
  assign y2204 = ~n15556 ;
  assign y2205 = n15557 ;
  assign y2206 = n15561 ;
  assign y2207 = ~n15562 ;
  assign y2208 = ~n15564 ;
  assign y2209 = ~n15566 ;
  assign y2210 = n15569 ;
  assign y2211 = n15572 ;
  assign y2212 = ~n15577 ;
  assign y2213 = ~n15581 ;
  assign y2214 = ~n15584 ;
  assign y2215 = ~n15588 ;
  assign y2216 = ~n15589 ;
  assign y2217 = ~n15591 ;
  assign y2218 = n15593 ;
  assign y2219 = n15596 ;
  assign y2220 = ~n15599 ;
  assign y2221 = n15600 ;
  assign y2222 = n15608 ;
  assign y2223 = n15610 ;
  assign y2224 = n15620 ;
  assign y2225 = ~n15622 ;
  assign y2226 = n15631 ;
  assign y2227 = ~n15632 ;
  assign y2228 = ~n15633 ;
  assign y2229 = n15637 ;
  assign y2230 = n15643 ;
  assign y2231 = n15647 ;
  assign y2232 = n15649 ;
  assign y2233 = n15651 ;
  assign y2234 = ~n15654 ;
  assign y2235 = n15658 ;
  assign y2236 = ~n15676 ;
  assign y2237 = ~n15679 ;
  assign y2238 = ~n15681 ;
  assign y2239 = ~n15684 ;
  assign y2240 = n15689 ;
  assign y2241 = n15699 ;
  assign y2242 = n15702 ;
  assign y2243 = ~n15703 ;
  assign y2244 = ~n15711 ;
  assign y2245 = ~n15720 ;
  assign y2246 = n15731 ;
  assign y2247 = n15735 ;
  assign y2248 = n15741 ;
  assign y2249 = ~n15745 ;
  assign y2250 = ~n15748 ;
  assign y2251 = ~n15750 ;
  assign y2252 = ~n15752 ;
  assign y2253 = ~n15762 ;
  assign y2254 = ~n15764 ;
  assign y2255 = ~n15766 ;
  assign y2256 = ~n15771 ;
  assign y2257 = ~n15774 ;
  assign y2258 = ~n15776 ;
  assign y2259 = ~n15782 ;
  assign y2260 = ~n15783 ;
  assign y2261 = n15784 ;
  assign y2262 = ~n15786 ;
  assign y2263 = n15788 ;
  assign y2264 = n15794 ;
  assign y2265 = n15799 ;
  assign y2266 = ~n15803 ;
  assign y2267 = ~n15804 ;
  assign y2268 = ~n15805 ;
  assign y2269 = n15810 ;
  assign y2270 = ~n15819 ;
  assign y2271 = n15824 ;
  assign y2272 = n15829 ;
  assign y2273 = ~n15837 ;
  assign y2274 = n15847 ;
  assign y2275 = ~n15858 ;
  assign y2276 = ~n15860 ;
  assign y2277 = ~n15866 ;
  assign y2278 = n15871 ;
  assign y2279 = n15882 ;
  assign y2280 = ~n15889 ;
  assign y2281 = n15891 ;
  assign y2282 = n15892 ;
  assign y2283 = n15902 ;
  assign y2284 = ~n15907 ;
  assign y2285 = n15911 ;
  assign y2286 = ~n15916 ;
  assign y2287 = ~n15918 ;
  assign y2288 = ~n15922 ;
  assign y2289 = ~n15932 ;
  assign y2290 = n15935 ;
  assign y2291 = n15937 ;
  assign y2292 = ~n15939 ;
  assign y2293 = ~n15941 ;
  assign y2294 = n15944 ;
  assign y2295 = ~n15948 ;
  assign y2296 = ~n15950 ;
  assign y2297 = ~n15958 ;
  assign y2298 = n15960 ;
  assign y2299 = ~n15961 ;
  assign y2300 = ~n15962 ;
  assign y2301 = ~n15963 ;
  assign y2302 = n15966 ;
  assign y2303 = n15977 ;
  assign y2304 = ~n15980 ;
  assign y2305 = ~n15981 ;
  assign y2306 = ~n15984 ;
  assign y2307 = ~n15985 ;
  assign y2308 = n15987 ;
  assign y2309 = n15992 ;
  assign y2310 = ~n15995 ;
  assign y2311 = ~n16000 ;
  assign y2312 = ~n16001 ;
  assign y2313 = n16004 ;
  assign y2314 = n16005 ;
  assign y2315 = n16009 ;
  assign y2316 = ~n16010 ;
  assign y2317 = n16011 ;
  assign y2318 = n16013 ;
  assign y2319 = ~n16017 ;
  assign y2320 = ~n16019 ;
  assign y2321 = ~n16021 ;
  assign y2322 = ~n16027 ;
  assign y2323 = ~n16030 ;
  assign y2324 = n16034 ;
  assign y2325 = n16037 ;
  assign y2326 = ~n16038 ;
  assign y2327 = n16039 ;
  assign y2328 = n16049 ;
  assign y2329 = ~n16051 ;
  assign y2330 = ~n16052 ;
  assign y2331 = n16054 ;
  assign y2332 = n16057 ;
  assign y2333 = ~n16062 ;
  assign y2334 = n16070 ;
  assign y2335 = n16074 ;
  assign y2336 = ~n16079 ;
  assign y2337 = n16080 ;
  assign y2338 = n16084 ;
  assign y2339 = ~n16087 ;
  assign y2340 = ~n16092 ;
  assign y2341 = n16094 ;
  assign y2342 = ~n16096 ;
  assign y2343 = ~n16097 ;
  assign y2344 = n16103 ;
  assign y2345 = ~n16108 ;
  assign y2346 = n16111 ;
  assign y2347 = n16114 ;
  assign y2348 = ~n16116 ;
  assign y2349 = ~n16118 ;
  assign y2350 = n16121 ;
  assign y2351 = n16123 ;
  assign y2352 = n16134 ;
  assign y2353 = n16138 ;
  assign y2354 = ~n16147 ;
  assign y2355 = n16157 ;
  assign y2356 = n16162 ;
  assign y2357 = ~n16166 ;
  assign y2358 = ~n16170 ;
  assign y2359 = ~n16172 ;
  assign y2360 = ~n16173 ;
  assign y2361 = n16176 ;
  assign y2362 = ~n16180 ;
  assign y2363 = ~n16185 ;
  assign y2364 = ~n16191 ;
  assign y2365 = n16192 ;
  assign y2366 = n16195 ;
  assign y2367 = n16196 ;
  assign y2368 = ~n16199 ;
  assign y2369 = ~n16200 ;
  assign y2370 = ~n16201 ;
  assign y2371 = ~n16203 ;
  assign y2372 = n16209 ;
  assign y2373 = n16210 ;
  assign y2374 = n16212 ;
  assign y2375 = ~n16215 ;
  assign y2376 = n16221 ;
  assign y2377 = ~n16234 ;
  assign y2378 = n16242 ;
  assign y2379 = n16245 ;
  assign y2380 = ~n16246 ;
  assign y2381 = n16250 ;
  assign y2382 = ~n16251 ;
  assign y2383 = n16260 ;
  assign y2384 = n16262 ;
  assign y2385 = ~n16263 ;
  assign y2386 = n16265 ;
  assign y2387 = n16267 ;
  assign y2388 = n16269 ;
  assign y2389 = ~n16273 ;
  assign y2390 = ~n16277 ;
  assign y2391 = n16279 ;
  assign y2392 = n16283 ;
  assign y2393 = ~n16295 ;
  assign y2394 = n16298 ;
  assign y2395 = n16305 ;
  assign y2396 = ~n16307 ;
  assign y2397 = n16309 ;
  assign y2398 = ~n16315 ;
  assign y2399 = ~n16317 ;
  assign y2400 = n16320 ;
  assign y2401 = n16321 ;
  assign y2402 = n16322 ;
  assign y2403 = ~n16324 ;
  assign y2404 = n16342 ;
  assign y2405 = n16344 ;
  assign y2406 = ~n16347 ;
  assign y2407 = ~n16350 ;
  assign y2408 = ~n16351 ;
  assign y2409 = n16360 ;
  assign y2410 = ~n16363 ;
  assign y2411 = ~n16365 ;
  assign y2412 = ~n16367 ;
  assign y2413 = n16375 ;
  assign y2414 = ~n16377 ;
  assign y2415 = n16380 ;
  assign y2416 = ~n16392 ;
  assign y2417 = ~n16395 ;
  assign y2418 = n16396 ;
  assign y2419 = n16399 ;
  assign y2420 = ~n16400 ;
  assign y2421 = n16405 ;
  assign y2422 = n16418 ;
  assign y2423 = n16424 ;
  assign y2424 = n16430 ;
  assign y2425 = n16441 ;
  assign y2426 = ~n16450 ;
  assign y2427 = n16452 ;
  assign y2428 = n16455 ;
  assign y2429 = n16457 ;
  assign y2430 = ~n16461 ;
  assign y2431 = n16465 ;
  assign y2432 = ~n16467 ;
  assign y2433 = ~n16470 ;
  assign y2434 = n16484 ;
  assign y2435 = n16494 ;
  assign y2436 = ~n16497 ;
  assign y2437 = n16503 ;
  assign y2438 = n16506 ;
  assign y2439 = ~n16508 ;
  assign y2440 = ~n16514 ;
  assign y2441 = n16522 ;
  assign y2442 = ~n16528 ;
  assign y2443 = n16529 ;
  assign y2444 = n16532 ;
  assign y2445 = ~n16536 ;
  assign y2446 = n16538 ;
  assign y2447 = n16541 ;
  assign y2448 = ~n16543 ;
  assign y2449 = n16547 ;
  assign y2450 = ~n16550 ;
  assign y2451 = n16556 ;
  assign y2452 = ~n16559 ;
  assign y2453 = ~n16560 ;
  assign y2454 = ~n16566 ;
  assign y2455 = ~n16567 ;
  assign y2456 = n16568 ;
  assign y2457 = n16569 ;
  assign y2458 = n16570 ;
  assign y2459 = n16575 ;
  assign y2460 = n16576 ;
  assign y2461 = ~n16579 ;
  assign y2462 = ~n16580 ;
  assign y2463 = n16582 ;
  assign y2464 = ~n16592 ;
  assign y2465 = ~n16594 ;
  assign y2466 = n16597 ;
  assign y2467 = ~n16602 ;
  assign y2468 = n16605 ;
  assign y2469 = n16607 ;
  assign y2470 = ~n16612 ;
  assign y2471 = ~n16615 ;
  assign y2472 = ~n16619 ;
  assign y2473 = n16624 ;
  assign y2474 = ~n16625 ;
  assign y2475 = n16629 ;
  assign y2476 = n16645 ;
  assign y2477 = n16649 ;
  assign y2478 = n16651 ;
  assign y2479 = n16653 ;
  assign y2480 = n16664 ;
  assign y2481 = ~n16673 ;
  assign y2482 = ~n16674 ;
  assign y2483 = ~n16675 ;
  assign y2484 = ~n16677 ;
  assign y2485 = ~n16678 ;
  assign y2486 = n16679 ;
  assign y2487 = ~n16680 ;
  assign y2488 = n16681 ;
  assign y2489 = n16683 ;
  assign y2490 = n16685 ;
  assign y2491 = n16688 ;
  assign y2492 = ~n16696 ;
  assign y2493 = n16697 ;
  assign y2494 = n16699 ;
  assign y2495 = n16701 ;
  assign y2496 = n16703 ;
  assign y2497 = ~n16707 ;
  assign y2498 = n16709 ;
  assign y2499 = ~n16715 ;
  assign y2500 = n16716 ;
  assign y2501 = n16723 ;
  assign y2502 = ~n16724 ;
  assign y2503 = n16725 ;
  assign y2504 = n16728 ;
  assign y2505 = ~n16729 ;
  assign y2506 = n16732 ;
  assign y2507 = ~n16737 ;
  assign y2508 = ~n16743 ;
  assign y2509 = n16745 ;
  assign y2510 = ~n16747 ;
  assign y2511 = n16748 ;
  assign y2512 = ~n16750 ;
  assign y2513 = ~n16756 ;
  assign y2514 = n16758 ;
  assign y2515 = n16762 ;
  assign y2516 = n16764 ;
  assign y2517 = ~n16765 ;
  assign y2518 = ~n16767 ;
  assign y2519 = n16769 ;
  assign y2520 = ~n16771 ;
  assign y2521 = n16776 ;
  assign y2522 = ~n16781 ;
  assign y2523 = ~n16784 ;
  assign y2524 = ~n16786 ;
  assign y2525 = ~n16788 ;
  assign y2526 = ~n16790 ;
  assign y2527 = ~n16792 ;
  assign y2528 = ~n16794 ;
  assign y2529 = ~n16795 ;
  assign y2530 = n16801 ;
  assign y2531 = n16804 ;
  assign y2532 = n16807 ;
  assign y2533 = n16808 ;
  assign y2534 = n16812 ;
  assign y2535 = ~n16818 ;
  assign y2536 = n16820 ;
  assign y2537 = ~n16826 ;
  assign y2538 = n16833 ;
  assign y2539 = n16835 ;
  assign y2540 = n16837 ;
  assign y2541 = n16839 ;
  assign y2542 = n16841 ;
  assign y2543 = n16843 ;
  assign y2544 = ~n16845 ;
  assign y2545 = ~n16847 ;
  assign y2546 = ~n16849 ;
  assign y2547 = n16857 ;
  assign y2548 = n16866 ;
  assign y2549 = n16872 ;
  assign y2550 = ~n16877 ;
  assign y2551 = n16879 ;
  assign y2552 = ~n16883 ;
  assign y2553 = n16887 ;
  assign y2554 = n16896 ;
  assign y2555 = n16899 ;
  assign y2556 = ~n16900 ;
  assign y2557 = ~n16903 ;
  assign y2558 = ~n16904 ;
  assign y2559 = ~n16909 ;
  assign y2560 = n16910 ;
  assign y2561 = n16922 ;
  assign y2562 = ~n16925 ;
  assign y2563 = n16928 ;
  assign y2564 = n16932 ;
  assign y2565 = n16933 ;
  assign y2566 = n16935 ;
  assign y2567 = n16937 ;
  assign y2568 = ~n16940 ;
  assign y2569 = ~n16945 ;
  assign y2570 = n16946 ;
  assign y2571 = ~n16948 ;
  assign y2572 = n16952 ;
  assign y2573 = n16953 ;
  assign y2574 = ~n16956 ;
  assign y2575 = n16960 ;
  assign y2576 = ~n16961 ;
  assign y2577 = n16962 ;
  assign y2578 = n16966 ;
  assign y2579 = ~n16971 ;
  assign y2580 = n16972 ;
  assign y2581 = ~n16974 ;
  assign y2582 = n16976 ;
  assign y2583 = n16978 ;
  assign y2584 = n16982 ;
  assign y2585 = n16985 ;
  assign y2586 = ~n16986 ;
  assign y2587 = n16992 ;
  assign y2588 = n16995 ;
  assign y2589 = ~n17000 ;
  assign y2590 = n17009 ;
  assign y2591 = ~n17012 ;
  assign y2592 = n17016 ;
  assign y2593 = ~n17020 ;
  assign y2594 = n17024 ;
  assign y2595 = ~n17028 ;
  assign y2596 = n17034 ;
  assign y2597 = ~n17036 ;
  assign y2598 = n17041 ;
  assign y2599 = n17052 ;
  assign y2600 = ~n17059 ;
  assign y2601 = n17060 ;
  assign y2602 = ~n17074 ;
  assign y2603 = n17078 ;
  assign y2604 = n17079 ;
  assign y2605 = n17085 ;
  assign y2606 = n17086 ;
  assign y2607 = ~n17087 ;
  assign y2608 = ~n17091 ;
  assign y2609 = ~n17095 ;
  assign y2610 = ~n17096 ;
  assign y2611 = ~n17097 ;
  assign y2612 = n17099 ;
  assign y2613 = n17101 ;
  assign y2614 = n17103 ;
  assign y2615 = ~n17109 ;
  assign y2616 = n17113 ;
  assign y2617 = ~n17117 ;
  assign y2618 = n17119 ;
  assign y2619 = n17120 ;
  assign y2620 = n17123 ;
  assign y2621 = ~n17128 ;
  assign y2622 = ~n17134 ;
  assign y2623 = ~n17141 ;
  assign y2624 = ~n17142 ;
  assign y2625 = n17145 ;
  assign y2626 = n17150 ;
  assign y2627 = ~n17156 ;
  assign y2628 = ~n17157 ;
  assign y2629 = n17162 ;
  assign y2630 = ~n17163 ;
  assign y2631 = ~n17171 ;
  assign y2632 = n17173 ;
  assign y2633 = ~n17178 ;
  assign y2634 = n17181 ;
  assign y2635 = ~n17182 ;
  assign y2636 = n17184 ;
  assign y2637 = n17185 ;
  assign y2638 = n17189 ;
  assign y2639 = n17192 ;
  assign y2640 = ~n17196 ;
  assign y2641 = n17198 ;
  assign y2642 = n17202 ;
  assign y2643 = n17205 ;
  assign y2644 = ~n17209 ;
  assign y2645 = n17210 ;
  assign y2646 = ~n17211 ;
  assign y2647 = n17212 ;
  assign y2648 = n17217 ;
  assign y2649 = n17222 ;
  assign y2650 = n17224 ;
  assign y2651 = n17225 ;
  assign y2652 = n17227 ;
  assign y2653 = ~n17229 ;
  assign y2654 = ~n17230 ;
  assign y2655 = ~n17233 ;
  assign y2656 = ~n17235 ;
  assign y2657 = n17236 ;
  assign y2658 = n17237 ;
  assign y2659 = ~n17238 ;
  assign y2660 = n17239 ;
  assign y2661 = ~n17242 ;
  assign y2662 = ~n17243 ;
  assign y2663 = ~n17246 ;
  assign y2664 = n17247 ;
  assign y2665 = n17254 ;
  assign y2666 = n17255 ;
  assign y2667 = ~n17261 ;
  assign y2668 = ~n17263 ;
  assign y2669 = ~n17265 ;
  assign y2670 = n17266 ;
  assign y2671 = ~n17274 ;
  assign y2672 = n17280 ;
  assign y2673 = ~n17283 ;
  assign y2674 = n17284 ;
  assign y2675 = ~n17285 ;
  assign y2676 = ~n17292 ;
  assign y2677 = n17295 ;
  assign y2678 = n17296 ;
  assign y2679 = n17300 ;
  assign y2680 = n17301 ;
  assign y2681 = ~n17303 ;
  assign y2682 = n17309 ;
  assign y2683 = ~n17311 ;
  assign y2684 = n17312 ;
  assign y2685 = n17313 ;
  assign y2686 = ~n17317 ;
  assign y2687 = ~n17320 ;
  assign y2688 = n17321 ;
  assign y2689 = n17324 ;
  assign y2690 = ~n17329 ;
  assign y2691 = n17330 ;
  assign y2692 = n17334 ;
  assign y2693 = n17336 ;
  assign y2694 = n17340 ;
  assign y2695 = n17342 ;
  assign y2696 = ~n17346 ;
  assign y2697 = ~n17350 ;
  assign y2698 = n17354 ;
  assign y2699 = ~n17355 ;
  assign y2700 = ~n17362 ;
  assign y2701 = n17367 ;
  assign y2702 = n17369 ;
  assign y2703 = ~n17377 ;
  assign y2704 = ~n17378 ;
  assign y2705 = n17380 ;
  assign y2706 = ~n17382 ;
  assign y2707 = ~n17384 ;
  assign y2708 = ~n17385 ;
  assign y2709 = ~n17388 ;
  assign y2710 = n17394 ;
  assign y2711 = n17396 ;
  assign y2712 = n17402 ;
  assign y2713 = ~n17404 ;
  assign y2714 = ~n17406 ;
  assign y2715 = ~n17413 ;
  assign y2716 = ~n17415 ;
  assign y2717 = n17417 ;
  assign y2718 = n17418 ;
  assign y2719 = ~n17420 ;
  assign y2720 = n17423 ;
  assign y2721 = ~n17424 ;
  assign y2722 = ~n17427 ;
  assign y2723 = ~n17433 ;
  assign y2724 = n17437 ;
  assign y2725 = n17438 ;
  assign y2726 = ~n17440 ;
  assign y2727 = n17445 ;
  assign y2728 = ~n17446 ;
  assign y2729 = n17450 ;
  assign y2730 = n17455 ;
  assign y2731 = n17457 ;
  assign y2732 = ~n17465 ;
  assign y2733 = n17469 ;
  assign y2734 = ~n17472 ;
  assign y2735 = ~n17477 ;
  assign y2736 = n17478 ;
  assign y2737 = n17480 ;
  assign y2738 = ~n17493 ;
  assign y2739 = ~n17499 ;
  assign y2740 = n17502 ;
  assign y2741 = ~n17505 ;
  assign y2742 = ~n17506 ;
  assign y2743 = ~n17509 ;
  assign y2744 = n17512 ;
  assign y2745 = n17514 ;
  assign y2746 = n17515 ;
  assign y2747 = n17516 ;
  assign y2748 = ~n17517 ;
  assign y2749 = ~n17519 ;
  assign y2750 = ~n17520 ;
  assign y2751 = n17527 ;
  assign y2752 = ~n17531 ;
  assign y2753 = n17542 ;
  assign y2754 = n17546 ;
  assign y2755 = n17550 ;
  assign y2756 = ~n17556 ;
  assign y2757 = ~n17560 ;
  assign y2758 = n17563 ;
  assign y2759 = n17565 ;
  assign y2760 = ~n17568 ;
  assign y2761 = n17572 ;
  assign y2762 = n17576 ;
  assign y2763 = n17587 ;
  assign y2764 = n17588 ;
  assign y2765 = ~n17590 ;
  assign y2766 = ~n17594 ;
  assign y2767 = n17599 ;
  assign y2768 = ~n17601 ;
  assign y2769 = ~n17605 ;
  assign y2770 = ~n17607 ;
  assign y2771 = ~n17608 ;
  assign y2772 = n17615 ;
  assign y2773 = ~n17617 ;
  assign y2774 = n17619 ;
  assign y2775 = ~n17639 ;
  assign y2776 = n17646 ;
  assign y2777 = n17650 ;
  assign y2778 = ~n17653 ;
  assign y2779 = n17657 ;
  assign y2780 = ~n17663 ;
  assign y2781 = n17665 ;
  assign y2782 = n17666 ;
  assign y2783 = n17667 ;
  assign y2784 = ~n17669 ;
  assign y2785 = ~n17670 ;
  assign y2786 = n17673 ;
  assign y2787 = ~n17675 ;
  assign y2788 = n17676 ;
  assign y2789 = ~n17677 ;
  assign y2790 = ~n17678 ;
  assign y2791 = n17679 ;
  assign y2792 = ~n17681 ;
  assign y2793 = n17684 ;
  assign y2794 = n17687 ;
  assign y2795 = n17689 ;
  assign y2796 = ~n17690 ;
  assign y2797 = ~n17692 ;
  assign y2798 = ~n17696 ;
  assign y2799 = ~n17698 ;
  assign y2800 = ~n17699 ;
  assign y2801 = n17701 ;
  assign y2802 = n17706 ;
  assign y2803 = ~n17711 ;
  assign y2804 = n17712 ;
  assign y2805 = n17713 ;
  assign y2806 = ~n17715 ;
  assign y2807 = ~n17719 ;
  assign y2808 = ~n17723 ;
  assign y2809 = ~n17725 ;
  assign y2810 = ~n17726 ;
  assign y2811 = ~n17728 ;
  assign y2812 = ~n17733 ;
  assign y2813 = ~n17735 ;
  assign y2814 = n17736 ;
  assign y2815 = ~n17737 ;
  assign y2816 = n17739 ;
  assign y2817 = ~n17742 ;
  assign y2818 = ~n17745 ;
  assign y2819 = ~n17748 ;
  assign y2820 = n17751 ;
  assign y2821 = ~n17752 ;
  assign y2822 = n17753 ;
  assign y2823 = ~n17755 ;
  assign y2824 = ~n17760 ;
  assign y2825 = ~n17763 ;
  assign y2826 = ~n17766 ;
  assign y2827 = n17768 ;
  assign y2828 = ~n17772 ;
  assign y2829 = ~n17774 ;
  assign y2830 = n17783 ;
  assign y2831 = ~n17788 ;
  assign y2832 = n17798 ;
  assign y2833 = ~n17805 ;
  assign y2834 = n17806 ;
  assign y2835 = n17810 ;
  assign y2836 = ~n17814 ;
  assign y2837 = ~n17821 ;
  assign y2838 = ~n17824 ;
  assign y2839 = n17825 ;
  assign y2840 = ~n17826 ;
  assign y2841 = n17834 ;
  assign y2842 = ~n17836 ;
  assign y2843 = ~n17837 ;
  assign y2844 = n17840 ;
  assign y2845 = n17843 ;
  assign y2846 = n17845 ;
  assign y2847 = n17847 ;
  assign y2848 = n17849 ;
  assign y2849 = n17852 ;
  assign y2850 = n17854 ;
  assign y2851 = n17856 ;
  assign y2852 = ~n17858 ;
  assign y2853 = ~n17862 ;
  assign y2854 = n17864 ;
  assign y2855 = n17867 ;
  assign y2856 = n17868 ;
  assign y2857 = n17869 ;
  assign y2858 = ~n17873 ;
  assign y2859 = n17875 ;
  assign y2860 = n17878 ;
  assign y2861 = n17881 ;
  assign y2862 = ~n17885 ;
  assign y2863 = n17888 ;
  assign y2864 = n17889 ;
  assign y2865 = ~n17891 ;
  assign y2866 = ~n17893 ;
  assign y2867 = ~n17896 ;
  assign y2868 = ~n17900 ;
  assign y2869 = n17902 ;
  assign y2870 = n17904 ;
  assign y2871 = n17905 ;
  assign y2872 = ~n17908 ;
  assign y2873 = n17910 ;
  assign y2874 = ~n17913 ;
  assign y2875 = n17916 ;
  assign y2876 = ~n17917 ;
  assign y2877 = n17919 ;
  assign y2878 = n17922 ;
  assign y2879 = ~n17924 ;
  assign y2880 = n17929 ;
  assign y2881 = n17936 ;
  assign y2882 = n17938 ;
  assign y2883 = ~n17940 ;
  assign y2884 = n17949 ;
  assign y2885 = n17953 ;
  assign y2886 = n17959 ;
  assign y2887 = n17967 ;
  assign y2888 = ~n17972 ;
  assign y2889 = ~n17975 ;
  assign y2890 = n17977 ;
  assign y2891 = ~n17983 ;
  assign y2892 = n17984 ;
  assign y2893 = ~n17992 ;
  assign y2894 = ~n17995 ;
  assign y2895 = ~n17997 ;
  assign y2896 = ~n18001 ;
  assign y2897 = ~n18003 ;
  assign y2898 = n18008 ;
  assign y2899 = n18009 ;
  assign y2900 = n18013 ;
  assign y2901 = n18015 ;
  assign y2902 = ~n18022 ;
  assign y2903 = n18025 ;
  assign y2904 = ~n18027 ;
  assign y2905 = n18028 ;
  assign y2906 = ~n18033 ;
  assign y2907 = ~n18035 ;
  assign y2908 = n18039 ;
  assign y2909 = n18042 ;
  assign y2910 = n18044 ;
  assign y2911 = ~n18045 ;
  assign y2912 = n18051 ;
  assign y2913 = n18057 ;
  assign y2914 = n18063 ;
  assign y2915 = n18065 ;
  assign y2916 = ~n18068 ;
  assign y2917 = ~n18071 ;
  assign y2918 = n18076 ;
  assign y2919 = n18077 ;
  assign y2920 = ~n18078 ;
  assign y2921 = n18088 ;
  assign y2922 = ~n18089 ;
  assign y2923 = ~n18091 ;
  assign y2924 = ~n18092 ;
  assign y2925 = ~n18093 ;
  assign y2926 = n18098 ;
  assign y2927 = ~n18102 ;
  assign y2928 = n18104 ;
  assign y2929 = n18107 ;
  assign y2930 = n18115 ;
  assign y2931 = ~n18119 ;
  assign y2932 = ~n18124 ;
  assign y2933 = ~n18126 ;
  assign y2934 = n18129 ;
  assign y2935 = ~n18130 ;
  assign y2936 = n18137 ;
  assign y2937 = n18143 ;
  assign y2938 = ~n18147 ;
  assign y2939 = ~n18155 ;
  assign y2940 = ~n18156 ;
  assign y2941 = ~n18158 ;
  assign y2942 = ~n18164 ;
  assign y2943 = ~n18169 ;
  assign y2944 = ~n18172 ;
  assign y2945 = n18174 ;
  assign y2946 = n18175 ;
  assign y2947 = n18176 ;
  assign y2948 = ~n18179 ;
  assign y2949 = n18182 ;
  assign y2950 = ~n18184 ;
  assign y2951 = ~n18186 ;
  assign y2952 = n18188 ;
  assign y2953 = n18190 ;
  assign y2954 = n18194 ;
  assign y2955 = ~n18199 ;
  assign y2956 = ~n18200 ;
  assign y2957 = n18203 ;
  assign y2958 = n18204 ;
  assign y2959 = n18206 ;
  assign y2960 = n18207 ;
  assign y2961 = n18213 ;
  assign y2962 = n18214 ;
  assign y2963 = ~n18216 ;
  assign y2964 = ~n18218 ;
  assign y2965 = ~n18223 ;
  assign y2966 = ~n18225 ;
  assign y2967 = n18238 ;
  assign y2968 = ~n18240 ;
  assign y2969 = n18241 ;
  assign y2970 = ~n18243 ;
  assign y2971 = n18245 ;
  assign y2972 = n18246 ;
  assign y2973 = ~n18248 ;
  assign y2974 = n18254 ;
  assign y2975 = ~n18255 ;
  assign y2976 = n18257 ;
  assign y2977 = n18259 ;
  assign y2978 = ~n18261 ;
  assign y2979 = n18266 ;
  assign y2980 = n18277 ;
  assign y2981 = ~n18278 ;
  assign y2982 = ~n18279 ;
  assign y2983 = n18280 ;
  assign y2984 = n18282 ;
  assign y2985 = ~n18284 ;
  assign y2986 = n18287 ;
  assign y2987 = ~n18294 ;
  assign y2988 = n18296 ;
  assign y2989 = ~n18297 ;
  assign y2990 = n18304 ;
  assign y2991 = n18305 ;
  assign y2992 = ~n18310 ;
  assign y2993 = ~n18312 ;
  assign y2994 = n18315 ;
  assign y2995 = ~n18323 ;
  assign y2996 = ~n18324 ;
  assign y2997 = ~n18333 ;
  assign y2998 = n18347 ;
  assign y2999 = ~n18352 ;
  assign y3000 = n18353 ;
  assign y3001 = n18359 ;
  assign y3002 = ~n18363 ;
  assign y3003 = n18370 ;
  assign y3004 = n18372 ;
  assign y3005 = n18374 ;
  assign y3006 = ~n18375 ;
  assign y3007 = n18379 ;
  assign y3008 = n18380 ;
  assign y3009 = n18381 ;
  assign y3010 = ~n18383 ;
  assign y3011 = ~n18390 ;
  assign y3012 = ~n18397 ;
  assign y3013 = ~n18407 ;
  assign y3014 = n18413 ;
  assign y3015 = ~n18415 ;
  assign y3016 = n18418 ;
  assign y3017 = n18426 ;
  assign y3018 = n18427 ;
  assign y3019 = n18430 ;
  assign y3020 = ~n18431 ;
  assign y3021 = n18433 ;
  assign y3022 = n18440 ;
  assign y3023 = ~n18448 ;
  assign y3024 = n18449 ;
  assign y3025 = n18450 ;
  assign y3026 = ~n18455 ;
  assign y3027 = ~n18459 ;
  assign y3028 = ~n18462 ;
  assign y3029 = n18465 ;
  assign y3030 = ~n18467 ;
  assign y3031 = ~n18468 ;
  assign y3032 = n18470 ;
  assign y3033 = ~n18471 ;
  assign y3034 = ~n18477 ;
  assign y3035 = ~n18481 ;
  assign y3036 = n18482 ;
  assign y3037 = n18485 ;
  assign y3038 = n18491 ;
  assign y3039 = ~n18494 ;
  assign y3040 = n18500 ;
  assign y3041 = n18501 ;
  assign y3042 = ~n18510 ;
  assign y3043 = n18513 ;
  assign y3044 = ~n18514 ;
  assign y3045 = ~n18520 ;
  assign y3046 = n18521 ;
  assign y3047 = n18532 ;
  assign y3048 = n18538 ;
  assign y3049 = n18540 ;
  assign y3050 = n18545 ;
  assign y3051 = ~n18547 ;
  assign y3052 = n18552 ;
  assign y3053 = n18554 ;
  assign y3054 = n18555 ;
  assign y3055 = ~n18558 ;
  assign y3056 = n18560 ;
  assign y3057 = ~n18562 ;
  assign y3058 = n18567 ;
  assign y3059 = n18569 ;
  assign y3060 = n18571 ;
  assign y3061 = n18573 ;
  assign y3062 = n18574 ;
  assign y3063 = ~n18576 ;
  assign y3064 = ~n18577 ;
  assign y3065 = ~n18580 ;
  assign y3066 = n18589 ;
  assign y3067 = n18594 ;
  assign y3068 = ~n18597 ;
  assign y3069 = ~n18598 ;
  assign y3070 = ~n18601 ;
  assign y3071 = n18607 ;
  assign y3072 = ~n18608 ;
  assign y3073 = n18611 ;
  assign y3074 = ~n18613 ;
  assign y3075 = n18614 ;
  assign y3076 = n18620 ;
  assign y3077 = ~n18622 ;
  assign y3078 = ~n18626 ;
  assign y3079 = ~n18627 ;
  assign y3080 = n18629 ;
  assign y3081 = n18636 ;
  assign y3082 = ~n18643 ;
  assign y3083 = ~n18645 ;
  assign y3084 = ~n18647 ;
  assign y3085 = ~n18649 ;
  assign y3086 = n18652 ;
  assign y3087 = ~n18656 ;
  assign y3088 = n18661 ;
  assign y3089 = ~n18664 ;
  assign y3090 = n18668 ;
  assign y3091 = ~n18669 ;
  assign y3092 = n18670 ;
  assign y3093 = ~n18672 ;
  assign y3094 = ~n18673 ;
  assign y3095 = n18678 ;
  assign y3096 = ~n18680 ;
  assign y3097 = ~n18681 ;
  assign y3098 = n18683 ;
  assign y3099 = n18686 ;
  assign y3100 = n18690 ;
  assign y3101 = n18698 ;
  assign y3102 = n18700 ;
  assign y3103 = n18706 ;
  assign y3104 = ~n18707 ;
  assign y3105 = ~n18709 ;
  assign y3106 = ~n18713 ;
  assign y3107 = ~n18715 ;
  assign y3108 = ~n18716 ;
  assign y3109 = n18718 ;
  assign y3110 = ~n18719 ;
  assign y3111 = ~n18723 ;
  assign y3112 = n18724 ;
  assign y3113 = ~n18726 ;
  assign y3114 = ~n18727 ;
  assign y3115 = ~n18733 ;
  assign y3116 = n18734 ;
  assign y3117 = n18741 ;
  assign y3118 = n18747 ;
  assign y3119 = ~n18748 ;
  assign y3120 = ~n18749 ;
  assign y3121 = n18758 ;
  assign y3122 = n18760 ;
  assign y3123 = ~n18763 ;
  assign y3124 = n18764 ;
  assign y3125 = n18767 ;
  assign y3126 = n18768 ;
  assign y3127 = n18771 ;
  assign y3128 = ~n18772 ;
  assign y3129 = ~n18775 ;
  assign y3130 = n18780 ;
  assign y3131 = n18784 ;
  assign y3132 = ~n18785 ;
  assign y3133 = ~n18788 ;
  assign y3134 = ~n18790 ;
  assign y3135 = ~n18791 ;
  assign y3136 = ~n18795 ;
  assign y3137 = n18796 ;
  assign y3138 = ~n18800 ;
  assign y3139 = n18804 ;
  assign y3140 = ~n18807 ;
  assign y3141 = n18812 ;
  assign y3142 = ~n18813 ;
  assign y3143 = n18815 ;
  assign y3144 = n18818 ;
  assign y3145 = n18822 ;
  assign y3146 = ~n18827 ;
  assign y3147 = ~n18828 ;
  assign y3148 = n18832 ;
  assign y3149 = ~n18835 ;
  assign y3150 = n18839 ;
  assign y3151 = n18848 ;
  assign y3152 = n18849 ;
  assign y3153 = ~n18856 ;
  assign y3154 = ~n18864 ;
  assign y3155 = n18874 ;
  assign y3156 = n18877 ;
  assign y3157 = n18880 ;
  assign y3158 = ~n18881 ;
  assign y3159 = n18886 ;
  assign y3160 = n18887 ;
  assign y3161 = n18889 ;
  assign y3162 = ~n18892 ;
  assign y3163 = n18897 ;
  assign y3164 = n18898 ;
  assign y3165 = n18900 ;
  assign y3166 = n18901 ;
  assign y3167 = ~n18903 ;
  assign y3168 = n18905 ;
  assign y3169 = ~n18911 ;
  assign y3170 = n18912 ;
  assign y3171 = ~n18914 ;
  assign y3172 = n18915 ;
  assign y3173 = n18919 ;
  assign y3174 = ~n18922 ;
  assign y3175 = ~n18923 ;
  assign y3176 = n18925 ;
  assign y3177 = ~n18926 ;
  assign y3178 = n18928 ;
  assign y3179 = ~n18933 ;
  assign y3180 = n18935 ;
  assign y3181 = ~n18941 ;
  assign y3182 = n18947 ;
  assign y3183 = n18950 ;
  assign y3184 = ~n18952 ;
  assign y3185 = ~n18965 ;
  assign y3186 = n18968 ;
  assign y3187 = n18971 ;
  assign y3188 = n18972 ;
  assign y3189 = n18975 ;
  assign y3190 = ~n18976 ;
  assign y3191 = n18982 ;
  assign y3192 = n18984 ;
  assign y3193 = ~n18987 ;
  assign y3194 = ~n18991 ;
  assign y3195 = ~n18992 ;
  assign y3196 = n18993 ;
  assign y3197 = n18998 ;
  assign y3198 = n19001 ;
  assign y3199 = ~n19004 ;
  assign y3200 = n19005 ;
  assign y3201 = ~n19006 ;
  assign y3202 = ~n19008 ;
  assign y3203 = n19009 ;
  assign y3204 = n19011 ;
  assign y3205 = n19015 ;
  assign y3206 = ~n19017 ;
  assign y3207 = n19019 ;
  assign y3208 = n19021 ;
  assign y3209 = ~n19024 ;
  assign y3210 = n19027 ;
  assign y3211 = n19030 ;
  assign y3212 = ~n19031 ;
  assign y3213 = ~n19032 ;
  assign y3214 = n19035 ;
  assign y3215 = n19042 ;
  assign y3216 = ~n19044 ;
  assign y3217 = n19051 ;
  assign y3218 = ~n19059 ;
  assign y3219 = n19061 ;
  assign y3220 = ~n19062 ;
  assign y3221 = ~n19067 ;
  assign y3222 = ~n19068 ;
  assign y3223 = n19070 ;
  assign y3224 = ~n19073 ;
  assign y3225 = n19074 ;
  assign y3226 = n19077 ;
  assign y3227 = ~n19084 ;
  assign y3228 = ~n19089 ;
  assign y3229 = n19090 ;
  assign y3230 = ~n19092 ;
  assign y3231 = ~n19093 ;
  assign y3232 = ~n19095 ;
  assign y3233 = ~n19098 ;
  assign y3234 = ~n19101 ;
  assign y3235 = n19102 ;
  assign y3236 = ~n19105 ;
  assign y3237 = n19114 ;
  assign y3238 = ~n19119 ;
  assign y3239 = ~n19121 ;
  assign y3240 = n19141 ;
  assign y3241 = ~n19145 ;
  assign y3242 = n19150 ;
  assign y3243 = n19158 ;
  assign y3244 = ~n19159 ;
  assign y3245 = ~n19167 ;
  assign y3246 = ~n19171 ;
  assign y3247 = n19173 ;
  assign y3248 = ~n19176 ;
  assign y3249 = ~n19177 ;
  assign y3250 = ~n19181 ;
  assign y3251 = ~n19185 ;
  assign y3252 = n19188 ;
  assign y3253 = n19189 ;
  assign y3254 = ~n19195 ;
  assign y3255 = n19203 ;
  assign y3256 = ~n19205 ;
  assign y3257 = n19206 ;
  assign y3258 = ~n19210 ;
  assign y3259 = ~n19212 ;
  assign y3260 = ~n19214 ;
  assign y3261 = n19215 ;
  assign y3262 = n19217 ;
  assign y3263 = n19219 ;
  assign y3264 = n19220 ;
  assign y3265 = n19229 ;
  assign y3266 = n19231 ;
  assign y3267 = ~n19233 ;
  assign y3268 = n19238 ;
  assign y3269 = n19239 ;
  assign y3270 = ~n19241 ;
  assign y3271 = ~n19244 ;
  assign y3272 = ~n19250 ;
  assign y3273 = ~n19251 ;
  assign y3274 = ~n19252 ;
  assign y3275 = n19256 ;
  assign y3276 = ~n19261 ;
  assign y3277 = n19264 ;
  assign y3278 = ~n19270 ;
  assign y3279 = n19271 ;
  assign y3280 = ~n19274 ;
  assign y3281 = n19281 ;
  assign y3282 = n19284 ;
  assign y3283 = n19286 ;
  assign y3284 = n19289 ;
  assign y3285 = ~n19292 ;
  assign y3286 = ~n19294 ;
  assign y3287 = ~n19300 ;
  assign y3288 = ~n19301 ;
  assign y3289 = n19311 ;
  assign y3290 = n19319 ;
  assign y3291 = n19323 ;
  assign y3292 = ~n19327 ;
  assign y3293 = ~n19329 ;
  assign y3294 = n19331 ;
  assign y3295 = ~n19332 ;
  assign y3296 = ~n19333 ;
  assign y3297 = ~n19336 ;
  assign y3298 = ~n19337 ;
  assign y3299 = n19340 ;
  assign y3300 = ~n19341 ;
  assign y3301 = n19345 ;
  assign y3302 = ~n19346 ;
  assign y3303 = n19348 ;
  assign y3304 = n19354 ;
  assign y3305 = ~n19356 ;
  assign y3306 = n19366 ;
  assign y3307 = n19367 ;
  assign y3308 = n19370 ;
  assign y3309 = ~n19375 ;
  assign y3310 = n19378 ;
  assign y3311 = n19384 ;
  assign y3312 = n19392 ;
  assign y3313 = ~n19393 ;
  assign y3314 = ~n19395 ;
  assign y3315 = ~n19396 ;
  assign y3316 = n19398 ;
  assign y3317 = n19399 ;
  assign y3318 = ~n19407 ;
  assign y3319 = n19408 ;
  assign y3320 = n19413 ;
  assign y3321 = ~n19416 ;
  assign y3322 = ~n19418 ;
  assign y3323 = ~n19421 ;
  assign y3324 = n19424 ;
  assign y3325 = ~n19433 ;
  assign y3326 = n19434 ;
  assign y3327 = ~n19437 ;
  assign y3328 = ~n19442 ;
  assign y3329 = ~n19446 ;
  assign y3330 = n19451 ;
  assign y3331 = n19458 ;
  assign y3332 = n19459 ;
  assign y3333 = n19460 ;
  assign y3334 = n19461 ;
  assign y3335 = ~n19462 ;
  assign y3336 = n19463 ;
  assign y3337 = n19464 ;
  assign y3338 = ~n19466 ;
  assign y3339 = n19470 ;
  assign y3340 = ~n19473 ;
  assign y3341 = ~n19474 ;
  assign y3342 = n19475 ;
  assign y3343 = ~n19479 ;
  assign y3344 = n19480 ;
  assign y3345 = n19483 ;
  assign y3346 = ~n19485 ;
  assign y3347 = n19487 ;
  assign y3348 = ~n19490 ;
  assign y3349 = ~n19496 ;
  assign y3350 = n19499 ;
  assign y3351 = ~n19504 ;
  assign y3352 = ~n19505 ;
  assign y3353 = ~n19515 ;
  assign y3354 = n19520 ;
  assign y3355 = n19521 ;
  assign y3356 = n19522 ;
  assign y3357 = ~n19523 ;
  assign y3358 = n19525 ;
  assign y3359 = n19526 ;
  assign y3360 = ~n19529 ;
  assign y3361 = n19532 ;
  assign y3362 = n19535 ;
  assign y3363 = n19537 ;
  assign y3364 = n19538 ;
  assign y3365 = ~n19541 ;
  assign y3366 = ~n19543 ;
  assign y3367 = n19544 ;
  assign y3368 = ~n19547 ;
  assign y3369 = n19551 ;
  assign y3370 = ~n19553 ;
  assign y3371 = n19555 ;
  assign y3372 = ~n19556 ;
  assign y3373 = n19558 ;
  assign y3374 = ~n19561 ;
  assign y3375 = n19564 ;
  assign y3376 = ~n19569 ;
  assign y3377 = ~n19576 ;
  assign y3378 = n19581 ;
  assign y3379 = ~n19582 ;
  assign y3380 = ~n19584 ;
  assign y3381 = n19585 ;
  assign y3382 = n19592 ;
  assign y3383 = n19594 ;
  assign y3384 = ~n19595 ;
  assign y3385 = n19598 ;
  assign y3386 = ~n19603 ;
  assign y3387 = ~n19606 ;
  assign y3388 = n19607 ;
  assign y3389 = n19617 ;
  assign y3390 = ~n19618 ;
  assign y3391 = n19621 ;
  assign y3392 = n19629 ;
  assign y3393 = n19630 ;
  assign y3394 = n19633 ;
  assign y3395 = n19635 ;
  assign y3396 = n19636 ;
  assign y3397 = ~n19645 ;
  assign y3398 = ~n19647 ;
  assign y3399 = ~n19648 ;
  assign y3400 = n19653 ;
  assign y3401 = n19655 ;
  assign y3402 = n19657 ;
  assign y3403 = n19662 ;
  assign y3404 = n19665 ;
  assign y3405 = n19670 ;
  assign y3406 = n19675 ;
  assign y3407 = n19676 ;
  assign y3408 = n19677 ;
  assign y3409 = n19683 ;
  assign y3410 = n19686 ;
  assign y3411 = n19688 ;
  assign y3412 = n19689 ;
  assign y3413 = n19690 ;
  assign y3414 = n19692 ;
  assign y3415 = ~n19699 ;
  assign y3416 = n19700 ;
  assign y3417 = ~n19703 ;
  assign y3418 = ~n19707 ;
  assign y3419 = n19711 ;
  assign y3420 = n19712 ;
  assign y3421 = ~n19716 ;
  assign y3422 = ~n19719 ;
  assign y3423 = n19723 ;
  assign y3424 = n19724 ;
  assign y3425 = n19732 ;
  assign y3426 = n19733 ;
  assign y3427 = n19736 ;
  assign y3428 = ~n19741 ;
  assign y3429 = n19746 ;
  assign y3430 = ~n19750 ;
  assign y3431 = n19751 ;
  assign y3432 = n19754 ;
  assign y3433 = n19755 ;
  assign y3434 = ~n19758 ;
  assign y3435 = n19760 ;
  assign y3436 = n19761 ;
  assign y3437 = ~n19763 ;
  assign y3438 = n19765 ;
  assign y3439 = ~n19768 ;
  assign y3440 = n19769 ;
  assign y3441 = n19770 ;
  assign y3442 = n19771 ;
  assign y3443 = n19775 ;
  assign y3444 = ~n19777 ;
  assign y3445 = ~n19783 ;
  assign y3446 = n19784 ;
  assign y3447 = n19787 ;
  assign y3448 = ~n19789 ;
  assign y3449 = ~n19793 ;
  assign y3450 = n19794 ;
  assign y3451 = ~n19795 ;
  assign y3452 = ~n19801 ;
  assign y3453 = ~n19804 ;
  assign y3454 = n19806 ;
  assign y3455 = ~n19809 ;
  assign y3456 = n19810 ;
  assign y3457 = n19812 ;
  assign y3458 = n19814 ;
  assign y3459 = n19817 ;
  assign y3460 = ~n19823 ;
  assign y3461 = ~n19826 ;
  assign y3462 = n19833 ;
  assign y3463 = ~n19839 ;
  assign y3464 = n19840 ;
  assign y3465 = n19842 ;
  assign y3466 = ~n19846 ;
  assign y3467 = n19847 ;
  assign y3468 = ~n19850 ;
  assign y3469 = ~n19853 ;
  assign y3470 = n19854 ;
  assign y3471 = n19856 ;
  assign y3472 = ~n19858 ;
  assign y3473 = n19861 ;
  assign y3474 = n19865 ;
  assign y3475 = n19870 ;
  assign y3476 = ~n19873 ;
  assign y3477 = ~n19874 ;
  assign y3478 = ~n19876 ;
  assign y3479 = n19878 ;
  assign y3480 = ~n19880 ;
  assign y3481 = n19881 ;
  assign y3482 = n19889 ;
  assign y3483 = n19890 ;
  assign y3484 = n19891 ;
  assign y3485 = ~n19894 ;
  assign y3486 = ~n19900 ;
  assign y3487 = n19902 ;
  assign y3488 = n19909 ;
  assign y3489 = n19910 ;
  assign y3490 = n19913 ;
  assign y3491 = n19914 ;
  assign y3492 = ~n19915 ;
  assign y3493 = n19921 ;
  assign y3494 = ~n19923 ;
  assign y3495 = n19927 ;
  assign y3496 = ~n19928 ;
  assign y3497 = n19933 ;
  assign y3498 = n19937 ;
  assign y3499 = n19943 ;
  assign y3500 = n19944 ;
  assign y3501 = ~n19948 ;
  assign y3502 = n19949 ;
  assign y3503 = ~n19950 ;
  assign y3504 = ~n19958 ;
  assign y3505 = ~n19959 ;
  assign y3506 = n19960 ;
  assign y3507 = ~n19968 ;
  assign y3508 = n19971 ;
  assign y3509 = ~n19974 ;
  assign y3510 = ~n19976 ;
  assign y3511 = n19984 ;
  assign y3512 = ~n19988 ;
  assign y3513 = ~n19992 ;
  assign y3514 = ~n19993 ;
  assign y3515 = ~n19997 ;
  assign y3516 = n19998 ;
  assign y3517 = ~n20001 ;
  assign y3518 = ~n20003 ;
  assign y3519 = ~n20009 ;
  assign y3520 = ~n20012 ;
  assign y3521 = n20014 ;
  assign y3522 = ~n20018 ;
  assign y3523 = n20022 ;
  assign y3524 = ~n20025 ;
  assign y3525 = n20034 ;
  assign y3526 = ~n20038 ;
  assign y3527 = n20039 ;
  assign y3528 = n20041 ;
  assign y3529 = n20046 ;
  assign y3530 = ~n20048 ;
  assign y3531 = n20050 ;
  assign y3532 = ~n20055 ;
  assign y3533 = ~n20058 ;
  assign y3534 = n20059 ;
  assign y3535 = ~n20066 ;
  assign y3536 = n20068 ;
  assign y3537 = n20072 ;
  assign y3538 = ~n20076 ;
  assign y3539 = ~n20078 ;
  assign y3540 = ~n20079 ;
  assign y3541 = n20082 ;
  assign y3542 = ~n20083 ;
  assign y3543 = ~n20084 ;
  assign y3544 = n20087 ;
  assign y3545 = n20088 ;
  assign y3546 = n20089 ;
  assign y3547 = ~n20090 ;
  assign y3548 = ~n20092 ;
  assign y3549 = ~n20093 ;
  assign y3550 = n20097 ;
  assign y3551 = n20108 ;
  assign y3552 = ~n20111 ;
  assign y3553 = ~n20115 ;
  assign y3554 = ~n20116 ;
  assign y3555 = ~n20117 ;
  assign y3556 = ~n20118 ;
  assign y3557 = n20123 ;
  assign y3558 = n20126 ;
  assign y3559 = ~n20129 ;
  assign y3560 = ~n20130 ;
  assign y3561 = ~n20131 ;
  assign y3562 = n20135 ;
  assign y3563 = n20137 ;
  assign y3564 = ~n20139 ;
  assign y3565 = ~n20142 ;
  assign y3566 = n20144 ;
  assign y3567 = n20145 ;
  assign y3568 = n20156 ;
  assign y3569 = ~n20161 ;
  assign y3570 = ~n20164 ;
  assign y3571 = n20166 ;
  assign y3572 = ~n20168 ;
  assign y3573 = n20171 ;
  assign y3574 = ~n20175 ;
  assign y3575 = ~n20190 ;
  assign y3576 = ~n20198 ;
  assign y3577 = ~n20200 ;
  assign y3578 = n20201 ;
  assign y3579 = n20203 ;
  assign y3580 = n20204 ;
  assign y3581 = n20205 ;
  assign y3582 = ~n20212 ;
  assign y3583 = n20214 ;
  assign y3584 = n20216 ;
  assign y3585 = n20222 ;
  assign y3586 = ~n20225 ;
  assign y3587 = ~n20232 ;
  assign y3588 = n20238 ;
  assign y3589 = n20244 ;
  assign y3590 = n20247 ;
  assign y3591 = n20248 ;
  assign y3592 = n20251 ;
  assign y3593 = ~n20257 ;
  assign y3594 = n20258 ;
  assign y3595 = n20260 ;
  assign y3596 = n20262 ;
  assign y3597 = ~n20266 ;
  assign y3598 = n20268 ;
  assign y3599 = ~n20269 ;
  assign y3600 = n20270 ;
  assign y3601 = n20273 ;
  assign y3602 = n20275 ;
  assign y3603 = n20277 ;
  assign y3604 = ~n20282 ;
  assign y3605 = n20287 ;
  assign y3606 = ~n20290 ;
  assign y3607 = ~n20291 ;
  assign y3608 = ~n20292 ;
  assign y3609 = n20296 ;
  assign y3610 = ~n20297 ;
  assign y3611 = ~n20300 ;
  assign y3612 = n20302 ;
  assign y3613 = n20307 ;
  assign y3614 = ~n20313 ;
  assign y3615 = ~n20315 ;
  assign y3616 = ~n20317 ;
  assign y3617 = n20319 ;
  assign y3618 = ~n20324 ;
  assign y3619 = n20330 ;
  assign y3620 = ~n20333 ;
  assign y3621 = n20341 ;
  assign y3622 = ~n20343 ;
  assign y3623 = n20345 ;
  assign y3624 = ~n20346 ;
  assign y3625 = n20348 ;
  assign y3626 = ~n20351 ;
  assign y3627 = ~n20352 ;
  assign y3628 = n20354 ;
  assign y3629 = n20359 ;
  assign y3630 = n20360 ;
  assign y3631 = n20362 ;
  assign y3632 = n20364 ;
  assign y3633 = n20365 ;
  assign y3634 = n20367 ;
  assign y3635 = n20371 ;
  assign y3636 = ~n20372 ;
  assign y3637 = n20373 ;
  assign y3638 = n20374 ;
  assign y3639 = ~n20378 ;
  assign y3640 = ~n20383 ;
  assign y3641 = ~n20386 ;
  assign y3642 = n20387 ;
  assign y3643 = n20388 ;
  assign y3644 = n20393 ;
  assign y3645 = n20394 ;
  assign y3646 = ~n20395 ;
  assign y3647 = n20397 ;
  assign y3648 = n20399 ;
  assign y3649 = n20404 ;
  assign y3650 = n20412 ;
  assign y3651 = ~n20413 ;
  assign y3652 = ~n20415 ;
  assign y3653 = ~n20418 ;
  assign y3654 = ~n20421 ;
  assign y3655 = n20423 ;
  assign y3656 = n20424 ;
  assign y3657 = n20427 ;
  assign y3658 = n20430 ;
  assign y3659 = ~n20432 ;
  assign y3660 = n20434 ;
  assign y3661 = ~n20436 ;
  assign y3662 = ~n20437 ;
  assign y3663 = ~n20440 ;
  assign y3664 = ~n20442 ;
  assign y3665 = ~n20443 ;
  assign y3666 = n20446 ;
  assign y3667 = ~n20449 ;
  assign y3668 = ~n20457 ;
  assign y3669 = n20459 ;
  assign y3670 = ~n20461 ;
  assign y3671 = n20464 ;
  assign y3672 = n20471 ;
  assign y3673 = n20473 ;
  assign y3674 = n20477 ;
  assign y3675 = ~n20481 ;
  assign y3676 = n20483 ;
  assign y3677 = n20484 ;
  assign y3678 = n20491 ;
  assign y3679 = ~n20492 ;
  assign y3680 = n20499 ;
  assign y3681 = ~n20500 ;
  assign y3682 = n20504 ;
  assign y3683 = ~n20507 ;
  assign y3684 = ~n20509 ;
  assign y3685 = n20513 ;
  assign y3686 = ~n20518 ;
  assign y3687 = n20522 ;
  assign y3688 = n20525 ;
  assign y3689 = n20527 ;
  assign y3690 = n20534 ;
  assign y3691 = n20536 ;
  assign y3692 = ~n20545 ;
  assign y3693 = ~n20548 ;
  assign y3694 = n20553 ;
  assign y3695 = ~n20555 ;
  assign y3696 = ~n20561 ;
  assign y3697 = n20585 ;
  assign y3698 = ~n20592 ;
  assign y3699 = ~n20593 ;
  assign y3700 = ~n20600 ;
  assign y3701 = ~n20602 ;
  assign y3702 = n20603 ;
  assign y3703 = ~n20607 ;
  assign y3704 = ~n20608 ;
  assign y3705 = n20610 ;
  assign y3706 = ~n20611 ;
  assign y3707 = n20615 ;
  assign y3708 = ~n20619 ;
  assign y3709 = n20622 ;
  assign y3710 = ~n20628 ;
  assign y3711 = ~n20630 ;
  assign y3712 = n20633 ;
  assign y3713 = ~n20636 ;
  assign y3714 = ~n20638 ;
  assign y3715 = ~n20644 ;
  assign y3716 = n20648 ;
  assign y3717 = ~n20649 ;
  assign y3718 = ~n20650 ;
  assign y3719 = n20655 ;
  assign y3720 = ~n20658 ;
  assign y3721 = ~n20662 ;
  assign y3722 = n20663 ;
  assign y3723 = n20664 ;
  assign y3724 = ~n20667 ;
  assign y3725 = ~n20668 ;
  assign y3726 = ~n20670 ;
  assign y3727 = n20672 ;
  assign y3728 = ~n20675 ;
  assign y3729 = ~n20676 ;
  assign y3730 = ~n20680 ;
  assign y3731 = ~n20682 ;
  assign y3732 = ~n20684 ;
  assign y3733 = ~n20685 ;
  assign y3734 = ~n20686 ;
  assign y3735 = n20688 ;
  assign y3736 = ~n20690 ;
  assign y3737 = n20692 ;
  assign y3738 = n20696 ;
  assign y3739 = ~n20697 ;
  assign y3740 = n20700 ;
  assign y3741 = n20702 ;
  assign y3742 = n20703 ;
  assign y3743 = n20706 ;
  assign y3744 = n20711 ;
  assign y3745 = n20716 ;
  assign y3746 = n20717 ;
  assign y3747 = ~n20719 ;
  assign y3748 = n20720 ;
  assign y3749 = n20736 ;
  assign y3750 = ~n20740 ;
  assign y3751 = ~n20742 ;
  assign y3752 = n20744 ;
  assign y3753 = ~n20747 ;
  assign y3754 = ~n20750 ;
  assign y3755 = ~n20752 ;
  assign y3756 = n20754 ;
  assign y3757 = ~n20758 ;
  assign y3758 = ~n20759 ;
  assign y3759 = n20763 ;
  assign y3760 = n20764 ;
  assign y3761 = ~n20766 ;
  assign y3762 = n20767 ;
  assign y3763 = n20768 ;
  assign y3764 = ~n20770 ;
  assign y3765 = n20773 ;
  assign y3766 = ~n20776 ;
  assign y3767 = n20777 ;
  assign y3768 = ~n20779 ;
  assign y3769 = ~n20780 ;
  assign y3770 = n20783 ;
  assign y3771 = ~n20785 ;
  assign y3772 = ~n20786 ;
  assign y3773 = n20787 ;
  assign y3774 = n20788 ;
  assign y3775 = ~n20789 ;
  assign y3776 = n20798 ;
  assign y3777 = n20799 ;
  assign y3778 = ~n20800 ;
  assign y3779 = n20806 ;
  assign y3780 = ~n20811 ;
  assign y3781 = ~n20812 ;
  assign y3782 = ~n20813 ;
  assign y3783 = n20814 ;
  assign y3784 = ~n20816 ;
  assign y3785 = n20819 ;
  assign y3786 = ~n20820 ;
  assign y3787 = ~n20822 ;
  assign y3788 = n20824 ;
  assign y3789 = ~n20826 ;
  assign y3790 = n20829 ;
  assign y3791 = n20830 ;
  assign y3792 = ~n20831 ;
  assign y3793 = n20835 ;
  assign y3794 = ~n20836 ;
  assign y3795 = ~n20838 ;
  assign y3796 = n20843 ;
  assign y3797 = ~n20846 ;
  assign y3798 = n20848 ;
  assign y3799 = ~n20849 ;
  assign y3800 = ~n20851 ;
  assign y3801 = ~n20857 ;
  assign y3802 = n20858 ;
  assign y3803 = n20861 ;
  assign y3804 = n20864 ;
  assign y3805 = ~n20867 ;
  assign y3806 = ~n20873 ;
  assign y3807 = n20876 ;
  assign y3808 = ~n20882 ;
  assign y3809 = n20883 ;
  assign y3810 = ~n20887 ;
  assign y3811 = n20892 ;
  assign y3812 = ~n20894 ;
  assign y3813 = ~n20896 ;
  assign y3814 = ~n20897 ;
  assign y3815 = ~n20900 ;
  assign y3816 = ~n20905 ;
  assign y3817 = n20910 ;
  assign y3818 = ~n20913 ;
  assign y3819 = ~n20918 ;
  assign y3820 = ~n20920 ;
  assign y3821 = n20921 ;
  assign y3822 = ~n20922 ;
  assign y3823 = ~n20926 ;
  assign y3824 = n20929 ;
  assign y3825 = ~n20930 ;
  assign y3826 = ~n20932 ;
  assign y3827 = n20933 ;
  assign y3828 = ~n20937 ;
  assign y3829 = ~n20938 ;
  assign y3830 = ~n20939 ;
  assign y3831 = ~n20940 ;
  assign y3832 = n20942 ;
  assign y3833 = ~n20947 ;
  assign y3834 = ~n20949 ;
  assign y3835 = n20950 ;
  assign y3836 = ~n20954 ;
  assign y3837 = ~n20955 ;
  assign y3838 = ~n20956 ;
  assign y3839 = ~n20958 ;
  assign y3840 = n20959 ;
  assign y3841 = ~n20963 ;
  assign y3842 = n20966 ;
  assign y3843 = n20968 ;
  assign y3844 = n20969 ;
  assign y3845 = n20971 ;
  assign y3846 = n20972 ;
  assign y3847 = ~n20974 ;
  assign y3848 = ~n20978 ;
  assign y3849 = ~n20979 ;
  assign y3850 = n20981 ;
  assign y3851 = ~n20982 ;
  assign y3852 = ~n20985 ;
  assign y3853 = n20986 ;
  assign y3854 = ~n20991 ;
  assign y3855 = ~n20992 ;
  assign y3856 = ~n20995 ;
  assign y3857 = n20999 ;
  assign y3858 = n21001 ;
  assign y3859 = ~n21004 ;
  assign y3860 = ~n21005 ;
  assign y3861 = n21009 ;
  assign y3862 = n21010 ;
  assign y3863 = n21011 ;
  assign y3864 = n21012 ;
  assign y3865 = n21015 ;
  assign y3866 = ~n21016 ;
  assign y3867 = ~n21017 ;
  assign y3868 = n21022 ;
  assign y3869 = ~n21025 ;
  assign y3870 = n21027 ;
  assign y3871 = n21031 ;
  assign y3872 = n21032 ;
  assign y3873 = n21034 ;
  assign y3874 = ~n21035 ;
  assign y3875 = n21040 ;
  assign y3876 = n21042 ;
  assign y3877 = ~n21043 ;
  assign y3878 = n21045 ;
  assign y3879 = n21048 ;
  assign y3880 = ~n21052 ;
  assign y3881 = n21053 ;
  assign y3882 = n21058 ;
  assign y3883 = ~n21061 ;
  assign y3884 = n21066 ;
  assign y3885 = n21074 ;
  assign y3886 = n21075 ;
  assign y3887 = ~n21077 ;
  assign y3888 = ~n21078 ;
  assign y3889 = ~n21079 ;
  assign y3890 = ~n21082 ;
  assign y3891 = n21083 ;
  assign y3892 = ~n21086 ;
  assign y3893 = n21090 ;
  assign y3894 = ~n21094 ;
  assign y3895 = n21100 ;
  assign y3896 = n21103 ;
  assign y3897 = ~n21105 ;
  assign y3898 = ~n21106 ;
  assign y3899 = ~n21112 ;
  assign y3900 = n21120 ;
  assign y3901 = ~n21121 ;
  assign y3902 = n21126 ;
  assign y3903 = n21129 ;
  assign y3904 = n21134 ;
  assign y3905 = ~n21135 ;
  assign y3906 = ~n21139 ;
  assign y3907 = n21140 ;
  assign y3908 = ~n21144 ;
  assign y3909 = n21145 ;
  assign y3910 = ~n21149 ;
  assign y3911 = n21151 ;
  assign y3912 = ~n21152 ;
  assign y3913 = ~n21154 ;
  assign y3914 = n21159 ;
  assign y3915 = ~n21163 ;
  assign y3916 = ~n21164 ;
  assign y3917 = ~n21169 ;
  assign y3918 = n21171 ;
  assign y3919 = n21176 ;
  assign y3920 = n21177 ;
  assign y3921 = n21178 ;
  assign y3922 = ~n21180 ;
  assign y3923 = ~n21183 ;
  assign y3924 = ~n21185 ;
  assign y3925 = n21187 ;
  assign y3926 = n21188 ;
  assign y3927 = n21189 ;
  assign y3928 = ~n21192 ;
  assign y3929 = ~n21193 ;
  assign y3930 = ~n21195 ;
  assign y3931 = n21197 ;
  assign y3932 = ~n21200 ;
  assign y3933 = n21208 ;
  assign y3934 = n21214 ;
  assign y3935 = ~n21215 ;
  assign y3936 = n21218 ;
  assign y3937 = n21221 ;
  assign y3938 = ~n21222 ;
  assign y3939 = ~n21224 ;
  assign y3940 = ~n21226 ;
  assign y3941 = n21228 ;
  assign y3942 = n21231 ;
  assign y3943 = n21233 ;
  assign y3944 = n21237 ;
  assign y3945 = ~n21238 ;
  assign y3946 = n21239 ;
  assign y3947 = n21240 ;
  assign y3948 = n21243 ;
  assign y3949 = ~n21244 ;
  assign y3950 = n21245 ;
  assign y3951 = ~n21247 ;
  assign y3952 = n21254 ;
  assign y3953 = ~n21255 ;
  assign y3954 = n21257 ;
  assign y3955 = n21263 ;
  assign y3956 = n21272 ;
  assign y3957 = n21276 ;
  assign y3958 = n21281 ;
  assign y3959 = n21286 ;
  assign y3960 = ~n21288 ;
  assign y3961 = ~n21290 ;
  assign y3962 = ~n21297 ;
  assign y3963 = ~n21303 ;
  assign y3964 = ~n21305 ;
  assign y3965 = n21306 ;
  assign y3966 = n21308 ;
  assign y3967 = n21309 ;
  assign y3968 = n21311 ;
  assign y3969 = n21317 ;
  assign y3970 = n21320 ;
  assign y3971 = ~n21322 ;
  assign y3972 = n21323 ;
  assign y3973 = n21324 ;
  assign y3974 = n21325 ;
  assign y3975 = ~n21328 ;
  assign y3976 = n21334 ;
  assign y3977 = ~n21339 ;
  assign y3978 = ~n21341 ;
  assign y3979 = n21343 ;
  assign y3980 = ~n21344 ;
  assign y3981 = ~n21345 ;
  assign y3982 = ~n21348 ;
  assign y3983 = ~n21350 ;
  assign y3984 = ~n21352 ;
  assign y3985 = n21355 ;
  assign y3986 = ~n21356 ;
  assign y3987 = ~n21358 ;
  assign y3988 = ~n21360 ;
  assign y3989 = n21362 ;
  assign y3990 = ~n21367 ;
  assign y3991 = ~n21371 ;
  assign y3992 = ~n21374 ;
  assign y3993 = n21376 ;
  assign y3994 = n21379 ;
  assign y3995 = ~n21381 ;
  assign y3996 = ~n21388 ;
  assign y3997 = n21389 ;
  assign y3998 = n21391 ;
  assign y3999 = n21394 ;
  assign y4000 = ~n21395 ;
  assign y4001 = ~n21399 ;
  assign y4002 = ~n21400 ;
  assign y4003 = ~n21404 ;
  assign y4004 = n21408 ;
  assign y4005 = ~n21412 ;
  assign y4006 = n21415 ;
  assign y4007 = ~n21420 ;
  assign y4008 = n21421 ;
  assign y4009 = ~n21423 ;
  assign y4010 = ~n21425 ;
  assign y4011 = n21426 ;
  assign y4012 = ~n21428 ;
  assign y4013 = n21431 ;
  assign y4014 = ~n21434 ;
  assign y4015 = n21438 ;
  assign y4016 = ~n21439 ;
  assign y4017 = n21443 ;
  assign y4018 = n21447 ;
  assign y4019 = n21448 ;
  assign y4020 = ~n21451 ;
  assign y4021 = n21453 ;
  assign y4022 = ~n21456 ;
  assign y4023 = ~n21457 ;
  assign y4024 = n21459 ;
  assign y4025 = ~n21468 ;
  assign y4026 = ~n21469 ;
  assign y4027 = ~n21472 ;
  assign y4028 = n21474 ;
  assign y4029 = n21477 ;
  assign y4030 = ~n21480 ;
  assign y4031 = n21482 ;
  assign y4032 = ~n21484 ;
  assign y4033 = ~n21485 ;
  assign y4034 = n21490 ;
  assign y4035 = n21491 ;
  assign y4036 = n21493 ;
  assign y4037 = n21495 ;
  assign y4038 = ~n21497 ;
  assign y4039 = n21505 ;
  assign y4040 = n21510 ;
  assign y4041 = n21512 ;
  assign y4042 = n21513 ;
  assign y4043 = ~n21515 ;
  assign y4044 = n21517 ;
  assign y4045 = n21520 ;
  assign y4046 = ~n21522 ;
  assign y4047 = n21526 ;
  assign y4048 = ~n21527 ;
  assign y4049 = ~n21529 ;
  assign y4050 = ~n21533 ;
  assign y4051 = n21536 ;
  assign y4052 = n21538 ;
  assign y4053 = ~n21539 ;
  assign y4054 = n21541 ;
  assign y4055 = n21542 ;
  assign y4056 = n21556 ;
  assign y4057 = ~n21557 ;
  assign y4058 = n21559 ;
  assign y4059 = n21563 ;
  assign y4060 = ~n21569 ;
  assign y4061 = ~n21574 ;
  assign y4062 = ~n21578 ;
  assign y4063 = n21580 ;
  assign y4064 = n21583 ;
  assign y4065 = n21584 ;
  assign y4066 = ~n21587 ;
  assign y4067 = n21592 ;
  assign y4068 = ~n21596 ;
  assign y4069 = ~n21597 ;
  assign y4070 = ~n21598 ;
  assign y4071 = n21614 ;
  assign y4072 = n21615 ;
  assign y4073 = n21622 ;
  assign y4074 = ~n21625 ;
  assign y4075 = ~n21631 ;
  assign y4076 = ~n21634 ;
  assign y4077 = ~n21635 ;
  assign y4078 = ~n21637 ;
  assign y4079 = ~n21639 ;
  assign y4080 = n21640 ;
  assign y4081 = n21641 ;
  assign y4082 = ~n21642 ;
  assign y4083 = ~n21650 ;
  assign y4084 = n21654 ;
  assign y4085 = ~n21658 ;
  assign y4086 = n21660 ;
  assign y4087 = ~n21666 ;
  assign y4088 = ~n21673 ;
  assign y4089 = n21675 ;
  assign y4090 = n21678 ;
  assign y4091 = n21679 ;
  assign y4092 = ~n21680 ;
  assign y4093 = ~n21683 ;
  assign y4094 = ~n21687 ;
  assign y4095 = n21691 ;
  assign y4096 = n21694 ;
  assign y4097 = ~n21696 ;
  assign y4098 = n21709 ;
  assign y4099 = n21710 ;
  assign y4100 = ~n21711 ;
  assign y4101 = n21712 ;
  assign y4102 = n21713 ;
  assign y4103 = n21715 ;
  assign y4104 = n21720 ;
  assign y4105 = n21726 ;
  assign y4106 = ~n21729 ;
  assign y4107 = ~n21733 ;
  assign y4108 = n21734 ;
  assign y4109 = ~n21736 ;
  assign y4110 = n21738 ;
  assign y4111 = ~n21740 ;
  assign y4112 = n21741 ;
  assign y4113 = ~n21747 ;
  assign y4114 = n21750 ;
  assign y4115 = ~n21751 ;
  assign y4116 = ~n21756 ;
  assign y4117 = n21759 ;
  assign y4118 = ~n21761 ;
  assign y4119 = n21765 ;
  assign y4120 = ~n21773 ;
  assign y4121 = n21775 ;
  assign y4122 = n21777 ;
  assign y4123 = n21778 ;
  assign y4124 = ~n21782 ;
  assign y4125 = n21785 ;
  assign y4126 = ~n21786 ;
  assign y4127 = ~n21789 ;
  assign y4128 = n21792 ;
  assign y4129 = n21795 ;
  assign y4130 = ~n21804 ;
  assign y4131 = ~n21805 ;
  assign y4132 = ~n21807 ;
  assign y4133 = n21809 ;
  assign y4134 = n21813 ;
  assign y4135 = ~n21816 ;
  assign y4136 = n21817 ;
  assign y4137 = ~n21819 ;
  assign y4138 = ~n21820 ;
  assign y4139 = n21821 ;
  assign y4140 = n21823 ;
  assign y4141 = ~n21830 ;
  assign y4142 = n21834 ;
  assign y4143 = ~n21835 ;
  assign y4144 = n21836 ;
  assign y4145 = ~n21840 ;
  assign y4146 = n21841 ;
  assign y4147 = ~n21844 ;
  assign y4148 = n21847 ;
  assign y4149 = ~n21849 ;
  assign y4150 = n21853 ;
  assign y4151 = n21857 ;
  assign y4152 = n21858 ;
  assign y4153 = n21860 ;
  assign y4154 = ~n21861 ;
  assign y4155 = n21862 ;
  assign y4156 = n21872 ;
  assign y4157 = n21874 ;
  assign y4158 = ~n21877 ;
  assign y4159 = ~n21881 ;
  assign y4160 = ~n21887 ;
  assign y4161 = n21893 ;
  assign y4162 = ~n21894 ;
  assign y4163 = ~n21898 ;
  assign y4164 = ~n21900 ;
  assign y4165 = n21903 ;
  assign y4166 = ~n21907 ;
  assign y4167 = ~n21908 ;
  assign y4168 = ~n21909 ;
  assign y4169 = n21913 ;
  assign y4170 = n21915 ;
  assign y4171 = n21916 ;
  assign y4172 = n21919 ;
  assign y4173 = ~n21920 ;
  assign y4174 = ~n21926 ;
  assign y4175 = ~n21927 ;
  assign y4176 = n21931 ;
  assign y4177 = ~n21937 ;
  assign y4178 = ~n21939 ;
  assign y4179 = ~n21940 ;
  assign y4180 = n21945 ;
  assign y4181 = n21946 ;
  assign y4182 = ~n21947 ;
  assign y4183 = n21950 ;
  assign y4184 = n21960 ;
  assign y4185 = ~n21961 ;
  assign y4186 = n21962 ;
  assign y4187 = n21968 ;
  assign y4188 = n21970 ;
  assign y4189 = ~n21972 ;
  assign y4190 = n21975 ;
  assign y4191 = ~n21977 ;
  assign y4192 = n21979 ;
  assign y4193 = n21984 ;
  assign y4194 = ~n21986 ;
  assign y4195 = ~n21988 ;
  assign y4196 = n21989 ;
  assign y4197 = n21990 ;
  assign y4198 = n21991 ;
  assign y4199 = ~n21992 ;
  assign y4200 = n21997 ;
  assign y4201 = n21998 ;
  assign y4202 = n21999 ;
  assign y4203 = ~n22000 ;
  assign y4204 = n22003 ;
  assign y4205 = ~n22007 ;
  assign y4206 = ~n22008 ;
  assign y4207 = n22009 ;
  assign y4208 = n22011 ;
  assign y4209 = ~n22012 ;
  assign y4210 = ~n22016 ;
  assign y4211 = n22020 ;
  assign y4212 = n22027 ;
  assign y4213 = ~n22037 ;
  assign y4214 = n22042 ;
  assign y4215 = n22047 ;
  assign y4216 = n22054 ;
  assign y4217 = n22058 ;
  assign y4218 = n22059 ;
  assign y4219 = n22061 ;
  assign y4220 = ~n22065 ;
  assign y4221 = n22067 ;
  assign y4222 = n22072 ;
  assign y4223 = n22074 ;
  assign y4224 = n22077 ;
  assign y4225 = n22082 ;
  assign y4226 = n22085 ;
  assign y4227 = n22091 ;
  assign y4228 = n22096 ;
  assign y4229 = ~n22100 ;
  assign y4230 = n22116 ;
  assign y4231 = n22120 ;
  assign y4232 = ~n22121 ;
  assign y4233 = n22122 ;
  assign y4234 = ~n22127 ;
  assign y4235 = n22129 ;
  assign y4236 = n22130 ;
  assign y4237 = ~n22135 ;
  assign y4238 = n22136 ;
  assign y4239 = ~n22142 ;
  assign y4240 = n22143 ;
  assign y4241 = n22144 ;
  assign y4242 = ~n22145 ;
  assign y4243 = ~n22146 ;
  assign y4244 = n22147 ;
  assign y4245 = n22149 ;
  assign y4246 = n22153 ;
  assign y4247 = ~n22155 ;
  assign y4248 = n22156 ;
  assign y4249 = ~n22158 ;
  assign y4250 = ~n22162 ;
  assign y4251 = n22165 ;
  assign y4252 = n22166 ;
  assign y4253 = n22170 ;
  assign y4254 = ~n22172 ;
  assign y4255 = ~n22174 ;
  assign y4256 = ~n22177 ;
  assign y4257 = ~n22178 ;
  assign y4258 = n22180 ;
  assign y4259 = ~n22181 ;
  assign y4260 = n22182 ;
  assign y4261 = n22184 ;
  assign y4262 = n22188 ;
  assign y4263 = n22196 ;
  assign y4264 = n22207 ;
  assign y4265 = n22210 ;
  assign y4266 = ~n22212 ;
  assign y4267 = n22214 ;
  assign y4268 = ~n22218 ;
  assign y4269 = n22221 ;
  assign y4270 = n22222 ;
  assign y4271 = n22227 ;
  assign y4272 = n22229 ;
  assign y4273 = n22235 ;
  assign y4274 = n22241 ;
  assign y4275 = n22242 ;
  assign y4276 = ~n22252 ;
  assign y4277 = ~n22257 ;
  assign y4278 = ~n22258 ;
  assign y4279 = n22261 ;
  assign y4280 = n22265 ;
  assign y4281 = n22271 ;
  assign y4282 = ~n22272 ;
  assign y4283 = ~n22278 ;
  assign y4284 = ~n22279 ;
  assign y4285 = ~n22283 ;
  assign y4286 = n22289 ;
  assign y4287 = n22295 ;
  assign y4288 = ~n22296 ;
  assign y4289 = n22301 ;
  assign y4290 = ~n22302 ;
  assign y4291 = n22303 ;
  assign y4292 = n22309 ;
  assign y4293 = n22311 ;
  assign y4294 = ~n22314 ;
  assign y4295 = n22316 ;
  assign y4296 = n22317 ;
  assign y4297 = n22320 ;
  assign y4298 = ~n22322 ;
  assign y4299 = ~n22323 ;
  assign y4300 = n22327 ;
  assign y4301 = n22330 ;
  assign y4302 = ~n22331 ;
  assign y4303 = ~n22333 ;
  assign y4304 = ~n22335 ;
  assign y4305 = n22338 ;
  assign y4306 = ~n22340 ;
  assign y4307 = ~n22342 ;
  assign y4308 = ~n22344 ;
  assign y4309 = n22345 ;
  assign y4310 = n22347 ;
  assign y4311 = ~n22348 ;
  assign y4312 = ~n22351 ;
  assign y4313 = ~n22354 ;
  assign y4314 = ~n22355 ;
  assign y4315 = ~n22356 ;
  assign y4316 = ~n22357 ;
  assign y4317 = ~n22361 ;
  assign y4318 = ~n22365 ;
  assign y4319 = ~n22366 ;
  assign y4320 = ~n22367 ;
  assign y4321 = ~n22368 ;
  assign y4322 = ~n22369 ;
  assign y4323 = ~n22371 ;
  assign y4324 = n22372 ;
  assign y4325 = n22374 ;
  assign y4326 = n22377 ;
  assign y4327 = n22378 ;
  assign y4328 = n22380 ;
  assign y4329 = ~n22381 ;
  assign y4330 = ~n22383 ;
  assign y4331 = ~n22384 ;
  assign y4332 = ~n22387 ;
  assign y4333 = ~n22389 ;
  assign y4334 = ~n22395 ;
  assign y4335 = n22401 ;
  assign y4336 = n22404 ;
  assign y4337 = n22405 ;
  assign y4338 = n22407 ;
  assign y4339 = ~n22408 ;
  assign y4340 = ~n22413 ;
  assign y4341 = n22418 ;
  assign y4342 = n22423 ;
  assign y4343 = n22427 ;
  assign y4344 = ~n22428 ;
  assign y4345 = ~n22429 ;
  assign y4346 = n22435 ;
  assign y4347 = n22436 ;
  assign y4348 = n22439 ;
  assign y4349 = n22443 ;
  assign y4350 = ~n22448 ;
  assign y4351 = ~n22449 ;
  assign y4352 = ~n22452 ;
  assign y4353 = ~n22454 ;
  assign y4354 = ~n22462 ;
  assign y4355 = n22466 ;
  assign y4356 = n22470 ;
  assign y4357 = ~n22472 ;
  assign y4358 = n22473 ;
  assign y4359 = ~n22475 ;
  assign y4360 = ~n22477 ;
  assign y4361 = ~n22479 ;
  assign y4362 = ~n22480 ;
  assign y4363 = n22483 ;
  assign y4364 = ~n22486 ;
  assign y4365 = ~n22490 ;
  assign y4366 = n22491 ;
  assign y4367 = n22494 ;
  assign y4368 = n22496 ;
  assign y4369 = n22500 ;
  assign y4370 = n22504 ;
  assign y4371 = n22505 ;
  assign y4372 = ~n22506 ;
  assign y4373 = ~n22508 ;
  assign y4374 = ~n22512 ;
  assign y4375 = ~n22514 ;
  assign y4376 = ~n22520 ;
  assign y4377 = ~n22521 ;
  assign y4378 = n22523 ;
  assign y4379 = n22525 ;
  assign y4380 = n22527 ;
  assign y4381 = ~n22528 ;
  assign y4382 = ~n22531 ;
  assign y4383 = n22533 ;
  assign y4384 = n22535 ;
  assign y4385 = ~n22536 ;
  assign y4386 = ~n22537 ;
  assign y4387 = n22539 ;
  assign y4388 = n22543 ;
  assign y4389 = ~n22544 ;
  assign y4390 = ~n22545 ;
  assign y4391 = n22549 ;
  assign y4392 = ~n22550 ;
  assign y4393 = n22555 ;
  assign y4394 = ~n22556 ;
  assign y4395 = n22558 ;
  assign y4396 = ~n22560 ;
  assign y4397 = n22562 ;
  assign y4398 = ~n22565 ;
  assign y4399 = n22569 ;
  assign y4400 = n22572 ;
  assign y4401 = n22575 ;
  assign y4402 = ~n22576 ;
  assign y4403 = n22579 ;
  assign y4404 = ~n22581 ;
  assign y4405 = ~n22584 ;
  assign y4406 = ~n22585 ;
  assign y4407 = ~n22587 ;
  assign y4408 = ~n22589 ;
  assign y4409 = ~n22590 ;
  assign y4410 = n22591 ;
  assign y4411 = n22593 ;
  assign y4412 = n22595 ;
  assign y4413 = ~n22596 ;
  assign y4414 = n22597 ;
  assign y4415 = n22600 ;
  assign y4416 = ~n22605 ;
  assign y4417 = ~n22606 ;
  assign y4418 = ~n22608 ;
  assign y4419 = n22609 ;
  assign y4420 = ~n22611 ;
  assign y4421 = n22612 ;
  assign y4422 = ~n22616 ;
  assign y4423 = n22617 ;
  assign y4424 = ~n22618 ;
  assign y4425 = ~n22621 ;
  assign y4426 = n22623 ;
  assign y4427 = ~n22625 ;
  assign y4428 = ~n22626 ;
  assign y4429 = n22627 ;
  assign y4430 = n22633 ;
  assign y4431 = n22635 ;
  assign y4432 = n22639 ;
  assign y4433 = ~n22643 ;
  assign y4434 = ~n22648 ;
  assign y4435 = ~n22651 ;
  assign y4436 = ~n22653 ;
  assign y4437 = ~n22655 ;
  assign y4438 = n22658 ;
  assign y4439 = n22659 ;
  assign y4440 = n22661 ;
  assign y4441 = n22665 ;
  assign y4442 = ~n22666 ;
  assign y4443 = ~n22669 ;
  assign y4444 = n22675 ;
  assign y4445 = ~n22676 ;
  assign y4446 = ~n22679 ;
  assign y4447 = n22680 ;
  assign y4448 = n22682 ;
  assign y4449 = n22683 ;
  assign y4450 = ~n22690 ;
  assign y4451 = ~n22693 ;
  assign y4452 = n22694 ;
  assign y4453 = n22695 ;
  assign y4454 = ~n22697 ;
  assign y4455 = ~n22700 ;
  assign y4456 = ~n22701 ;
  assign y4457 = ~n22703 ;
  assign y4458 = n22704 ;
  assign y4459 = n22705 ;
  assign y4460 = n22709 ;
  assign y4461 = n22713 ;
  assign y4462 = n22714 ;
  assign y4463 = n22716 ;
  assign y4464 = n22721 ;
  assign y4465 = n22727 ;
  assign y4466 = ~n22729 ;
  assign y4467 = ~n22734 ;
  assign y4468 = n22735 ;
  assign y4469 = n22741 ;
  assign y4470 = n22742 ;
  assign y4471 = ~n22743 ;
  assign y4472 = n22744 ;
  assign y4473 = n22750 ;
  assign y4474 = ~n22753 ;
  assign y4475 = n22755 ;
  assign y4476 = n22756 ;
  assign y4477 = ~n22757 ;
  assign y4478 = n22761 ;
  assign y4479 = ~n22763 ;
  assign y4480 = n22765 ;
  assign y4481 = ~n22768 ;
  assign y4482 = n22775 ;
  assign y4483 = n22777 ;
  assign y4484 = n22780 ;
  assign y4485 = n22786 ;
  assign y4486 = n22787 ;
  assign y4487 = n22789 ;
  assign y4488 = ~n22791 ;
  assign y4489 = ~n22795 ;
  assign y4490 = ~n22797 ;
  assign y4491 = n22798 ;
  assign y4492 = ~n22801 ;
  assign y4493 = ~n22803 ;
  assign y4494 = ~n22805 ;
  assign y4495 = ~n22807 ;
  assign y4496 = ~n22808 ;
  assign y4497 = n22809 ;
  assign y4498 = n22810 ;
  assign y4499 = ~n22811 ;
  assign y4500 = ~n22815 ;
  assign y4501 = ~n22822 ;
  assign y4502 = n22824 ;
  assign y4503 = ~n22826 ;
  assign y4504 = n22829 ;
  assign y4505 = n22830 ;
  assign y4506 = ~n22831 ;
  assign y4507 = ~n22832 ;
  assign y4508 = ~n22833 ;
  assign y4509 = n22837 ;
  assign y4510 = n22841 ;
  assign y4511 = ~n22844 ;
  assign y4512 = n22845 ;
  assign y4513 = ~n22846 ;
  assign y4514 = ~n22848 ;
  assign y4515 = n22851 ;
  assign y4516 = ~n22854 ;
  assign y4517 = ~n22855 ;
  assign y4518 = ~n22856 ;
  assign y4519 = n22863 ;
  assign y4520 = n22864 ;
  assign y4521 = n22866 ;
  assign y4522 = n22869 ;
  assign y4523 = ~n22874 ;
  assign y4524 = ~n22876 ;
  assign y4525 = n22878 ;
  assign y4526 = ~n22880 ;
  assign y4527 = n22882 ;
  assign y4528 = ~n22883 ;
  assign y4529 = ~n22884 ;
  assign y4530 = n22885 ;
  assign y4531 = ~n22886 ;
  assign y4532 = n22889 ;
  assign y4533 = n22892 ;
  assign y4534 = n22895 ;
  assign y4535 = n22897 ;
  assign y4536 = n22900 ;
  assign y4537 = n22901 ;
  assign y4538 = ~n22902 ;
  assign y4539 = n22904 ;
  assign y4540 = n22913 ;
  assign y4541 = ~n22918 ;
  assign y4542 = n22921 ;
  assign y4543 = ~n22922 ;
  assign y4544 = ~n22923 ;
  assign y4545 = n22924 ;
  assign y4546 = ~n22928 ;
  assign y4547 = n22929 ;
  assign y4548 = ~n22931 ;
  assign y4549 = n22932 ;
  assign y4550 = ~n22933 ;
  assign y4551 = ~n22936 ;
  assign y4552 = n22937 ;
  assign y4553 = ~n22940 ;
  assign y4554 = n22943 ;
  assign y4555 = n22951 ;
  assign y4556 = n22952 ;
  assign y4557 = n22953 ;
  assign y4558 = n22954 ;
  assign y4559 = n22957 ;
  assign y4560 = n22958 ;
  assign y4561 = n22964 ;
  assign y4562 = ~n22966 ;
  assign y4563 = n22967 ;
  assign y4564 = n22977 ;
  assign y4565 = ~n22978 ;
  assign y4566 = ~n22982 ;
  assign y4567 = ~n22983 ;
  assign y4568 = ~n22984 ;
  assign y4569 = ~n22985 ;
  assign y4570 = ~n22988 ;
  assign y4571 = n22989 ;
  assign y4572 = ~n22991 ;
  assign y4573 = ~n22993 ;
  assign y4574 = ~n22994 ;
  assign y4575 = n22997 ;
  assign y4576 = n22999 ;
  assign y4577 = ~n23002 ;
  assign y4578 = ~n23004 ;
  assign y4579 = n23005 ;
  assign y4580 = ~n23007 ;
  assign y4581 = ~n23009 ;
  assign y4582 = n23014 ;
  assign y4583 = n23021 ;
  assign y4584 = n23025 ;
  assign y4585 = n23027 ;
  assign y4586 = ~n23030 ;
  assign y4587 = n23034 ;
  assign y4588 = ~n23039 ;
  assign y4589 = n23040 ;
  assign y4590 = n23044 ;
  assign y4591 = ~n23046 ;
  assign y4592 = n23047 ;
  assign y4593 = ~n23054 ;
  assign y4594 = ~n23056 ;
  assign y4595 = ~n23064 ;
  assign y4596 = ~n23065 ;
  assign y4597 = ~n23069 ;
  assign y4598 = n23072 ;
  assign y4599 = n23074 ;
  assign y4600 = ~n23075 ;
  assign y4601 = n23077 ;
  assign y4602 = ~n23081 ;
  assign y4603 = ~n23083 ;
  assign y4604 = ~n23090 ;
  assign y4605 = ~n23093 ;
  assign y4606 = ~n23094 ;
  assign y4607 = ~n23096 ;
  assign y4608 = ~n23098 ;
  assign y4609 = n23099 ;
  assign y4610 = ~n23101 ;
  assign y4611 = ~n23104 ;
  assign y4612 = n23106 ;
  assign y4613 = n23108 ;
  assign y4614 = n23109 ;
  assign y4615 = ~n23112 ;
  assign y4616 = n23113 ;
  assign y4617 = ~n23116 ;
  assign y4618 = ~n23118 ;
  assign y4619 = ~n23122 ;
  assign y4620 = ~n23126 ;
  assign y4621 = n23134 ;
  assign y4622 = ~n23135 ;
  assign y4623 = n23146 ;
  assign y4624 = ~n23147 ;
  assign y4625 = n23154 ;
  assign y4626 = n23156 ;
  assign y4627 = n23158 ;
  assign y4628 = n23162 ;
  assign y4629 = n23163 ;
  assign y4630 = n23165 ;
  assign y4631 = ~n23166 ;
  assign y4632 = ~n23168 ;
  assign y4633 = n23176 ;
  assign y4634 = n23178 ;
  assign y4635 = n23179 ;
  assign y4636 = n23181 ;
  assign y4637 = n23183 ;
  assign y4638 = ~n23188 ;
  assign y4639 = n23190 ;
  assign y4640 = n23201 ;
  assign y4641 = ~n23202 ;
  assign y4642 = ~n23203 ;
  assign y4643 = ~n23205 ;
  assign y4644 = n23208 ;
  assign y4645 = ~n23209 ;
  assign y4646 = n23211 ;
  assign y4647 = ~n23212 ;
  assign y4648 = ~n23214 ;
  assign y4649 = n23215 ;
  assign y4650 = ~n23218 ;
  assign y4651 = n23219 ;
  assign y4652 = ~n23221 ;
  assign y4653 = n23223 ;
  assign y4654 = ~n23228 ;
  assign y4655 = n23229 ;
  assign y4656 = n23230 ;
  assign y4657 = n23231 ;
  assign y4658 = ~n23232 ;
  assign y4659 = ~n23235 ;
  assign y4660 = ~n23237 ;
  assign y4661 = ~n23249 ;
  assign y4662 = ~n23254 ;
  assign y4663 = n23258 ;
  assign y4664 = n23262 ;
  assign y4665 = n23264 ;
  assign y4666 = n23267 ;
  assign y4667 = ~n23270 ;
  assign y4668 = ~n23274 ;
  assign y4669 = n23277 ;
  assign y4670 = ~n23279 ;
  assign y4671 = n23281 ;
  assign y4672 = ~n23283 ;
  assign y4673 = n23284 ;
  assign y4674 = n23285 ;
  assign y4675 = n23294 ;
  assign y4676 = n23295 ;
  assign y4677 = ~n23297 ;
  assign y4678 = n23301 ;
  assign y4679 = ~n23302 ;
  assign y4680 = ~n23305 ;
  assign y4681 = n23306 ;
  assign y4682 = ~n23307 ;
  assign y4683 = ~n23309 ;
  assign y4684 = n23317 ;
  assign y4685 = ~n23318 ;
  assign y4686 = n23319 ;
  assign y4687 = ~n23327 ;
  assign y4688 = ~n23328 ;
  assign y4689 = n23332 ;
  assign y4690 = n23337 ;
  assign y4691 = n23343 ;
  assign y4692 = ~n23344 ;
  assign y4693 = n23346 ;
  assign y4694 = n23352 ;
  assign y4695 = ~n23353 ;
  assign y4696 = ~n23358 ;
  assign y4697 = ~n23361 ;
  assign y4698 = n23364 ;
  assign y4699 = n23366 ;
  assign y4700 = n23367 ;
  assign y4701 = n23369 ;
  assign y4702 = ~n23372 ;
  assign y4703 = ~n23374 ;
  assign y4704 = ~n23377 ;
  assign y4705 = ~n23380 ;
  assign y4706 = ~n23382 ;
  assign y4707 = n23384 ;
  assign y4708 = n23385 ;
  assign y4709 = ~n23386 ;
  assign y4710 = n23391 ;
  assign y4711 = n23397 ;
  assign y4712 = ~n23398 ;
  assign y4713 = ~n23402 ;
  assign y4714 = n23403 ;
  assign y4715 = n23410 ;
  assign y4716 = n23412 ;
  assign y4717 = ~n23413 ;
  assign y4718 = ~n23414 ;
  assign y4719 = ~n23416 ;
  assign y4720 = ~n23417 ;
  assign y4721 = ~n23425 ;
  assign y4722 = ~n23427 ;
  assign y4723 = ~n23429 ;
  assign y4724 = ~n23430 ;
  assign y4725 = n23432 ;
  assign y4726 = n23436 ;
  assign y4727 = ~n23437 ;
  assign y4728 = ~n23440 ;
  assign y4729 = ~n23442 ;
  assign y4730 = n23445 ;
  assign y4731 = n23446 ;
  assign y4732 = n23450 ;
  assign y4733 = ~n23455 ;
  assign y4734 = n23461 ;
  assign y4735 = n23471 ;
  assign y4736 = ~n23475 ;
  assign y4737 = n23476 ;
  assign y4738 = ~n23477 ;
  assign y4739 = ~n23479 ;
  assign y4740 = ~n23480 ;
  assign y4741 = ~n23482 ;
  assign y4742 = ~n23486 ;
  assign y4743 = ~n23487 ;
  assign y4744 = ~n23488 ;
  assign y4745 = ~n23491 ;
  assign y4746 = n23493 ;
  assign y4747 = n23496 ;
  assign y4748 = n23501 ;
  assign y4749 = ~n23503 ;
  assign y4750 = ~n23504 ;
  assign y4751 = n23507 ;
  assign y4752 = n23508 ;
  assign y4753 = ~n23509 ;
  assign y4754 = n23512 ;
  assign y4755 = n23513 ;
  assign y4756 = n23514 ;
  assign y4757 = ~n23517 ;
  assign y4758 = n23518 ;
  assign y4759 = n23524 ;
  assign y4760 = n23527 ;
  assign y4761 = n23528 ;
  assign y4762 = n23529 ;
  assign y4763 = ~n23535 ;
  assign y4764 = n23538 ;
  assign y4765 = n23542 ;
  assign y4766 = ~n23544 ;
  assign y4767 = ~n23546 ;
  assign y4768 = ~n23547 ;
  assign y4769 = n23548 ;
  assign y4770 = n23551 ;
  assign y4771 = ~n23553 ;
  assign y4772 = ~n23555 ;
  assign y4773 = ~n23556 ;
  assign y4774 = n23560 ;
  assign y4775 = ~n23565 ;
  assign y4776 = ~n23567 ;
  assign y4777 = n23571 ;
  assign y4778 = ~n23574 ;
  assign y4779 = n23578 ;
  assign y4780 = ~n23581 ;
  assign y4781 = n23583 ;
  assign y4782 = ~n23585 ;
  assign y4783 = ~n23588 ;
  assign y4784 = ~n23591 ;
  assign y4785 = n23593 ;
  assign y4786 = n23594 ;
  assign y4787 = n23601 ;
  assign y4788 = ~n23603 ;
  assign y4789 = n23606 ;
  assign y4790 = ~n23610 ;
  assign y4791 = ~n23612 ;
  assign y4792 = n23613 ;
  assign y4793 = ~n23614 ;
  assign y4794 = ~n23616 ;
  assign y4795 = n23620 ;
  assign y4796 = ~n23626 ;
  assign y4797 = ~n23627 ;
  assign y4798 = ~n23632 ;
  assign y4799 = n23636 ;
  assign y4800 = ~n23637 ;
  assign y4801 = n23638 ;
  assign y4802 = ~n23639 ;
  assign y4803 = n23643 ;
  assign y4804 = ~n23645 ;
  assign y4805 = n23647 ;
  assign y4806 = n23648 ;
  assign y4807 = ~n23650 ;
  assign y4808 = n23652 ;
  assign y4809 = ~n23653 ;
  assign y4810 = ~n23655 ;
  assign y4811 = ~n23656 ;
  assign y4812 = n23657 ;
  assign y4813 = n23658 ;
  assign y4814 = ~n23665 ;
  assign y4815 = ~n23668 ;
  assign y4816 = n23671 ;
  assign y4817 = ~n23674 ;
  assign y4818 = ~n23676 ;
  assign y4819 = ~n23679 ;
  assign y4820 = n23680 ;
  assign y4821 = ~n23682 ;
  assign y4822 = ~n23683 ;
  assign y4823 = ~n23685 ;
  assign y4824 = ~n23692 ;
  assign y4825 = ~n23695 ;
  assign y4826 = ~n23701 ;
  assign y4827 = n23702 ;
  assign y4828 = n23707 ;
  assign y4829 = ~n23708 ;
  assign y4830 = ~n23710 ;
  assign y4831 = n23711 ;
  assign y4832 = n23712 ;
  assign y4833 = ~n23713 ;
  assign y4834 = n23714 ;
  assign y4835 = n23716 ;
  assign y4836 = ~n23720 ;
  assign y4837 = ~n23723 ;
  assign y4838 = n23727 ;
  assign y4839 = n23728 ;
  assign y4840 = n23732 ;
  assign y4841 = ~n23740 ;
  assign y4842 = n23744 ;
  assign y4843 = ~n23745 ;
  assign y4844 = n23752 ;
  assign y4845 = ~n23754 ;
  assign y4846 = n23760 ;
  assign y4847 = n23762 ;
  assign y4848 = n23767 ;
  assign y4849 = ~n23771 ;
  assign y4850 = ~n23772 ;
  assign y4851 = ~n23774 ;
  assign y4852 = ~n23780 ;
  assign y4853 = n23782 ;
  assign y4854 = n23785 ;
  assign y4855 = n23788 ;
  assign y4856 = n23789 ;
  assign y4857 = n23792 ;
  assign y4858 = n23796 ;
  assign y4859 = ~n23798 ;
  assign y4860 = ~n23800 ;
  assign y4861 = ~n23804 ;
  assign y4862 = ~n23806 ;
  assign y4863 = ~n23807 ;
  assign y4864 = n23811 ;
  assign y4865 = n23812 ;
  assign y4866 = ~n23813 ;
  assign y4867 = n23814 ;
  assign y4868 = ~n23815 ;
  assign y4869 = n23819 ;
  assign y4870 = ~n23823 ;
  assign y4871 = ~n23832 ;
  assign y4872 = ~n23833 ;
  assign y4873 = ~n23834 ;
  assign y4874 = n23836 ;
  assign y4875 = n23838 ;
  assign y4876 = n23844 ;
  assign y4877 = ~n23845 ;
  assign y4878 = ~n23847 ;
  assign y4879 = n23850 ;
  assign y4880 = ~n23853 ;
  assign y4881 = n23856 ;
  assign y4882 = n23857 ;
  assign y4883 = ~n23858 ;
  assign y4884 = ~n23859 ;
  assign y4885 = ~n23862 ;
  assign y4886 = n23864 ;
  assign y4887 = n23866 ;
  assign y4888 = ~n23869 ;
  assign y4889 = n23870 ;
  assign y4890 = ~n23872 ;
  assign y4891 = n23879 ;
  assign y4892 = n23883 ;
  assign y4893 = ~n23885 ;
  assign y4894 = ~n23886 ;
  assign y4895 = n23889 ;
  assign y4896 = ~n23890 ;
  assign y4897 = ~n23894 ;
  assign y4898 = ~n23896 ;
  assign y4899 = n23897 ;
  assign y4900 = n23898 ;
  assign y4901 = ~n23905 ;
  assign y4902 = ~n23910 ;
  assign y4903 = ~n23911 ;
  assign y4904 = ~n23913 ;
  assign y4905 = n23914 ;
  assign y4906 = n23915 ;
  assign y4907 = ~n23918 ;
  assign y4908 = ~n23921 ;
  assign y4909 = ~n23925 ;
  assign y4910 = n23927 ;
  assign y4911 = ~n23928 ;
  assign y4912 = n23929 ;
  assign y4913 = ~n23930 ;
  assign y4914 = n23931 ;
  assign y4915 = ~n23932 ;
  assign y4916 = ~n23934 ;
  assign y4917 = n23936 ;
  assign y4918 = n23941 ;
  assign y4919 = ~n23942 ;
  assign y4920 = n23951 ;
  assign y4921 = ~n23952 ;
  assign y4922 = n23958 ;
  assign y4923 = ~n23963 ;
  assign y4924 = ~n23968 ;
  assign y4925 = n23969 ;
  assign y4926 = ~n23975 ;
  assign y4927 = ~n23979 ;
  assign y4928 = ~n23982 ;
  assign y4929 = n23985 ;
  assign y4930 = ~n23987 ;
  assign y4931 = n23989 ;
  assign y4932 = ~n23991 ;
  assign y4933 = ~n23992 ;
  assign y4934 = ~n23996 ;
  assign y4935 = ~n23998 ;
  assign y4936 = ~n24000 ;
  assign y4937 = ~n24001 ;
  assign y4938 = n24005 ;
  assign y4939 = ~n24009 ;
  assign y4940 = n24011 ;
  assign y4941 = ~n24015 ;
  assign y4942 = ~n24018 ;
  assign y4943 = n24021 ;
  assign y4944 = n24023 ;
  assign y4945 = ~n24024 ;
  assign y4946 = n24025 ;
  assign y4947 = n24027 ;
  assign y4948 = ~n24031 ;
  assign y4949 = n24034 ;
  assign y4950 = n24040 ;
  assign y4951 = ~n24041 ;
  assign y4952 = ~n24044 ;
  assign y4953 = ~n24045 ;
  assign y4954 = n24048 ;
  assign y4955 = n24051 ;
  assign y4956 = n24052 ;
  assign y4957 = ~n24057 ;
  assign y4958 = ~n24061 ;
  assign y4959 = ~n24063 ;
  assign y4960 = ~n24065 ;
  assign y4961 = n24066 ;
  assign y4962 = ~n24070 ;
  assign y4963 = n24072 ;
  assign y4964 = n24081 ;
  assign y4965 = n24085 ;
  assign y4966 = ~n24089 ;
  assign y4967 = ~n24093 ;
  assign y4968 = n24096 ;
  assign y4969 = n24100 ;
  assign y4970 = ~n24102 ;
  assign y4971 = n24105 ;
  assign y4972 = n24112 ;
  assign y4973 = n24114 ;
  assign y4974 = n24116 ;
  assign y4975 = ~n24117 ;
  assign y4976 = ~n24119 ;
  assign y4977 = ~n24122 ;
  assign y4978 = ~n24124 ;
  assign y4979 = n24128 ;
  assign y4980 = n24130 ;
  assign y4981 = ~n24131 ;
  assign y4982 = ~n24133 ;
  assign y4983 = n24137 ;
  assign y4984 = ~n24138 ;
  assign y4985 = ~n24139 ;
  assign y4986 = n24142 ;
  assign y4987 = n24143 ;
  assign y4988 = ~n24144 ;
  assign y4989 = ~n24146 ;
  assign y4990 = n24147 ;
  assign y4991 = ~n24148 ;
  assign y4992 = n24150 ;
  assign y4993 = n24152 ;
  assign y4994 = ~n24153 ;
  assign y4995 = n24158 ;
  assign y4996 = ~n24165 ;
  assign y4997 = n24168 ;
  assign y4998 = ~n24169 ;
  assign y4999 = n24170 ;
  assign y5000 = n24172 ;
  assign y5001 = ~n24174 ;
  assign y5002 = n24177 ;
  assign y5003 = n24179 ;
  assign y5004 = n24182 ;
  assign y5005 = ~n24183 ;
  assign y5006 = n24184 ;
  assign y5007 = ~n24185 ;
  assign y5008 = n24186 ;
  assign y5009 = ~n24188 ;
  assign y5010 = ~n24191 ;
  assign y5011 = n24192 ;
  assign y5012 = n24194 ;
  assign y5013 = ~n24202 ;
  assign y5014 = ~n24208 ;
  assign y5015 = n24209 ;
  assign y5016 = n24210 ;
  assign y5017 = n24212 ;
  assign y5018 = n24218 ;
  assign y5019 = n24220 ;
  assign y5020 = ~n24223 ;
  assign y5021 = n24224 ;
  assign y5022 = ~n24226 ;
  assign y5023 = ~n24227 ;
  assign y5024 = n24228 ;
  assign y5025 = n24229 ;
  assign y5026 = n24235 ;
  assign y5027 = n24237 ;
  assign y5028 = ~n24239 ;
  assign y5029 = n24243 ;
  assign y5030 = n24246 ;
  assign y5031 = ~n24247 ;
  assign y5032 = ~n24249 ;
  assign y5033 = ~n24256 ;
  assign y5034 = ~n24259 ;
  assign y5035 = n24261 ;
  assign y5036 = ~n24263 ;
  assign y5037 = n24265 ;
  assign y5038 = ~n24266 ;
  assign y5039 = n24267 ;
  assign y5040 = ~n24272 ;
  assign y5041 = n24277 ;
  assign y5042 = ~n24278 ;
  assign y5043 = n24279 ;
  assign y5044 = n24281 ;
  assign y5045 = n24286 ;
  assign y5046 = ~n24290 ;
  assign y5047 = n24293 ;
  assign y5048 = n24298 ;
  assign y5049 = ~n24301 ;
  assign y5050 = n24303 ;
  assign y5051 = n24306 ;
  assign y5052 = n24309 ;
  assign y5053 = n24310 ;
  assign y5054 = ~n24311 ;
  assign y5055 = n24314 ;
  assign y5056 = n24317 ;
  assign y5057 = n24322 ;
  assign y5058 = n24324 ;
  assign y5059 = n24325 ;
  assign y5060 = ~n24326 ;
  assign y5061 = ~n24327 ;
  assign y5062 = ~n24328 ;
  assign y5063 = ~n24329 ;
  assign y5064 = ~n24331 ;
  assign y5065 = n24332 ;
  assign y5066 = ~n24333 ;
  assign y5067 = n24334 ;
  assign y5068 = ~n24337 ;
  assign y5069 = ~n24338 ;
  assign y5070 = ~n24341 ;
  assign y5071 = n24342 ;
  assign y5072 = n24345 ;
  assign y5073 = ~n24346 ;
  assign y5074 = n24349 ;
  assign y5075 = n24359 ;
  assign y5076 = n24365 ;
  assign y5077 = ~n24367 ;
  assign y5078 = ~n24369 ;
  assign y5079 = ~n24372 ;
  assign y5080 = n24373 ;
  assign y5081 = n24375 ;
  assign y5082 = ~n24376 ;
  assign y5083 = n24379 ;
  assign y5084 = ~n24382 ;
  assign y5085 = ~n24383 ;
  assign y5086 = n24385 ;
  assign y5087 = ~n24389 ;
  assign y5088 = n24392 ;
  assign y5089 = ~n24393 ;
  assign y5090 = ~n24395 ;
  assign y5091 = ~n24400 ;
  assign y5092 = n24401 ;
  assign y5093 = ~n24404 ;
  assign y5094 = ~n24405 ;
  assign y5095 = ~n24406 ;
  assign y5096 = ~n24407 ;
  assign y5097 = ~n24410 ;
  assign y5098 = n24413 ;
  assign y5099 = n24418 ;
  assign y5100 = n24419 ;
  assign y5101 = n24422 ;
  assign y5102 = ~n24427 ;
  assign y5103 = ~n24432 ;
  assign y5104 = n24434 ;
  assign y5105 = ~n24438 ;
  assign y5106 = n24441 ;
  assign y5107 = ~n24442 ;
  assign y5108 = ~n24443 ;
  assign y5109 = n24448 ;
  assign y5110 = ~n24451 ;
  assign y5111 = n24452 ;
  assign y5112 = n24454 ;
  assign y5113 = ~n24456 ;
  assign y5114 = ~n24460 ;
  assign y5115 = n24464 ;
  assign y5116 = n24466 ;
  assign y5117 = ~n24467 ;
  assign y5118 = ~n24471 ;
  assign y5119 = ~n24475 ;
  assign y5120 = ~n24476 ;
  assign y5121 = ~n24480 ;
  assign y5122 = ~n24481 ;
  assign y5123 = ~n24483 ;
  assign y5124 = ~n24485 ;
  assign y5125 = n24486 ;
  assign y5126 = ~n24487 ;
  assign y5127 = ~n24493 ;
  assign y5128 = ~n24494 ;
  assign y5129 = n24498 ;
  assign y5130 = n24500 ;
  assign y5131 = n24502 ;
  assign y5132 = ~n24506 ;
  assign y5133 = n24510 ;
  assign y5134 = n24511 ;
  assign y5135 = n24512 ;
  assign y5136 = n24514 ;
  assign y5137 = ~n24519 ;
  assign y5138 = ~n24523 ;
  assign y5139 = ~n24524 ;
  assign y5140 = ~n24526 ;
  assign y5141 = ~n24530 ;
  assign y5142 = ~n24531 ;
  assign y5143 = n24532 ;
  assign y5144 = n24533 ;
  assign y5145 = ~n24535 ;
  assign y5146 = ~n24537 ;
  assign y5147 = ~n24539 ;
  assign y5148 = n24542 ;
  assign y5149 = n24543 ;
  assign y5150 = ~n24544 ;
  assign y5151 = n24545 ;
  assign y5152 = n24548 ;
  assign y5153 = n24549 ;
  assign y5154 = ~n24553 ;
  assign y5155 = n24559 ;
  assign y5156 = n24562 ;
  assign y5157 = ~n24568 ;
  assign y5158 = n24571 ;
  assign y5159 = ~n24573 ;
  assign y5160 = ~n24574 ;
  assign y5161 = n24575 ;
  assign y5162 = ~n24579 ;
  assign y5163 = ~n24580 ;
  assign y5164 = n24582 ;
  assign y5165 = ~n24587 ;
  assign y5166 = ~n24588 ;
  assign y5167 = ~n24590 ;
  assign y5168 = n24592 ;
  assign y5169 = n24594 ;
  assign y5170 = ~n24595 ;
  assign y5171 = n24596 ;
  assign y5172 = ~n24599 ;
  assign y5173 = ~n24600 ;
  assign y5174 = n24603 ;
  assign y5175 = ~n24606 ;
  assign y5176 = ~n24612 ;
  assign y5177 = ~n24615 ;
  assign y5178 = n24618 ;
  assign y5179 = ~n24620 ;
  assign y5180 = n24621 ;
  assign y5181 = ~n24623 ;
  assign y5182 = ~n24625 ;
  assign y5183 = n24632 ;
  assign y5184 = ~n24633 ;
  assign y5185 = ~n24634 ;
  assign y5186 = n24637 ;
  assign y5187 = ~n24638 ;
  assign y5188 = n24641 ;
  assign y5189 = n24642 ;
  assign y5190 = n24646 ;
  assign y5191 = n24648 ;
  assign y5192 = n24649 ;
  assign y5193 = n24652 ;
  assign y5194 = n24654 ;
  assign y5195 = ~n24657 ;
  assign y5196 = ~n24661 ;
  assign y5197 = ~n24665 ;
  assign y5198 = n24669 ;
  assign y5199 = n24670 ;
  assign y5200 = ~n24672 ;
  assign y5201 = n24673 ;
  assign y5202 = ~n24674 ;
  assign y5203 = n24676 ;
  assign y5204 = n24677 ;
  assign y5205 = ~n24678 ;
  assign y5206 = ~n24680 ;
  assign y5207 = ~n24683 ;
  assign y5208 = ~n24686 ;
  assign y5209 = n24687 ;
  assign y5210 = ~n24689 ;
  assign y5211 = ~n24692 ;
  assign y5212 = n24694 ;
  assign y5213 = n24695 ;
  assign y5214 = ~n24698 ;
  assign y5215 = n24699 ;
  assign y5216 = n24700 ;
  assign y5217 = n24703 ;
  assign y5218 = ~n24709 ;
  assign y5219 = ~n24712 ;
  assign y5220 = ~n24713 ;
  assign y5221 = n24719 ;
  assign y5222 = n24722 ;
  assign y5223 = ~n24727 ;
  assign y5224 = n24728 ;
  assign y5225 = ~n24735 ;
  assign y5226 = n24739 ;
  assign y5227 = ~n24741 ;
  assign y5228 = ~n24742 ;
  assign y5229 = ~n24745 ;
  assign y5230 = n24747 ;
  assign y5231 = n24749 ;
  assign y5232 = n24750 ;
  assign y5233 = n24751 ;
  assign y5234 = n24752 ;
  assign y5235 = ~n24755 ;
  assign y5236 = ~n24758 ;
  assign y5237 = n24759 ;
  assign y5238 = n24760 ;
  assign y5239 = ~n24762 ;
  assign y5240 = n24767 ;
  assign y5241 = ~n24771 ;
  assign y5242 = n24772 ;
  assign y5243 = ~n24774 ;
  assign y5244 = ~n24777 ;
  assign y5245 = ~n24782 ;
  assign y5246 = ~n24785 ;
  assign y5247 = ~n24787 ;
  assign y5248 = n24791 ;
  assign y5249 = ~n24794 ;
  assign y5250 = n24796 ;
  assign y5251 = ~n24799 ;
  assign y5252 = ~n24815 ;
  assign y5253 = ~n24818 ;
  assign y5254 = n24821 ;
  assign y5255 = ~n24822 ;
  assign y5256 = ~n24825 ;
  assign y5257 = ~n24827 ;
  assign y5258 = n24834 ;
  assign y5259 = ~n24837 ;
  assign y5260 = ~n24840 ;
  assign y5261 = n24842 ;
  assign y5262 = ~n24844 ;
  assign y5263 = n24845 ;
  assign y5264 = n24847 ;
  assign y5265 = n24848 ;
  assign y5266 = ~n24849 ;
  assign y5267 = n24850 ;
  assign y5268 = n24855 ;
  assign y5269 = n24857 ;
  assign y5270 = n24860 ;
  assign y5271 = n24861 ;
  assign y5272 = n24862 ;
  assign y5273 = ~n24864 ;
  assign y5274 = ~n24865 ;
  assign y5275 = n24866 ;
  assign y5276 = n24871 ;
  assign y5277 = ~n24872 ;
  assign y5278 = ~n24873 ;
  assign y5279 = ~n24876 ;
  assign y5280 = n24878 ;
  assign y5281 = ~n24880 ;
  assign y5282 = n24881 ;
  assign y5283 = ~n24886 ;
  assign y5284 = n24889 ;
  assign y5285 = n24890 ;
  assign y5286 = ~n24892 ;
  assign y5287 = ~n24893 ;
  assign y5288 = n24894 ;
  assign y5289 = n24895 ;
  assign y5290 = ~n24898 ;
  assign y5291 = n24902 ;
  assign y5292 = n24904 ;
  assign y5293 = n24906 ;
  assign y5294 = ~n24907 ;
  assign y5295 = n24908 ;
  assign y5296 = ~n24909 ;
  assign y5297 = ~n24911 ;
  assign y5298 = ~n24915 ;
  assign y5299 = ~n24916 ;
  assign y5300 = n24917 ;
  assign y5301 = n24918 ;
  assign y5302 = n24920 ;
  assign y5303 = n24923 ;
  assign y5304 = n24925 ;
  assign y5305 = n24929 ;
  assign y5306 = ~n24932 ;
  assign y5307 = n24933 ;
  assign y5308 = ~n24935 ;
  assign y5309 = n24939 ;
  assign y5310 = n24945 ;
  assign y5311 = ~n24947 ;
  assign y5312 = n24952 ;
  assign y5313 = ~n24955 ;
  assign y5314 = ~n24957 ;
  assign y5315 = ~n24959 ;
  assign y5316 = n24960 ;
  assign y5317 = n24961 ;
  assign y5318 = ~n24963 ;
  assign y5319 = ~n24964 ;
  assign y5320 = n24965 ;
  assign y5321 = n24966 ;
  assign y5322 = n24973 ;
  assign y5323 = ~n24974 ;
  assign y5324 = n24976 ;
  assign y5325 = ~n24979 ;
  assign y5326 = n24980 ;
  assign y5327 = ~n24981 ;
  assign y5328 = ~n24983 ;
  assign y5329 = ~n24984 ;
  assign y5330 = ~n24985 ;
  assign y5331 = ~n24988 ;
  assign y5332 = n24992 ;
  assign y5333 = n24993 ;
  assign y5334 = n24994 ;
  assign y5335 = ~n24995 ;
  assign y5336 = n24997 ;
  assign y5337 = n24999 ;
  assign y5338 = n25004 ;
  assign y5339 = ~n25009 ;
  assign y5340 = n25012 ;
  assign y5341 = ~n25013 ;
  assign y5342 = n25015 ;
  assign y5343 = ~n25016 ;
  assign y5344 = ~n25017 ;
  assign y5345 = ~n25018 ;
  assign y5346 = ~n25019 ;
  assign y5347 = n25021 ;
  assign y5348 = n25023 ;
  assign y5349 = n25025 ;
  assign y5350 = n25029 ;
  assign y5351 = n25030 ;
  assign y5352 = ~n25037 ;
  assign y5353 = n25038 ;
  assign y5354 = ~n25040 ;
  assign y5355 = n25043 ;
  assign y5356 = n25046 ;
  assign y5357 = ~n25049 ;
  assign y5358 = ~n25051 ;
  assign y5359 = n25054 ;
  assign y5360 = n25055 ;
  assign y5361 = n25057 ;
  assign y5362 = n25058 ;
  assign y5363 = ~n25059 ;
  assign y5364 = ~n25061 ;
  assign y5365 = n25065 ;
  assign y5366 = n25068 ;
  assign y5367 = ~n25076 ;
  assign y5368 = n25077 ;
  assign y5369 = n25078 ;
  assign y5370 = ~n25079 ;
  assign y5371 = n25080 ;
  assign y5372 = n25084 ;
  assign y5373 = ~n25087 ;
  assign y5374 = n25088 ;
  assign y5375 = n25089 ;
  assign y5376 = n25090 ;
  assign y5377 = ~n25091 ;
  assign y5378 = ~n25096 ;
  assign y5379 = ~n25099 ;
  assign y5380 = ~n25100 ;
  assign y5381 = ~n25103 ;
  assign y5382 = ~n25104 ;
  assign y5383 = n25108 ;
  assign y5384 = n25115 ;
  assign y5385 = ~n25117 ;
  assign y5386 = n25119 ;
  assign y5387 = ~n25120 ;
  assign y5388 = ~n25121 ;
  assign y5389 = n25122 ;
  assign y5390 = n25124 ;
  assign y5391 = n25127 ;
  assign y5392 = n25128 ;
  assign y5393 = n25129 ;
  assign y5394 = ~n25131 ;
  assign y5395 = n25134 ;
  assign y5396 = n25135 ;
  assign y5397 = ~n25136 ;
  assign y5398 = ~n25142 ;
  assign y5399 = ~n25145 ;
  assign y5400 = ~n25149 ;
  assign y5401 = ~n25150 ;
  assign y5402 = n25151 ;
  assign y5403 = ~n25156 ;
  assign y5404 = ~n25157 ;
  assign y5405 = n25164 ;
  assign y5406 = ~n25166 ;
  assign y5407 = n25168 ;
  assign y5408 = ~n25169 ;
  assign y5409 = ~n25170 ;
  assign y5410 = ~n25171 ;
  assign y5411 = n25174 ;
  assign y5412 = n25183 ;
  assign y5413 = ~n25187 ;
  assign y5414 = n25189 ;
  assign y5415 = ~n25190 ;
  assign y5416 = n25191 ;
  assign y5417 = n25192 ;
  assign y5418 = n25198 ;
  assign y5419 = ~n25203 ;
  assign y5420 = n25204 ;
  assign y5421 = n25206 ;
  assign y5422 = ~n25208 ;
  assign y5423 = ~n25216 ;
  assign y5424 = ~n25217 ;
  assign y5425 = n25218 ;
  assign y5426 = ~n25222 ;
  assign y5427 = n25223 ;
  assign y5428 = ~n25225 ;
  assign y5429 = n25227 ;
  assign y5430 = ~n25229 ;
  assign y5431 = ~n25231 ;
  assign y5432 = ~n25233 ;
  assign y5433 = n25234 ;
  assign y5434 = ~n25235 ;
  assign y5435 = ~n25237 ;
  assign y5436 = n25242 ;
  assign y5437 = ~n25243 ;
  assign y5438 = ~n25245 ;
  assign y5439 = ~n25249 ;
  assign y5440 = n25250 ;
  assign y5441 = n25251 ;
  assign y5442 = ~n25256 ;
  assign y5443 = ~n25260 ;
  assign y5444 = n25261 ;
  assign y5445 = ~n25265 ;
  assign y5446 = ~n25266 ;
  assign y5447 = n25269 ;
  assign y5448 = n25270 ;
  assign y5449 = n25271 ;
  assign y5450 = ~n25272 ;
  assign y5451 = n25274 ;
  assign y5452 = n25276 ;
  assign y5453 = ~n25277 ;
  assign y5454 = n25278 ;
  assign y5455 = n25282 ;
  assign y5456 = n25289 ;
  assign y5457 = n25291 ;
  assign y5458 = ~n25293 ;
  assign y5459 = ~n25300 ;
  assign y5460 = n25301 ;
  assign y5461 = n25303 ;
  assign y5462 = ~n25304 ;
  assign y5463 = n25305 ;
  assign y5464 = n25306 ;
  assign y5465 = n25307 ;
  assign y5466 = n25309 ;
  assign y5467 = ~n25310 ;
  assign y5468 = n25315 ;
  assign y5469 = ~n25316 ;
  assign y5470 = n25317 ;
  assign y5471 = ~n25318 ;
  assign y5472 = n25319 ;
  assign y5473 = n25322 ;
  assign y5474 = ~n25323 ;
  assign y5475 = ~n25325 ;
  assign y5476 = ~n25331 ;
  assign y5477 = ~n25334 ;
  assign y5478 = ~n25335 ;
  assign y5479 = ~n25336 ;
  assign y5480 = ~n25344 ;
  assign y5481 = n25345 ;
  assign y5482 = n25347 ;
  assign y5483 = n25349 ;
  assign y5484 = n25358 ;
  assign y5485 = n25359 ;
  assign y5486 = n25360 ;
  assign y5487 = ~n25364 ;
  assign y5488 = ~n25365 ;
  assign y5489 = ~n25375 ;
  assign y5490 = ~n25382 ;
  assign y5491 = ~n25383 ;
  assign y5492 = n25385 ;
  assign y5493 = n25387 ;
  assign y5494 = ~n25393 ;
  assign y5495 = ~n25394 ;
  assign y5496 = n25395 ;
  assign y5497 = ~n25397 ;
  assign y5498 = n25399 ;
  assign y5499 = n25402 ;
  assign y5500 = n25408 ;
  assign y5501 = n25410 ;
  assign y5502 = n25411 ;
  assign y5503 = ~n25413 ;
  assign y5504 = n25417 ;
  assign y5505 = n25419 ;
  assign y5506 = n25420 ;
  assign y5507 = n25421 ;
  assign y5508 = n25423 ;
  assign y5509 = ~n25425 ;
  assign y5510 = n25430 ;
  assign y5511 = n25434 ;
  assign y5512 = n25437 ;
  assign y5513 = n25439 ;
  assign y5514 = n25441 ;
  assign y5515 = ~n25445 ;
  assign y5516 = n25448 ;
  assign y5517 = ~n25449 ;
  assign y5518 = ~n25451 ;
  assign y5519 = ~n25452 ;
  assign y5520 = n25454 ;
  assign y5521 = n25456 ;
  assign y5522 = n25458 ;
  assign y5523 = n25462 ;
  assign y5524 = n25464 ;
  assign y5525 = ~n25466 ;
  assign y5526 = ~n25469 ;
  assign y5527 = ~n25471 ;
  assign y5528 = n25476 ;
  assign y5529 = n25477 ;
  assign y5530 = n25479 ;
  assign y5531 = ~n25480 ;
  assign y5532 = ~n25481 ;
  assign y5533 = n25485 ;
  assign y5534 = n25488 ;
  assign y5535 = ~n25489 ;
  assign y5536 = ~n25491 ;
  assign y5537 = ~n25493 ;
  assign y5538 = ~n25496 ;
  assign y5539 = ~n25497 ;
  assign y5540 = n25501 ;
  assign y5541 = n25506 ;
  assign y5542 = n25510 ;
  assign y5543 = n25512 ;
  assign y5544 = n25521 ;
  assign y5545 = ~n25524 ;
  assign y5546 = ~n25526 ;
  assign y5547 = ~n25527 ;
  assign y5548 = ~n25528 ;
  assign y5549 = n25530 ;
  assign y5550 = n25532 ;
  assign y5551 = ~n25533 ;
  assign y5552 = n25535 ;
  assign y5553 = n25537 ;
  assign y5554 = n25540 ;
  assign y5555 = ~n25541 ;
  assign y5556 = ~n25543 ;
  assign y5557 = n25544 ;
  assign y5558 = ~n25545 ;
  assign y5559 = n25548 ;
  assign y5560 = ~n25551 ;
  assign y5561 = ~n25555 ;
  assign y5562 = ~n25556 ;
  assign y5563 = ~n25557 ;
  assign y5564 = n25562 ;
  assign y5565 = ~n25565 ;
  assign y5566 = ~n25571 ;
  assign y5567 = ~n25575 ;
  assign y5568 = n25579 ;
  assign y5569 = n25583 ;
  assign y5570 = n25587 ;
  assign y5571 = n25594 ;
  assign y5572 = n25598 ;
  assign y5573 = n25600 ;
  assign y5574 = ~n25603 ;
  assign y5575 = ~n25606 ;
  assign y5576 = n25607 ;
  assign y5577 = ~n25610 ;
  assign y5578 = n25613 ;
  assign y5579 = ~n25615 ;
  assign y5580 = ~n25618 ;
  assign y5581 = n25620 ;
  assign y5582 = n25626 ;
  assign y5583 = ~n25627 ;
  assign y5584 = n25629 ;
  assign y5585 = ~n25635 ;
  assign y5586 = ~n25638 ;
  assign y5587 = ~n25643 ;
  assign y5588 = n25644 ;
  assign y5589 = n25648 ;
  assign y5590 = n25650 ;
  assign y5591 = ~n25651 ;
  assign y5592 = ~n25659 ;
  assign y5593 = ~n25660 ;
  assign y5594 = ~n25663 ;
  assign y5595 = ~n25666 ;
  assign y5596 = ~n25668 ;
  assign y5597 = ~n25670 ;
  assign y5598 = ~n25672 ;
  assign y5599 = n25673 ;
  assign y5600 = n25675 ;
  assign y5601 = n25676 ;
  assign y5602 = ~n25677 ;
  assign y5603 = ~n25678 ;
  assign y5604 = ~n25679 ;
  assign y5605 = n25681 ;
  assign y5606 = n25684 ;
  assign y5607 = n25687 ;
  assign y5608 = ~n25688 ;
  assign y5609 = n25691 ;
  assign y5610 = n25694 ;
  assign y5611 = n25697 ;
  assign y5612 = ~n25707 ;
  assign y5613 = ~n25708 ;
  assign y5614 = n25713 ;
  assign y5615 = ~n25715 ;
  assign y5616 = n25719 ;
  assign y5617 = ~n25721 ;
  assign y5618 = n25722 ;
  assign y5619 = n25723 ;
  assign y5620 = ~n25728 ;
  assign y5621 = n25730 ;
  assign y5622 = n25731 ;
  assign y5623 = n25732 ;
  assign y5624 = ~n25734 ;
  assign y5625 = n25735 ;
  assign y5626 = ~n25739 ;
  assign y5627 = ~n25740 ;
  assign y5628 = ~n25742 ;
  assign y5629 = n25743 ;
  assign y5630 = ~n25744 ;
  assign y5631 = ~n25745 ;
  assign y5632 = n25749 ;
  assign y5633 = n25753 ;
  assign y5634 = ~n25756 ;
  assign y5635 = n25757 ;
  assign y5636 = n25759 ;
  assign y5637 = ~n25760 ;
  assign y5638 = ~n25762 ;
  assign y5639 = n25764 ;
  assign y5640 = n25766 ;
  assign y5641 = ~n25770 ;
  assign y5642 = ~n25774 ;
  assign y5643 = ~n25775 ;
  assign y5644 = n25776 ;
  assign y5645 = n25779 ;
  assign y5646 = ~n25782 ;
  assign y5647 = n25791 ;
  assign y5648 = n25792 ;
  assign y5649 = ~n25793 ;
  assign y5650 = ~n25796 ;
  assign y5651 = ~n25798 ;
  assign y5652 = ~n25801 ;
  assign y5653 = ~n25802 ;
  assign y5654 = n25806 ;
  assign y5655 = n25808 ;
  assign y5656 = ~n25810 ;
  assign y5657 = ~n25814 ;
  assign y5658 = ~n25816 ;
  assign y5659 = n25818 ;
  assign y5660 = n25822 ;
  assign y5661 = ~n25823 ;
  assign y5662 = ~n25825 ;
  assign y5663 = ~n25828 ;
  assign y5664 = n25831 ;
  assign y5665 = n25832 ;
  assign y5666 = n25833 ;
  assign y5667 = n25835 ;
  assign y5668 = n25841 ;
  assign y5669 = n25844 ;
  assign y5670 = ~n25847 ;
  assign y5671 = ~n25850 ;
  assign y5672 = n25854 ;
  assign y5673 = ~n25859 ;
  assign y5674 = n25861 ;
  assign y5675 = n25863 ;
  assign y5676 = n25868 ;
  assign y5677 = n25869 ;
  assign y5678 = n25872 ;
  assign y5679 = n25873 ;
  assign y5680 = n25874 ;
  assign y5681 = ~n25877 ;
  assign y5682 = n25880 ;
  assign y5683 = ~n25882 ;
  assign y5684 = n25885 ;
  assign y5685 = ~n25887 ;
  assign y5686 = n25890 ;
  assign y5687 = ~n25891 ;
  assign y5688 = ~n25893 ;
  assign y5689 = ~n25899 ;
  assign y5690 = ~n25900 ;
  assign y5691 = ~n25905 ;
  assign y5692 = ~n25908 ;
  assign y5693 = ~n25912 ;
  assign y5694 = n25914 ;
  assign y5695 = ~n25915 ;
  assign y5696 = n25917 ;
  assign y5697 = ~n25918 ;
  assign y5698 = n25922 ;
  assign y5699 = ~n25924 ;
  assign y5700 = n25928 ;
  assign y5701 = ~n25929 ;
  assign y5702 = n25930 ;
  assign y5703 = ~n25931 ;
  assign y5704 = ~n25937 ;
  assign y5705 = n25946 ;
  assign y5706 = ~n25947 ;
  assign y5707 = n25949 ;
  assign y5708 = ~n25951 ;
  assign y5709 = ~n25956 ;
  assign y5710 = n25958 ;
  assign y5711 = n25959 ;
  assign y5712 = ~n25963 ;
  assign y5713 = ~n25965 ;
  assign y5714 = n25966 ;
  assign y5715 = n25967 ;
  assign y5716 = ~n25969 ;
  assign y5717 = n25971 ;
  assign y5718 = n25972 ;
  assign y5719 = ~n25974 ;
  assign y5720 = ~n25975 ;
  assign y5721 = ~n25976 ;
  assign y5722 = n25978 ;
  assign y5723 = ~n25980 ;
  assign y5724 = n25986 ;
  assign y5725 = ~n25988 ;
  assign y5726 = n25991 ;
  assign y5727 = n25992 ;
  assign y5728 = ~n25997 ;
  assign y5729 = ~n26003 ;
  assign y5730 = ~n26004 ;
  assign y5731 = n26008 ;
  assign y5732 = ~n26009 ;
  assign y5733 = ~n26011 ;
  assign y5734 = ~n26016 ;
  assign y5735 = ~n26022 ;
  assign y5736 = n26025 ;
  assign y5737 = ~n26028 ;
  assign y5738 = n26030 ;
  assign y5739 = n26032 ;
  assign y5740 = n26034 ;
  assign y5741 = n26040 ;
  assign y5742 = n26047 ;
  assign y5743 = ~n26051 ;
  assign y5744 = ~n26053 ;
  assign y5745 = ~n26054 ;
  assign y5746 = ~n26055 ;
  assign y5747 = n26058 ;
  assign y5748 = ~n26063 ;
  assign y5749 = ~n26066 ;
  assign y5750 = ~n26071 ;
  assign y5751 = n26072 ;
  assign y5752 = n26078 ;
  assign y5753 = n26079 ;
  assign y5754 = n26080 ;
  assign y5755 = n26082 ;
  assign y5756 = n26085 ;
  assign y5757 = ~n26090 ;
  assign y5758 = ~n26094 ;
  assign y5759 = n26096 ;
  assign y5760 = n26100 ;
  assign y5761 = ~n26101 ;
  assign y5762 = n26109 ;
  assign y5763 = ~n26111 ;
  assign y5764 = ~n26113 ;
  assign y5765 = n26117 ;
  assign y5766 = n26120 ;
  assign y5767 = ~n26121 ;
  assign y5768 = ~n26128 ;
  assign y5769 = ~n26133 ;
  assign y5770 = n26135 ;
  assign y5771 = ~n26137 ;
  assign y5772 = ~n26140 ;
  assign y5773 = ~n26141 ;
  assign y5774 = n26146 ;
  assign y5775 = n26147 ;
  assign y5776 = ~n26148 ;
  assign y5777 = ~n26149 ;
  assign y5778 = n26150 ;
  assign y5779 = ~n26151 ;
  assign y5780 = n26153 ;
  assign y5781 = ~n26154 ;
  assign y5782 = n26155 ;
  assign y5783 = n26157 ;
  assign y5784 = ~n26158 ;
  assign y5785 = ~n26161 ;
  assign y5786 = ~n26163 ;
  assign y5787 = n26165 ;
  assign y5788 = n26169 ;
  assign y5789 = ~n26174 ;
  assign y5790 = ~n26175 ;
  assign y5791 = n26176 ;
  assign y5792 = ~n26181 ;
  assign y5793 = ~n26183 ;
  assign y5794 = ~n26184 ;
  assign y5795 = n26185 ;
  assign y5796 = n26187 ;
  assign y5797 = ~n26188 ;
  assign y5798 = ~n26189 ;
  assign y5799 = ~n26191 ;
  assign y5800 = n26196 ;
  assign y5801 = n26199 ;
  assign y5802 = ~n26201 ;
  assign y5803 = n26202 ;
  assign y5804 = ~n26205 ;
  assign y5805 = ~n26206 ;
  assign y5806 = ~n26208 ;
  assign y5807 = n26210 ;
  assign y5808 = n26211 ;
  assign y5809 = ~n26217 ;
  assign y5810 = n26218 ;
  assign y5811 = n26221 ;
  assign y5812 = ~n26222 ;
  assign y5813 = ~n26226 ;
  assign y5814 = ~n26229 ;
  assign y5815 = n26230 ;
  assign y5816 = n26231 ;
  assign y5817 = n26232 ;
  assign y5818 = ~n26233 ;
  assign y5819 = n26235 ;
  assign y5820 = n26241 ;
  assign y5821 = ~n26244 ;
  assign y5822 = ~n26247 ;
  assign y5823 = n26248 ;
  assign y5824 = ~n26249 ;
  assign y5825 = n26251 ;
  assign y5826 = ~n26252 ;
  assign y5827 = ~n26253 ;
  assign y5828 = ~n26255 ;
  assign y5829 = n26256 ;
  assign y5830 = n26257 ;
  assign y5831 = n26258 ;
  assign y5832 = n26259 ;
  assign y5833 = ~n26263 ;
  assign y5834 = n26266 ;
  assign y5835 = ~n26269 ;
  assign y5836 = ~n26273 ;
  assign y5837 = n26275 ;
  assign y5838 = n26276 ;
  assign y5839 = ~n26277 ;
  assign y5840 = ~n26279 ;
  assign y5841 = n26281 ;
  assign y5842 = ~n26284 ;
  assign y5843 = ~n26285 ;
  assign y5844 = n26287 ;
  assign y5845 = ~n26288 ;
  assign y5846 = n26290 ;
  assign y5847 = n26293 ;
  assign y5848 = n26294 ;
  assign y5849 = n26298 ;
  assign y5850 = ~n26299 ;
  assign y5851 = n26300 ;
  assign y5852 = n26302 ;
  assign y5853 = ~n26304 ;
  assign y5854 = ~n26305 ;
  assign y5855 = ~n26306 ;
  assign y5856 = n26309 ;
  assign y5857 = n26313 ;
  assign y5858 = ~n26314 ;
  assign y5859 = n26315 ;
  assign y5860 = n26316 ;
  assign y5861 = ~n26324 ;
  assign y5862 = n26326 ;
  assign y5863 = n26327 ;
  assign y5864 = n26329 ;
  assign y5865 = n26332 ;
  assign y5866 = ~n26333 ;
  assign y5867 = n26335 ;
  assign y5868 = n26336 ;
  assign y5869 = ~n26337 ;
  assign y5870 = ~n26340 ;
  assign y5871 = n26346 ;
  assign y5872 = ~n26347 ;
  assign y5873 = ~n26350 ;
  assign y5874 = ~n26353 ;
  assign y5875 = ~n26355 ;
  assign y5876 = n26358 ;
  assign y5877 = n26361 ;
  assign y5878 = ~n26362 ;
  assign y5879 = ~n26366 ;
  assign y5880 = ~n26367 ;
  assign y5881 = ~n26369 ;
  assign y5882 = n26371 ;
  assign y5883 = n26374 ;
  assign y5884 = ~n26376 ;
  assign y5885 = n26378 ;
  assign y5886 = ~n26382 ;
  assign y5887 = n26388 ;
  assign y5888 = n26390 ;
  assign y5889 = n26392 ;
  assign y5890 = ~n26396 ;
  assign y5891 = ~n26400 ;
  assign y5892 = n26405 ;
  assign y5893 = ~n26408 ;
  assign y5894 = n26410 ;
  assign y5895 = n26411 ;
  assign y5896 = n26413 ;
  assign y5897 = n26414 ;
  assign y5898 = ~n26417 ;
  assign y5899 = ~n26418 ;
  assign y5900 = ~n26420 ;
  assign y5901 = n26424 ;
  assign y5902 = ~n26425 ;
  assign y5903 = ~n26428 ;
  assign y5904 = ~n26430 ;
  assign y5905 = ~n26434 ;
  assign y5906 = n26435 ;
  assign y5907 = n26437 ;
  assign y5908 = ~n26440 ;
  assign y5909 = ~n26441 ;
  assign y5910 = n26445 ;
  assign y5911 = ~n26447 ;
  assign y5912 = ~n26449 ;
  assign y5913 = n26456 ;
  assign y5914 = ~n26457 ;
  assign y5915 = n26458 ;
  assign y5916 = n26462 ;
  assign y5917 = ~n26463 ;
  assign y5918 = n26465 ;
  assign y5919 = ~n26469 ;
  assign y5920 = n26472 ;
  assign y5921 = ~n26475 ;
  assign y5922 = n26478 ;
  assign y5923 = ~n26481 ;
  assign y5924 = ~n26482 ;
  assign y5925 = ~n26485 ;
  assign y5926 = ~n26486 ;
  assign y5927 = ~n26487 ;
  assign y5928 = ~n26490 ;
  assign y5929 = n26496 ;
  assign y5930 = n26498 ;
  assign y5931 = ~n26500 ;
  assign y5932 = n26501 ;
  assign y5933 = n26502 ;
  assign y5934 = ~n26504 ;
  assign y5935 = ~n26507 ;
  assign y5936 = n26508 ;
  assign y5937 = ~n26510 ;
  assign y5938 = ~n26515 ;
  assign y5939 = ~n26519 ;
  assign y5940 = n26521 ;
  assign y5941 = n26522 ;
  assign y5942 = ~n26524 ;
  assign y5943 = ~n26525 ;
  assign y5944 = ~n26526 ;
  assign y5945 = n26527 ;
  assign y5946 = ~n26530 ;
  assign y5947 = ~n26532 ;
  assign y5948 = n26534 ;
  assign y5949 = ~n26536 ;
  assign y5950 = ~n26545 ;
  assign y5951 = n26549 ;
  assign y5952 = ~n26550 ;
  assign y5953 = n26551 ;
  assign y5954 = n26552 ;
  assign y5955 = n26554 ;
  assign y5956 = n26556 ;
  assign y5957 = n26558 ;
  assign y5958 = ~n26559 ;
  assign y5959 = n26561 ;
  assign y5960 = ~n26562 ;
  assign y5961 = n26563 ;
  assign y5962 = ~n26564 ;
  assign y5963 = n26566 ;
  assign y5964 = n26570 ;
  assign y5965 = n26574 ;
  assign y5966 = ~n26579 ;
  assign y5967 = ~n26581 ;
  assign y5968 = ~n26582 ;
  assign y5969 = ~n26588 ;
  assign y5970 = n26589 ;
  assign y5971 = ~n26590 ;
  assign y5972 = n26593 ;
  assign y5973 = n26594 ;
  assign y5974 = n26595 ;
  assign y5975 = n26597 ;
  assign y5976 = ~n26598 ;
  assign y5977 = n26602 ;
  assign y5978 = n26605 ;
  assign y5979 = ~n26607 ;
  assign y5980 = n26608 ;
  assign y5981 = ~n26613 ;
  assign y5982 = ~n26615 ;
  assign y5983 = ~n26616 ;
  assign y5984 = n26618 ;
  assign y5985 = n26620 ;
  assign y5986 = n26622 ;
  assign y5987 = ~n26624 ;
  assign y5988 = n26625 ;
  assign y5989 = ~n26626 ;
  assign y5990 = ~n26628 ;
  assign y5991 = ~n26630 ;
  assign y5992 = n26635 ;
  assign y5993 = n26636 ;
  assign y5994 = ~n26648 ;
  assign y5995 = n26649 ;
  assign y5996 = ~n26652 ;
  assign y5997 = n26654 ;
  assign y5998 = n26656 ;
  assign y5999 = ~n26659 ;
  assign y6000 = ~n26661 ;
  assign y6001 = ~n26662 ;
  assign y6002 = n26663 ;
  assign y6003 = ~n26664 ;
  assign y6004 = n26669 ;
  assign y6005 = ~n26671 ;
  assign y6006 = n26675 ;
  assign y6007 = ~n26677 ;
  assign y6008 = n26678 ;
  assign y6009 = n26680 ;
  assign y6010 = n26681 ;
  assign y6011 = n26683 ;
  assign y6012 = n26686 ;
  assign y6013 = n26687 ;
  assign y6014 = n26688 ;
  assign y6015 = n26689 ;
  assign y6016 = ~n26691 ;
  assign y6017 = ~n26692 ;
  assign y6018 = n26695 ;
  assign y6019 = ~n26696 ;
  assign y6020 = ~n26701 ;
  assign y6021 = n26703 ;
  assign y6022 = n26705 ;
  assign y6023 = ~n26709 ;
  assign y6024 = n26715 ;
  assign y6025 = ~n26717 ;
  assign y6026 = ~n26720 ;
  assign y6027 = n26722 ;
  assign y6028 = n26723 ;
  assign y6029 = n26726 ;
  assign y6030 = n26727 ;
  assign y6031 = n26730 ;
  assign y6032 = n26731 ;
  assign y6033 = ~n26732 ;
  assign y6034 = n26733 ;
  assign y6035 = ~n26736 ;
  assign y6036 = ~n26737 ;
  assign y6037 = n26738 ;
  assign y6038 = ~n26739 ;
  assign y6039 = ~n26740 ;
  assign y6040 = ~n26743 ;
  assign y6041 = ~n26745 ;
  assign y6042 = n26746 ;
  assign y6043 = n26749 ;
  assign y6044 = n26752 ;
  assign y6045 = ~n26753 ;
  assign y6046 = n26754 ;
  assign y6047 = ~n26755 ;
  assign y6048 = ~n26757 ;
  assign y6049 = n26758 ;
  assign y6050 = ~n26760 ;
  assign y6051 = ~n26764 ;
  assign y6052 = ~n26765 ;
  assign y6053 = n26767 ;
  assign y6054 = n26768 ;
  assign y6055 = ~n26769 ;
  assign y6056 = n26774 ;
  assign y6057 = n26776 ;
  assign y6058 = ~n26780 ;
  assign y6059 = n26782 ;
  assign y6060 = ~n26785 ;
  assign y6061 = n26791 ;
  assign y6062 = n26792 ;
  assign y6063 = n26793 ;
  assign y6064 = n26795 ;
  assign y6065 = n26796 ;
  assign y6066 = n26800 ;
  assign y6067 = ~n26801 ;
  assign y6068 = n26803 ;
  assign y6069 = n26810 ;
  assign y6070 = ~n26813 ;
  assign y6071 = n26815 ;
  assign y6072 = n26817 ;
  assign y6073 = ~n26819 ;
  assign y6074 = n26823 ;
  assign y6075 = n26826 ;
  assign y6076 = ~n26828 ;
  assign y6077 = ~n26830 ;
  assign y6078 = n26833 ;
  assign y6079 = ~n26835 ;
  assign y6080 = ~n26837 ;
  assign y6081 = n26842 ;
  assign y6082 = ~n26843 ;
  assign y6083 = ~n26844 ;
  assign y6084 = ~n26848 ;
  assign y6085 = ~n26851 ;
  assign y6086 = n26853 ;
  assign y6087 = n26855 ;
  assign y6088 = ~n26857 ;
  assign y6089 = n26861 ;
  assign y6090 = ~n26863 ;
  assign y6091 = n26865 ;
  assign y6092 = n26868 ;
  assign y6093 = n26873 ;
  assign y6094 = n26877 ;
  assign y6095 = ~n26878 ;
  assign y6096 = ~n26880 ;
  assign y6097 = n26882 ;
  assign y6098 = ~n26885 ;
  assign y6099 = n26886 ;
  assign y6100 = n26891 ;
  assign y6101 = n26892 ;
  assign y6102 = ~n26894 ;
  assign y6103 = n26895 ;
  assign y6104 = ~n26896 ;
  assign y6105 = ~n26897 ;
  assign y6106 = n26900 ;
  assign y6107 = ~n26906 ;
  assign y6108 = ~n26911 ;
  assign y6109 = n26912 ;
  assign y6110 = n26914 ;
  assign y6111 = ~n26915 ;
  assign y6112 = ~n26916 ;
  assign y6113 = n26917 ;
  assign y6114 = ~n26918 ;
  assign y6115 = n26921 ;
  assign y6116 = ~n26922 ;
  assign y6117 = ~n26926 ;
  assign y6118 = n26927 ;
  assign y6119 = n26930 ;
  assign y6120 = n26933 ;
  assign y6121 = ~n26935 ;
  assign y6122 = n26938 ;
  assign y6123 = ~n26942 ;
  assign y6124 = ~n26943 ;
  assign y6125 = ~n26944 ;
  assign y6126 = ~n26946 ;
  assign y6127 = n26949 ;
  assign y6128 = n26951 ;
  assign y6129 = ~n26953 ;
  assign y6130 = n26954 ;
  assign y6131 = n26958 ;
  assign y6132 = n26963 ;
  assign y6133 = ~n26965 ;
  assign y6134 = ~n26967 ;
  assign y6135 = n26968 ;
  assign y6136 = ~n26971 ;
  assign y6137 = ~n26972 ;
  assign y6138 = ~n26973 ;
  assign y6139 = n26975 ;
  assign y6140 = ~n26976 ;
  assign y6141 = ~n26978 ;
  assign y6142 = ~n26979 ;
  assign y6143 = n26981 ;
  assign y6144 = ~n26983 ;
  assign y6145 = n26986 ;
  assign y6146 = n26989 ;
  assign y6147 = ~n26990 ;
  assign y6148 = ~n26993 ;
  assign y6149 = n26994 ;
  assign y6150 = ~n26997 ;
  assign y6151 = ~n26999 ;
  assign y6152 = ~n27002 ;
  assign y6153 = n27007 ;
  assign y6154 = n27008 ;
  assign y6155 = n27011 ;
  assign y6156 = n27014 ;
  assign y6157 = ~n27015 ;
  assign y6158 = n27016 ;
  assign y6159 = ~n27017 ;
  assign y6160 = ~n27018 ;
  assign y6161 = ~n27022 ;
  assign y6162 = ~n27023 ;
  assign y6163 = n27026 ;
  assign y6164 = ~n27027 ;
  assign y6165 = n27029 ;
  assign y6166 = n27033 ;
  assign y6167 = ~n27035 ;
  assign y6168 = n27040 ;
  assign y6169 = ~n27044 ;
  assign y6170 = ~n27045 ;
  assign y6171 = n27048 ;
  assign y6172 = n27050 ;
  assign y6173 = n27054 ;
  assign y6174 = ~n27055 ;
  assign y6175 = n27060 ;
  assign y6176 = ~n27064 ;
  assign y6177 = n27066 ;
  assign y6178 = n27068 ;
  assign y6179 = ~n27072 ;
  assign y6180 = n27074 ;
  assign y6181 = ~n27075 ;
  assign y6182 = n27078 ;
  assign y6183 = ~n27080 ;
  assign y6184 = n27082 ;
  assign y6185 = ~n27083 ;
  assign y6186 = n27084 ;
  assign y6187 = ~n27086 ;
  assign y6188 = n27091 ;
  assign y6189 = ~n27092 ;
  assign y6190 = ~n27093 ;
  assign y6191 = n27095 ;
  assign y6192 = n27099 ;
  assign y6193 = n27102 ;
  assign y6194 = n27103 ;
  assign y6195 = ~n27104 ;
  assign y6196 = ~n27106 ;
  assign y6197 = n27107 ;
  assign y6198 = n27109 ;
  assign y6199 = n27111 ;
  assign y6200 = ~n27112 ;
  assign y6201 = n27116 ;
  assign y6202 = n27117 ;
  assign y6203 = n27118 ;
  assign y6204 = ~n27119 ;
  assign y6205 = n27122 ;
  assign y6206 = ~n27124 ;
  assign y6207 = ~n27127 ;
  assign y6208 = n27131 ;
  assign y6209 = ~n27132 ;
  assign y6210 = ~n27134 ;
  assign y6211 = n27137 ;
  assign y6212 = n27139 ;
  assign y6213 = n27140 ;
  assign y6214 = n27141 ;
  assign y6215 = n27142 ;
  assign y6216 = n27143 ;
  assign y6217 = ~n27144 ;
  assign y6218 = ~n27147 ;
  assign y6219 = ~n27148 ;
  assign y6220 = ~n27149 ;
  assign y6221 = n27150 ;
  assign y6222 = n27154 ;
  assign y6223 = n27160 ;
  assign y6224 = n27161 ;
  assign y6225 = n27163 ;
  assign y6226 = ~n27166 ;
  assign y6227 = n27169 ;
  assign y6228 = ~n27171 ;
  assign y6229 = ~n27172 ;
  assign y6230 = ~n27173 ;
  assign y6231 = ~n27176 ;
  assign y6232 = ~n27178 ;
  assign y6233 = ~n27179 ;
  assign y6234 = ~n27180 ;
  assign y6235 = ~n27184 ;
  assign y6236 = n27186 ;
  assign y6237 = n27187 ;
  assign y6238 = ~n27188 ;
  assign y6239 = n27190 ;
  assign y6240 = n27194 ;
  assign y6241 = n27195 ;
  assign y6242 = ~n27197 ;
  assign y6243 = ~n27201 ;
  assign y6244 = n27208 ;
  assign y6245 = ~n27213 ;
  assign y6246 = n27218 ;
  assign y6247 = n27219 ;
  assign y6248 = n27220 ;
  assign y6249 = n27222 ;
  assign y6250 = n27223 ;
  assign y6251 = ~n27225 ;
  assign y6252 = n27226 ;
  assign y6253 = n27229 ;
  assign y6254 = ~n27230 ;
  assign y6255 = ~n27232 ;
  assign y6256 = n27233 ;
  assign y6257 = n27237 ;
  assign y6258 = ~n27241 ;
  assign y6259 = ~n27242 ;
  assign y6260 = n27248 ;
  assign y6261 = ~n27253 ;
  assign y6262 = ~n27257 ;
  assign y6263 = n27259 ;
  assign y6264 = n27260 ;
  assign y6265 = n27261 ;
  assign y6266 = n27263 ;
  assign y6267 = ~n27266 ;
  assign y6268 = n27270 ;
  assign y6269 = ~n27272 ;
  assign y6270 = n27275 ;
  assign y6271 = ~n27278 ;
  assign y6272 = n27281 ;
  assign y6273 = n27282 ;
  assign y6274 = n27283 ;
  assign y6275 = n27285 ;
  assign y6276 = n27286 ;
  assign y6277 = n27287 ;
  assign y6278 = n27288 ;
  assign y6279 = n27289 ;
  assign y6280 = ~n27291 ;
  assign y6281 = n27293 ;
  assign y6282 = ~n27298 ;
  assign y6283 = ~n27300 ;
  assign y6284 = ~n27301 ;
  assign y6285 = n27303 ;
  assign y6286 = ~n27306 ;
  assign y6287 = n27307 ;
  assign y6288 = ~n27312 ;
  assign y6289 = ~n27313 ;
  assign y6290 = n27315 ;
  assign y6291 = n27318 ;
  assign y6292 = n27319 ;
  assign y6293 = n27320 ;
  assign y6294 = ~n27322 ;
  assign y6295 = ~n27323 ;
  assign y6296 = ~n27326 ;
  assign y6297 = ~n27328 ;
  assign y6298 = n27329 ;
  assign y6299 = n27332 ;
  assign y6300 = ~n27333 ;
  assign y6301 = n27334 ;
  assign y6302 = n27337 ;
  assign y6303 = n27339 ;
  assign y6304 = ~n27340 ;
  assign y6305 = ~n27341 ;
  assign y6306 = ~n27342 ;
  assign y6307 = ~n27344 ;
  assign y6308 = ~n27346 ;
  assign y6309 = n27348 ;
  assign y6310 = n27349 ;
  assign y6311 = ~n27350 ;
  assign y6312 = ~n27352 ;
  assign y6313 = n27353 ;
  assign y6314 = ~n27354 ;
  assign y6315 = ~n27356 ;
  assign y6316 = n27357 ;
  assign y6317 = n27363 ;
  assign y6318 = ~n27366 ;
  assign y6319 = n27368 ;
  assign y6320 = n27369 ;
  assign y6321 = n27373 ;
  assign y6322 = ~n27374 ;
  assign y6323 = ~n27375 ;
  assign y6324 = n27376 ;
  assign y6325 = ~n27377 ;
  assign y6326 = n27379 ;
  assign y6327 = n27380 ;
  assign y6328 = ~n27382 ;
  assign y6329 = n27385 ;
  assign y6330 = n27388 ;
  assign y6331 = ~n27390 ;
  assign y6332 = n27394 ;
  assign y6333 = ~n27395 ;
  assign y6334 = ~n27396 ;
  assign y6335 = ~n27397 ;
  assign y6336 = n27400 ;
  assign y6337 = n27403 ;
  assign y6338 = ~n27404 ;
  assign y6339 = n27405 ;
  assign y6340 = ~n27406 ;
  assign y6341 = n27410 ;
  assign y6342 = ~n27412 ;
  assign y6343 = ~n27416 ;
  assign y6344 = ~n27419 ;
  assign y6345 = n27420 ;
  assign y6346 = n27423 ;
  assign y6347 = ~n27426 ;
  assign y6348 = ~n27428 ;
  assign y6349 = n27431 ;
  assign y6350 = n27434 ;
  assign y6351 = n27437 ;
  assign y6352 = n27440 ;
  assign y6353 = ~n27445 ;
  assign y6354 = ~n27446 ;
  assign y6355 = n27447 ;
  assign y6356 = ~n27448 ;
  assign y6357 = n27449 ;
  assign y6358 = ~n27453 ;
  assign y6359 = ~n27454 ;
  assign y6360 = ~n27457 ;
  assign y6361 = ~n27458 ;
  assign y6362 = ~n27459 ;
  assign y6363 = n27460 ;
  assign y6364 = n27462 ;
  assign y6365 = ~n27463 ;
  assign y6366 = n27465 ;
  assign y6367 = n27466 ;
  assign y6368 = ~n27467 ;
  assign y6369 = ~n27469 ;
  assign y6370 = n27470 ;
  assign y6371 = ~n27472 ;
  assign y6372 = n27474 ;
  assign y6373 = ~n27476 ;
  assign y6374 = ~n27477 ;
  assign y6375 = ~n27478 ;
  assign y6376 = ~n27480 ;
  assign y6377 = ~n27481 ;
  assign y6378 = n27483 ;
  assign y6379 = n27487 ;
  assign y6380 = ~n27488 ;
  assign y6381 = n27490 ;
  assign y6382 = ~n27492 ;
  assign y6383 = ~n27493 ;
  assign y6384 = ~n27497 ;
  assign y6385 = ~n27499 ;
  assign y6386 = n27500 ;
  assign y6387 = ~n27501 ;
  assign y6388 = ~n27503 ;
  assign y6389 = ~n27506 ;
  assign y6390 = n27508 ;
  assign y6391 = n27509 ;
  assign y6392 = ~n27510 ;
  assign y6393 = ~n27512 ;
  assign y6394 = n27514 ;
  assign y6395 = n27518 ;
  assign y6396 = ~n27519 ;
  assign y6397 = n27522 ;
  assign y6398 = ~n27528 ;
  assign y6399 = ~n27532 ;
  assign y6400 = ~n27535 ;
  assign y6401 = n27536 ;
  assign y6402 = ~n27539 ;
  assign y6403 = n27543 ;
  assign y6404 = n27544 ;
  assign y6405 = ~n27545 ;
  assign y6406 = n27546 ;
  assign y6407 = n27547 ;
  assign y6408 = ~n27551 ;
  assign y6409 = ~n27552 ;
  assign y6410 = ~n27554 ;
  assign y6411 = ~n27556 ;
  assign y6412 = ~n27557 ;
  assign y6413 = ~n27563 ;
  assign y6414 = n27564 ;
  assign y6415 = n27565 ;
  assign y6416 = ~n27569 ;
  assign y6417 = ~n27570 ;
  assign y6418 = ~n27571 ;
  assign y6419 = ~n27573 ;
  assign y6420 = n27574 ;
  assign y6421 = ~n27576 ;
  assign y6422 = ~n27580 ;
  assign y6423 = n27581 ;
  assign y6424 = ~n27584 ;
  assign y6425 = ~n27585 ;
  assign y6426 = n27587 ;
  assign y6427 = ~n27589 ;
  assign y6428 = ~n27591 ;
  assign y6429 = ~n27592 ;
  assign y6430 = n27594 ;
  assign y6431 = n27599 ;
  assign y6432 = ~n27602 ;
  assign y6433 = ~n27609 ;
  assign y6434 = ~n27612 ;
  assign y6435 = n27615 ;
  assign y6436 = n27616 ;
  assign y6437 = ~n27620 ;
  assign y6438 = ~n27622 ;
  assign y6439 = n27623 ;
  assign y6440 = ~n27624 ;
  assign y6441 = ~n27625 ;
  assign y6442 = n27627 ;
  assign y6443 = ~n27631 ;
  assign y6444 = n27634 ;
  assign y6445 = ~n27636 ;
  assign y6446 = n27637 ;
  assign y6447 = n27638 ;
  assign y6448 = n27641 ;
  assign y6449 = n27645 ;
  assign y6450 = ~n27646 ;
  assign y6451 = ~n27647 ;
  assign y6452 = ~n27649 ;
  assign y6453 = ~n27650 ;
  assign y6454 = n27651 ;
  assign y6455 = n27653 ;
  assign y6456 = ~n27654 ;
  assign y6457 = n27655 ;
  assign y6458 = ~n27659 ;
  assign y6459 = ~n27664 ;
  assign y6460 = n27666 ;
  assign y6461 = n27670 ;
  assign y6462 = ~n27673 ;
  assign y6463 = n27675 ;
  assign y6464 = n27682 ;
  assign y6465 = n27683 ;
  assign y6466 = n27684 ;
  assign y6467 = n27687 ;
  assign y6468 = ~n27688 ;
  assign y6469 = n27690 ;
  assign y6470 = ~n27692 ;
  assign y6471 = ~n27694 ;
  assign y6472 = ~n27698 ;
  assign y6473 = n27699 ;
  assign y6474 = ~n27701 ;
  assign y6475 = ~n27702 ;
  assign y6476 = ~n27704 ;
  assign y6477 = ~n27710 ;
  assign y6478 = ~n27712 ;
  assign y6479 = ~n27714 ;
  assign y6480 = n27717 ;
  assign y6481 = n27718 ;
  assign y6482 = n27719 ;
  assign y6483 = ~n27720 ;
  assign y6484 = ~n27722 ;
  assign y6485 = n27727 ;
  assign y6486 = ~n27730 ;
  assign y6487 = n27736 ;
  assign y6488 = ~n27737 ;
  assign y6489 = ~n27738 ;
  assign y6490 = n27739 ;
  assign y6491 = n27741 ;
  assign y6492 = n27743 ;
  assign y6493 = n27745 ;
  assign y6494 = ~n27746 ;
  assign y6495 = ~n27747 ;
  assign y6496 = n27748 ;
  assign y6497 = n27750 ;
  assign y6498 = ~n27751 ;
  assign y6499 = ~n27752 ;
  assign y6500 = n27757 ;
  assign y6501 = n27761 ;
  assign y6502 = n27763 ;
  assign y6503 = n27767 ;
  assign y6504 = n27768 ;
  assign y6505 = n27769 ;
  assign y6506 = n27772 ;
  assign y6507 = ~n27774 ;
  assign y6508 = n27775 ;
  assign y6509 = ~n27784 ;
  assign y6510 = n27785 ;
  assign y6511 = n27789 ;
  assign y6512 = n27790 ;
  assign y6513 = ~n27791 ;
  assign y6514 = n27792 ;
  assign y6515 = n27795 ;
  assign y6516 = ~n27802 ;
  assign y6517 = ~n27804 ;
  assign y6518 = ~n27805 ;
  assign y6519 = ~n27806 ;
  assign y6520 = n27808 ;
  assign y6521 = ~n27809 ;
  assign y6522 = n27810 ;
  assign y6523 = n27814 ;
  assign y6524 = ~n27816 ;
  assign y6525 = n27819 ;
  assign y6526 = n27821 ;
  assign y6527 = ~n27822 ;
  assign y6528 = n27826 ;
  assign y6529 = n27829 ;
  assign y6530 = ~n27830 ;
  assign y6531 = ~n27832 ;
  assign y6532 = n27834 ;
  assign y6533 = n27836 ;
  assign y6534 = ~n27837 ;
  assign y6535 = ~n27838 ;
  assign y6536 = n27839 ;
  assign y6537 = ~n27840 ;
  assign y6538 = ~n27844 ;
  assign y6539 = n27846 ;
  assign y6540 = ~n27848 ;
  assign y6541 = ~n27858 ;
  assign y6542 = n27859 ;
  assign y6543 = n27861 ;
  assign y6544 = n27863 ;
  assign y6545 = n27864 ;
  assign y6546 = ~n27866 ;
  assign y6547 = ~n27867 ;
  assign y6548 = ~n27873 ;
  assign y6549 = ~n27875 ;
  assign y6550 = ~n27879 ;
  assign y6551 = ~n27880 ;
  assign y6552 = n27885 ;
  assign y6553 = ~n27889 ;
  assign y6554 = ~n27890 ;
  assign y6555 = ~n27894 ;
  assign y6556 = n27895 ;
  assign y6557 = n27900 ;
  assign y6558 = n27901 ;
  assign y6559 = n27903 ;
  assign y6560 = n27905 ;
  assign y6561 = ~n27911 ;
  assign y6562 = n27912 ;
  assign y6563 = ~n27914 ;
  assign y6564 = ~n27915 ;
  assign y6565 = ~n27922 ;
  assign y6566 = n27925 ;
  assign y6567 = ~n27930 ;
  assign y6568 = ~n27931 ;
  assign y6569 = ~n27932 ;
  assign y6570 = n27934 ;
  assign y6571 = n27936 ;
  assign y6572 = ~n27937 ;
  assign y6573 = n27939 ;
  assign y6574 = ~n27941 ;
  assign y6575 = n27944 ;
  assign y6576 = n27945 ;
  assign y6577 = n27947 ;
  assign y6578 = ~n27950 ;
  assign y6579 = ~n27951 ;
  assign y6580 = n27952 ;
  assign y6581 = n27955 ;
  assign y6582 = ~n27956 ;
  assign y6583 = ~n27958 ;
  assign y6584 = n27959 ;
  assign y6585 = ~n27960 ;
  assign y6586 = ~n27962 ;
  assign y6587 = ~n27966 ;
  assign y6588 = ~n27967 ;
  assign y6589 = n27969 ;
  assign y6590 = ~n27970 ;
  assign y6591 = n27972 ;
  assign y6592 = ~n27976 ;
  assign y6593 = n27979 ;
  assign y6594 = n27981 ;
  assign y6595 = ~n27982 ;
  assign y6596 = ~n27987 ;
  assign y6597 = ~n27988 ;
  assign y6598 = ~n27992 ;
  assign y6599 = n27993 ;
  assign y6600 = ~n27995 ;
  assign y6601 = n28000 ;
  assign y6602 = ~n28001 ;
  assign y6603 = n28004 ;
  assign y6604 = n28008 ;
  assign y6605 = ~n28010 ;
  assign y6606 = n28015 ;
  assign y6607 = n28016 ;
  assign y6608 = n28017 ;
  assign y6609 = n28021 ;
  assign y6610 = ~n28022 ;
  assign y6611 = n28024 ;
  assign y6612 = ~n28026 ;
  assign y6613 = ~n28031 ;
  assign y6614 = n28033 ;
  assign y6615 = n28034 ;
  assign y6616 = n28040 ;
  assign y6617 = n28042 ;
  assign y6618 = n28043 ;
  assign y6619 = n28047 ;
  assign y6620 = n28051 ;
  assign y6621 = n28054 ;
  assign y6622 = ~n28055 ;
  assign y6623 = ~n28056 ;
  assign y6624 = n28060 ;
  assign y6625 = n28067 ;
  assign y6626 = ~n28070 ;
  assign y6627 = n28071 ;
  assign y6628 = n28072 ;
  assign y6629 = n28073 ;
  assign y6630 = ~n28074 ;
  assign y6631 = ~n28076 ;
  assign y6632 = n28079 ;
  assign y6633 = ~n28080 ;
  assign y6634 = n28082 ;
  assign y6635 = ~n28084 ;
  assign y6636 = ~n28087 ;
  assign y6637 = n28091 ;
  assign y6638 = ~n28093 ;
  assign y6639 = ~n28094 ;
  assign y6640 = n28095 ;
  assign y6641 = n28096 ;
  assign y6642 = n28098 ;
  assign y6643 = ~n28099 ;
  assign y6644 = ~n28100 ;
  assign y6645 = n28101 ;
  assign y6646 = ~n28102 ;
  assign y6647 = n28103 ;
  assign y6648 = n28107 ;
  assign y6649 = n28108 ;
  assign y6650 = ~n28115 ;
  assign y6651 = n28116 ;
  assign y6652 = n28118 ;
  assign y6653 = ~n28119 ;
  assign y6654 = ~n28122 ;
  assign y6655 = ~n28124 ;
  assign y6656 = ~n28128 ;
  assign y6657 = ~n28130 ;
  assign y6658 = ~n28132 ;
  assign y6659 = n28135 ;
  assign y6660 = ~n28140 ;
  assign y6661 = ~n28143 ;
  assign y6662 = n28147 ;
  assign y6663 = n28149 ;
  assign y6664 = n28156 ;
  assign y6665 = ~n28157 ;
  assign y6666 = ~n28163 ;
  assign y6667 = ~n28166 ;
  assign y6668 = ~n28168 ;
  assign y6669 = ~n28170 ;
  assign y6670 = ~n28171 ;
  assign y6671 = n28175 ;
  assign y6672 = n28178 ;
  assign y6673 = n28179 ;
  assign y6674 = n28181 ;
  assign y6675 = n28183 ;
  assign y6676 = ~n28184 ;
  assign y6677 = n28185 ;
  assign y6678 = n28186 ;
  assign y6679 = n28187 ;
  assign y6680 = n28189 ;
  assign y6681 = n28191 ;
  assign y6682 = n28194 ;
  assign y6683 = ~n28196 ;
  assign y6684 = ~n28201 ;
  assign y6685 = n28202 ;
  assign y6686 = ~n28204 ;
  assign y6687 = n28205 ;
  assign y6688 = n28207 ;
  assign y6689 = ~n28209 ;
  assign y6690 = n28210 ;
  assign y6691 = n28211 ;
  assign y6692 = ~n28212 ;
  assign y6693 = n28213 ;
  assign y6694 = ~n28214 ;
  assign y6695 = n28215 ;
  assign y6696 = ~n28217 ;
  assign y6697 = n28218 ;
  assign y6698 = ~n28220 ;
  assign y6699 = n28223 ;
  assign y6700 = ~n28226 ;
  assign y6701 = ~n28227 ;
  assign y6702 = n28231 ;
  assign y6703 = ~n28236 ;
  assign y6704 = ~n28240 ;
  assign y6705 = ~n28244 ;
  assign y6706 = ~n28245 ;
  assign y6707 = n28247 ;
  assign y6708 = n28249 ;
  assign y6709 = ~n28250 ;
  assign y6710 = n28252 ;
  assign y6711 = n28254 ;
  assign y6712 = n28257 ;
  assign y6713 = ~n28260 ;
  assign y6714 = ~n28263 ;
  assign y6715 = n28267 ;
  assign y6716 = n28269 ;
  assign y6717 = ~n28273 ;
  assign y6718 = ~n28277 ;
  assign y6719 = n28278 ;
  assign y6720 = n28279 ;
  assign y6721 = n28280 ;
  assign y6722 = n28284 ;
  assign y6723 = ~n28285 ;
  assign y6724 = n28286 ;
  assign y6725 = n28290 ;
  assign y6726 = n28291 ;
  assign y6727 = n28293 ;
  assign y6728 = n28296 ;
  assign y6729 = ~n28297 ;
  assign y6730 = n28298 ;
  assign y6731 = n28299 ;
  assign y6732 = ~n28300 ;
  assign y6733 = n28301 ;
  assign y6734 = ~n28305 ;
  assign y6735 = ~n28309 ;
  assign y6736 = n28311 ;
  assign y6737 = ~n28312 ;
  assign y6738 = n28315 ;
  assign y6739 = ~n28317 ;
  assign y6740 = ~n28320 ;
  assign y6741 = ~n28324 ;
  assign y6742 = n28325 ;
  assign y6743 = ~n28327 ;
  assign y6744 = ~n28329 ;
  assign y6745 = ~n28330 ;
  assign y6746 = ~n28331 ;
  assign y6747 = ~n28333 ;
  assign y6748 = ~n28335 ;
  assign y6749 = ~n28337 ;
  assign y6750 = ~n28338 ;
  assign y6751 = n28339 ;
  assign y6752 = n28340 ;
  assign y6753 = n28341 ;
  assign y6754 = n28342 ;
  assign y6755 = n28343 ;
  assign y6756 = n28345 ;
  assign y6757 = n28348 ;
  assign y6758 = n28349 ;
  assign y6759 = ~n28352 ;
  assign y6760 = n28353 ;
  assign y6761 = n28355 ;
  assign y6762 = n28357 ;
  assign y6763 = n28359 ;
  assign y6764 = ~n28361 ;
  assign y6765 = n28362 ;
  assign y6766 = n28364 ;
  assign y6767 = ~n28367 ;
  assign y6768 = n28371 ;
  assign y6769 = n28373 ;
  assign y6770 = n28375 ;
  assign y6771 = n28376 ;
  assign y6772 = ~n28377 ;
  assign y6773 = ~n28381 ;
  assign y6774 = n28382 ;
  assign y6775 = ~n28384 ;
  assign y6776 = ~n28388 ;
  assign y6777 = ~n28389 ;
  assign y6778 = n28392 ;
  assign y6779 = ~n28394 ;
  assign y6780 = n28395 ;
  assign y6781 = ~n28396 ;
  assign y6782 = ~n28398 ;
  assign y6783 = n28399 ;
  assign y6784 = n28400 ;
  assign y6785 = ~n28403 ;
  assign y6786 = ~n28404 ;
  assign y6787 = ~n28407 ;
  assign y6788 = n28409 ;
  assign y6789 = ~n28413 ;
  assign y6790 = n28416 ;
  assign y6791 = n28420 ;
  assign y6792 = ~n28422 ;
  assign y6793 = ~n28427 ;
  assign y6794 = n28428 ;
  assign y6795 = ~n28430 ;
  assign y6796 = n28432 ;
  assign y6797 = n28436 ;
  assign y6798 = n28441 ;
  assign y6799 = ~n28443 ;
  assign y6800 = n28445 ;
  assign y6801 = ~n28447 ;
  assign y6802 = ~n28452 ;
  assign y6803 = n28455 ;
  assign y6804 = n28457 ;
  assign y6805 = n28458 ;
  assign y6806 = ~n28459 ;
  assign y6807 = ~n28461 ;
  assign y6808 = ~n28462 ;
  assign y6809 = n28463 ;
  assign y6810 = n28465 ;
  assign y6811 = n28466 ;
  assign y6812 = n28471 ;
  assign y6813 = n28473 ;
  assign y6814 = n28474 ;
  assign y6815 = ~n28476 ;
  assign y6816 = ~n28477 ;
  assign y6817 = ~n28480 ;
  assign y6818 = n28485 ;
  assign y6819 = n28486 ;
  assign y6820 = ~n28491 ;
  assign y6821 = n28495 ;
  assign y6822 = ~n28500 ;
  assign y6823 = ~n28502 ;
  assign y6824 = ~n28503 ;
  assign y6825 = ~n28507 ;
  assign y6826 = ~n28511 ;
  assign y6827 = ~n28514 ;
  assign y6828 = ~n28519 ;
  assign y6829 = n28521 ;
  assign y6830 = ~n28527 ;
  assign y6831 = n28528 ;
  assign y6832 = n28529 ;
  assign y6833 = n28531 ;
  assign y6834 = n28534 ;
  assign y6835 = n28535 ;
  assign y6836 = ~n28537 ;
  assign y6837 = ~n28542 ;
  assign y6838 = ~n28543 ;
  assign y6839 = ~n28549 ;
  assign y6840 = n28551 ;
  assign y6841 = ~n28553 ;
  assign y6842 = n28556 ;
  assign y6843 = n28558 ;
  assign y6844 = n28560 ;
  assign y6845 = ~n28561 ;
  assign y6846 = ~n28565 ;
  assign y6847 = n28567 ;
  assign y6848 = ~n28569 ;
  assign y6849 = ~n28571 ;
  assign y6850 = ~n28572 ;
  assign y6851 = n28573 ;
  assign y6852 = ~n28574 ;
  assign y6853 = ~n28576 ;
  assign y6854 = ~n28578 ;
  assign y6855 = n28581 ;
  assign y6856 = n28582 ;
  assign y6857 = ~n28583 ;
  assign y6858 = ~n28584 ;
  assign y6859 = ~n28585 ;
  assign y6860 = n28588 ;
  assign y6861 = n28589 ;
  assign y6862 = n28595 ;
  assign y6863 = n28602 ;
  assign y6864 = n28603 ;
  assign y6865 = n28604 ;
  assign y6866 = n28607 ;
  assign y6867 = ~n28608 ;
  assign y6868 = n28609 ;
  assign y6869 = ~n28610 ;
  assign y6870 = ~n28613 ;
  assign y6871 = n28615 ;
  assign y6872 = n28616 ;
  assign y6873 = ~n28617 ;
  assign y6874 = ~n28618 ;
  assign y6875 = n28619 ;
  assign y6876 = n28621 ;
  assign y6877 = ~n28623 ;
  assign y6878 = ~n28624 ;
  assign y6879 = n28627 ;
  assign y6880 = n28629 ;
  assign y6881 = ~n28631 ;
  assign y6882 = ~n28632 ;
  assign y6883 = n28635 ;
  assign y6884 = ~n28641 ;
  assign y6885 = ~n28643 ;
  assign y6886 = ~n28647 ;
  assign y6887 = n28651 ;
  assign y6888 = ~n28652 ;
  assign y6889 = ~n28654 ;
  assign y6890 = n28655 ;
  assign y6891 = n28656 ;
  assign y6892 = ~n28657 ;
  assign y6893 = ~n28660 ;
  assign y6894 = n28662 ;
  assign y6895 = n28663 ;
  assign y6896 = ~n28664 ;
  assign y6897 = n28665 ;
  assign y6898 = n28669 ;
  assign y6899 = n28671 ;
  assign y6900 = n28672 ;
  assign y6901 = n28675 ;
  assign y6902 = n28678 ;
  assign y6903 = ~n28680 ;
  assign y6904 = ~n28684 ;
  assign y6905 = n28685 ;
  assign y6906 = ~n28690 ;
  assign y6907 = ~n28691 ;
  assign y6908 = ~n28697 ;
  assign y6909 = ~n28700 ;
  assign y6910 = ~n28701 ;
  assign y6911 = ~n28702 ;
  assign y6912 = ~n28703 ;
  assign y6913 = ~n28704 ;
  assign y6914 = ~n28705 ;
  assign y6915 = n28708 ;
  assign y6916 = n28709 ;
  assign y6917 = n28711 ;
  assign y6918 = n28712 ;
  assign y6919 = n28714 ;
  assign y6920 = ~n28719 ;
  assign y6921 = n28721 ;
  assign y6922 = n28722 ;
  assign y6923 = ~n28723 ;
  assign y6924 = n28724 ;
  assign y6925 = ~n28725 ;
  assign y6926 = ~n28727 ;
  assign y6927 = n28730 ;
  assign y6928 = ~n28736 ;
  assign y6929 = n28739 ;
  assign y6930 = ~n28741 ;
  assign y6931 = ~n28743 ;
  assign y6932 = n28744 ;
  assign y6933 = ~n28745 ;
  assign y6934 = ~n28746 ;
  assign y6935 = ~n28747 ;
  assign y6936 = ~n28748 ;
  assign y6937 = ~n28751 ;
  assign y6938 = n28756 ;
  assign y6939 = n28757 ;
  assign y6940 = n28760 ;
  assign y6941 = ~n28761 ;
  assign y6942 = ~n28764 ;
  assign y6943 = n28766 ;
  assign y6944 = ~n28769 ;
  assign y6945 = ~n28771 ;
  assign y6946 = ~n28772 ;
  assign y6947 = ~n28774 ;
  assign y6948 = n28776 ;
  assign y6949 = n28780 ;
  assign y6950 = ~n28783 ;
  assign y6951 = ~n28784 ;
  assign y6952 = ~n28785 ;
  assign y6953 = n28787 ;
  assign y6954 = n28789 ;
  assign y6955 = ~n28794 ;
  assign y6956 = n28795 ;
  assign y6957 = n28799 ;
  assign y6958 = n28802 ;
  assign y6959 = n28803 ;
  assign y6960 = n28804 ;
  assign y6961 = n28805 ;
  assign y6962 = ~n28807 ;
  assign y6963 = n28809 ;
  assign y6964 = ~n28811 ;
  assign y6965 = ~n28812 ;
  assign y6966 = ~n28815 ;
  assign y6967 = ~n28818 ;
  assign y6968 = n28821 ;
  assign y6969 = n28823 ;
  assign y6970 = n28829 ;
  assign y6971 = n28830 ;
  assign y6972 = ~n28833 ;
  assign y6973 = n28837 ;
  assign y6974 = ~n28840 ;
  assign y6975 = n28841 ;
  assign y6976 = n28844 ;
  assign y6977 = ~n28847 ;
  assign y6978 = n28855 ;
  assign y6979 = ~n28857 ;
  assign y6980 = n28858 ;
  assign y6981 = n28859 ;
  assign y6982 = ~n28860 ;
  assign y6983 = n28861 ;
  assign y6984 = n28863 ;
  assign y6985 = n28864 ;
  assign y6986 = ~n28868 ;
  assign y6987 = n28869 ;
  assign y6988 = ~n28871 ;
  assign y6989 = n28872 ;
  assign y6990 = n28876 ;
  assign y6991 = ~n28885 ;
  assign y6992 = n28887 ;
  assign y6993 = ~n28888 ;
  assign y6994 = n28893 ;
  assign y6995 = ~n28895 ;
  assign y6996 = n28897 ;
  assign y6997 = n28902 ;
  assign y6998 = n28904 ;
  assign y6999 = ~n28905 ;
  assign y7000 = ~n28906 ;
  assign y7001 = n28907 ;
  assign y7002 = n28912 ;
  assign y7003 = n28913 ;
  assign y7004 = n28916 ;
  assign y7005 = ~n28917 ;
  assign y7006 = n28920 ;
  assign y7007 = n28921 ;
  assign y7008 = ~n28923 ;
  assign y7009 = ~n28924 ;
  assign y7010 = n28925 ;
  assign y7011 = n28932 ;
  assign y7012 = ~n28933 ;
  assign y7013 = n28934 ;
  assign y7014 = ~n28936 ;
  assign y7015 = ~n28940 ;
  assign y7016 = n28943 ;
  assign y7017 = n28945 ;
  assign y7018 = ~n28951 ;
  assign y7019 = n28954 ;
  assign y7020 = ~n28957 ;
  assign y7021 = n28960 ;
  assign y7022 = ~n28961 ;
  assign y7023 = n28962 ;
  assign y7024 = ~n28963 ;
  assign y7025 = n28965 ;
  assign y7026 = n28967 ;
  assign y7027 = n28969 ;
  assign y7028 = n28970 ;
  assign y7029 = ~n28975 ;
  assign y7030 = ~n28977 ;
  assign y7031 = n28978 ;
  assign y7032 = n28980 ;
  assign y7033 = ~n28982 ;
  assign y7034 = ~n28983 ;
  assign y7035 = ~n28984 ;
  assign y7036 = ~n28985 ;
  assign y7037 = n28986 ;
  assign y7038 = n28987 ;
  assign y7039 = ~n28988 ;
  assign y7040 = n28990 ;
  assign y7041 = n28998 ;
  assign y7042 = n29000 ;
  assign y7043 = n29001 ;
  assign y7044 = n29005 ;
  assign y7045 = n29007 ;
  assign y7046 = n29013 ;
  assign y7047 = n29017 ;
  assign y7048 = n29020 ;
  assign y7049 = ~n29021 ;
  assign y7050 = n29022 ;
  assign y7051 = n29024 ;
  assign y7052 = n29025 ;
  assign y7053 = ~n29026 ;
  assign y7054 = n29027 ;
  assign y7055 = n29028 ;
  assign y7056 = ~n29029 ;
  assign y7057 = ~n29030 ;
  assign y7058 = n29032 ;
  assign y7059 = ~n29034 ;
  assign y7060 = ~n29035 ;
  assign y7061 = ~n29036 ;
  assign y7062 = n29038 ;
  assign y7063 = ~n29039 ;
  assign y7064 = ~n29042 ;
  assign y7065 = n29044 ;
  assign y7066 = n29045 ;
  assign y7067 = n29046 ;
  assign y7068 = ~n29047 ;
  assign y7069 = ~n29048 ;
  assign y7070 = n29051 ;
  assign y7071 = n29052 ;
  assign y7072 = n29055 ;
  assign y7073 = n29056 ;
  assign y7074 = ~n29057 ;
  assign y7075 = ~n29059 ;
  assign y7076 = ~n29060 ;
  assign y7077 = ~n29063 ;
  assign y7078 = ~n29064 ;
  assign y7079 = ~n29065 ;
  assign y7080 = ~n29069 ;
  assign y7081 = n29073 ;
  assign y7082 = n29079 ;
  assign y7083 = n29081 ;
  assign y7084 = n29082 ;
  assign y7085 = n29083 ;
  assign y7086 = ~n29084 ;
  assign y7087 = n29088 ;
  assign y7088 = ~n29091 ;
  assign y7089 = ~n29092 ;
  assign y7090 = n29094 ;
  assign y7091 = n29101 ;
  assign y7092 = n29105 ;
  assign y7093 = ~n29107 ;
  assign y7094 = n29109 ;
  assign y7095 = ~n29113 ;
  assign y7096 = ~n29114 ;
  assign y7097 = n29116 ;
  assign y7098 = ~n29120 ;
  assign y7099 = ~n29121 ;
  assign y7100 = ~n29122 ;
  assign y7101 = n29123 ;
  assign y7102 = n29125 ;
  assign y7103 = n29128 ;
  assign y7104 = n29134 ;
  assign y7105 = n29139 ;
  assign y7106 = n29140 ;
  assign y7107 = ~n29143 ;
  assign y7108 = ~n29144 ;
  assign y7109 = ~n29147 ;
  assign y7110 = n29148 ;
  assign y7111 = ~n29149 ;
  assign y7112 = n29150 ;
  assign y7113 = ~n29152 ;
  assign y7114 = n29153 ;
  assign y7115 = n29155 ;
  assign y7116 = n29157 ;
  assign y7117 = n29159 ;
  assign y7118 = n29161 ;
  assign y7119 = n29165 ;
  assign y7120 = n29170 ;
  assign y7121 = n29171 ;
  assign y7122 = ~n29174 ;
  assign y7123 = ~n29176 ;
  assign y7124 = ~n29178 ;
  assign y7125 = ~n29181 ;
  assign y7126 = ~n29184 ;
  assign y7127 = ~n29185 ;
  assign y7128 = n29186 ;
  assign y7129 = n29187 ;
  assign y7130 = n29189 ;
  assign y7131 = n29190 ;
  assign y7132 = n29191 ;
  assign y7133 = n29192 ;
  assign y7134 = ~n29195 ;
  assign y7135 = ~n29198 ;
  assign y7136 = n29199 ;
  assign y7137 = ~n29202 ;
  assign y7138 = n29203 ;
  assign y7139 = ~n29204 ;
  assign y7140 = ~n29207 ;
  assign y7141 = ~n29208 ;
  assign y7142 = n29213 ;
  assign y7143 = ~n29215 ;
  assign y7144 = n29219 ;
  assign y7145 = n29221 ;
  assign y7146 = n29222 ;
  assign y7147 = n29225 ;
  assign y7148 = ~n29229 ;
  assign y7149 = n29230 ;
  assign y7150 = ~n29233 ;
  assign y7151 = n29234 ;
  assign y7152 = n29236 ;
  assign y7153 = ~n29241 ;
  assign y7154 = ~n29242 ;
  assign y7155 = n29247 ;
  assign y7156 = ~n29248 ;
  assign y7157 = ~n29249 ;
  assign y7158 = ~n29253 ;
  assign y7159 = ~n29257 ;
  assign y7160 = ~n29258 ;
  assign y7161 = n29259 ;
  assign y7162 = n29260 ;
  assign y7163 = n29263 ;
  assign y7164 = ~n29265 ;
  assign y7165 = n29267 ;
  assign y7166 = n29269 ;
  assign y7167 = n29270 ;
  assign y7168 = ~n29272 ;
  assign y7169 = n29273 ;
  assign y7170 = ~n29274 ;
  assign y7171 = ~n29276 ;
  assign y7172 = n29279 ;
  assign y7173 = n29280 ;
  assign y7174 = ~n29282 ;
  assign y7175 = n29285 ;
  assign y7176 = n29287 ;
  assign y7177 = ~n29290 ;
  assign y7178 = ~n29294 ;
  assign y7179 = n29295 ;
  assign y7180 = n29297 ;
  assign y7181 = n29299 ;
  assign y7182 = n29302 ;
  assign y7183 = n29304 ;
  assign y7184 = n29305 ;
  assign y7185 = ~n29309 ;
  assign y7186 = ~n29311 ;
  assign y7187 = ~n29312 ;
  assign y7188 = ~n29316 ;
  assign y7189 = ~n29318 ;
  assign y7190 = ~n29320 ;
  assign y7191 = n29322 ;
  assign y7192 = ~n29324 ;
  assign y7193 = ~n29330 ;
  assign y7194 = n29331 ;
  assign y7195 = ~n29333 ;
  assign y7196 = ~n29335 ;
  assign y7197 = n29337 ;
  assign y7198 = n29338 ;
  assign y7199 = n29341 ;
  assign y7200 = ~n29343 ;
  assign y7201 = ~n29347 ;
  assign y7202 = n29350 ;
  assign y7203 = n29351 ;
  assign y7204 = n29352 ;
  assign y7205 = ~n29357 ;
  assign y7206 = n29358 ;
  assign y7207 = ~n29359 ;
  assign y7208 = ~n29360 ;
  assign y7209 = n29361 ;
  assign y7210 = ~n29363 ;
  assign y7211 = ~n29366 ;
  assign y7212 = n29369 ;
  assign y7213 = n29373 ;
  assign y7214 = ~n29379 ;
  assign y7215 = n29380 ;
  assign y7216 = ~n29381 ;
  assign y7217 = n29382 ;
  assign y7218 = ~n29386 ;
  assign y7219 = n29388 ;
  assign y7220 = ~n29389 ;
  assign y7221 = n29390 ;
  assign y7222 = n29391 ;
  assign y7223 = ~n29394 ;
  assign y7224 = n29396 ;
  assign y7225 = ~n29399 ;
  assign y7226 = ~n29400 ;
  assign y7227 = n29401 ;
  assign y7228 = n29405 ;
  assign y7229 = n29408 ;
  assign y7230 = ~n29409 ;
  assign y7231 = n29411 ;
  assign y7232 = n29412 ;
  assign y7233 = ~n29413 ;
  assign y7234 = n29415 ;
  assign y7235 = ~n29416 ;
  assign y7236 = n29417 ;
  assign y7237 = ~n29418 ;
  assign y7238 = n29420 ;
  assign y7239 = n29426 ;
  assign y7240 = n29427 ;
  assign y7241 = n29429 ;
  assign y7242 = n29434 ;
  assign y7243 = ~n29435 ;
  assign y7244 = ~n29436 ;
  assign y7245 = n29438 ;
  assign y7246 = ~n29439 ;
  assign y7247 = ~n29441 ;
  assign y7248 = n29444 ;
  assign y7249 = n29446 ;
  assign y7250 = n29447 ;
  assign y7251 = ~n29449 ;
  assign y7252 = n29451 ;
  assign y7253 = ~n29453 ;
  assign y7254 = ~n29454 ;
  assign y7255 = ~n29458 ;
  assign y7256 = n29459 ;
  assign y7257 = n29461 ;
  assign y7258 = ~n29462 ;
  assign y7259 = n29465 ;
  assign y7260 = ~n29467 ;
  assign y7261 = n29469 ;
  assign y7262 = ~n29471 ;
  assign y7263 = n29472 ;
  assign y7264 = ~n29474 ;
  assign y7265 = n29475 ;
  assign y7266 = n29477 ;
  assign y7267 = ~n29478 ;
  assign y7268 = n29480 ;
  assign y7269 = n29481 ;
  assign y7270 = ~n29483 ;
  assign y7271 = ~n29486 ;
  assign y7272 = n29487 ;
  assign y7273 = n29489 ;
  assign y7274 = ~n29490 ;
  assign y7275 = n29492 ;
  assign y7276 = ~n29494 ;
  assign y7277 = ~n29497 ;
  assign y7278 = n29498 ;
  assign y7279 = n29500 ;
  assign y7280 = n29502 ;
  assign y7281 = n29503 ;
  assign y7282 = ~n29504 ;
  assign y7283 = ~n29506 ;
  assign y7284 = ~n29509 ;
  assign y7285 = n29511 ;
  assign y7286 = ~n29512 ;
  assign y7287 = n29515 ;
  assign y7288 = n29517 ;
  assign y7289 = n29519 ;
  assign y7290 = n29522 ;
  assign y7291 = n29523 ;
  assign y7292 = n29525 ;
  assign y7293 = n29527 ;
  assign y7294 = ~n29528 ;
  assign y7295 = ~n29529 ;
  assign y7296 = n29531 ;
  assign y7297 = n29535 ;
  assign y7298 = ~n29537 ;
  assign y7299 = ~n29541 ;
  assign y7300 = ~n29544 ;
  assign y7301 = ~n29547 ;
  assign y7302 = ~n29550 ;
  assign y7303 = n29551 ;
  assign y7304 = ~n29552 ;
  assign y7305 = ~n29555 ;
  assign y7306 = ~n29557 ;
  assign y7307 = n29562 ;
  assign y7308 = ~n29563 ;
  assign y7309 = ~n29565 ;
  assign y7310 = ~n29567 ;
  assign y7311 = n29569 ;
  assign y7312 = n29570 ;
  assign y7313 = n29571 ;
  assign y7314 = n29573 ;
  assign y7315 = n29575 ;
  assign y7316 = ~n29580 ;
  assign y7317 = n29583 ;
  assign y7318 = n29585 ;
  assign y7319 = n29587 ;
  assign y7320 = n29590 ;
  assign y7321 = n29595 ;
  assign y7322 = n29597 ;
  assign y7323 = ~n29598 ;
  assign y7324 = n29601 ;
  assign y7325 = ~n29603 ;
  assign y7326 = ~n29604 ;
  assign y7327 = ~n29605 ;
  assign y7328 = ~n29611 ;
  assign y7329 = ~n29614 ;
  assign y7330 = ~n29615 ;
  assign y7331 = n29618 ;
  assign y7332 = n29619 ;
  assign y7333 = ~n29621 ;
  assign y7334 = n29623 ;
  assign y7335 = ~n29624 ;
  assign y7336 = n29625 ;
  assign y7337 = ~n29627 ;
  assign y7338 = ~n29628 ;
  assign y7339 = n29633 ;
  assign y7340 = ~n29634 ;
  assign y7341 = ~n29636 ;
  assign y7342 = ~n29638 ;
  assign y7343 = ~n29639 ;
  assign y7344 = n29642 ;
  assign y7345 = ~n29644 ;
  assign y7346 = ~n29645 ;
  assign y7347 = n29649 ;
  assign y7348 = ~n29650 ;
  assign y7349 = ~n29651 ;
  assign y7350 = n29652 ;
  assign y7351 = ~n29656 ;
  assign y7352 = ~n29657 ;
  assign y7353 = n29658 ;
  assign y7354 = ~n29659 ;
  assign y7355 = ~n29660 ;
  assign y7356 = ~n29661 ;
  assign y7357 = n29667 ;
  assign y7358 = ~n29668 ;
  assign y7359 = n29669 ;
  assign y7360 = ~n29672 ;
  assign y7361 = ~n29673 ;
  assign y7362 = n29675 ;
  assign y7363 = n29680 ;
  assign y7364 = ~n29681 ;
  assign y7365 = n29682 ;
  assign y7366 = ~n29685 ;
  assign y7367 = n29686 ;
  assign y7368 = ~n29688 ;
  assign y7369 = ~n29689 ;
  assign y7370 = n29696 ;
  assign y7371 = ~n29703 ;
  assign y7372 = n29706 ;
  assign y7373 = ~n29709 ;
  assign y7374 = ~n29710 ;
  assign y7375 = ~n29711 ;
  assign y7376 = n29712 ;
  assign y7377 = ~n29713 ;
  assign y7378 = n29716 ;
  assign y7379 = ~n29717 ;
  assign y7380 = n29726 ;
  assign y7381 = n29727 ;
  assign y7382 = n29728 ;
  assign y7383 = n29729 ;
  assign y7384 = n29731 ;
  assign y7385 = ~n29734 ;
  assign y7386 = n29737 ;
  assign y7387 = ~n29738 ;
  assign y7388 = n29739 ;
  assign y7389 = ~n29740 ;
  assign y7390 = n29742 ;
  assign y7391 = n29745 ;
  assign y7392 = n29746 ;
  assign y7393 = n29747 ;
  assign y7394 = ~n29749 ;
  assign y7395 = ~n29751 ;
  assign y7396 = ~n29752 ;
  assign y7397 = n29753 ;
  assign y7398 = ~n29754 ;
  assign y7399 = n29757 ;
  assign y7400 = n29758 ;
  assign y7401 = n29759 ;
  assign y7402 = n29760 ;
  assign y7403 = ~n29762 ;
  assign y7404 = n29763 ;
  assign y7405 = n29767 ;
  assign y7406 = ~n29773 ;
  assign y7407 = n29775 ;
  assign y7408 = ~n29778 ;
  assign y7409 = n29779 ;
  assign y7410 = ~n29781 ;
  assign y7411 = ~n29785 ;
  assign y7412 = ~n29787 ;
  assign y7413 = ~n29790 ;
  assign y7414 = n29795 ;
  assign y7415 = n29796 ;
  assign y7416 = n29798 ;
  assign y7417 = ~n29801 ;
  assign y7418 = ~n29802 ;
  assign y7419 = ~n29804 ;
  assign y7420 = n29805 ;
  assign y7421 = ~n29807 ;
  assign y7422 = n29810 ;
  assign y7423 = ~n29812 ;
  assign y7424 = n29817 ;
  assign y7425 = n29820 ;
  assign y7426 = n29824 ;
  assign y7427 = ~n29826 ;
  assign y7428 = n29827 ;
  assign y7429 = ~n29828 ;
  assign y7430 = n29829 ;
  assign y7431 = ~n29830 ;
  assign y7432 = n29835 ;
  assign y7433 = ~n29837 ;
  assign y7434 = ~n29840 ;
  assign y7435 = ~n29842 ;
  assign y7436 = n29843 ;
  assign y7437 = ~n29844 ;
  assign y7438 = n29846 ;
  assign y7439 = ~n29849 ;
  assign y7440 = ~n29851 ;
  assign y7441 = n29853 ;
  assign y7442 = n29855 ;
  assign y7443 = ~n29856 ;
  assign y7444 = n29858 ;
  assign y7445 = ~n29859 ;
  assign y7446 = n29860 ;
  assign y7447 = ~n29867 ;
  assign y7448 = n29873 ;
  assign y7449 = n29875 ;
  assign y7450 = ~n29876 ;
  assign y7451 = ~n29878 ;
  assign y7452 = ~n29881 ;
  assign y7453 = ~n29883 ;
  assign y7454 = n29884 ;
  assign y7455 = ~n29890 ;
  assign y7456 = n29891 ;
  assign y7457 = ~n29892 ;
  assign y7458 = n29893 ;
  assign y7459 = ~n29896 ;
  assign y7460 = ~n29898 ;
  assign y7461 = ~n29899 ;
  assign y7462 = n29902 ;
  assign y7463 = ~n29903 ;
  assign y7464 = n29905 ;
  assign y7465 = ~n29906 ;
  assign y7466 = n29908 ;
  assign y7467 = n29909 ;
  assign y7468 = ~n29911 ;
  assign y7469 = n29912 ;
  assign y7470 = ~n29913 ;
  assign y7471 = n29914 ;
  assign y7472 = ~n29919 ;
  assign y7473 = n29924 ;
  assign y7474 = ~n29928 ;
  assign y7475 = n29929 ;
  assign y7476 = ~n29930 ;
  assign y7477 = n29931 ;
  assign y7478 = n29933 ;
  assign y7479 = ~n29934 ;
  assign y7480 = ~n29935 ;
  assign y7481 = n29936 ;
  assign y7482 = n29938 ;
  assign y7483 = ~n29940 ;
  assign y7484 = n29945 ;
  assign y7485 = n29947 ;
  assign y7486 = n29949 ;
  assign y7487 = n29951 ;
  assign y7488 = ~n29953 ;
  assign y7489 = ~n29954 ;
  assign y7490 = n29956 ;
  assign y7491 = n29961 ;
  assign y7492 = ~n29962 ;
  assign y7493 = n29964 ;
  assign y7494 = ~n29966 ;
  assign y7495 = ~n29968 ;
  assign y7496 = ~n29971 ;
  assign y7497 = ~n29972 ;
  assign y7498 = n29974 ;
  assign y7499 = n29976 ;
  assign y7500 = ~n29977 ;
  assign y7501 = ~n29978 ;
  assign y7502 = n29980 ;
  assign y7503 = n29981 ;
  assign y7504 = ~n29984 ;
  assign y7505 = ~n29985 ;
  assign y7506 = n29987 ;
  assign y7507 = ~n29988 ;
  assign y7508 = n29990 ;
  assign y7509 = ~n29993 ;
  assign y7510 = ~n29996 ;
  assign y7511 = n29998 ;
  assign y7512 = n29999 ;
  assign y7513 = ~n30001 ;
  assign y7514 = n30002 ;
  assign y7515 = ~n30004 ;
  assign y7516 = ~n30005 ;
  assign y7517 = n30008 ;
  assign y7518 = ~n30010 ;
  assign y7519 = ~n30011 ;
  assign y7520 = n30012 ;
  assign y7521 = n30016 ;
  assign y7522 = ~n30019 ;
  assign y7523 = ~n30021 ;
  assign y7524 = ~n30024 ;
  assign y7525 = ~n30026 ;
  assign y7526 = ~n30027 ;
  assign y7527 = ~n30029 ;
  assign y7528 = n30034 ;
  assign y7529 = n30035 ;
  assign y7530 = n30038 ;
  assign y7531 = n30040 ;
  assign y7532 = ~n30041 ;
  assign y7533 = n30047 ;
  assign y7534 = ~n30049 ;
  assign y7535 = n30050 ;
  assign y7536 = ~n30052 ;
  assign y7537 = ~n30053 ;
  assign y7538 = n30056 ;
  assign y7539 = ~n30057 ;
  assign y7540 = n30058 ;
  assign y7541 = n30059 ;
  assign y7542 = n30062 ;
  assign y7543 = n30065 ;
  assign y7544 = ~n30068 ;
  assign y7545 = ~n30070 ;
  assign y7546 = n30072 ;
  assign y7547 = n30074 ;
  assign y7548 = n30075 ;
  assign y7549 = n30077 ;
  assign y7550 = n30080 ;
  assign y7551 = ~n30081 ;
  assign y7552 = n30082 ;
  assign y7553 = ~n30086 ;
  assign y7554 = n30087 ;
  assign y7555 = n30089 ;
  assign y7556 = n30092 ;
  assign y7557 = n30096 ;
  assign y7558 = ~n30099 ;
  assign y7559 = ~n30101 ;
  assign y7560 = ~n30104 ;
  assign y7561 = ~n30107 ;
  assign y7562 = n30108 ;
  assign y7563 = ~n30112 ;
  assign y7564 = n30119 ;
  assign y7565 = ~n30120 ;
  assign y7566 = n30122 ;
  assign y7567 = n30123 ;
  assign y7568 = n30126 ;
  assign y7569 = n30128 ;
  assign y7570 = ~n30132 ;
  assign y7571 = ~n30140 ;
  assign y7572 = ~n30143 ;
  assign y7573 = n30144 ;
  assign y7574 = n30148 ;
  assign y7575 = ~n30150 ;
  assign y7576 = n30151 ;
  assign y7577 = ~n30153 ;
  assign y7578 = n30154 ;
  assign y7579 = n30155 ;
  assign y7580 = n30157 ;
  assign y7581 = ~n30159 ;
  assign y7582 = ~n30160 ;
  assign y7583 = ~n30161 ;
  assign y7584 = ~n30164 ;
  assign y7585 = ~n30168 ;
  assign y7586 = ~n30169 ;
  assign y7587 = ~n30170 ;
  assign y7588 = ~n30173 ;
  assign y7589 = ~n30176 ;
  assign y7590 = ~n30181 ;
  assign y7591 = ~n30182 ;
  assign y7592 = n30183 ;
  assign y7593 = ~n30184 ;
  assign y7594 = ~n30187 ;
  assign y7595 = ~n30188 ;
  assign y7596 = ~n30192 ;
  assign y7597 = n30194 ;
  assign y7598 = ~n30195 ;
  assign y7599 = n30196 ;
  assign y7600 = ~n30200 ;
  assign y7601 = ~n30202 ;
  assign y7602 = ~n30204 ;
  assign y7603 = ~n30207 ;
  assign y7604 = n30208 ;
  assign y7605 = n30211 ;
  assign y7606 = ~n30213 ;
  assign y7607 = n30214 ;
  assign y7608 = n30216 ;
  assign y7609 = n30219 ;
  assign y7610 = n30222 ;
  assign y7611 = n30224 ;
  assign y7612 = ~n30225 ;
  assign y7613 = ~n30226 ;
  assign y7614 = n30227 ;
  assign y7615 = ~n30228 ;
  assign y7616 = n30229 ;
  assign y7617 = ~n30230 ;
  assign y7618 = ~n30231 ;
  assign y7619 = n30234 ;
  assign y7620 = ~n30238 ;
  assign y7621 = n30243 ;
  assign y7622 = ~n30245 ;
  assign y7623 = n30248 ;
  assign y7624 = n30249 ;
  assign y7625 = ~n30251 ;
  assign y7626 = n30252 ;
  assign y7627 = ~n30253 ;
  assign y7628 = ~n30255 ;
  assign y7629 = n30256 ;
  assign y7630 = n30258 ;
endmodule
