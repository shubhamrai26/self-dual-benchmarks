module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n149 , n150 , n151 , n153 , n154 , n155 , n157 , n158 , n159 , n161 , n162 , n163 , n165 , n166 , n167 , n169 , n170 , n171 , n173 , n174 , n175 , n177 , n178 , n179 , n181 , n182 , n183 , n185 , n186 , n187 , n189 , n190 , n191 , n193 , n194 , n195 , n198 , n199 , n200 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3241 , n3242 , n3243 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3277 , n3278 , n3279 , n3280 , n3281 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3297 , n3298 , n3299 , n3300 , n3301 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3323 , n3324 , n3325 , n3326 , n3327 , n3329 , n3330 , n3331 , n3332 , n3333 , n3335 , n3336 , n3337 , n3338 , n3339 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3359 , n3360 , n3361 ;
  assign n149 = x108 & x147 ;
  assign n150 = x108 & ~x147 ;
  assign n151 = ~n149 & ~n150 ;
  assign n153 = x83 & x148 ;
  assign n154 = x83 & ~x148 ;
  assign n155 = ~n153 & ~n154 ;
  assign n157 = x104 & x149 ;
  assign n158 = x104 & ~x149 ;
  assign n159 = ~n157 & ~n158 ;
  assign n161 = x103 & x150 ;
  assign n162 = x103 & ~x150 ;
  assign n163 = ~n161 & ~n162 ;
  assign n165 = x102 & x151 ;
  assign n166 = x102 & ~x151 ;
  assign n167 = ~n165 & ~n166 ;
  assign n169 = x105 & x152 ;
  assign n170 = x105 & ~x152 ;
  assign n171 = ~n169 & ~n170 ;
  assign n173 = x107 & x153 ;
  assign n174 = x107 & ~x153 ;
  assign n175 = ~n173 & ~n174 ;
  assign n177 = x101 & x154 ;
  assign n178 = x101 & ~x154 ;
  assign n179 = ~n177 & ~n178 ;
  assign n181 = x126 & x155 ;
  assign n182 = x126 & ~x155 ;
  assign n183 = ~n181 & ~n182 ;
  assign n185 = x121 & x156 ;
  assign n186 = x121 & ~x156 ;
  assign n187 = ~n185 & ~n186 ;
  assign n189 = x1 & x157 ;
  assign n190 = x1 & ~x157 ;
  assign n191 = ~n189 & ~n190 ;
  assign n193 = x0 & x158 ;
  assign n194 = x0 & ~x158 ;
  assign n195 = ~n193 & ~n194 ;
  assign n198 = x130 & x160 ;
  assign n199 = x130 & ~x160 ;
  assign n200 = ~n198 & ~n199 ;
  assign n202 = x128 & x161 ;
  assign n203 = x128 & ~x161 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = ~x13 & ~x14 ;
  assign n206 = ~x6 & ~x7 ;
  assign n207 = n205 & n206 ;
  assign n208 = ~x17 & ~x21 ;
  assign n209 = ~x8 & n208 ;
  assign n210 = ~x12 & n209 ;
  assign n211 = n207 & n210 ;
  assign n212 = ~x18 & ~x19 ;
  assign n213 = ~x4 & ~x16 ;
  assign n214 = n212 & n213 ;
  assign n215 = ~x5 & ~x22 ;
  assign n216 = ~x9 & ~x11 ;
  assign n217 = n215 & n216 ;
  assign n218 = n214 & n217 ;
  assign n219 = n211 & n218 ;
  assign n220 = x54 & ~n219 ;
  assign n221 = ~x0 & ~n220 ;
  assign n222 = n215 & ~n216 ;
  assign n223 = ~x56 & n222 ;
  assign n224 = ~x56 & ~n215 ;
  assign n225 = ~x8 & ~x21 ;
  assign n226 = ~x7 & x13 ;
  assign n227 = n225 & n226 ;
  assign n228 = ~x7 & n225 ;
  assign n229 = x7 & ~n225 ;
  assign n230 = ~n228 & ~n229 ;
  assign n231 = x8 & x21 ;
  assign n232 = ~x13 & ~n231 ;
  assign n233 = n230 & n232 ;
  assign n234 = ~n227 & ~n233 ;
  assign n235 = ~x14 & ~n234 ;
  assign n236 = ~x13 & x14 ;
  assign n237 = n228 & n236 ;
  assign n238 = ~n235 & ~n237 ;
  assign n239 = ~x10 & ~n238 ;
  assign n240 = x10 & n205 ;
  assign n241 = n228 & n240 ;
  assign n242 = ~n239 & ~n241 ;
  assign n243 = n215 & ~n242 ;
  assign n244 = n214 & n243 ;
  assign n245 = ~x17 & n244 ;
  assign n246 = ~x6 & ~x12 ;
  assign n247 = n245 & n246 ;
  assign n248 = ~n224 & ~n247 ;
  assign n249 = n216 & ~n248 ;
  assign n250 = ~n223 & ~n249 ;
  assign n251 = x54 & ~n250 ;
  assign n252 = ~n221 & ~n251 ;
  assign n253 = ~x129 & ~n252 ;
  assign n254 = ~x3 & n253 ;
  assign n304 = ~n254 & x162 ;
  assign n255 = x13 & x14 ;
  assign n256 = x6 & x7 ;
  assign n257 = n255 & n256 ;
  assign n258 = x17 & x21 ;
  assign n259 = x8 & n258 ;
  assign n260 = x12 & n259 ;
  assign n261 = n257 & n260 ;
  assign n262 = x18 & x19 ;
  assign n263 = x4 & x16 ;
  assign n264 = n262 & n263 ;
  assign n265 = x5 & x22 ;
  assign n266 = x9 & x11 ;
  assign n267 = n265 & n266 ;
  assign n268 = n264 & n267 ;
  assign n269 = n261 & n268 ;
  assign n270 = ~x54 & ~n269 ;
  assign n271 = x0 & ~n270 ;
  assign n272 = n265 & ~n266 ;
  assign n273 = x56 & n272 ;
  assign n274 = x56 & ~n265 ;
  assign n275 = x7 & ~x13 ;
  assign n276 = n231 & n275 ;
  assign n277 = x7 & n231 ;
  assign n278 = ~x7 & ~n231 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = x13 & ~n225 ;
  assign n281 = n279 & n280 ;
  assign n282 = ~n276 & ~n281 ;
  assign n283 = x14 & ~n282 ;
  assign n284 = x13 & ~x14 ;
  assign n285 = n277 & n284 ;
  assign n286 = ~n283 & ~n285 ;
  assign n287 = x10 & ~n286 ;
  assign n288 = ~x10 & n255 ;
  assign n289 = n277 & n288 ;
  assign n290 = ~n287 & ~n289 ;
  assign n291 = n265 & ~n290 ;
  assign n292 = n264 & n291 ;
  assign n293 = x17 & n292 ;
  assign n294 = x6 & x12 ;
  assign n295 = n293 & n294 ;
  assign n296 = ~n274 & ~n295 ;
  assign n297 = n266 & ~n296 ;
  assign n298 = ~n273 & ~n297 ;
  assign n299 = ~x54 & ~n298 ;
  assign n300 = ~n271 & ~n299 ;
  assign n301 = x129 & ~n300 ;
  assign n302 = x3 & n301 ;
  assign n305 = n302 & ~x162 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = ~x11 & ~x12 ;
  assign n308 = n225 & n307 ;
  assign n309 = n214 & n308 ;
  assign n310 = ~x10 & ~x22 ;
  assign n311 = ~x7 & ~x13 ;
  assign n312 = ~x5 & ~x6 ;
  assign n313 = n311 & n312 ;
  assign n314 = ~x14 & n313 ;
  assign n315 = n310 & n314 ;
  assign n316 = n309 & n315 ;
  assign n317 = ~x17 & x54 ;
  assign n318 = ~n316 & n317 ;
  assign n319 = ~x1 & ~n318 ;
  assign n320 = ~x14 & x54 ;
  assign n321 = ~x8 & ~x11 ;
  assign n322 = n208 & n321 ;
  assign n323 = ~x5 & n246 ;
  assign n324 = x5 & ~n246 ;
  assign n325 = ~n323 & ~n324 ;
  assign n326 = ~x7 & ~n294 ;
  assign n327 = n325 & n326 ;
  assign n328 = x7 & n323 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = ~x13 & ~n329 ;
  assign n331 = n226 & n323 ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = ~x9 & ~n332 ;
  assign n334 = n311 & n323 ;
  assign n335 = x9 & n334 ;
  assign n336 = ~n333 & ~n335 ;
  assign n337 = n214 & ~n336 ;
  assign n338 = n322 & n337 ;
  assign n339 = n320 & n338 ;
  assign n340 = n310 & n339 ;
  assign n341 = ~n319 & ~n340 ;
  assign n342 = ~x129 & ~n341 ;
  assign n343 = ~x3 & n342 ;
  assign n382 = ~n343 & x163 ;
  assign n344 = x11 & x12 ;
  assign n345 = n231 & n344 ;
  assign n346 = n264 & n345 ;
  assign n347 = x10 & x22 ;
  assign n348 = x7 & x13 ;
  assign n349 = x5 & x6 ;
  assign n350 = n348 & n349 ;
  assign n351 = x14 & n350 ;
  assign n352 = n347 & n351 ;
  assign n353 = n346 & n352 ;
  assign n354 = x17 & ~x54 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = x1 & ~n355 ;
  assign n357 = x14 & ~x54 ;
  assign n358 = x8 & x11 ;
  assign n359 = n258 & n358 ;
  assign n360 = x5 & n294 ;
  assign n361 = ~x5 & ~n294 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = x7 & ~n246 ;
  assign n364 = n362 & n363 ;
  assign n365 = ~x7 & n360 ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = x13 & ~n366 ;
  assign n368 = n275 & n360 ;
  assign n369 = ~n367 & ~n368 ;
  assign n370 = x9 & ~n369 ;
  assign n371 = n348 & n360 ;
  assign n372 = ~x9 & n371 ;
  assign n373 = ~n370 & ~n372 ;
  assign n374 = n264 & ~n373 ;
  assign n375 = n359 & n374 ;
  assign n376 = n357 & n375 ;
  assign n377 = n347 & n376 ;
  assign n378 = ~n356 & ~n377 ;
  assign n379 = x129 & ~n378 ;
  assign n380 = x3 & n379 ;
  assign n383 = n380 & ~x163 ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = x122 & x127 ;
  assign n386 = ~x45 & ~x48 ;
  assign n387 = ~x43 & ~x47 ;
  assign n388 = n386 & n387 ;
  assign n389 = ~x15 & ~x20 ;
  assign n390 = ~x24 & ~x49 ;
  assign n391 = n389 & n390 ;
  assign n392 = n388 & n391 ;
  assign n393 = ~x41 & ~x46 ;
  assign n394 = ~x38 & ~x50 ;
  assign n395 = n393 & n394 ;
  assign n396 = ~x42 & ~x44 ;
  assign n397 = ~x40 & n396 ;
  assign n398 = ~x2 & n397 ;
  assign n399 = n395 & n398 ;
  assign n400 = n392 & n399 ;
  assign n401 = x82 & ~n400 ;
  assign n402 = ~n385 & ~n401 ;
  assign n403 = ~x65 & n402 ;
  assign n404 = ~x24 & ~x45 ;
  assign n405 = ~x47 & ~x48 ;
  assign n406 = n404 & n405 ;
  assign n407 = ~x49 & n389 ;
  assign n408 = n406 & n407 ;
  assign n409 = ~x38 & ~x40 ;
  assign n410 = n396 & n409 ;
  assign n411 = ~x46 & ~x50 ;
  assign n412 = ~x41 & n411 ;
  assign n413 = n410 & n412 ;
  assign n414 = ~x43 & n413 ;
  assign n415 = n408 & n414 ;
  assign n416 = x82 & ~n415 ;
  assign n417 = ~x82 & n385 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = x2 & ~n418 ;
  assign n420 = ~n403 & ~n419 ;
  assign n421 = ~x129 & ~n420 ;
  assign n460 = n421 & x164 ;
  assign n422 = ~x122 & ~x127 ;
  assign n423 = x45 & x48 ;
  assign n424 = x43 & x47 ;
  assign n425 = n423 & n424 ;
  assign n426 = x15 & x20 ;
  assign n427 = x24 & x49 ;
  assign n428 = n426 & n427 ;
  assign n429 = n425 & n428 ;
  assign n430 = x41 & x46 ;
  assign n431 = x38 & x50 ;
  assign n432 = n430 & n431 ;
  assign n433 = x42 & x44 ;
  assign n434 = x40 & n433 ;
  assign n435 = x2 & n434 ;
  assign n436 = n432 & n435 ;
  assign n437 = n429 & n436 ;
  assign n438 = ~x82 & ~n437 ;
  assign n439 = ~n422 & ~n438 ;
  assign n440 = x65 & n439 ;
  assign n441 = x24 & x45 ;
  assign n442 = x47 & x48 ;
  assign n443 = n441 & n442 ;
  assign n444 = x49 & n426 ;
  assign n445 = n443 & n444 ;
  assign n446 = x38 & x40 ;
  assign n447 = n433 & n446 ;
  assign n448 = x46 & x50 ;
  assign n449 = x41 & n448 ;
  assign n450 = n447 & n449 ;
  assign n451 = x43 & n450 ;
  assign n452 = n445 & n451 ;
  assign n453 = ~x82 & ~n452 ;
  assign n454 = x82 & n422 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = ~x2 & ~n455 ;
  assign n457 = ~n440 & ~n456 ;
  assign n458 = x129 & ~n457 ;
  assign n461 = ~n458 & ~x164 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~x9 & ~x14 ;
  assign n464 = n310 & n463 ;
  assign n465 = n313 & n464 ;
  assign n466 = ~x8 & ~x17 ;
  assign n467 = n307 & n466 ;
  assign n468 = ~x21 & n214 ;
  assign n469 = n467 & n468 ;
  assign n470 = n465 & n469 ;
  assign n471 = ~x61 & ~x118 ;
  assign n472 = ~n470 & n471 ;
  assign n473 = x0 & ~x123 ;
  assign n474 = ~x113 & n473 ;
  assign n475 = ~n472 & ~n474 ;
  assign n476 = ~x129 & ~n475 ;
  assign n492 = n476 & x165 ;
  assign n477 = x9 & x14 ;
  assign n478 = n347 & n477 ;
  assign n479 = n350 & n478 ;
  assign n480 = x8 & x17 ;
  assign n481 = n344 & n480 ;
  assign n482 = x21 & n264 ;
  assign n483 = n481 & n482 ;
  assign n484 = n479 & n483 ;
  assign n485 = x61 & x118 ;
  assign n486 = ~n484 & n485 ;
  assign n487 = ~x0 & x123 ;
  assign n488 = x113 & n487 ;
  assign n489 = ~n486 & ~n488 ;
  assign n490 = x129 & ~n489 ;
  assign n493 = ~n490 & ~x165 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = x10 & ~x22 ;
  assign n496 = n463 & n495 ;
  assign n497 = n334 & n496 ;
  assign n498 = x54 & n214 ;
  assign n499 = n322 & n498 ;
  assign n500 = n497 & n499 ;
  assign n501 = x4 & ~x54 ;
  assign n502 = ~n500 & ~n501 ;
  assign n503 = ~x129 & ~n502 ;
  assign n504 = ~x3 & n503 ;
  assign n516 = n504 & x166 ;
  assign n505 = ~x10 & x22 ;
  assign n506 = n477 & n505 ;
  assign n507 = n371 & n506 ;
  assign n508 = ~x54 & n264 ;
  assign n509 = n359 & n508 ;
  assign n510 = n507 & n509 ;
  assign n511 = ~x4 & x54 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = x129 & ~n512 ;
  assign n514 = x3 & n513 ;
  assign n517 = ~n514 & ~x166 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = x5 & ~x54 ;
  assign n520 = ~x7 & n246 ;
  assign n521 = ~x25 & ~x29 ;
  assign n522 = x28 & n521 ;
  assign n523 = n520 & n522 ;
  assign n524 = ~x13 & n464 ;
  assign n525 = n523 & n524 ;
  assign n526 = ~x59 & n322 ;
  assign n527 = ~x16 & x54 ;
  assign n528 = ~x4 & ~x19 ;
  assign n529 = ~x18 & n528 ;
  assign n530 = ~x5 & n529 ;
  assign n531 = n527 & n530 ;
  assign n532 = n526 & n531 ;
  assign n533 = n525 & n532 ;
  assign n534 = ~n519 & ~n533 ;
  assign n535 = ~x129 & ~n534 ;
  assign n536 = ~x3 & n535 ;
  assign n556 = n536 & x167 ;
  assign n537 = ~x5 & x54 ;
  assign n538 = x7 & n294 ;
  assign n539 = x25 & x29 ;
  assign n540 = ~x28 & n539 ;
  assign n541 = n538 & n540 ;
  assign n542 = x13 & n478 ;
  assign n543 = n541 & n542 ;
  assign n544 = x59 & n359 ;
  assign n545 = x16 & ~x54 ;
  assign n546 = x4 & x19 ;
  assign n547 = x18 & n546 ;
  assign n548 = x5 & n547 ;
  assign n549 = n545 & n548 ;
  assign n550 = n544 & n549 ;
  assign n551 = n543 & n550 ;
  assign n552 = ~n537 & ~n551 ;
  assign n553 = x129 & ~n552 ;
  assign n554 = x3 & n553 ;
  assign n557 = ~n554 & ~x167 ;
  assign n558 = ~n556 & ~n557 ;
  assign n559 = x6 & ~x54 ;
  assign n560 = ~x5 & ~x7 ;
  assign n561 = x25 & ~x29 ;
  assign n562 = ~x28 & n561 ;
  assign n563 = ~x12 & n562 ;
  assign n564 = n560 & n563 ;
  assign n565 = n524 & n564 ;
  assign n566 = ~x6 & n529 ;
  assign n567 = n527 & n566 ;
  assign n568 = n526 & n567 ;
  assign n569 = n565 & n568 ;
  assign n570 = ~n559 & ~n569 ;
  assign n571 = ~x129 & ~n570 ;
  assign n572 = ~x3 & n571 ;
  assign n588 = n572 & x168 ;
  assign n573 = ~x6 & x54 ;
  assign n574 = x5 & x7 ;
  assign n575 = ~x25 & x29 ;
  assign n576 = x28 & n575 ;
  assign n577 = x12 & n576 ;
  assign n578 = n574 & n577 ;
  assign n579 = n542 & n578 ;
  assign n580 = x6 & n547 ;
  assign n581 = n545 & n580 ;
  assign n582 = n544 & n581 ;
  assign n583 = n579 & n582 ;
  assign n584 = ~n573 & ~n583 ;
  assign n585 = x129 & ~n584 ;
  assign n586 = x3 & n585 ;
  assign n589 = ~n586 & ~x168 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = x7 & ~x54 ;
  assign n592 = ~x18 & ~x21 ;
  assign n593 = x8 & ~x17 ;
  assign n594 = n592 & n593 ;
  assign n595 = ~x7 & n528 ;
  assign n596 = n527 & n595 ;
  assign n597 = n594 & n596 ;
  assign n598 = ~x6 & n307 ;
  assign n599 = ~x5 & n598 ;
  assign n600 = n524 & n599 ;
  assign n601 = n597 & n600 ;
  assign n602 = ~n591 & ~n601 ;
  assign n603 = ~x129 & ~n602 ;
  assign n604 = ~x3 & n603 ;
  assign n620 = n604 & x169 ;
  assign n605 = ~x7 & x54 ;
  assign n606 = x18 & x21 ;
  assign n607 = ~x8 & x17 ;
  assign n608 = n606 & n607 ;
  assign n609 = x7 & n546 ;
  assign n610 = n545 & n609 ;
  assign n611 = n608 & n610 ;
  assign n612 = x6 & n344 ;
  assign n613 = x5 & n612 ;
  assign n614 = n542 & n613 ;
  assign n615 = n611 & n614 ;
  assign n616 = ~n605 & ~n615 ;
  assign n617 = x129 & ~n616 ;
  assign n618 = x3 & n617 ;
  assign n621 = ~n618 & ~x169 ;
  assign n622 = ~n620 & ~n621 ;
  assign n623 = x8 & ~x54 ;
  assign n624 = n334 & n464 ;
  assign n625 = ~x17 & ~x18 ;
  assign n626 = ~x11 & x21 ;
  assign n627 = n625 & n626 ;
  assign n628 = ~x8 & n528 ;
  assign n629 = n527 & n628 ;
  assign n630 = n627 & n629 ;
  assign n631 = n624 & n630 ;
  assign n632 = ~n623 & ~n631 ;
  assign n633 = ~x129 & ~n632 ;
  assign n634 = ~x3 & n633 ;
  assign n648 = n634 & x170 ;
  assign n635 = ~x8 & x54 ;
  assign n636 = n371 & n478 ;
  assign n637 = x17 & x18 ;
  assign n638 = x11 & ~x21 ;
  assign n639 = n637 & n638 ;
  assign n640 = x8 & n546 ;
  assign n641 = n545 & n640 ;
  assign n642 = n639 & n641 ;
  assign n643 = n636 & n642 ;
  assign n644 = ~n635 & ~n643 ;
  assign n645 = x129 & ~n644 ;
  assign n646 = x3 & n645 ;
  assign n649 = ~n646 & ~x170 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = x9 & ~x54 ;
  assign n652 = n205 & n310 ;
  assign n653 = x11 & n560 ;
  assign n654 = n246 & n653 ;
  assign n655 = n652 & n654 ;
  assign n656 = n466 & n592 ;
  assign n657 = ~x9 & n528 ;
  assign n658 = n527 & n657 ;
  assign n659 = n656 & n658 ;
  assign n660 = n655 & n659 ;
  assign n661 = ~n651 & ~n660 ;
  assign n662 = ~x129 & ~n661 ;
  assign n663 = ~x3 & n662 ;
  assign n678 = n663 & x171 ;
  assign n664 = ~x9 & x54 ;
  assign n665 = n255 & n347 ;
  assign n666 = ~x11 & n574 ;
  assign n667 = n294 & n666 ;
  assign n668 = n665 & n667 ;
  assign n669 = n480 & n606 ;
  assign n670 = x9 & n546 ;
  assign n671 = n545 & n670 ;
  assign n672 = n669 & n671 ;
  assign n673 = n668 & n672 ;
  assign n674 = ~n664 & ~n673 ;
  assign n675 = x129 & ~n674 ;
  assign n676 = x3 & n675 ;
  assign n679 = ~n676 & ~x171 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = x10 & ~x54 ;
  assign n682 = ~x10 & n528 ;
  assign n683 = n527 & n682 ;
  assign n684 = n656 & n683 ;
  assign n685 = n560 & n598 ;
  assign n686 = ~x9 & ~x22 ;
  assign n687 = n236 & n686 ;
  assign n688 = n685 & n687 ;
  assign n689 = n684 & n688 ;
  assign n690 = ~n681 & ~n689 ;
  assign n691 = ~x129 & ~n690 ;
  assign n692 = ~x3 & n691 ;
  assign n706 = n692 & x172 ;
  assign n693 = ~x10 & x54 ;
  assign n694 = x10 & n546 ;
  assign n695 = n545 & n694 ;
  assign n696 = n669 & n695 ;
  assign n697 = n574 & n612 ;
  assign n698 = x9 & x22 ;
  assign n699 = n284 & n698 ;
  assign n700 = n697 & n699 ;
  assign n701 = n696 & n700 ;
  assign n702 = ~n693 & ~n701 ;
  assign n703 = x129 & ~n702 ;
  assign n704 = x3 & n703 ;
  assign n707 = ~n704 & ~x172 ;
  assign n708 = ~n706 & ~n707 ;
  assign n709 = x11 & ~x54 ;
  assign n710 = ~x11 & n528 ;
  assign n711 = n527 & n710 ;
  assign n712 = n656 & n711 ;
  assign n713 = n463 & n505 ;
  assign n714 = n334 & n713 ;
  assign n715 = n712 & n714 ;
  assign n716 = ~n709 & ~n715 ;
  assign n717 = ~x129 & ~n716 ;
  assign n718 = ~x3 & n717 ;
  assign n730 = n718 & x173 ;
  assign n719 = ~x11 & x54 ;
  assign n720 = x11 & n546 ;
  assign n721 = n545 & n720 ;
  assign n722 = n669 & n721 ;
  assign n723 = n477 & n495 ;
  assign n724 = n371 & n723 ;
  assign n725 = n722 & n724 ;
  assign n726 = ~n719 & ~n725 ;
  assign n727 = x129 & ~n726 ;
  assign n728 = x3 & n727 ;
  assign n731 = ~n728 & ~x173 ;
  assign n732 = ~n730 & ~n731 ;
  assign n733 = x12 & ~x54 ;
  assign n734 = ~x12 & n528 ;
  assign n735 = n527 & n734 ;
  assign n736 = x18 & n209 ;
  assign n737 = n735 & n736 ;
  assign n738 = ~x11 & n465 ;
  assign n739 = n737 & n738 ;
  assign n740 = ~n733 & ~n739 ;
  assign n741 = ~x129 & ~n740 ;
  assign n742 = ~x3 & n741 ;
  assign n754 = n742 & x174 ;
  assign n743 = ~x12 & x54 ;
  assign n744 = x12 & n546 ;
  assign n745 = n545 & n744 ;
  assign n746 = ~x18 & n259 ;
  assign n747 = n745 & n746 ;
  assign n748 = x11 & n479 ;
  assign n749 = n747 & n748 ;
  assign n750 = ~n743 & ~n749 ;
  assign n751 = x129 & ~n750 ;
  assign n752 = x3 & n751 ;
  assign n755 = ~n752 & ~x174 ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = x13 & ~x54 ;
  assign n758 = ~x13 & n529 ;
  assign n759 = n527 & n758 ;
  assign n760 = n526 & n759 ;
  assign n761 = ~x28 & n575 ;
  assign n762 = n323 & n761 ;
  assign n763 = ~x7 & n464 ;
  assign n764 = n762 & n763 ;
  assign n765 = n760 & n764 ;
  assign n766 = ~n757 & ~n765 ;
  assign n767 = ~x129 & ~n766 ;
  assign n768 = ~x3 & n767 ;
  assign n782 = n768 & x175 ;
  assign n769 = ~x13 & x54 ;
  assign n770 = x13 & n547 ;
  assign n771 = n545 & n770 ;
  assign n772 = n544 & n771 ;
  assign n773 = x28 & n561 ;
  assign n774 = n360 & n773 ;
  assign n775 = x7 & n478 ;
  assign n776 = n774 & n775 ;
  assign n777 = n772 & n776 ;
  assign n778 = ~n769 & ~n777 ;
  assign n779 = x129 & ~n778 ;
  assign n780 = x3 & n779 ;
  assign n783 = ~n780 & ~x175 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~x16 & n320 ;
  assign n786 = n528 & n785 ;
  assign n787 = n656 & n786 ;
  assign n788 = ~x9 & x13 ;
  assign n789 = n310 & n788 ;
  assign n790 = n685 & n789 ;
  assign n791 = n787 & n790 ;
  assign n792 = ~n357 & ~n791 ;
  assign n793 = ~x129 & ~n792 ;
  assign n794 = ~x3 & n793 ;
  assign n806 = n794 & x176 ;
  assign n795 = x16 & n357 ;
  assign n796 = n546 & n795 ;
  assign n797 = n669 & n796 ;
  assign n798 = x9 & ~x13 ;
  assign n799 = n347 & n798 ;
  assign n800 = n697 & n799 ;
  assign n801 = n797 & n800 ;
  assign n802 = ~n320 & ~n801 ;
  assign n803 = x129 & ~n802 ;
  assign n804 = x3 & n803 ;
  assign n807 = ~n804 & ~x176 ;
  assign n808 = ~n806 & ~n807 ;
  assign n809 = ~x41 & ~x43 ;
  assign n810 = n405 & n809 ;
  assign n811 = ~x45 & n390 ;
  assign n812 = n810 & n811 ;
  assign n813 = ~x46 & n394 ;
  assign n814 = n397 & n813 ;
  assign n815 = ~x15 & n814 ;
  assign n816 = n812 & n815 ;
  assign n817 = x82 & ~n816 ;
  assign n818 = ~n385 & ~n817 ;
  assign n819 = ~x70 & n818 ;
  assign n820 = ~x48 & n387 ;
  assign n821 = n811 & n820 ;
  assign n822 = n413 & n821 ;
  assign n823 = x15 & ~n822 ;
  assign n824 = ~x45 & n405 ;
  assign n825 = ~x2 & ~x20 ;
  assign n826 = ~x15 & ~n825 ;
  assign n827 = n414 & n826 ;
  assign n828 = n390 & n827 ;
  assign n829 = n824 & n828 ;
  assign n830 = ~n823 & ~n829 ;
  assign n831 = x82 & ~n830 ;
  assign n832 = x15 & n417 ;
  assign n833 = ~n831 & ~n832 ;
  assign n834 = ~n819 & n833 ;
  assign n835 = ~x129 & ~n834 ;
  assign n864 = n835 & x177 ;
  assign n836 = x41 & x43 ;
  assign n837 = n442 & n836 ;
  assign n838 = x45 & n427 ;
  assign n839 = n837 & n838 ;
  assign n840 = x46 & n431 ;
  assign n841 = n434 & n840 ;
  assign n842 = x15 & n841 ;
  assign n843 = n839 & n842 ;
  assign n844 = ~x82 & ~n843 ;
  assign n845 = ~n422 & ~n844 ;
  assign n846 = x70 & n845 ;
  assign n847 = x48 & n424 ;
  assign n848 = n838 & n847 ;
  assign n849 = n450 & n848 ;
  assign n850 = ~x15 & ~n849 ;
  assign n851 = x45 & n442 ;
  assign n852 = x2 & x20 ;
  assign n853 = x15 & ~n852 ;
  assign n854 = n451 & n853 ;
  assign n855 = n427 & n854 ;
  assign n856 = n851 & n855 ;
  assign n857 = ~n850 & ~n856 ;
  assign n858 = ~x82 & ~n857 ;
  assign n859 = ~x15 & n454 ;
  assign n860 = ~n858 & ~n859 ;
  assign n861 = ~n846 & n860 ;
  assign n862 = x129 & ~n861 ;
  assign n865 = ~n862 & ~x177 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = x6 & ~x12 ;
  assign n868 = ~x5 & n867 ;
  assign n869 = n311 & n868 ;
  assign n870 = n464 & n869 ;
  assign n871 = n499 & n870 ;
  assign n872 = ~n545 & ~n871 ;
  assign n873 = ~x129 & ~n872 ;
  assign n874 = ~x3 & n873 ;
  assign n884 = n874 & x178 ;
  assign n875 = ~x6 & x12 ;
  assign n876 = x5 & n875 ;
  assign n877 = n348 & n876 ;
  assign n878 = n478 & n877 ;
  assign n879 = n509 & n878 ;
  assign n880 = ~n527 & ~n879 ;
  assign n881 = x129 & ~n880 ;
  assign n882 = x3 & n881 ;
  assign n885 = ~n882 & ~x178 ;
  assign n886 = ~n884 & ~n885 ;
  assign n887 = ~x7 & n312 ;
  assign n888 = ~x25 & ~x28 ;
  assign n889 = ~x12 & n888 ;
  assign n890 = n887 & n889 ;
  assign n891 = n524 & n890 ;
  assign n892 = ~x16 & n317 ;
  assign n893 = n529 & n892 ;
  assign n894 = ~x11 & n225 ;
  assign n895 = ~x29 & x59 ;
  assign n896 = n894 & n895 ;
  assign n897 = n893 & n896 ;
  assign n898 = n891 & n897 ;
  assign n899 = ~n354 & ~n898 ;
  assign n900 = ~x129 & ~n899 ;
  assign n901 = ~x3 & n900 ;
  assign n918 = n901 & x179 ;
  assign n902 = x7 & n349 ;
  assign n903 = x25 & x28 ;
  assign n904 = x12 & n903 ;
  assign n905 = n902 & n904 ;
  assign n906 = n542 & n905 ;
  assign n907 = x16 & n354 ;
  assign n908 = n547 & n907 ;
  assign n909 = x11 & n231 ;
  assign n910 = x29 & ~x59 ;
  assign n911 = n909 & n910 ;
  assign n912 = n908 & n911 ;
  assign n913 = n906 & n912 ;
  assign n914 = ~n317 & ~n913 ;
  assign n915 = x129 & ~n914 ;
  assign n916 = x3 & n915 ;
  assign n919 = ~n916 & ~x179 ;
  assign n920 = ~n918 & ~n919 ;
  assign n921 = x18 & ~x54 ;
  assign n922 = x16 & x54 ;
  assign n923 = n529 & n922 ;
  assign n924 = n322 & n923 ;
  assign n925 = n624 & n924 ;
  assign n926 = ~n921 & ~n925 ;
  assign n927 = ~x129 & ~n926 ;
  assign n928 = ~x3 & n927 ;
  assign n938 = n928 & x180 ;
  assign n929 = ~x18 & x54 ;
  assign n930 = ~x16 & ~x54 ;
  assign n931 = n547 & n930 ;
  assign n932 = n359 & n931 ;
  assign n933 = n636 & n932 ;
  assign n934 = ~n929 & ~n933 ;
  assign n935 = x129 & ~n934 ;
  assign n936 = x3 & n935 ;
  assign n939 = ~n936 & ~x180 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = x19 & ~x54 ;
  assign n942 = x17 & n894 ;
  assign n943 = ~x4 & ~x18 ;
  assign n944 = ~x19 & n943 ;
  assign n945 = n527 & n944 ;
  assign n946 = n942 & n945 ;
  assign n947 = n624 & n946 ;
  assign n948 = ~n941 & ~n947 ;
  assign n949 = ~x129 & ~n948 ;
  assign n950 = ~x3 & n949 ;
  assign n962 = n950 & x181 ;
  assign n951 = ~x19 & x54 ;
  assign n952 = ~x17 & n909 ;
  assign n953 = x4 & x18 ;
  assign n954 = x19 & n953 ;
  assign n955 = n545 & n954 ;
  assign n956 = n952 & n955 ;
  assign n957 = n636 & n956 ;
  assign n958 = ~n951 & ~n957 ;
  assign n959 = x129 & ~n958 ;
  assign n960 = x3 & n959 ;
  assign n963 = ~n960 & ~x181 ;
  assign n964 = ~n962 & ~n963 ;
  assign n965 = n387 & n393 ;
  assign n966 = ~x24 & n386 ;
  assign n967 = n965 & n966 ;
  assign n968 = ~x40 & ~x42 ;
  assign n969 = n394 & n968 ;
  assign n970 = ~x44 & n407 ;
  assign n971 = n969 & n970 ;
  assign n972 = n967 & n971 ;
  assign n973 = x82 & ~n972 ;
  assign n974 = ~n385 & ~n973 ;
  assign n975 = ~x71 & n974 ;
  assign n976 = ~x50 & n409 ;
  assign n977 = ~x15 & ~x49 ;
  assign n978 = n396 & n977 ;
  assign n979 = n976 & n978 ;
  assign n980 = n967 & n979 ;
  assign n981 = x20 & ~n980 ;
  assign n982 = x2 & n972 ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = x82 & ~n983 ;
  assign n985 = x20 & n417 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~n975 & n986 ;
  assign n988 = ~x129 & ~n987 ;
  assign n1014 = n988 & x182 ;
  assign n989 = n424 & n430 ;
  assign n990 = x24 & n423 ;
  assign n991 = n989 & n990 ;
  assign n992 = x40 & x42 ;
  assign n993 = n431 & n992 ;
  assign n994 = x44 & n444 ;
  assign n995 = n993 & n994 ;
  assign n996 = n991 & n995 ;
  assign n997 = ~x82 & ~n996 ;
  assign n998 = ~n422 & ~n997 ;
  assign n999 = x71 & n998 ;
  assign n1000 = x50 & n446 ;
  assign n1001 = x15 & x49 ;
  assign n1002 = n433 & n1001 ;
  assign n1003 = n1000 & n1002 ;
  assign n1004 = n991 & n1003 ;
  assign n1005 = ~x20 & ~n1004 ;
  assign n1006 = ~x2 & n996 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = ~x82 & ~n1007 ;
  assign n1009 = ~x20 & n454 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = ~n999 & n1010 ;
  assign n1012 = x129 & ~n1011 ;
  assign n1015 = ~n1012 & ~x182 ;
  assign n1016 = ~n1014 & ~n1015 ;
  assign n1017 = x21 & ~x54 ;
  assign n1018 = n321 & n625 ;
  assign n1019 = ~x21 & x54 ;
  assign n1020 = x19 & n1019 ;
  assign n1021 = n213 & n1020 ;
  assign n1022 = n1018 & n1021 ;
  assign n1023 = n624 & n1022 ;
  assign n1024 = ~n1017 & ~n1023 ;
  assign n1025 = ~x129 & ~n1024 ;
  assign n1026 = ~x3 & n1025 ;
  assign n1036 = n1026 & x183 ;
  assign n1027 = n358 & n637 ;
  assign n1028 = ~x19 & n1017 ;
  assign n1029 = n263 & n1028 ;
  assign n1030 = n1027 & n1029 ;
  assign n1031 = n636 & n1030 ;
  assign n1032 = ~n1019 & ~n1031 ;
  assign n1033 = x129 & ~n1032 ;
  assign n1034 = x3 & n1033 ;
  assign n1037 = ~n1034 & ~x183 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = x22 & ~x54 ;
  assign n1040 = ~x22 & n528 ;
  assign n1041 = n527 & n1040 ;
  assign n1042 = n656 & n1041 ;
  assign n1043 = ~x9 & ~x10 ;
  assign n1044 = n205 & n1043 ;
  assign n1045 = x5 & ~x7 ;
  assign n1046 = n598 & n1045 ;
  assign n1047 = n1044 & n1046 ;
  assign n1048 = n1042 & n1047 ;
  assign n1049 = ~n1039 & ~n1048 ;
  assign n1050 = ~x129 & ~n1049 ;
  assign n1051 = ~x3 & n1050 ;
  assign n1066 = n1051 & x184 ;
  assign n1052 = ~x22 & x54 ;
  assign n1053 = x22 & n546 ;
  assign n1054 = n545 & n1053 ;
  assign n1055 = n669 & n1054 ;
  assign n1056 = x9 & x10 ;
  assign n1057 = n255 & n1056 ;
  assign n1058 = ~x5 & x7 ;
  assign n1059 = n612 & n1058 ;
  assign n1060 = n1057 & n1059 ;
  assign n1061 = n1055 & n1060 ;
  assign n1062 = ~n1052 & ~n1061 ;
  assign n1063 = x129 & ~n1062 ;
  assign n1064 = x3 & n1063 ;
  assign n1067 = ~n1064 & ~x184 ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1069 = ~x23 & x55 ;
  assign n1070 = ~x129 & ~n1069 ;
  assign n1071 = x61 & n1070 ;
  assign n1076 = n1071 & x185 ;
  assign n1072 = x23 & ~x55 ;
  assign n1073 = x129 & ~n1072 ;
  assign n1074 = ~x61 & n1073 ;
  assign n1077 = ~n1074 & ~x185 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1079 = ~x47 & n809 ;
  assign n1080 = n386 & n1079 ;
  assign n1081 = n814 & n1080 ;
  assign n1082 = x82 & ~n1081 ;
  assign n1083 = n825 & n977 ;
  assign n1084 = x82 & ~n1083 ;
  assign n1085 = n385 & ~n1084 ;
  assign n1086 = ~n1082 & ~n1085 ;
  assign n1087 = ~x24 & ~n1086 ;
  assign n1088 = ~x2 & ~x45 ;
  assign n1089 = n405 & n1088 ;
  assign n1090 = n407 & n1089 ;
  assign n1091 = n414 & n1090 ;
  assign n1092 = x82 & ~n1091 ;
  assign n1093 = ~n385 & ~n1092 ;
  assign n1094 = x63 & n1093 ;
  assign n1095 = ~x43 & n393 ;
  assign n1096 = n824 & n1095 ;
  assign n1097 = x24 & x82 ;
  assign n1098 = n396 & n1097 ;
  assign n1099 = n976 & n1098 ;
  assign n1100 = n1096 & n1099 ;
  assign n1101 = ~x129 & ~n1100 ;
  assign n1102 = ~n1094 & n1101 ;
  assign n1103 = ~n1087 & n1102 ;
  assign n1130 = n1103 & x186 ;
  assign n1104 = x47 & n836 ;
  assign n1105 = n423 & n1104 ;
  assign n1106 = n841 & n1105 ;
  assign n1107 = ~x82 & ~n1106 ;
  assign n1108 = n852 & n1001 ;
  assign n1109 = ~x82 & ~n1108 ;
  assign n1110 = n422 & ~n1109 ;
  assign n1111 = ~n1107 & ~n1110 ;
  assign n1112 = x24 & ~n1111 ;
  assign n1113 = x2 & x45 ;
  assign n1114 = n442 & n1113 ;
  assign n1115 = n444 & n1114 ;
  assign n1116 = n451 & n1115 ;
  assign n1117 = ~x82 & ~n1116 ;
  assign n1118 = ~n422 & ~n1117 ;
  assign n1119 = ~x63 & n1118 ;
  assign n1120 = x43 & n430 ;
  assign n1121 = n851 & n1120 ;
  assign n1122 = ~x24 & ~x82 ;
  assign n1123 = n433 & n1122 ;
  assign n1124 = n1000 & n1123 ;
  assign n1125 = n1121 & n1124 ;
  assign n1126 = x129 & ~n1125 ;
  assign n1127 = ~n1119 & n1126 ;
  assign n1128 = ~n1112 & n1127 ;
  assign n1131 = ~n1128 & ~x186 ;
  assign n1132 = ~n1130 & ~n1131 ;
  assign n1133 = x85 & x116 ;
  assign n1134 = ~x85 & ~x110 ;
  assign n1135 = ~x96 & n1134 ;
  assign n1136 = ~n1133 & ~n1135 ;
  assign n1137 = x100 & ~n1136 ;
  assign n1138 = x25 & ~x116 ;
  assign n1139 = x85 & n1138 ;
  assign n1140 = ~n1137 & ~n1139 ;
  assign n1141 = ~x26 & ~n1140 ;
  assign n1142 = ~x51 & ~x52 ;
  assign n1143 = ~x39 & n1142 ;
  assign n1144 = ~x95 & ~x100 ;
  assign n1145 = ~x97 & n1144 ;
  assign n1146 = ~x110 & ~n1145 ;
  assign n1147 = x25 & ~n1146 ;
  assign n1148 = x26 & x116 ;
  assign n1149 = ~n1147 & ~n1148 ;
  assign n1150 = ~n1143 & ~n1149 ;
  assign n1151 = x26 & n1138 ;
  assign n1152 = ~n1150 & ~n1151 ;
  assign n1153 = ~x85 & ~n1152 ;
  assign n1154 = ~n1141 & ~n1153 ;
  assign n1155 = ~x27 & ~n1154 ;
  assign n1156 = ~x39 & ~x52 ;
  assign n1157 = ~x51 & n1156 ;
  assign n1158 = x116 & n1157 ;
  assign n1159 = ~n1138 & ~n1158 ;
  assign n1160 = x27 & ~n1159 ;
  assign n1161 = n1143 & n1147 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~x26 & ~x85 ;
  assign n1164 = ~n1162 & n1163 ;
  assign n1165 = ~n1155 & ~n1164 ;
  assign n1166 = ~x53 & ~n1165 ;
  assign n1167 = x25 & ~x26 ;
  assign n1168 = ~x116 & n1167 ;
  assign n1169 = x53 & ~x85 ;
  assign n1170 = ~x27 & n1169 ;
  assign n1171 = n1168 & n1170 ;
  assign n1172 = ~n1166 & ~n1171 ;
  assign n1173 = ~x58 & ~n1172 ;
  assign n1174 = ~x27 & ~x85 ;
  assign n1175 = ~x53 & x58 ;
  assign n1176 = n1174 & n1175 ;
  assign n1177 = n1168 & n1176 ;
  assign n1178 = ~n1173 & ~n1177 ;
  assign n1179 = ~x129 & ~n1178 ;
  assign n1180 = ~x3 & n1179 ;
  assign n1230 = n1180 & x187 ;
  assign n1181 = ~x85 & ~x116 ;
  assign n1182 = x85 & x110 ;
  assign n1183 = x96 & n1182 ;
  assign n1184 = ~n1181 & ~n1183 ;
  assign n1185 = ~x100 & ~n1184 ;
  assign n1186 = ~x25 & x116 ;
  assign n1187 = ~x85 & n1186 ;
  assign n1188 = ~n1185 & ~n1187 ;
  assign n1189 = x26 & ~n1188 ;
  assign n1190 = x51 & x52 ;
  assign n1191 = x39 & n1190 ;
  assign n1192 = x95 & x100 ;
  assign n1193 = x97 & n1192 ;
  assign n1194 = x110 & ~n1193 ;
  assign n1195 = ~x25 & ~n1194 ;
  assign n1196 = ~x26 & ~x116 ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = ~n1191 & ~n1197 ;
  assign n1199 = ~x26 & n1186 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1201 = x85 & ~n1200 ;
  assign n1202 = ~n1189 & ~n1201 ;
  assign n1203 = x27 & ~n1202 ;
  assign n1204 = x39 & x52 ;
  assign n1205 = x51 & n1204 ;
  assign n1206 = ~x116 & n1205 ;
  assign n1207 = ~n1186 & ~n1206 ;
  assign n1208 = ~x27 & ~n1207 ;
  assign n1209 = n1191 & n1195 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = x26 & x85 ;
  assign n1212 = ~n1210 & n1211 ;
  assign n1213 = ~n1203 & ~n1212 ;
  assign n1214 = x53 & ~n1213 ;
  assign n1215 = ~x25 & x26 ;
  assign n1216 = x116 & n1215 ;
  assign n1217 = ~x53 & x85 ;
  assign n1218 = x27 & n1217 ;
  assign n1219 = n1216 & n1218 ;
  assign n1220 = ~n1214 & ~n1219 ;
  assign n1221 = x58 & ~n1220 ;
  assign n1222 = x27 & x85 ;
  assign n1223 = x53 & ~x58 ;
  assign n1224 = n1222 & n1223 ;
  assign n1225 = n1216 & n1224 ;
  assign n1226 = ~n1221 & ~n1225 ;
  assign n1227 = x129 & ~n1226 ;
  assign n1228 = x3 & n1227 ;
  assign n1231 = ~n1228 & ~x187 ;
  assign n1232 = ~n1230 & ~n1231 ;
  assign n1233 = x85 & ~x116 ;
  assign n1234 = ~x110 & ~n1233 ;
  assign n1235 = ~n1148 & n1234 ;
  assign n1236 = ~x96 & n1235 ;
  assign n1237 = ~x26 & n1133 ;
  assign n1238 = ~n1236 & ~n1237 ;
  assign n1239 = x100 & ~n1238 ;
  assign n1240 = ~x85 & ~n1158 ;
  assign n1241 = x26 & n1240 ;
  assign n1242 = ~n1239 & ~n1241 ;
  assign n1243 = ~x129 & ~n1242 ;
  assign n1244 = ~x3 & n1243 ;
  assign n1245 = ~x27 & ~x53 ;
  assign n1246 = ~x58 & n1245 ;
  assign n1247 = n1244 & n1246 ;
  assign n1264 = n1247 & x188 ;
  assign n1248 = ~x85 & x116 ;
  assign n1249 = x110 & ~n1248 ;
  assign n1250 = ~n1196 & n1249 ;
  assign n1251 = x96 & n1250 ;
  assign n1252 = x26 & n1181 ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = ~x100 & ~n1253 ;
  assign n1255 = x85 & ~n1206 ;
  assign n1256 = ~x26 & n1255 ;
  assign n1257 = ~n1254 & ~n1256 ;
  assign n1258 = x129 & ~n1257 ;
  assign n1259 = x3 & n1258 ;
  assign n1260 = x27 & x53 ;
  assign n1261 = x58 & n1260 ;
  assign n1262 = n1259 & n1261 ;
  assign n1265 = ~n1262 & ~x188 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = x95 & ~x96 ;
  assign n1268 = x27 & x116 ;
  assign n1269 = n1234 & ~n1268 ;
  assign n1270 = n1267 & n1269 ;
  assign n1271 = ~x27 & n1133 ;
  assign n1272 = ~n1270 & ~n1271 ;
  assign n1273 = ~x100 & ~n1272 ;
  assign n1274 = x27 & n1240 ;
  assign n1275 = ~n1273 & ~n1274 ;
  assign n1276 = ~x129 & ~n1275 ;
  assign n1277 = ~x3 & n1276 ;
  assign n1278 = ~x53 & ~x58 ;
  assign n1279 = ~x26 & n1278 ;
  assign n1280 = n1277 & n1279 ;
  assign n1296 = n1280 & x189 ;
  assign n1281 = ~x95 & x96 ;
  assign n1282 = ~x27 & ~x116 ;
  assign n1283 = n1249 & ~n1282 ;
  assign n1284 = n1281 & n1283 ;
  assign n1285 = x27 & n1181 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = x100 & ~n1286 ;
  assign n1288 = ~x27 & n1255 ;
  assign n1289 = ~n1287 & ~n1288 ;
  assign n1290 = x129 & ~n1289 ;
  assign n1291 = x3 & n1290 ;
  assign n1292 = x53 & x58 ;
  assign n1293 = x26 & n1292 ;
  assign n1294 = n1291 & n1293 ;
  assign n1297 = ~n1294 & ~x189 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = ~x26 & ~n1143 ;
  assign n1300 = ~x27 & n1157 ;
  assign n1301 = ~n1299 & ~n1300 ;
  assign n1302 = ~n1146 & ~n1301 ;
  assign n1303 = x26 & ~x27 ;
  assign n1304 = ~x26 & x27 ;
  assign n1305 = ~n1303 & ~n1304 ;
  assign n1306 = ~x116 & ~n1305 ;
  assign n1307 = ~n1302 & ~n1306 ;
  assign n1308 = x28 & ~n1307 ;
  assign n1309 = ~x26 & ~x100 ;
  assign n1310 = ~x110 & n1309 ;
  assign n1311 = n1267 & n1310 ;
  assign n1312 = n1148 & n1157 ;
  assign n1313 = ~n1311 & ~n1312 ;
  assign n1314 = ~x27 & ~n1313 ;
  assign n1315 = n1268 & n1299 ;
  assign n1316 = ~n1314 & ~n1315 ;
  assign n1317 = ~n1308 & n1316 ;
  assign n1318 = ~x85 & ~n1317 ;
  assign n1319 = x28 & ~x116 ;
  assign n1320 = ~x100 & x116 ;
  assign n1321 = ~n1319 & ~n1320 ;
  assign n1322 = x85 & ~n1321 ;
  assign n1323 = ~x26 & ~x27 ;
  assign n1324 = n1322 & n1323 ;
  assign n1325 = ~n1318 & ~n1324 ;
  assign n1326 = ~x53 & ~n1325 ;
  assign n1327 = ~x27 & x28 ;
  assign n1328 = ~x116 & n1327 ;
  assign n1329 = ~x26 & n1169 ;
  assign n1330 = n1328 & n1329 ;
  assign n1331 = ~n1326 & ~n1330 ;
  assign n1332 = ~x58 & ~n1331 ;
  assign n1333 = n1163 & n1175 ;
  assign n1334 = n1328 & n1333 ;
  assign n1335 = ~n1332 & ~n1334 ;
  assign n1336 = ~x129 & ~n1335 ;
  assign n1337 = ~x3 & n1336 ;
  assign n1375 = n1337 & x190 ;
  assign n1338 = x26 & ~n1191 ;
  assign n1339 = x27 & n1205 ;
  assign n1340 = ~n1338 & ~n1339 ;
  assign n1341 = ~n1194 & ~n1340 ;
  assign n1342 = x116 & ~n1305 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = ~x28 & ~n1343 ;
  assign n1345 = x26 & x100 ;
  assign n1346 = x110 & n1345 ;
  assign n1347 = n1281 & n1346 ;
  assign n1348 = n1196 & n1205 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = x27 & ~n1349 ;
  assign n1351 = n1282 & n1338 ;
  assign n1352 = ~n1350 & ~n1351 ;
  assign n1353 = ~n1344 & n1352 ;
  assign n1354 = x85 & ~n1353 ;
  assign n1355 = ~x28 & x116 ;
  assign n1356 = x100 & ~x116 ;
  assign n1357 = ~n1355 & ~n1356 ;
  assign n1358 = ~x85 & ~n1357 ;
  assign n1359 = x26 & x27 ;
  assign n1360 = n1358 & n1359 ;
  assign n1361 = ~n1354 & ~n1360 ;
  assign n1362 = x53 & ~n1361 ;
  assign n1363 = x27 & ~x28 ;
  assign n1364 = x116 & n1363 ;
  assign n1365 = x26 & n1217 ;
  assign n1366 = n1364 & n1365 ;
  assign n1367 = ~n1362 & ~n1366 ;
  assign n1368 = x58 & ~n1367 ;
  assign n1369 = n1211 & n1223 ;
  assign n1370 = n1364 & n1369 ;
  assign n1371 = ~n1368 & ~n1370 ;
  assign n1372 = x129 & ~n1371 ;
  assign n1373 = x3 & n1372 ;
  assign n1376 = ~n1373 & ~x190 ;
  assign n1377 = ~n1375 & ~n1376 ;
  assign n1378 = x29 & x110 ;
  assign n1379 = x97 & ~x110 ;
  assign n1380 = ~x96 & n1379 ;
  assign n1381 = x29 & ~x97 ;
  assign n1382 = ~n1380 & ~n1381 ;
  assign n1383 = n1144 & ~n1382 ;
  assign n1384 = ~n1378 & ~n1383 ;
  assign n1385 = ~x58 & ~n1384 ;
  assign n1386 = x97 & x116 ;
  assign n1387 = x29 & ~x116 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = x58 & ~n1388 ;
  assign n1390 = ~n1385 & ~n1389 ;
  assign n1391 = ~x53 & ~n1390 ;
  assign n1392 = n1223 & n1387 ;
  assign n1393 = ~n1391 & ~n1392 ;
  assign n1394 = ~x27 & ~n1393 ;
  assign n1395 = x27 & n1387 ;
  assign n1396 = n1278 & n1395 ;
  assign n1397 = ~n1394 & ~n1396 ;
  assign n1398 = ~x85 & ~n1397 ;
  assign n1399 = x85 & n1246 ;
  assign n1400 = n1387 & n1399 ;
  assign n1401 = ~n1398 & ~n1400 ;
  assign n1402 = ~x26 & ~n1401 ;
  assign n1403 = n1174 & n1278 ;
  assign n1404 = x26 & n1403 ;
  assign n1405 = n1387 & n1404 ;
  assign n1406 = ~n1402 & ~n1405 ;
  assign n1407 = ~x129 & ~n1406 ;
  assign n1408 = ~x3 & n1407 ;
  assign n1441 = n1408 & x191 ;
  assign n1409 = ~x29 & ~x110 ;
  assign n1410 = ~x97 & x110 ;
  assign n1411 = x96 & n1410 ;
  assign n1412 = ~x29 & x97 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = n1192 & ~n1413 ;
  assign n1415 = ~n1409 & ~n1414 ;
  assign n1416 = x58 & ~n1415 ;
  assign n1417 = ~x97 & ~x116 ;
  assign n1418 = ~x29 & x116 ;
  assign n1419 = ~n1417 & ~n1418 ;
  assign n1420 = ~x58 & ~n1419 ;
  assign n1421 = ~n1416 & ~n1420 ;
  assign n1422 = x53 & ~n1421 ;
  assign n1423 = n1175 & n1418 ;
  assign n1424 = ~n1422 & ~n1423 ;
  assign n1425 = x27 & ~n1424 ;
  assign n1426 = ~x27 & n1418 ;
  assign n1427 = n1292 & n1426 ;
  assign n1428 = ~n1425 & ~n1427 ;
  assign n1429 = x85 & ~n1428 ;
  assign n1430 = ~x85 & n1261 ;
  assign n1431 = n1418 & n1430 ;
  assign n1432 = ~n1429 & ~n1431 ;
  assign n1433 = x26 & ~n1432 ;
  assign n1434 = n1222 & n1292 ;
  assign n1435 = ~x26 & n1434 ;
  assign n1436 = n1418 & n1435 ;
  assign n1437 = ~n1433 & ~n1436 ;
  assign n1438 = x129 & ~n1437 ;
  assign n1439 = x3 & n1438 ;
  assign n1442 = ~n1439 & ~x191 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = x30 & ~x109 ;
  assign n1445 = x60 & x109 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = ~x106 & ~n1446 ;
  assign n1448 = x88 & x106 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1450 = ~x129 & ~n1449 ;
  assign n1459 = n1450 & x192 ;
  assign n1451 = ~x30 & x109 ;
  assign n1452 = ~x60 & ~x109 ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = x106 & ~n1453 ;
  assign n1455 = ~x88 & ~x106 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = x129 & ~n1456 ;
  assign n1460 = ~n1457 & ~x192 ;
  assign n1461 = ~n1459 & ~n1460 ;
  assign n1462 = x89 & x106 ;
  assign n1463 = x30 & x109 ;
  assign n1464 = x31 & ~x109 ;
  assign n1465 = ~n1463 & ~n1464 ;
  assign n1466 = ~x106 & ~n1465 ;
  assign n1467 = ~n1462 & ~n1466 ;
  assign n1468 = ~x129 & ~n1467 ;
  assign n1477 = n1468 & x193 ;
  assign n1469 = ~x89 & ~x106 ;
  assign n1470 = ~x30 & ~x109 ;
  assign n1471 = ~x31 & x109 ;
  assign n1472 = ~n1470 & ~n1471 ;
  assign n1473 = x106 & ~n1472 ;
  assign n1474 = ~n1469 & ~n1473 ;
  assign n1475 = x129 & ~n1474 ;
  assign n1478 = ~n1475 & ~x193 ;
  assign n1479 = ~n1477 & ~n1478 ;
  assign n1480 = x99 & x106 ;
  assign n1481 = x31 & x109 ;
  assign n1482 = x32 & ~x109 ;
  assign n1483 = ~n1481 & ~n1482 ;
  assign n1484 = ~x106 & ~n1483 ;
  assign n1485 = ~n1480 & ~n1484 ;
  assign n1486 = ~x129 & ~n1485 ;
  assign n1495 = n1486 & x194 ;
  assign n1487 = ~x99 & ~x106 ;
  assign n1488 = ~x31 & ~x109 ;
  assign n1489 = ~x32 & x109 ;
  assign n1490 = ~n1488 & ~n1489 ;
  assign n1491 = x106 & ~n1490 ;
  assign n1492 = ~n1487 & ~n1491 ;
  assign n1493 = x129 & ~n1492 ;
  assign n1496 = ~n1493 & ~x194 ;
  assign n1497 = ~n1495 & ~n1496 ;
  assign n1498 = x90 & x106 ;
  assign n1499 = x32 & x109 ;
  assign n1500 = x33 & ~x109 ;
  assign n1501 = ~n1499 & ~n1500 ;
  assign n1502 = ~x106 & ~n1501 ;
  assign n1503 = ~n1498 & ~n1502 ;
  assign n1504 = ~x129 & ~n1503 ;
  assign n1513 = n1504 & x195 ;
  assign n1505 = ~x90 & ~x106 ;
  assign n1506 = ~x32 & ~x109 ;
  assign n1507 = ~x33 & x109 ;
  assign n1508 = ~n1506 & ~n1507 ;
  assign n1509 = x106 & ~n1508 ;
  assign n1510 = ~n1505 & ~n1509 ;
  assign n1511 = x129 & ~n1510 ;
  assign n1514 = ~n1511 & ~x195 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = x91 & x106 ;
  assign n1517 = x33 & x109 ;
  assign n1518 = x34 & ~x109 ;
  assign n1519 = ~n1517 & ~n1518 ;
  assign n1520 = ~x106 & ~n1519 ;
  assign n1521 = ~n1516 & ~n1520 ;
  assign n1522 = ~x129 & ~n1521 ;
  assign n1531 = n1522 & x196 ;
  assign n1523 = ~x91 & ~x106 ;
  assign n1524 = ~x33 & ~x109 ;
  assign n1525 = ~x34 & x109 ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = x106 & ~n1526 ;
  assign n1528 = ~n1523 & ~n1527 ;
  assign n1529 = x129 & ~n1528 ;
  assign n1532 = ~n1529 & ~x196 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = x92 & x106 ;
  assign n1535 = x34 & x109 ;
  assign n1536 = x35 & ~x109 ;
  assign n1537 = ~n1535 & ~n1536 ;
  assign n1538 = ~x106 & ~n1537 ;
  assign n1539 = ~n1534 & ~n1538 ;
  assign n1540 = ~x129 & ~n1539 ;
  assign n1549 = n1540 & x197 ;
  assign n1541 = ~x92 & ~x106 ;
  assign n1542 = ~x34 & ~x109 ;
  assign n1543 = ~x35 & x109 ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1545 = x106 & ~n1544 ;
  assign n1546 = ~n1541 & ~n1545 ;
  assign n1547 = x129 & ~n1546 ;
  assign n1550 = ~n1547 & ~x197 ;
  assign n1551 = ~n1549 & ~n1550 ;
  assign n1552 = x98 & x106 ;
  assign n1553 = x35 & x109 ;
  assign n1554 = x36 & ~x109 ;
  assign n1555 = ~n1553 & ~n1554 ;
  assign n1556 = ~x106 & ~n1555 ;
  assign n1557 = ~n1552 & ~n1556 ;
  assign n1558 = ~x129 & ~n1557 ;
  assign n1567 = n1558 & x198 ;
  assign n1559 = ~x98 & ~x106 ;
  assign n1560 = ~x35 & ~x109 ;
  assign n1561 = ~x36 & x109 ;
  assign n1562 = ~n1560 & ~n1561 ;
  assign n1563 = x106 & ~n1562 ;
  assign n1564 = ~n1559 & ~n1563 ;
  assign n1565 = x129 & ~n1564 ;
  assign n1568 = ~n1565 & ~x198 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = x93 & x106 ;
  assign n1571 = x36 & x109 ;
  assign n1572 = x37 & ~x109 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = ~x106 & ~n1573 ;
  assign n1575 = ~n1570 & ~n1574 ;
  assign n1576 = ~x129 & ~n1575 ;
  assign n1585 = n1576 & x199 ;
  assign n1577 = ~x93 & ~x106 ;
  assign n1578 = ~x36 & ~x109 ;
  assign n1579 = ~x37 & x109 ;
  assign n1580 = ~n1578 & ~n1579 ;
  assign n1581 = x106 & ~n1580 ;
  assign n1582 = ~n1577 & ~n1581 ;
  assign n1583 = x129 & ~n1582 ;
  assign n1586 = ~n1583 & ~x199 ;
  assign n1587 = ~n1585 & ~n1586 ;
  assign n1588 = x82 & ~n397 ;
  assign n1589 = n412 & n820 ;
  assign n1590 = n391 & n1088 ;
  assign n1591 = n1589 & n1590 ;
  assign n1592 = x82 & ~n1591 ;
  assign n1593 = n385 & ~n1592 ;
  assign n1594 = ~n1588 & ~n1593 ;
  assign n1595 = ~x38 & ~n1594 ;
  assign n1596 = ~x2 & ~x48 ;
  assign n1597 = n404 & n1596 ;
  assign n1598 = n407 & n1597 ;
  assign n1599 = ~x50 & n397 ;
  assign n1600 = n965 & n1599 ;
  assign n1601 = n1598 & n1600 ;
  assign n1602 = x82 & ~n1601 ;
  assign n1603 = ~n385 & ~n1602 ;
  assign n1604 = x74 & n1603 ;
  assign n1605 = ~x44 & x82 ;
  assign n1606 = x38 & n968 ;
  assign n1607 = n1605 & n1606 ;
  assign n1608 = ~x129 & ~n1607 ;
  assign n1609 = ~n1604 & n1608 ;
  assign n1610 = ~n1595 & n1609 ;
  assign n1635 = n1610 & x200 ;
  assign n1611 = ~x82 & ~n434 ;
  assign n1612 = n449 & n847 ;
  assign n1613 = n428 & n1113 ;
  assign n1614 = n1612 & n1613 ;
  assign n1615 = ~x82 & ~n1614 ;
  assign n1616 = n422 & ~n1615 ;
  assign n1617 = ~n1611 & ~n1616 ;
  assign n1618 = x38 & ~n1617 ;
  assign n1619 = x2 & x48 ;
  assign n1620 = n441 & n1619 ;
  assign n1621 = n444 & n1620 ;
  assign n1622 = x50 & n434 ;
  assign n1623 = n989 & n1622 ;
  assign n1624 = n1621 & n1623 ;
  assign n1625 = ~x82 & ~n1624 ;
  assign n1626 = ~n422 & ~n1625 ;
  assign n1627 = ~x74 & n1626 ;
  assign n1628 = x44 & ~x82 ;
  assign n1629 = ~x38 & n992 ;
  assign n1630 = n1628 & n1629 ;
  assign n1631 = x129 & ~n1630 ;
  assign n1632 = ~n1627 & n1631 ;
  assign n1633 = ~n1618 & n1632 ;
  assign n1636 = ~n1633 & ~x200 ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = ~x51 & x109 ;
  assign n1639 = n1156 & n1638 ;
  assign n1640 = ~x106 & ~n1639 ;
  assign n1641 = x109 & n1142 ;
  assign n1642 = x39 & ~n1641 ;
  assign n1643 = n1640 & ~n1642 ;
  assign n1644 = ~x129 & ~n1643 ;
  assign n1653 = n1644 & x201 ;
  assign n1645 = x51 & ~x109 ;
  assign n1646 = n1204 & n1645 ;
  assign n1647 = x106 & ~n1646 ;
  assign n1648 = ~x109 & n1190 ;
  assign n1649 = ~x39 & ~n1648 ;
  assign n1650 = n1647 & ~n1649 ;
  assign n1651 = x129 & ~n1650 ;
  assign n1654 = ~n1651 & ~x201 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = x82 & ~n396 ;
  assign n1657 = n820 & n1590 ;
  assign n1658 = n395 & n1657 ;
  assign n1659 = x82 & ~n1658 ;
  assign n1660 = n385 & ~n1659 ;
  assign n1661 = ~n1656 & ~n1660 ;
  assign n1662 = ~x40 & ~n1661 ;
  assign n1663 = n394 & n396 ;
  assign n1664 = n965 & n1663 ;
  assign n1665 = n1598 & n1664 ;
  assign n1666 = x82 & ~n1665 ;
  assign n1667 = ~n385 & ~n1666 ;
  assign n1668 = x73 & n1667 ;
  assign n1669 = x40 & x82 ;
  assign n1670 = n396 & n1669 ;
  assign n1671 = ~x129 & ~n1670 ;
  assign n1672 = ~n1668 & n1671 ;
  assign n1673 = ~n1662 & n1672 ;
  assign n1693 = n1673 & x202 ;
  assign n1674 = ~x82 & ~n433 ;
  assign n1675 = n847 & n1613 ;
  assign n1676 = n432 & n1675 ;
  assign n1677 = ~x82 & ~n1676 ;
  assign n1678 = n422 & ~n1677 ;
  assign n1679 = ~n1674 & ~n1678 ;
  assign n1680 = x40 & ~n1679 ;
  assign n1681 = n431 & n433 ;
  assign n1682 = n989 & n1681 ;
  assign n1683 = n1621 & n1682 ;
  assign n1684 = ~x82 & ~n1683 ;
  assign n1685 = ~n422 & ~n1684 ;
  assign n1686 = ~x73 & n1685 ;
  assign n1687 = ~x40 & ~x82 ;
  assign n1688 = n433 & n1687 ;
  assign n1689 = x129 & ~n1688 ;
  assign n1690 = ~n1686 & n1689 ;
  assign n1691 = ~n1680 & n1690 ;
  assign n1694 = ~n1691 & ~x202 ;
  assign n1695 = ~n1693 & ~n1694 ;
  assign n1696 = x82 & ~n814 ;
  assign n1697 = x82 & ~n1657 ;
  assign n1698 = n385 & ~n1697 ;
  assign n1699 = ~n1696 & ~n1698 ;
  assign n1700 = ~x41 & ~n1699 ;
  assign n1701 = n387 & n411 ;
  assign n1702 = n410 & n1701 ;
  assign n1703 = n1598 & n1702 ;
  assign n1704 = x82 & ~n1703 ;
  assign n1705 = ~n385 & ~n1704 ;
  assign n1706 = x76 & n1705 ;
  assign n1707 = n409 & n411 ;
  assign n1708 = x41 & x82 ;
  assign n1709 = n396 & n1708 ;
  assign n1710 = n1707 & n1709 ;
  assign n1711 = ~x129 & ~n1710 ;
  assign n1712 = ~n1706 & n1711 ;
  assign n1713 = ~n1700 & n1712 ;
  assign n1733 = n1713 & x203 ;
  assign n1714 = ~x82 & ~n841 ;
  assign n1715 = ~x82 & ~n1675 ;
  assign n1716 = n422 & ~n1715 ;
  assign n1717 = ~n1714 & ~n1716 ;
  assign n1718 = x41 & ~n1717 ;
  assign n1719 = n424 & n448 ;
  assign n1720 = n447 & n1719 ;
  assign n1721 = n1621 & n1720 ;
  assign n1722 = ~x82 & ~n1721 ;
  assign n1723 = ~n422 & ~n1722 ;
  assign n1724 = ~x76 & n1723 ;
  assign n1725 = n446 & n448 ;
  assign n1726 = ~x41 & ~x82 ;
  assign n1727 = n433 & n1726 ;
  assign n1728 = n1725 & n1727 ;
  assign n1729 = x129 & ~n1728 ;
  assign n1730 = ~n1724 & n1729 ;
  assign n1731 = ~n1718 & n1730 ;
  assign n1734 = ~n1731 & ~x203 ;
  assign n1735 = ~n1733 & ~n1734 ;
  assign n1736 = x44 & x82 ;
  assign n1737 = n1079 & n1707 ;
  assign n1738 = n1598 & n1737 ;
  assign n1739 = x82 & ~n1738 ;
  assign n1740 = n385 & ~n1739 ;
  assign n1741 = ~n1736 & ~n1740 ;
  assign n1742 = ~x42 & ~n1741 ;
  assign n1743 = ~x44 & n976 ;
  assign n1744 = n965 & n1743 ;
  assign n1745 = n1598 & n1744 ;
  assign n1746 = x82 & ~n1745 ;
  assign n1747 = ~n385 & ~n1746 ;
  assign n1748 = x72 & n1747 ;
  assign n1749 = x42 & n1605 ;
  assign n1750 = ~x129 & ~n1749 ;
  assign n1751 = ~n1748 & n1750 ;
  assign n1752 = ~n1742 & n1751 ;
  assign n1771 = n1752 & x204 ;
  assign n1753 = ~x44 & ~x82 ;
  assign n1754 = n1104 & n1725 ;
  assign n1755 = n1621 & n1754 ;
  assign n1756 = ~x82 & ~n1755 ;
  assign n1757 = n422 & ~n1756 ;
  assign n1758 = ~n1753 & ~n1757 ;
  assign n1759 = x42 & ~n1758 ;
  assign n1760 = x44 & n1000 ;
  assign n1761 = n989 & n1760 ;
  assign n1762 = n1621 & n1761 ;
  assign n1763 = ~x82 & ~n1762 ;
  assign n1764 = ~n422 & ~n1763 ;
  assign n1765 = ~x72 & n1764 ;
  assign n1766 = ~x42 & n1628 ;
  assign n1767 = x129 & ~n1766 ;
  assign n1768 = ~n1765 & n1767 ;
  assign n1769 = ~n1759 & n1768 ;
  assign n1772 = ~n1769 & ~x204 ;
  assign n1773 = ~n1771 & ~n1772 ;
  assign n1774 = x82 & ~n413 ;
  assign n1775 = n391 & n1089 ;
  assign n1776 = x82 & ~n1775 ;
  assign n1777 = n385 & ~n1776 ;
  assign n1778 = ~n1774 & ~n1777 ;
  assign n1779 = ~x43 & ~n1778 ;
  assign n1780 = ~x47 & n413 ;
  assign n1781 = n1598 & n1780 ;
  assign n1782 = x82 & ~n1781 ;
  assign n1783 = ~n385 & ~n1782 ;
  assign n1784 = x77 & n1783 ;
  assign n1785 = x43 & n968 ;
  assign n1786 = n1605 & n1785 ;
  assign n1787 = n395 & n1786 ;
  assign n1788 = ~x129 & ~n1787 ;
  assign n1789 = ~n1784 & n1788 ;
  assign n1790 = ~n1779 & n1789 ;
  assign n1809 = n1790 & x205 ;
  assign n1791 = ~x82 & ~n450 ;
  assign n1792 = n428 & n1114 ;
  assign n1793 = ~x82 & ~n1792 ;
  assign n1794 = n422 & ~n1793 ;
  assign n1795 = ~n1791 & ~n1794 ;
  assign n1796 = x43 & ~n1795 ;
  assign n1797 = x47 & n450 ;
  assign n1798 = n1621 & n1797 ;
  assign n1799 = ~x82 & ~n1798 ;
  assign n1800 = ~n422 & ~n1799 ;
  assign n1801 = ~x77 & n1800 ;
  assign n1802 = ~x43 & n992 ;
  assign n1803 = n1628 & n1802 ;
  assign n1804 = n432 & n1803 ;
  assign n1805 = x129 & ~n1804 ;
  assign n1806 = ~n1801 & n1805 ;
  assign n1807 = ~n1796 & n1806 ;
  assign n1810 = ~n1807 & ~x205 ;
  assign n1811 = ~n1809 & ~n1810 ;
  assign n1812 = n965 & n969 ;
  assign n1813 = n1598 & n1812 ;
  assign n1814 = x82 & ~n1813 ;
  assign n1815 = x67 & ~n385 ;
  assign n1816 = ~x44 & n385 ;
  assign n1817 = ~n1815 & ~n1816 ;
  assign n1818 = ~n1814 & ~n1817 ;
  assign n1819 = ~x129 & ~n1736 ;
  assign n1820 = ~n1818 & n1819 ;
  assign n1831 = n1820 & x206 ;
  assign n1821 = n989 & n993 ;
  assign n1822 = n1621 & n1821 ;
  assign n1823 = ~x82 & ~n1822 ;
  assign n1824 = ~x67 & ~n422 ;
  assign n1825 = x44 & n422 ;
  assign n1826 = ~n1824 & ~n1825 ;
  assign n1827 = ~n1823 & ~n1826 ;
  assign n1828 = x129 & ~n1753 ;
  assign n1829 = ~n1827 & n1828 ;
  assign n1832 = ~n1829 & ~x206 ;
  assign n1833 = ~n1831 & ~n1832 ;
  assign n1834 = n405 & n1095 ;
  assign n1835 = n394 & n397 ;
  assign n1836 = n1834 & n1835 ;
  assign n1837 = x82 & ~n1836 ;
  assign n1838 = ~x24 & n1083 ;
  assign n1839 = x82 & ~n1838 ;
  assign n1840 = n385 & ~n1839 ;
  assign n1841 = ~n1837 & ~n1840 ;
  assign n1842 = ~x45 & ~n1841 ;
  assign n1843 = ~x2 & n405 ;
  assign n1844 = n391 & n1843 ;
  assign n1845 = n414 & n1844 ;
  assign n1846 = x82 & ~n1845 ;
  assign n1847 = ~n385 & ~n1846 ;
  assign n1848 = x68 & n1847 ;
  assign n1849 = ~x38 & n968 ;
  assign n1850 = x45 & n1849 ;
  assign n1851 = n1605 & n1850 ;
  assign n1852 = n1589 & n1851 ;
  assign n1853 = ~x129 & ~n1852 ;
  assign n1854 = ~n1848 & n1853 ;
  assign n1855 = ~n1842 & n1854 ;
  assign n1879 = n1855 & x207 ;
  assign n1856 = n442 & n1120 ;
  assign n1857 = n431 & n434 ;
  assign n1858 = n1856 & n1857 ;
  assign n1859 = ~x82 & ~n1858 ;
  assign n1860 = x24 & n1108 ;
  assign n1861 = ~x82 & ~n1860 ;
  assign n1862 = n422 & ~n1861 ;
  assign n1863 = ~n1859 & ~n1862 ;
  assign n1864 = x45 & ~n1863 ;
  assign n1865 = x2 & n442 ;
  assign n1866 = n428 & n1865 ;
  assign n1867 = n451 & n1866 ;
  assign n1868 = ~x82 & ~n1867 ;
  assign n1869 = ~n422 & ~n1868 ;
  assign n1870 = ~x68 & n1869 ;
  assign n1871 = x38 & n992 ;
  assign n1872 = ~x45 & n1871 ;
  assign n1873 = n1628 & n1872 ;
  assign n1874 = n1612 & n1873 ;
  assign n1875 = x129 & ~n1874 ;
  assign n1876 = ~n1870 & n1875 ;
  assign n1877 = ~n1864 & n1876 ;
  assign n1880 = ~n1877 & ~x207 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = x82 & ~n1835 ;
  assign n1883 = n1079 & n1598 ;
  assign n1884 = x82 & ~n1883 ;
  assign n1885 = n385 & ~n1884 ;
  assign n1886 = ~n1882 & ~n1885 ;
  assign n1887 = ~x46 & ~n1886 ;
  assign n1888 = ~x50 & n410 ;
  assign n1889 = n1883 & n1888 ;
  assign n1890 = x82 & ~n1889 ;
  assign n1891 = ~n385 & ~n1890 ;
  assign n1892 = x75 & n1891 ;
  assign n1893 = x46 & x82 ;
  assign n1894 = n1888 & n1893 ;
  assign n1895 = ~x129 & ~n1894 ;
  assign n1896 = ~n1892 & n1895 ;
  assign n1897 = ~n1887 & n1896 ;
  assign n1915 = n1897 & x208 ;
  assign n1898 = ~x82 & ~n1857 ;
  assign n1899 = n1104 & n1621 ;
  assign n1900 = ~x82 & ~n1899 ;
  assign n1901 = n422 & ~n1900 ;
  assign n1902 = ~n1898 & ~n1901 ;
  assign n1903 = x46 & ~n1902 ;
  assign n1904 = x50 & n447 ;
  assign n1905 = n1899 & n1904 ;
  assign n1906 = ~x82 & ~n1905 ;
  assign n1907 = ~n422 & ~n1906 ;
  assign n1908 = ~x75 & n1907 ;
  assign n1909 = ~x46 & ~x82 ;
  assign n1910 = n1904 & n1909 ;
  assign n1911 = x129 & ~n1910 ;
  assign n1912 = ~n1908 & n1911 ;
  assign n1913 = ~n1903 & n1912 ;
  assign n1916 = ~n1913 & ~x208 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = x82 & ~n414 ;
  assign n1919 = x82 & ~n1598 ;
  assign n1920 = n385 & ~n1919 ;
  assign n1921 = ~n1918 & ~n1920 ;
  assign n1922 = ~x47 & ~n1921 ;
  assign n1923 = n414 & n1598 ;
  assign n1924 = x82 & ~n1923 ;
  assign n1925 = ~n385 & ~n1924 ;
  assign n1926 = x64 & n1925 ;
  assign n1927 = n809 & n813 ;
  assign n1928 = x47 & n968 ;
  assign n1929 = n1605 & n1928 ;
  assign n1930 = n1927 & n1929 ;
  assign n1931 = ~x129 & ~n1930 ;
  assign n1932 = ~n1926 & n1931 ;
  assign n1933 = ~n1922 & n1932 ;
  assign n1951 = n1933 & x209 ;
  assign n1934 = ~x82 & ~n451 ;
  assign n1935 = ~x82 & ~n1621 ;
  assign n1936 = n422 & ~n1935 ;
  assign n1937 = ~n1934 & ~n1936 ;
  assign n1938 = x47 & ~n1937 ;
  assign n1939 = n451 & n1621 ;
  assign n1940 = ~x82 & ~n1939 ;
  assign n1941 = ~n422 & ~n1940 ;
  assign n1942 = ~x64 & n1941 ;
  assign n1943 = n836 & n840 ;
  assign n1944 = ~x47 & n992 ;
  assign n1945 = n1628 & n1944 ;
  assign n1946 = n1943 & n1945 ;
  assign n1947 = x129 & ~n1946 ;
  assign n1948 = ~n1942 & n1947 ;
  assign n1949 = ~n1938 & n1948 ;
  assign n1952 = ~n1949 & ~x209 ;
  assign n1953 = ~n1951 & ~n1952 ;
  assign n1954 = n965 & n1835 ;
  assign n1955 = x82 & ~n1954 ;
  assign n1956 = x82 & ~n1590 ;
  assign n1957 = n385 & ~n1956 ;
  assign n1958 = ~n1955 & ~n1957 ;
  assign n1959 = ~x48 & ~n1958 ;
  assign n1960 = ~x2 & ~x47 ;
  assign n1961 = n404 & n407 ;
  assign n1962 = n1960 & n1961 ;
  assign n1963 = n414 & n1962 ;
  assign n1964 = x82 & ~n1963 ;
  assign n1965 = ~n385 & ~n1964 ;
  assign n1966 = x62 & n1965 ;
  assign n1967 = n387 & n412 ;
  assign n1968 = x48 & n1849 ;
  assign n1969 = n1605 & n1968 ;
  assign n1970 = n1967 & n1969 ;
  assign n1971 = ~x129 & ~n1970 ;
  assign n1972 = ~n1966 & n1971 ;
  assign n1973 = ~n1959 & n1972 ;
  assign n1995 = n1973 & x210 ;
  assign n1974 = n989 & n1857 ;
  assign n1975 = ~x82 & ~n1974 ;
  assign n1976 = ~x82 & ~n1613 ;
  assign n1977 = n422 & ~n1976 ;
  assign n1978 = ~n1975 & ~n1977 ;
  assign n1979 = x48 & ~n1978 ;
  assign n1980 = x2 & x47 ;
  assign n1981 = n441 & n444 ;
  assign n1982 = n1980 & n1981 ;
  assign n1983 = n451 & n1982 ;
  assign n1984 = ~x82 & ~n1983 ;
  assign n1985 = ~n422 & ~n1984 ;
  assign n1986 = ~x62 & n1985 ;
  assign n1987 = n424 & n449 ;
  assign n1988 = ~x48 & n1871 ;
  assign n1989 = n1628 & n1988 ;
  assign n1990 = n1987 & n1989 ;
  assign n1991 = x129 & ~n1990 ;
  assign n1992 = ~n1986 & n1991 ;
  assign n1993 = ~n1979 & n1992 ;
  assign n1996 = ~n1993 & ~x210 ;
  assign n1997 = ~n1995 & ~n1996 ;
  assign n1998 = n390 & n1888 ;
  assign n1999 = n1096 & n1998 ;
  assign n2000 = x82 & ~n1999 ;
  assign n2001 = ~n385 & ~n2000 ;
  assign n2002 = ~x69 & n2001 ;
  assign n2003 = ~x24 & ~x42 ;
  assign n2004 = n1743 & n2003 ;
  assign n2005 = n1096 & n2004 ;
  assign n2006 = x49 & ~n2005 ;
  assign n2007 = ~x2 & n389 ;
  assign n2008 = n1998 & ~n2007 ;
  assign n2009 = n965 & n2008 ;
  assign n2010 = n386 & n2009 ;
  assign n2011 = ~n2006 & ~n2010 ;
  assign n2012 = x82 & ~n2011 ;
  assign n2013 = x49 & n417 ;
  assign n2014 = ~n2012 & ~n2013 ;
  assign n2015 = ~n2002 & n2014 ;
  assign n2016 = ~x129 & ~n2015 ;
  assign n2037 = n2016 & x211 ;
  assign n2017 = n427 & n1904 ;
  assign n2018 = n1121 & n2017 ;
  assign n2019 = ~x82 & ~n2018 ;
  assign n2020 = ~n422 & ~n2019 ;
  assign n2021 = x69 & n2020 ;
  assign n2022 = x24 & x42 ;
  assign n2023 = n1760 & n2022 ;
  assign n2024 = n1121 & n2023 ;
  assign n2025 = ~x49 & ~n2024 ;
  assign n2026 = x2 & n426 ;
  assign n2027 = n2017 & ~n2026 ;
  assign n2028 = n989 & n2027 ;
  assign n2029 = n423 & n2028 ;
  assign n2030 = ~n2025 & ~n2029 ;
  assign n2031 = ~x82 & ~n2030 ;
  assign n2032 = ~x49 & n454 ;
  assign n2033 = ~n2031 & ~n2032 ;
  assign n2034 = ~n2021 & n2033 ;
  assign n2035 = x129 & ~n2034 ;
  assign n2038 = ~n2035 & ~x211 ;
  assign n2039 = ~n2037 & ~n2038 ;
  assign n2040 = x82 & ~n410 ;
  assign n2041 = n1095 & n1843 ;
  assign n2042 = n1961 & n2041 ;
  assign n2043 = x82 & ~n2042 ;
  assign n2044 = n385 & ~n2043 ;
  assign n2045 = ~n2040 & ~n2044 ;
  assign n2046 = ~x50 & ~n2045 ;
  assign n2047 = n410 & n965 ;
  assign n2048 = n1598 & n2047 ;
  assign n2049 = x82 & ~n2048 ;
  assign n2050 = ~n385 & ~n2049 ;
  assign n2051 = x66 & n2050 ;
  assign n2052 = x50 & n1849 ;
  assign n2053 = n1605 & n2052 ;
  assign n2054 = ~x129 & ~n2053 ;
  assign n2055 = ~n2051 & n2054 ;
  assign n2056 = ~n2046 & n2055 ;
  assign n2075 = n2056 & x212 ;
  assign n2057 = ~x82 & ~n447 ;
  assign n2058 = n1120 & n1865 ;
  assign n2059 = n1981 & n2058 ;
  assign n2060 = ~x82 & ~n2059 ;
  assign n2061 = n422 & ~n2060 ;
  assign n2062 = ~n2057 & ~n2061 ;
  assign n2063 = x50 & ~n2062 ;
  assign n2064 = n447 & n989 ;
  assign n2065 = n1621 & n2064 ;
  assign n2066 = ~x82 & ~n2065 ;
  assign n2067 = ~n422 & ~n2066 ;
  assign n2068 = ~x66 & n2067 ;
  assign n2069 = ~x50 & n1871 ;
  assign n2070 = n1628 & n2069 ;
  assign n2071 = x129 & ~n2070 ;
  assign n2072 = ~n2068 & n2071 ;
  assign n2073 = ~n2063 & n2072 ;
  assign n2076 = ~n2073 & ~x212 ;
  assign n2077 = ~n2075 & ~n2076 ;
  assign n2078 = ~n1638 & ~n1645 ;
  assign n2079 = ~x106 & n2078 ;
  assign n2080 = ~x129 & ~n2079 ;
  assign n2084 = n2080 & x213 ;
  assign n2081 = x106 & n2078 ;
  assign n2082 = x129 & ~n2081 ;
  assign n2085 = ~n2082 & ~x213 ;
  assign n2086 = ~n2084 & ~n2085 ;
  assign n2087 = x52 & ~n1638 ;
  assign n2088 = ~x106 & ~n1641 ;
  assign n2089 = ~n2087 & n2088 ;
  assign n2090 = ~x129 & ~n2089 ;
  assign n2096 = n2090 & x214 ;
  assign n2091 = ~x52 & ~n1645 ;
  assign n2092 = x106 & ~n1648 ;
  assign n2093 = ~n2091 & n2092 ;
  assign n2094 = x129 & ~n2093 ;
  assign n2097 = ~n2094 & ~x214 ;
  assign n2098 = ~n2096 & ~n2097 ;
  assign n2099 = x58 & x116 ;
  assign n2100 = ~x58 & ~x110 ;
  assign n2101 = ~x96 & n2100 ;
  assign n2102 = n1144 & n2101 ;
  assign n2103 = ~n2099 & ~n2102 ;
  assign n2104 = ~x53 & ~n2103 ;
  assign n2105 = x97 & n2104 ;
  assign n2106 = ~x116 & n1223 ;
  assign n2107 = ~n2105 & ~n2106 ;
  assign n2108 = ~x129 & ~n2107 ;
  assign n2109 = ~x3 & n2108 ;
  assign n2110 = n1174 & n2109 ;
  assign n2111 = ~x26 & n2110 ;
  assign n2126 = n2111 & x215 ;
  assign n2112 = ~x58 & ~x116 ;
  assign n2113 = x58 & x110 ;
  assign n2114 = x96 & n2113 ;
  assign n2115 = n1192 & n2114 ;
  assign n2116 = ~n2112 & ~n2115 ;
  assign n2117 = x53 & ~n2116 ;
  assign n2118 = ~x97 & n2117 ;
  assign n2119 = x116 & n1175 ;
  assign n2120 = ~n2118 & ~n2119 ;
  assign n2121 = x129 & ~n2120 ;
  assign n2122 = x3 & n2121 ;
  assign n2123 = n1222 & n2122 ;
  assign n2124 = x26 & n2123 ;
  assign n2127 = ~n2124 & ~x215 ;
  assign n2128 = ~n2126 & ~n2127 ;
  assign n2129 = n414 & n1775 ;
  assign n2130 = x82 & ~n2129 ;
  assign n2131 = ~n385 & ~n2130 ;
  assign n2132 = ~x129 & ~n2131 ;
  assign n2138 = ~n2132 & x216 ;
  assign n2133 = n451 & n1792 ;
  assign n2134 = ~x82 & ~n2133 ;
  assign n2135 = ~n422 & ~n2134 ;
  assign n2136 = x129 & ~n2135 ;
  assign n2139 = n2136 & ~x216 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = ~x123 & ~x129 ;
  assign n2142 = x114 & ~x122 ;
  assign n2143 = n2141 & n2142 ;
  assign n2148 = n2143 & x217 ;
  assign n2144 = x123 & x129 ;
  assign n2145 = ~x114 & x122 ;
  assign n2146 = n2144 & n2145 ;
  assign n2149 = ~n2146 & ~x217 ;
  assign n2150 = ~n2148 & ~n2149 ;
  assign n2151 = ~x26 & x58 ;
  assign n2152 = x26 & ~x58 ;
  assign n2153 = x116 & n2152 ;
  assign n2154 = ~n2151 & ~n2153 ;
  assign n2155 = x94 & ~n2154 ;
  assign n2156 = x58 & ~x116 ;
  assign n2157 = x37 & ~x116 ;
  assign n2158 = ~n2151 & ~n2157 ;
  assign n2159 = ~n2156 & ~n2158 ;
  assign n2160 = ~n2155 & ~n2159 ;
  assign n2161 = ~x53 & ~n2160 ;
  assign n2162 = ~x26 & x37 ;
  assign n2163 = ~x58 & n2162 ;
  assign n2164 = ~n2161 & ~n2163 ;
  assign n2165 = ~x85 & ~n2164 ;
  assign n2166 = n1278 & n2162 ;
  assign n2167 = ~n2165 & ~n2166 ;
  assign n2168 = ~x27 & ~n2167 ;
  assign n2169 = ~x85 & n1278 ;
  assign n2170 = n2162 & n2169 ;
  assign n2171 = ~n2168 & ~n2170 ;
  assign n2172 = ~x129 & ~n2171 ;
  assign n2173 = ~x3 & n2172 ;
  assign n2196 = n2173 & x218 ;
  assign n2174 = ~x116 & n2151 ;
  assign n2175 = ~n2152 & ~n2174 ;
  assign n2176 = ~x94 & ~n2175 ;
  assign n2177 = ~x58 & x116 ;
  assign n2178 = ~x37 & x116 ;
  assign n2179 = ~n2152 & ~n2178 ;
  assign n2180 = ~n2177 & ~n2179 ;
  assign n2181 = ~n2176 & ~n2180 ;
  assign n2182 = x53 & ~n2181 ;
  assign n2183 = x26 & ~x37 ;
  assign n2184 = x58 & n2183 ;
  assign n2185 = ~n2182 & ~n2184 ;
  assign n2186 = x85 & ~n2185 ;
  assign n2187 = n1292 & n2183 ;
  assign n2188 = ~n2186 & ~n2187 ;
  assign n2189 = x27 & ~n2188 ;
  assign n2190 = x85 & n1292 ;
  assign n2191 = n2183 & n2190 ;
  assign n2192 = ~n2189 & ~n2191 ;
  assign n2193 = x129 & ~n2192 ;
  assign n2194 = x3 & n2193 ;
  assign n2197 = ~n2194 & ~x218 ;
  assign n2198 = ~n2196 & ~n2197 ;
  assign n2199 = ~x26 & ~x53 ;
  assign n2200 = x26 & x53 ;
  assign n2201 = ~x85 & ~n2200 ;
  assign n2202 = ~n2199 & ~n2201 ;
  assign n2203 = ~x58 & ~n2202 ;
  assign n2204 = ~x85 & n2199 ;
  assign n2205 = ~x116 & n2204 ;
  assign n2206 = ~n2203 & ~n2205 ;
  assign n2207 = x57 & ~n2206 ;
  assign n2208 = x60 & n2099 ;
  assign n2209 = n2204 & n2208 ;
  assign n2210 = ~n2207 & ~n2209 ;
  assign n2211 = ~x27 & ~n2210 ;
  assign n2212 = x57 & ~x58 ;
  assign n2213 = n2204 & n2212 ;
  assign n2214 = ~n2211 & ~n2213 ;
  assign n2215 = ~x129 & ~n2214 ;
  assign n2216 = ~x3 & n2215 ;
  assign n2234 = n2216 & x219 ;
  assign n2217 = x85 & ~n2199 ;
  assign n2218 = ~n2200 & ~n2217 ;
  assign n2219 = x58 & ~n2218 ;
  assign n2220 = x85 & n2200 ;
  assign n2221 = x116 & n2220 ;
  assign n2222 = ~n2219 & ~n2221 ;
  assign n2223 = ~x57 & ~n2222 ;
  assign n2224 = ~x60 & n2112 ;
  assign n2225 = n2220 & n2224 ;
  assign n2226 = ~n2223 & ~n2225 ;
  assign n2227 = x27 & ~n2226 ;
  assign n2228 = ~x57 & x58 ;
  assign n2229 = n2220 & n2228 ;
  assign n2230 = ~n2227 & ~n2229 ;
  assign n2231 = x129 & ~n2230 ;
  assign n2232 = x3 & n2231 ;
  assign n2235 = ~n2232 & ~x219 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = n1323 & n2156 ;
  assign n2238 = ~x58 & n1342 ;
  assign n2239 = n1157 & n2238 ;
  assign n2240 = ~n2237 & ~n2239 ;
  assign n2241 = ~x129 & ~n2240 ;
  assign n2242 = ~x3 & n2241 ;
  assign n2243 = ~x53 & n2242 ;
  assign n2244 = ~x85 & n2243 ;
  assign n2254 = n2244 & x220 ;
  assign n2245 = n1359 & n2177 ;
  assign n2246 = x58 & n1306 ;
  assign n2247 = n1205 & n2246 ;
  assign n2248 = ~n2245 & ~n2247 ;
  assign n2249 = x129 & ~n2248 ;
  assign n2250 = x3 & n2249 ;
  assign n2251 = x53 & n2250 ;
  assign n2252 = x85 & n2251 ;
  assign n2255 = ~n2252 & ~x220 ;
  assign n2256 = ~n2254 & ~n2255 ;
  assign n2257 = ~n1175 & ~n1223 ;
  assign n2258 = ~x116 & ~n2257 ;
  assign n2259 = ~n1146 & n1278 ;
  assign n2260 = ~n2258 & ~n2259 ;
  assign n2261 = x59 & ~n2260 ;
  assign n2262 = n1146 & n1278 ;
  assign n2263 = x96 & n2262 ;
  assign n2264 = ~n2261 & ~n2263 ;
  assign n2265 = ~x85 & ~n2264 ;
  assign n2266 = x59 & ~x116 ;
  assign n2267 = x85 & n1278 ;
  assign n2268 = n2266 & n2267 ;
  assign n2269 = ~n2265 & ~n2268 ;
  assign n2270 = ~x27 & ~n2269 ;
  assign n2271 = x27 & n2169 ;
  assign n2272 = n2266 & n2271 ;
  assign n2273 = ~n2270 & ~n2272 ;
  assign n2274 = ~x26 & ~n2273 ;
  assign n2275 = n1404 & n2266 ;
  assign n2276 = ~n2274 & ~n2275 ;
  assign n2277 = ~x129 & ~n2276 ;
  assign n2278 = ~x3 & n2277 ;
  assign n2301 = n2278 & x221 ;
  assign n2279 = x116 & ~n2257 ;
  assign n2280 = ~n1194 & n1292 ;
  assign n2281 = ~n2279 & ~n2280 ;
  assign n2282 = ~x59 & ~n2281 ;
  assign n2283 = n1194 & n1292 ;
  assign n2284 = ~x96 & n2283 ;
  assign n2285 = ~n2282 & ~n2284 ;
  assign n2286 = x85 & ~n2285 ;
  assign n2287 = ~x59 & x116 ;
  assign n2288 = ~x85 & n1292 ;
  assign n2289 = n2287 & n2288 ;
  assign n2290 = ~n2286 & ~n2289 ;
  assign n2291 = x27 & ~n2290 ;
  assign n2292 = ~x27 & n2190 ;
  assign n2293 = n2287 & n2292 ;
  assign n2294 = ~n2291 & ~n2293 ;
  assign n2295 = x26 & ~n2294 ;
  assign n2296 = n1435 & n2287 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2298 = x129 & ~n2297 ;
  assign n2299 = x3 & n2298 ;
  assign n2302 = ~n2299 & ~x221 ;
  assign n2303 = ~n2301 & ~n2302 ;
  assign n2304 = ~x117 & ~x122 ;
  assign n2305 = x60 & ~n2304 ;
  assign n2306 = x123 & n2304 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2313 = ~n2307 & x222 ;
  assign n2308 = x117 & x122 ;
  assign n2309 = ~x60 & ~n2308 ;
  assign n2310 = ~x123 & n2308 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2314 = n2311 & ~x222 ;
  assign n2315 = ~n2313 & ~n2314 ;
  assign n2316 = ~x114 & x123 ;
  assign n2317 = ~x122 & n2316 ;
  assign n2318 = ~x129 & n2317 ;
  assign n2323 = n2318 & x223 ;
  assign n2319 = x114 & ~x123 ;
  assign n2320 = x122 & n2319 ;
  assign n2321 = x129 & n2320 ;
  assign n2324 = ~n2321 & ~x223 ;
  assign n2325 = ~n2323 & ~n2324 ;
  assign n2326 = ~x137 & ~x138 ;
  assign n2327 = x136 & n2326 ;
  assign n2328 = x132 & x133 ;
  assign n2329 = x131 & n2328 ;
  assign n2330 = n2327 & n2329 ;
  assign n2331 = x62 & ~n2330 ;
  assign n2332 = x136 & ~x137 ;
  assign n2333 = ~x140 & n2332 ;
  assign n2334 = ~x138 & n2329 ;
  assign n2335 = n2333 & n2334 ;
  assign n2336 = ~n2331 & ~n2335 ;
  assign n2337 = ~x129 & ~n2336 ;
  assign n2351 = ~n2337 & x224 ;
  assign n2338 = x137 & x138 ;
  assign n2339 = ~x136 & n2338 ;
  assign n2340 = ~x132 & ~x133 ;
  assign n2341 = ~x131 & n2340 ;
  assign n2342 = n2339 & n2341 ;
  assign n2343 = ~x62 & ~n2342 ;
  assign n2344 = ~x136 & x137 ;
  assign n2345 = x140 & n2344 ;
  assign n2346 = x138 & n2341 ;
  assign n2347 = n2345 & n2346 ;
  assign n2348 = ~n2343 & ~n2347 ;
  assign n2349 = x129 & ~n2348 ;
  assign n2352 = n2349 & ~x224 ;
  assign n2353 = ~n2351 & ~n2352 ;
  assign n2354 = x63 & ~n2330 ;
  assign n2355 = ~x142 & n2332 ;
  assign n2356 = n2334 & n2355 ;
  assign n2357 = ~n2354 & ~n2356 ;
  assign n2358 = ~x129 & ~n2357 ;
  assign n2365 = ~n2358 & x225 ;
  assign n2359 = ~x63 & ~n2342 ;
  assign n2360 = x142 & n2344 ;
  assign n2361 = n2346 & n2360 ;
  assign n2362 = ~n2359 & ~n2361 ;
  assign n2363 = x129 & ~n2362 ;
  assign n2366 = n2363 & ~x225 ;
  assign n2367 = ~n2365 & ~n2366 ;
  assign n2368 = x64 & ~n2330 ;
  assign n2369 = ~x139 & n2332 ;
  assign n2370 = n2334 & n2369 ;
  assign n2371 = ~n2368 & ~n2370 ;
  assign n2372 = ~x129 & ~n2371 ;
  assign n2379 = ~n2372 & x226 ;
  assign n2373 = ~x64 & ~n2342 ;
  assign n2374 = x139 & n2344 ;
  assign n2375 = n2346 & n2374 ;
  assign n2376 = ~n2373 & ~n2375 ;
  assign n2377 = x129 & ~n2376 ;
  assign n2380 = n2377 & ~x226 ;
  assign n2381 = ~n2379 & ~n2380 ;
  assign n2382 = x65 & ~n2330 ;
  assign n2383 = ~x146 & n2332 ;
  assign n2384 = n2334 & n2383 ;
  assign n2385 = ~n2382 & ~n2384 ;
  assign n2386 = ~x129 & ~n2385 ;
  assign n2393 = ~n2386 & x227 ;
  assign n2387 = ~x65 & ~n2342 ;
  assign n2388 = x146 & n2344 ;
  assign n2389 = n2346 & n2388 ;
  assign n2390 = ~n2387 & ~n2389 ;
  assign n2391 = x129 & ~n2390 ;
  assign n2394 = n2391 & ~x227 ;
  assign n2395 = ~n2393 & ~n2394 ;
  assign n2396 = ~x136 & ~x137 ;
  assign n2397 = n2334 & n2396 ;
  assign n2398 = x66 & ~n2397 ;
  assign n2399 = ~x143 & n2397 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = ~x129 & ~n2400 ;
  assign n2409 = ~n2401 & x228 ;
  assign n2402 = x136 & x137 ;
  assign n2403 = n2346 & n2402 ;
  assign n2404 = ~x66 & ~n2403 ;
  assign n2405 = x143 & n2403 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = x129 & ~n2406 ;
  assign n2410 = n2407 & ~x228 ;
  assign n2411 = ~n2409 & ~n2410 ;
  assign n2412 = x67 & ~n2397 ;
  assign n2413 = ~x139 & n2397 ;
  assign n2414 = ~n2412 & ~n2413 ;
  assign n2415 = ~x129 & ~n2414 ;
  assign n2421 = ~n2415 & x229 ;
  assign n2416 = ~x67 & ~n2403 ;
  assign n2417 = x139 & n2403 ;
  assign n2418 = ~n2416 & ~n2417 ;
  assign n2419 = x129 & ~n2418 ;
  assign n2422 = n2419 & ~x229 ;
  assign n2423 = ~n2421 & ~n2422 ;
  assign n2424 = x68 & ~n2330 ;
  assign n2425 = ~x141 & n2332 ;
  assign n2426 = n2334 & n2425 ;
  assign n2427 = ~n2424 & ~n2426 ;
  assign n2428 = ~x129 & ~n2427 ;
  assign n2435 = ~n2428 & x230 ;
  assign n2429 = ~x68 & ~n2342 ;
  assign n2430 = x141 & n2344 ;
  assign n2431 = n2346 & n2430 ;
  assign n2432 = ~n2429 & ~n2431 ;
  assign n2433 = x129 & ~n2432 ;
  assign n2436 = n2433 & ~x230 ;
  assign n2437 = ~n2435 & ~n2436 ;
  assign n2438 = x69 & ~n2330 ;
  assign n2439 = ~x143 & n2332 ;
  assign n2440 = n2334 & n2439 ;
  assign n2441 = ~n2438 & ~n2440 ;
  assign n2442 = ~x129 & ~n2441 ;
  assign n2449 = ~n2442 & x231 ;
  assign n2443 = ~x69 & ~n2342 ;
  assign n2444 = x143 & n2344 ;
  assign n2445 = n2346 & n2444 ;
  assign n2446 = ~n2443 & ~n2445 ;
  assign n2447 = x129 & ~n2446 ;
  assign n2450 = n2447 & ~x231 ;
  assign n2451 = ~n2449 & ~n2450 ;
  assign n2452 = x70 & ~n2330 ;
  assign n2453 = ~x144 & n2332 ;
  assign n2454 = n2334 & n2453 ;
  assign n2455 = ~n2452 & ~n2454 ;
  assign n2456 = ~x129 & ~n2455 ;
  assign n2463 = ~n2456 & x232 ;
  assign n2457 = ~x70 & ~n2342 ;
  assign n2458 = x144 & n2344 ;
  assign n2459 = n2346 & n2458 ;
  assign n2460 = ~n2457 & ~n2459 ;
  assign n2461 = x129 & ~n2460 ;
  assign n2464 = n2461 & ~x232 ;
  assign n2465 = ~n2463 & ~n2464 ;
  assign n2466 = x71 & ~n2330 ;
  assign n2467 = ~x145 & n2332 ;
  assign n2468 = n2334 & n2467 ;
  assign n2469 = ~n2466 & ~n2468 ;
  assign n2470 = ~x129 & ~n2469 ;
  assign n2477 = ~n2470 & x233 ;
  assign n2471 = ~x71 & ~n2342 ;
  assign n2472 = x145 & n2344 ;
  assign n2473 = n2346 & n2472 ;
  assign n2474 = ~n2471 & ~n2473 ;
  assign n2475 = x129 & ~n2474 ;
  assign n2478 = n2475 & ~x233 ;
  assign n2479 = ~n2477 & ~n2478 ;
  assign n2480 = x72 & ~n2397 ;
  assign n2481 = ~x140 & n2397 ;
  assign n2482 = ~n2480 & ~n2481 ;
  assign n2483 = ~x129 & ~n2482 ;
  assign n2489 = ~n2483 & x234 ;
  assign n2484 = ~x72 & ~n2403 ;
  assign n2485 = x140 & n2403 ;
  assign n2486 = ~n2484 & ~n2485 ;
  assign n2487 = x129 & ~n2486 ;
  assign n2490 = n2487 & ~x234 ;
  assign n2491 = ~n2489 & ~n2490 ;
  assign n2492 = x73 & ~n2397 ;
  assign n2493 = ~x141 & n2397 ;
  assign n2494 = ~n2492 & ~n2493 ;
  assign n2495 = ~x129 & ~n2494 ;
  assign n2501 = ~n2495 & x235 ;
  assign n2496 = ~x73 & ~n2403 ;
  assign n2497 = x141 & n2403 ;
  assign n2498 = ~n2496 & ~n2497 ;
  assign n2499 = x129 & ~n2498 ;
  assign n2502 = n2499 & ~x235 ;
  assign n2503 = ~n2501 & ~n2502 ;
  assign n2504 = x74 & ~n2397 ;
  assign n2505 = ~x142 & n2397 ;
  assign n2506 = ~n2504 & ~n2505 ;
  assign n2507 = ~x129 & ~n2506 ;
  assign n2513 = ~n2507 & x236 ;
  assign n2508 = ~x74 & ~n2403 ;
  assign n2509 = x142 & n2403 ;
  assign n2510 = ~n2508 & ~n2509 ;
  assign n2511 = x129 & ~n2510 ;
  assign n2514 = n2511 & ~x236 ;
  assign n2515 = ~n2513 & ~n2514 ;
  assign n2516 = x75 & ~n2397 ;
  assign n2517 = ~x144 & n2397 ;
  assign n2518 = ~n2516 & ~n2517 ;
  assign n2519 = ~x129 & ~n2518 ;
  assign n2525 = ~n2519 & x237 ;
  assign n2520 = ~x75 & ~n2403 ;
  assign n2521 = x144 & n2403 ;
  assign n2522 = ~n2520 & ~n2521 ;
  assign n2523 = x129 & ~n2522 ;
  assign n2526 = n2523 & ~x237 ;
  assign n2527 = ~n2525 & ~n2526 ;
  assign n2528 = x76 & ~n2397 ;
  assign n2529 = ~x145 & n2397 ;
  assign n2530 = ~n2528 & ~n2529 ;
  assign n2531 = ~x129 & ~n2530 ;
  assign n2537 = ~n2531 & x238 ;
  assign n2532 = ~x76 & ~n2403 ;
  assign n2533 = x145 & n2403 ;
  assign n2534 = ~n2532 & ~n2533 ;
  assign n2535 = x129 & ~n2534 ;
  assign n2538 = n2535 & ~x238 ;
  assign n2539 = ~n2537 & ~n2538 ;
  assign n2540 = x77 & ~n2397 ;
  assign n2541 = ~x146 & n2397 ;
  assign n2542 = ~n2540 & ~n2541 ;
  assign n2543 = ~x129 & ~n2542 ;
  assign n2549 = ~n2543 & x239 ;
  assign n2544 = ~x77 & ~n2403 ;
  assign n2545 = x146 & n2403 ;
  assign n2546 = ~n2544 & ~n2545 ;
  assign n2547 = x129 & ~n2546 ;
  assign n2550 = n2547 & ~x239 ;
  assign n2551 = ~n2549 & ~n2550 ;
  assign n2552 = n2334 & n2344 ;
  assign n2553 = x78 & ~n2552 ;
  assign n2554 = x142 & n2552 ;
  assign n2555 = ~n2553 & ~n2554 ;
  assign n2556 = ~x129 & ~n2555 ;
  assign n2563 = n2556 & x240 ;
  assign n2557 = n2332 & n2346 ;
  assign n2558 = ~x78 & ~n2557 ;
  assign n2559 = ~x142 & n2557 ;
  assign n2560 = ~n2558 & ~n2559 ;
  assign n2561 = x129 & ~n2560 ;
  assign n2564 = ~n2561 & ~x240 ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = x79 & ~n2552 ;
  assign n2567 = x143 & n2552 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = ~x129 & ~n2568 ;
  assign n2575 = n2569 & x241 ;
  assign n2570 = ~x79 & ~n2557 ;
  assign n2571 = ~x143 & n2557 ;
  assign n2572 = ~n2570 & ~n2571 ;
  assign n2573 = x129 & ~n2572 ;
  assign n2576 = ~n2573 & ~x241 ;
  assign n2577 = ~n2575 & ~n2576 ;
  assign n2578 = x80 & ~n2552 ;
  assign n2579 = x144 & n2552 ;
  assign n2580 = ~n2578 & ~n2579 ;
  assign n2581 = ~x129 & ~n2580 ;
  assign n2587 = n2581 & x242 ;
  assign n2582 = ~x80 & ~n2557 ;
  assign n2583 = ~x144 & n2557 ;
  assign n2584 = ~n2582 & ~n2583 ;
  assign n2585 = x129 & ~n2584 ;
  assign n2588 = ~n2585 & ~x242 ;
  assign n2589 = ~n2587 & ~n2588 ;
  assign n2590 = x81 & ~n2552 ;
  assign n2591 = x145 & n2552 ;
  assign n2592 = ~n2590 & ~n2591 ;
  assign n2593 = ~x129 & ~n2592 ;
  assign n2599 = n2593 & x243 ;
  assign n2594 = ~x81 & ~n2557 ;
  assign n2595 = ~x145 & n2557 ;
  assign n2596 = ~n2594 & ~n2595 ;
  assign n2597 = x129 & ~n2596 ;
  assign n2600 = ~n2597 & ~x243 ;
  assign n2601 = ~n2599 & ~n2600 ;
  assign n2602 = x82 & ~n2552 ;
  assign n2603 = x146 & n2552 ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = ~x129 & ~n2604 ;
  assign n2611 = n2605 & x244 ;
  assign n2606 = ~x82 & ~n2557 ;
  assign n2607 = ~x146 & n2557 ;
  assign n2608 = ~n2606 & ~n2607 ;
  assign n2609 = x129 & ~n2608 ;
  assign n2612 = ~n2609 & ~x244 ;
  assign n2613 = ~n2611 & ~n2612 ;
  assign n2614 = x89 & x138 ;
  assign n2615 = ~x62 & ~x138 ;
  assign n2616 = ~n2614 & ~n2615 ;
  assign n2617 = x136 & ~n2616 ;
  assign n2618 = x119 & x138 ;
  assign n2619 = ~x72 & ~x138 ;
  assign n2620 = ~n2618 & ~n2619 ;
  assign n2621 = ~x136 & ~n2620 ;
  assign n2622 = ~n2617 & ~n2621 ;
  assign n2623 = ~x137 & ~n2622 ;
  assign n2624 = ~x115 & x138 ;
  assign n2625 = x87 & ~x138 ;
  assign n2626 = ~n2624 & ~n2625 ;
  assign n2627 = ~x136 & ~n2626 ;
  assign n2628 = x136 & ~x138 ;
  assign n2629 = x31 & n2628 ;
  assign n2630 = ~n2627 & ~n2629 ;
  assign n2631 = x137 & ~n2630 ;
  assign n2632 = ~n2623 & ~n2631 ;
  assign n2653 = ~n2632 & x245 ;
  assign n2633 = ~x89 & ~x138 ;
  assign n2634 = x62 & x138 ;
  assign n2635 = ~n2633 & ~n2634 ;
  assign n2636 = ~x136 & ~n2635 ;
  assign n2637 = ~x119 & ~x138 ;
  assign n2638 = x72 & x138 ;
  assign n2639 = ~n2637 & ~n2638 ;
  assign n2640 = x136 & ~n2639 ;
  assign n2641 = ~n2636 & ~n2640 ;
  assign n2642 = x137 & ~n2641 ;
  assign n2643 = x115 & ~x138 ;
  assign n2644 = ~x87 & x138 ;
  assign n2645 = ~n2643 & ~n2644 ;
  assign n2646 = x136 & ~n2645 ;
  assign n2647 = ~x136 & x138 ;
  assign n2648 = ~x31 & n2647 ;
  assign n2649 = ~n2646 & ~n2648 ;
  assign n2650 = ~x137 & ~n2649 ;
  assign n2651 = ~n2642 & ~n2650 ;
  assign n2654 = n2651 & ~x245 ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = x84 & ~n2552 ;
  assign n2657 = x141 & n2552 ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = ~x129 & ~n2658 ;
  assign n2665 = n2659 & x246 ;
  assign n2660 = ~x84 & ~n2557 ;
  assign n2661 = ~x141 & n2557 ;
  assign n2662 = ~n2660 & ~n2661 ;
  assign n2663 = x129 & ~n2662 ;
  assign n2666 = ~n2663 & ~x246 ;
  assign n2667 = ~n2665 & ~n2666 ;
  assign n2668 = ~x85 & ~n1145 ;
  assign n2669 = ~x110 & n2668 ;
  assign n2670 = x96 & n2669 ;
  assign n2671 = ~n1233 & ~n2670 ;
  assign n2672 = ~x129 & ~n2671 ;
  assign n2673 = ~x3 & n2672 ;
  assign n2674 = n1246 & n2673 ;
  assign n2675 = ~x26 & n2674 ;
  assign n2685 = n2675 & x247 ;
  assign n2676 = x85 & ~n1193 ;
  assign n2677 = x110 & n2676 ;
  assign n2678 = ~x96 & n2677 ;
  assign n2679 = ~n1248 & ~n2678 ;
  assign n2680 = x129 & ~n2679 ;
  assign n2681 = x3 & n2680 ;
  assign n2682 = n1261 & n2681 ;
  assign n2683 = x26 & n2682 ;
  assign n2686 = ~n2683 & ~x247 ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = x86 & ~n2552 ;
  assign n2689 = x139 & n2552 ;
  assign n2690 = ~n2688 & ~n2689 ;
  assign n2691 = ~x129 & ~n2690 ;
  assign n2697 = n2691 & x248 ;
  assign n2692 = ~x86 & ~n2557 ;
  assign n2693 = ~x139 & n2557 ;
  assign n2694 = ~n2692 & ~n2693 ;
  assign n2695 = x129 & ~n2694 ;
  assign n2698 = ~n2695 & ~x248 ;
  assign n2699 = ~n2697 & ~n2698 ;
  assign n2700 = x87 & ~n2552 ;
  assign n2701 = x140 & n2552 ;
  assign n2702 = ~n2700 & ~n2701 ;
  assign n2703 = ~x129 & ~n2702 ;
  assign n2709 = n2703 & x249 ;
  assign n2704 = ~x87 & ~n2557 ;
  assign n2705 = ~x140 & n2557 ;
  assign n2706 = ~n2704 & ~n2705 ;
  assign n2707 = x129 & ~n2706 ;
  assign n2710 = ~n2707 & ~x249 ;
  assign n2711 = ~n2709 & ~n2710 ;
  assign n2712 = n2334 & n2402 ;
  assign n2713 = x88 & ~n2712 ;
  assign n2714 = x139 & n2712 ;
  assign n2715 = ~n2713 & ~n2714 ;
  assign n2716 = ~x129 & ~n2715 ;
  assign n2723 = n2716 & x250 ;
  assign n2717 = n2346 & n2396 ;
  assign n2718 = ~x88 & ~n2717 ;
  assign n2719 = ~x139 & n2717 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2721 = x129 & ~n2720 ;
  assign n2724 = ~n2721 & ~x250 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = x89 & ~n2712 ;
  assign n2727 = x140 & n2712 ;
  assign n2728 = ~n2726 & ~n2727 ;
  assign n2729 = ~x129 & ~n2728 ;
  assign n2735 = n2729 & x251 ;
  assign n2730 = ~x89 & ~n2717 ;
  assign n2731 = ~x140 & n2717 ;
  assign n2732 = ~n2730 & ~n2731 ;
  assign n2733 = x129 & ~n2732 ;
  assign n2736 = ~n2733 & ~x251 ;
  assign n2737 = ~n2735 & ~n2736 ;
  assign n2738 = x90 & ~n2712 ;
  assign n2739 = x142 & n2712 ;
  assign n2740 = ~n2738 & ~n2739 ;
  assign n2741 = ~x129 & ~n2740 ;
  assign n2747 = n2741 & x252 ;
  assign n2742 = ~x90 & ~n2717 ;
  assign n2743 = ~x142 & n2717 ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = x129 & ~n2744 ;
  assign n2748 = ~n2745 & ~x252 ;
  assign n2749 = ~n2747 & ~n2748 ;
  assign n2750 = x91 & ~n2712 ;
  assign n2751 = x143 & n2712 ;
  assign n2752 = ~n2750 & ~n2751 ;
  assign n2753 = ~x129 & ~n2752 ;
  assign n2759 = n2753 & x253 ;
  assign n2754 = ~x91 & ~n2717 ;
  assign n2755 = ~x143 & n2717 ;
  assign n2756 = ~n2754 & ~n2755 ;
  assign n2757 = x129 & ~n2756 ;
  assign n2760 = ~n2757 & ~x253 ;
  assign n2761 = ~n2759 & ~n2760 ;
  assign n2762 = x92 & ~n2712 ;
  assign n2763 = x144 & n2712 ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = ~x129 & ~n2764 ;
  assign n2771 = n2765 & x254 ;
  assign n2766 = ~x92 & ~n2717 ;
  assign n2767 = ~x144 & n2717 ;
  assign n2768 = ~n2766 & ~n2767 ;
  assign n2769 = x129 & ~n2768 ;
  assign n2772 = ~n2769 & ~x254 ;
  assign n2773 = ~n2771 & ~n2772 ;
  assign n2774 = x93 & ~n2712 ;
  assign n2775 = x146 & n2712 ;
  assign n2776 = ~n2774 & ~n2775 ;
  assign n2777 = ~x129 & ~n2776 ;
  assign n2783 = n2777 & x255 ;
  assign n2778 = ~x93 & ~n2717 ;
  assign n2779 = ~x146 & n2717 ;
  assign n2780 = ~n2778 & ~n2779 ;
  assign n2781 = x129 & ~n2780 ;
  assign n2784 = ~n2781 & ~x255 ;
  assign n2785 = ~n2783 & ~n2784 ;
  assign n2786 = x82 & ~x137 ;
  assign n2787 = ~x136 & n2786 ;
  assign n2788 = x138 & n2329 ;
  assign n2789 = n2787 & n2788 ;
  assign n2790 = x94 & ~n2789 ;
  assign n2791 = x142 & n2789 ;
  assign n2792 = ~n2790 & ~n2791 ;
  assign n2793 = ~x129 & ~n2792 ;
  assign n2803 = n2793 & x256 ;
  assign n2794 = ~x82 & x137 ;
  assign n2795 = x136 & n2794 ;
  assign n2796 = ~x138 & n2341 ;
  assign n2797 = n2795 & n2796 ;
  assign n2798 = ~x94 & ~n2797 ;
  assign n2799 = ~x142 & n2797 ;
  assign n2800 = ~n2798 & ~n2799 ;
  assign n2801 = x129 & ~n2800 ;
  assign n2804 = ~n2801 & ~x256 ;
  assign n2805 = ~n2803 & ~n2804 ;
  assign n2806 = ~x3 & ~n2329 ;
  assign n2807 = ~x110 & n2806 ;
  assign n2808 = x138 & n2787 ;
  assign n2809 = n2329 & ~n2808 ;
  assign n2810 = ~n2807 & ~n2809 ;
  assign n2811 = x95 & ~n2810 ;
  assign n2812 = x143 & n2789 ;
  assign n2813 = ~n2811 & ~n2812 ;
  assign n2814 = ~x129 & ~n2813 ;
  assign n2825 = n2814 & x257 ;
  assign n2815 = x3 & ~n2341 ;
  assign n2816 = x110 & n2815 ;
  assign n2817 = ~x138 & n2795 ;
  assign n2818 = n2341 & ~n2817 ;
  assign n2819 = ~n2816 & ~n2818 ;
  assign n2820 = ~x95 & ~n2819 ;
  assign n2821 = ~x143 & n2797 ;
  assign n2822 = ~n2820 & ~n2821 ;
  assign n2823 = x129 & ~n2822 ;
  assign n2826 = ~n2823 & ~x257 ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = x96 & ~n2810 ;
  assign n2829 = x146 & n2789 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = ~x129 & ~n2830 ;
  assign n2837 = n2831 & x258 ;
  assign n2832 = ~x96 & ~n2819 ;
  assign n2833 = ~x146 & n2797 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = x129 & ~n2834 ;
  assign n2838 = ~n2835 & ~x258 ;
  assign n2839 = ~n2837 & ~n2838 ;
  assign n2840 = x97 & ~n2810 ;
  assign n2841 = x145 & n2789 ;
  assign n2842 = ~n2840 & ~n2841 ;
  assign n2843 = ~x129 & ~n2842 ;
  assign n2849 = n2843 & x259 ;
  assign n2844 = ~x97 & ~n2819 ;
  assign n2845 = ~x145 & n2797 ;
  assign n2846 = ~n2844 & ~n2845 ;
  assign n2847 = x129 & ~n2846 ;
  assign n2850 = ~n2847 & ~x259 ;
  assign n2851 = ~n2849 & ~n2850 ;
  assign n2852 = x98 & ~n2712 ;
  assign n2853 = x145 & n2712 ;
  assign n2854 = ~n2852 & ~n2853 ;
  assign n2855 = ~x129 & ~n2854 ;
  assign n2861 = n2855 & x260 ;
  assign n2856 = ~x98 & ~n2717 ;
  assign n2857 = ~x145 & n2717 ;
  assign n2858 = ~n2856 & ~n2857 ;
  assign n2859 = x129 & ~n2858 ;
  assign n2862 = ~n2859 & ~x260 ;
  assign n2863 = ~n2861 & ~n2862 ;
  assign n2864 = x99 & ~n2712 ;
  assign n2865 = x141 & n2712 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = ~x129 & ~n2866 ;
  assign n2873 = n2867 & x261 ;
  assign n2868 = ~x99 & ~n2717 ;
  assign n2869 = ~x141 & n2717 ;
  assign n2870 = ~n2868 & ~n2869 ;
  assign n2871 = x129 & ~n2870 ;
  assign n2874 = ~n2871 & ~x261 ;
  assign n2875 = ~n2873 & ~n2874 ;
  assign n2876 = x100 & ~n2810 ;
  assign n2877 = x144 & n2789 ;
  assign n2878 = ~n2876 & ~n2877 ;
  assign n2879 = ~x129 & ~n2878 ;
  assign n2885 = n2879 & x262 ;
  assign n2880 = ~x100 & ~n2819 ;
  assign n2881 = ~x144 & n2797 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = x129 & ~n2882 ;
  assign n2886 = ~n2883 & ~x262 ;
  assign n2887 = ~n2885 & ~n2886 ;
  assign n2888 = x124 & x138 ;
  assign n2889 = ~x77 & ~x138 ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n2891 = ~x136 & ~n2890 ;
  assign n2892 = ~x65 & ~x138 ;
  assign n2893 = x93 & x138 ;
  assign n2894 = ~n2892 & ~n2893 ;
  assign n2895 = x136 & ~n2894 ;
  assign n2896 = ~n2891 & ~n2895 ;
  assign n2897 = ~x137 & ~n2896 ;
  assign n2898 = x37 & n2628 ;
  assign n2899 = x96 & x138 ;
  assign n2900 = x82 & ~x138 ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = ~x136 & ~n2901 ;
  assign n2903 = ~n2898 & ~n2902 ;
  assign n2904 = x137 & ~n2903 ;
  assign n2905 = ~n2897 & ~n2904 ;
  assign n2925 = ~n2905 & x263 ;
  assign n2906 = ~x124 & ~x138 ;
  assign n2907 = x77 & x138 ;
  assign n2908 = ~n2906 & ~n2907 ;
  assign n2909 = x136 & ~n2908 ;
  assign n2910 = x65 & x138 ;
  assign n2911 = ~x93 & ~x138 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = ~x136 & ~n2912 ;
  assign n2914 = ~n2909 & ~n2913 ;
  assign n2915 = x137 & ~n2914 ;
  assign n2916 = ~x37 & n2647 ;
  assign n2917 = ~x96 & ~x138 ;
  assign n2918 = ~x82 & x138 ;
  assign n2919 = ~n2917 & ~n2918 ;
  assign n2920 = x136 & ~n2919 ;
  assign n2921 = ~n2916 & ~n2920 ;
  assign n2922 = ~x137 & ~n2921 ;
  assign n2923 = ~n2915 & ~n2922 ;
  assign n2926 = n2923 & ~x263 ;
  assign n2927 = ~n2925 & ~n2926 ;
  assign n2928 = x91 & n2332 ;
  assign n2929 = x95 & n2344 ;
  assign n2930 = ~n2928 & ~n2929 ;
  assign n2931 = x138 & ~n2930 ;
  assign n2932 = x79 & ~x136 ;
  assign n2933 = x34 & x136 ;
  assign n2934 = ~n2932 & ~n2933 ;
  assign n2935 = x137 & ~n2934 ;
  assign n2936 = ~x69 & x136 ;
  assign n2937 = ~x66 & ~x136 ;
  assign n2938 = ~n2936 & ~n2937 ;
  assign n2939 = ~x137 & ~n2938 ;
  assign n2940 = ~n2935 & ~n2939 ;
  assign n2941 = ~x138 & ~n2940 ;
  assign n2942 = ~n2931 & ~n2941 ;
  assign n2959 = ~n2942 & x264 ;
  assign n2943 = ~x91 & n2344 ;
  assign n2944 = ~x95 & n2332 ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = ~x138 & ~n2945 ;
  assign n2947 = ~x79 & x136 ;
  assign n2948 = ~x34 & ~x136 ;
  assign n2949 = ~n2947 & ~n2948 ;
  assign n2950 = ~x137 & ~n2949 ;
  assign n2951 = x69 & ~x136 ;
  assign n2952 = x66 & x136 ;
  assign n2953 = ~n2951 & ~n2952 ;
  assign n2954 = x137 & ~n2953 ;
  assign n2955 = ~n2950 & ~n2954 ;
  assign n2956 = x138 & ~n2955 ;
  assign n2957 = ~n2946 & ~n2956 ;
  assign n2960 = n2957 & ~x264 ;
  assign n2961 = ~n2959 & ~n2960 ;
  assign n2962 = x90 & n2332 ;
  assign n2963 = x94 & n2344 ;
  assign n2964 = ~n2962 & ~n2963 ;
  assign n2965 = x138 & ~n2964 ;
  assign n2966 = x78 & ~x136 ;
  assign n2967 = x33 & x136 ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = x137 & ~n2968 ;
  assign n2970 = ~x63 & x136 ;
  assign n2971 = ~x74 & ~x136 ;
  assign n2972 = ~n2970 & ~n2971 ;
  assign n2973 = ~x137 & ~n2972 ;
  assign n2974 = ~n2969 & ~n2973 ;
  assign n2975 = ~x138 & ~n2974 ;
  assign n2976 = ~n2965 & ~n2975 ;
  assign n2993 = ~n2976 & x265 ;
  assign n2977 = ~x90 & n2344 ;
  assign n2978 = ~x94 & n2332 ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = ~x138 & ~n2979 ;
  assign n2981 = ~x78 & x136 ;
  assign n2982 = ~x33 & ~x136 ;
  assign n2983 = ~n2981 & ~n2982 ;
  assign n2984 = ~x137 & ~n2983 ;
  assign n2985 = x63 & ~x136 ;
  assign n2986 = x74 & x136 ;
  assign n2987 = ~n2985 & ~n2986 ;
  assign n2988 = x137 & ~n2987 ;
  assign n2989 = ~n2984 & ~n2988 ;
  assign n2990 = x138 & ~n2989 ;
  assign n2991 = ~n2980 & ~n2990 ;
  assign n2994 = n2991 & ~x265 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = x99 & n2332 ;
  assign n2997 = ~x112 & n2344 ;
  assign n2998 = ~n2996 & ~n2997 ;
  assign n2999 = x138 & ~n2998 ;
  assign n3000 = ~x68 & x136 ;
  assign n3001 = ~x73 & ~x136 ;
  assign n3002 = ~n3000 & ~n3001 ;
  assign n3003 = ~x137 & ~n3002 ;
  assign n3004 = x84 & ~x136 ;
  assign n3005 = x32 & x136 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = x137 & ~n3006 ;
  assign n3008 = ~n3003 & ~n3007 ;
  assign n3009 = ~x138 & ~n3008 ;
  assign n3010 = ~n2999 & ~n3009 ;
  assign n3027 = ~n3010 & x266 ;
  assign n3011 = ~x99 & n2344 ;
  assign n3012 = x112 & n2332 ;
  assign n3013 = ~n3011 & ~n3012 ;
  assign n3014 = ~x138 & ~n3013 ;
  assign n3015 = x68 & ~x136 ;
  assign n3016 = x73 & x136 ;
  assign n3017 = ~n3015 & ~n3016 ;
  assign n3018 = x137 & ~n3017 ;
  assign n3019 = ~x84 & x136 ;
  assign n3020 = ~x32 & ~x136 ;
  assign n3021 = ~n3019 & ~n3020 ;
  assign n3022 = ~x137 & ~n3021 ;
  assign n3023 = ~n3018 & ~n3022 ;
  assign n3024 = x138 & ~n3023 ;
  assign n3025 = ~n3014 & ~n3024 ;
  assign n3028 = n3025 & ~x266 ;
  assign n3029 = ~n3027 & ~n3028 ;
  assign n3030 = x92 & x138 ;
  assign n3031 = ~x70 & ~x138 ;
  assign n3032 = ~n3030 & ~n3031 ;
  assign n3033 = x136 & ~n3032 ;
  assign n3034 = x125 & x138 ;
  assign n3035 = ~x75 & ~x138 ;
  assign n3036 = ~n3034 & ~n3035 ;
  assign n3037 = ~x136 & ~n3036 ;
  assign n3038 = ~n3033 & ~n3037 ;
  assign n3039 = ~x137 & ~n3038 ;
  assign n3040 = x80 & ~x138 ;
  assign n3041 = x100 & x138 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = ~x136 & ~n3042 ;
  assign n3044 = x35 & n2628 ;
  assign n3045 = ~n3043 & ~n3044 ;
  assign n3046 = x137 & ~n3045 ;
  assign n3047 = ~n3039 & ~n3046 ;
  assign n3067 = ~n3047 & x267 ;
  assign n3048 = ~x92 & ~x138 ;
  assign n3049 = x70 & x138 ;
  assign n3050 = ~n3048 & ~n3049 ;
  assign n3051 = ~x136 & ~n3050 ;
  assign n3052 = ~x125 & ~x138 ;
  assign n3053 = x75 & x138 ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = x136 & ~n3054 ;
  assign n3056 = ~n3051 & ~n3055 ;
  assign n3057 = x137 & ~n3056 ;
  assign n3058 = ~x80 & x138 ;
  assign n3059 = ~x100 & ~x138 ;
  assign n3060 = ~n3058 & ~n3059 ;
  assign n3061 = x136 & ~n3060 ;
  assign n3062 = ~x35 & n2647 ;
  assign n3063 = ~n3061 & ~n3062 ;
  assign n3064 = ~x137 & ~n3063 ;
  assign n3065 = ~n3057 & ~n3064 ;
  assign n3068 = n3065 & ~x267 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = n1279 & n2669 ;
  assign n3071 = ~x27 & n3070 ;
  assign n3072 = ~n1133 & ~n3071 ;
  assign n3073 = ~x129 & ~n3072 ;
  assign n3074 = ~x3 & n3073 ;
  assign n3081 = n3074 & x268 ;
  assign n3075 = n1293 & n2677 ;
  assign n3076 = x27 & n3075 ;
  assign n3077 = ~n1181 & ~n3076 ;
  assign n3078 = x129 & ~n3077 ;
  assign n3079 = x3 & n3078 ;
  assign n3082 = ~n3079 & ~x268 ;
  assign n3083 = ~n3081 & ~n3082 ;
  assign n3084 = x98 & x138 ;
  assign n3085 = ~x71 & ~x138 ;
  assign n3086 = ~n3084 & ~n3085 ;
  assign n3087 = x136 & ~n3086 ;
  assign n3088 = ~x76 & ~x138 ;
  assign n3089 = x23 & x138 ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = ~x136 & ~n3090 ;
  assign n3092 = ~n3087 & ~n3091 ;
  assign n3093 = ~x137 & ~n3092 ;
  assign n3094 = x36 & n2628 ;
  assign n3095 = x81 & ~x138 ;
  assign n3096 = x97 & x138 ;
  assign n3097 = ~n3095 & ~n3096 ;
  assign n3098 = ~x136 & ~n3097 ;
  assign n3099 = ~n3094 & ~n3098 ;
  assign n3100 = x137 & ~n3099 ;
  assign n3101 = ~n3093 & ~n3100 ;
  assign n3121 = ~n3101 & x269 ;
  assign n3102 = ~x98 & ~x138 ;
  assign n3103 = x71 & x138 ;
  assign n3104 = ~n3102 & ~n3103 ;
  assign n3105 = ~x136 & ~n3104 ;
  assign n3106 = x76 & x138 ;
  assign n3107 = ~x23 & ~x138 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = x136 & ~n3108 ;
  assign n3110 = ~n3105 & ~n3109 ;
  assign n3111 = x137 & ~n3110 ;
  assign n3112 = ~x36 & n2647 ;
  assign n3113 = ~x81 & x138 ;
  assign n3114 = ~x97 & ~x138 ;
  assign n3115 = ~n3113 & ~n3114 ;
  assign n3116 = x136 & ~n3115 ;
  assign n3117 = ~n3112 & ~n3116 ;
  assign n3118 = ~x137 & ~n3117 ;
  assign n3119 = ~n3111 & ~n3118 ;
  assign n3122 = n3119 & ~x269 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = x88 & x138 ;
  assign n3125 = ~x64 & ~x138 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = x136 & ~n3126 ;
  assign n3128 = x120 & x138 ;
  assign n3129 = ~x67 & ~x138 ;
  assign n3130 = ~n3128 & ~n3129 ;
  assign n3131 = ~x136 & ~n3130 ;
  assign n3132 = ~n3127 & ~n3131 ;
  assign n3133 = ~x137 & ~n3132 ;
  assign n3134 = x86 & ~x138 ;
  assign n3135 = x111 & x138 ;
  assign n3136 = ~n3134 & ~n3135 ;
  assign n3137 = ~x136 & ~n3136 ;
  assign n3138 = x30 & n2628 ;
  assign n3139 = ~n3137 & ~n3138 ;
  assign n3140 = x137 & ~n3139 ;
  assign n3141 = ~n3133 & ~n3140 ;
  assign n3161 = ~n3141 & x270 ;
  assign n3142 = ~x88 & ~x138 ;
  assign n3143 = x64 & x138 ;
  assign n3144 = ~n3142 & ~n3143 ;
  assign n3145 = ~x136 & ~n3144 ;
  assign n3146 = ~x120 & ~x138 ;
  assign n3147 = x67 & x138 ;
  assign n3148 = ~n3146 & ~n3147 ;
  assign n3149 = x136 & ~n3148 ;
  assign n3150 = ~n3145 & ~n3149 ;
  assign n3151 = x137 & ~n3150 ;
  assign n3152 = ~x86 & x138 ;
  assign n3153 = ~x111 & ~x138 ;
  assign n3154 = ~n3152 & ~n3153 ;
  assign n3155 = x136 & ~n3154 ;
  assign n3156 = ~x30 & n2647 ;
  assign n3157 = ~n3155 & ~n3156 ;
  assign n3158 = ~x137 & ~n3157 ;
  assign n3159 = ~n3151 & ~n3158 ;
  assign n3162 = n3159 & ~x270 ;
  assign n3163 = ~n3161 & ~n3162 ;
  assign n3164 = ~n1157 & n1304 ;
  assign n3165 = ~n1303 & ~n3164 ;
  assign n3166 = ~x129 & ~n3165 ;
  assign n3167 = ~x3 & n3166 ;
  assign n3168 = x116 & n3167 ;
  assign n3175 = n3168 & x271 ;
  assign n3169 = ~n1205 & n1303 ;
  assign n3170 = ~n1304 & ~n3169 ;
  assign n3171 = x129 & ~n3170 ;
  assign n3172 = x3 & n3171 ;
  assign n3173 = ~x116 & n3172 ;
  assign n3176 = ~n3173 & ~x271 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = ~x97 & n1175 ;
  assign n3179 = ~n1223 & ~n3178 ;
  assign n3180 = ~x129 & ~n3179 ;
  assign n3181 = ~x3 & n3180 ;
  assign n3182 = x116 & n3181 ;
  assign n3189 = n3182 & x272 ;
  assign n3183 = x97 & n1223 ;
  assign n3184 = ~n1175 & ~n3183 ;
  assign n3185 = x129 & ~n3184 ;
  assign n3186 = x3 & n3185 ;
  assign n3187 = ~x116 & n3186 ;
  assign n3190 = ~n3187 & ~x272 ;
  assign n3191 = ~n3189 & ~n3190 ;
  assign n3192 = x111 & ~n2808 ;
  assign n3193 = ~x136 & x139 ;
  assign n3194 = ~x137 & x138 ;
  assign n3195 = x82 & n3194 ;
  assign n3196 = n3193 & n3195 ;
  assign n3197 = ~n3192 & ~n3196 ;
  assign n3198 = n2329 & ~n3197 ;
  assign n3199 = ~x129 & n3198 ;
  assign n3209 = n3199 & x273 ;
  assign n3200 = ~x111 & ~n2817 ;
  assign n3201 = x136 & ~x139 ;
  assign n3202 = x137 & ~x138 ;
  assign n3203 = ~x82 & n3202 ;
  assign n3204 = n3201 & n3203 ;
  assign n3205 = ~n3200 & ~n3204 ;
  assign n3206 = n2341 & ~n3205 ;
  assign n3207 = x129 & n3206 ;
  assign n3210 = ~n3207 & ~x273 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = ~x136 & x141 ;
  assign n3213 = n3195 & n3212 ;
  assign n3214 = ~x112 & ~n2808 ;
  assign n3215 = ~n3213 & ~n3214 ;
  assign n3216 = n2329 & ~n3215 ;
  assign n3217 = ~x129 & n3216 ;
  assign n3225 = n3217 & x274 ;
  assign n3218 = x136 & ~x141 ;
  assign n3219 = n3203 & n3218 ;
  assign n3220 = x112 & ~n2817 ;
  assign n3221 = ~n3219 & ~n3220 ;
  assign n3222 = n2341 & ~n3221 ;
  assign n3223 = x129 & n3222 ;
  assign n3226 = ~n3223 & ~x274 ;
  assign n3227 = ~n3225 & ~n3226 ;
  assign n3228 = ~x54 & ~x113 ;
  assign n3229 = ~x11 & ~x22 ;
  assign n3230 = x54 & ~n3229 ;
  assign n3231 = ~n3228 & ~n3230 ;
  assign n3232 = ~x129 & ~n3231 ;
  assign n3233 = ~x3 & n3232 ;
  assign n3241 = n3233 & x275 ;
  assign n3234 = x54 & x113 ;
  assign n3235 = x11 & x22 ;
  assign n3236 = ~x54 & ~n3235 ;
  assign n3237 = ~n3234 & ~n3236 ;
  assign n3238 = x129 & ~n3237 ;
  assign n3239 = x3 & n3238 ;
  assign n3242 = ~n3239 & ~x275 ;
  assign n3243 = ~n3241 & ~n3242 ;
  assign n3245 = ~n2141 & x276 ;
  assign n3246 = n2144 & ~x276 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = ~x136 & x140 ;
  assign n3249 = n3195 & n3248 ;
  assign n3250 = ~x115 & ~n2808 ;
  assign n3251 = ~n3249 & ~n3250 ;
  assign n3252 = n2329 & ~n3251 ;
  assign n3253 = ~x129 & n3252 ;
  assign n3261 = n3253 & x277 ;
  assign n3254 = x136 & ~x140 ;
  assign n3255 = n3203 & n3254 ;
  assign n3256 = x115 & ~n2817 ;
  assign n3257 = ~n3255 & ~n3256 ;
  assign n3258 = n2341 & ~n3257 ;
  assign n3259 = x129 & n3258 ;
  assign n3262 = ~n3259 & ~x277 ;
  assign n3263 = ~n3261 & ~n3262 ;
  assign n3264 = ~x4 & ~x12 ;
  assign n3265 = ~x7 & ~x9 ;
  assign n3266 = n3264 & n3265 ;
  assign n3267 = ~x129 & ~n3266 ;
  assign n3268 = ~x3 & n3267 ;
  assign n3269 = x54 & n3268 ;
  assign n3277 = n3269 & x278 ;
  assign n3270 = x4 & x12 ;
  assign n3271 = x7 & x9 ;
  assign n3272 = n3270 & n3271 ;
  assign n3273 = x129 & ~n3272 ;
  assign n3274 = x3 & n3273 ;
  assign n3275 = ~x54 & n3274 ;
  assign n3278 = ~n3275 & ~x278 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = x122 & ~x129 ;
  assign n3283 = ~n3280 & x279 ;
  assign n3281 = ~x122 & x129 ;
  assign n3284 = n3281 & ~x279 ;
  assign n3285 = ~n3283 & ~n3284 ;
  assign n3286 = ~x54 & x118 ;
  assign n3287 = x54 & ~x59 ;
  assign n3288 = n761 & n3287 ;
  assign n3289 = ~n3286 & ~n3288 ;
  assign n3290 = ~x129 & ~n3289 ;
  assign n3297 = n3290 & x280 ;
  assign n3291 = x54 & ~x118 ;
  assign n3292 = ~x54 & x59 ;
  assign n3293 = n773 & n3292 ;
  assign n3294 = ~n3291 & ~n3293 ;
  assign n3295 = x129 & ~n3294 ;
  assign n3298 = ~n3295 & ~x280 ;
  assign n3299 = ~n3297 & ~n3298 ;
  assign n3300 = ~x129 & ~n1144 ;
  assign n3303 = n3300 & x281 ;
  assign n3301 = x129 & ~n1192 ;
  assign n3304 = ~n3301 & ~x281 ;
  assign n3305 = ~n3303 & ~n3304 ;
  assign n3306 = ~x110 & ~x120 ;
  assign n3307 = ~x3 & n3306 ;
  assign n3308 = ~x129 & ~n3307 ;
  assign n3309 = ~x111 & n3308 ;
  assign n3315 = n3309 & x282 ;
  assign n3310 = x110 & x120 ;
  assign n3311 = x3 & n3310 ;
  assign n3312 = x129 & ~n3311 ;
  assign n3313 = x111 & n3312 ;
  assign n3316 = ~n3313 & ~x282 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = x81 & x120 ;
  assign n3319 = ~x129 & n3318 ;
  assign n3323 = n3319 & x283 ;
  assign n3320 = ~x81 & ~x120 ;
  assign n3321 = x129 & n3320 ;
  assign n3324 = ~n3321 & ~x283 ;
  assign n3325 = ~n3323 & ~n3324 ;
  assign n3326 = ~x129 & ~x134 ;
  assign n3329 = ~n3326 & x284 ;
  assign n3327 = x129 & x134 ;
  assign n3330 = n3327 & ~x284 ;
  assign n3331 = ~n3329 & ~n3330 ;
  assign n3332 = ~x129 & ~x135 ;
  assign n3335 = ~n3332 & x285 ;
  assign n3333 = x129 & x135 ;
  assign n3336 = n3333 & ~x285 ;
  assign n3337 = ~n3335 & ~n3336 ;
  assign n3338 = x57 & ~x129 ;
  assign n3341 = n3338 & x286 ;
  assign n3339 = ~x57 & x129 ;
  assign n3342 = ~n3339 & ~x286 ;
  assign n3343 = ~n3341 & ~n3342 ;
  assign n3344 = ~x96 & x125 ;
  assign n3345 = ~x3 & ~n3344 ;
  assign n3346 = ~x129 & ~n3345 ;
  assign n3351 = n3346 & x287 ;
  assign n3347 = x96 & ~x125 ;
  assign n3348 = x3 & ~n3347 ;
  assign n3349 = x129 & ~n3348 ;
  assign n3352 = ~n3349 & ~x287 ;
  assign n3353 = ~n3351 & ~n3352 ;
  assign n3354 = ~x126 & x132 ;
  assign n3355 = x133 & n3354 ;
  assign n3359 = n3355 & x288 ;
  assign n3356 = x126 & ~x132 ;
  assign n3357 = ~x133 & n3356 ;
  assign n3360 = ~n3357 & ~x288 ;
  assign n3361 = ~n3359 & ~n3360 ;
  assign y0 = ~n151 ;
  assign y1 = ~n155 ;
  assign y2 = ~n159 ;
  assign y3 = ~n163 ;
  assign y4 = ~n167 ;
  assign y5 = ~n171 ;
  assign y6 = ~n175 ;
  assign y7 = ~n179 ;
  assign y8 = ~n183 ;
  assign y9 = ~n187 ;
  assign y10 = ~n191 ;
  assign y11 = ~n195 ;
  assign y12 = x159 ;
  assign y13 = ~n200 ;
  assign y14 = ~n204 ;
  assign y15 = ~n306 ;
  assign y16 = ~n384 ;
  assign y17 = ~n462 ;
  assign y18 = ~n494 ;
  assign y19 = ~n518 ;
  assign y20 = ~n558 ;
  assign y21 = ~n590 ;
  assign y22 = ~n622 ;
  assign y23 = ~n650 ;
  assign y24 = ~n680 ;
  assign y25 = ~n708 ;
  assign y26 = ~n732 ;
  assign y27 = ~n756 ;
  assign y28 = ~n784 ;
  assign y29 = ~n808 ;
  assign y30 = ~n866 ;
  assign y31 = ~n886 ;
  assign y32 = ~n920 ;
  assign y33 = ~n940 ;
  assign y34 = ~n964 ;
  assign y35 = ~n1016 ;
  assign y36 = ~n1038 ;
  assign y37 = ~n1068 ;
  assign y38 = ~n1078 ;
  assign y39 = ~n1132 ;
  assign y40 = ~n1232 ;
  assign y41 = ~n1266 ;
  assign y42 = ~n1298 ;
  assign y43 = ~n1377 ;
  assign y44 = ~n1443 ;
  assign y45 = ~n1461 ;
  assign y46 = ~n1479 ;
  assign y47 = ~n1497 ;
  assign y48 = ~n1515 ;
  assign y49 = ~n1533 ;
  assign y50 = ~n1551 ;
  assign y51 = ~n1569 ;
  assign y52 = ~n1587 ;
  assign y53 = ~n1637 ;
  assign y54 = ~n1655 ;
  assign y55 = ~n1695 ;
  assign y56 = ~n1735 ;
  assign y57 = ~n1773 ;
  assign y58 = ~n1811 ;
  assign y59 = ~n1833 ;
  assign y60 = ~n1881 ;
  assign y61 = ~n1917 ;
  assign y62 = ~n1953 ;
  assign y63 = ~n1997 ;
  assign y64 = ~n2039 ;
  assign y65 = ~n2077 ;
  assign y66 = ~n2086 ;
  assign y67 = ~n2098 ;
  assign y68 = ~n2128 ;
  assign y69 = ~n2140 ;
  assign y70 = ~n2150 ;
  assign y71 = ~n2198 ;
  assign y72 = ~n2236 ;
  assign y73 = ~n2256 ;
  assign y74 = ~n2303 ;
  assign y75 = ~n2315 ;
  assign y76 = ~n2325 ;
  assign y77 = ~n2353 ;
  assign y78 = ~n2367 ;
  assign y79 = ~n2381 ;
  assign y80 = ~n2395 ;
  assign y81 = ~n2411 ;
  assign y82 = ~n2423 ;
  assign y83 = ~n2437 ;
  assign y84 = ~n2451 ;
  assign y85 = ~n2465 ;
  assign y86 = ~n2479 ;
  assign y87 = ~n2491 ;
  assign y88 = ~n2503 ;
  assign y89 = ~n2515 ;
  assign y90 = ~n2527 ;
  assign y91 = ~n2539 ;
  assign y92 = ~n2551 ;
  assign y93 = ~n2565 ;
  assign y94 = ~n2577 ;
  assign y95 = ~n2589 ;
  assign y96 = ~n2601 ;
  assign y97 = ~n2613 ;
  assign y98 = ~n2655 ;
  assign y99 = ~n2667 ;
  assign y100 = ~n2687 ;
  assign y101 = ~n2699 ;
  assign y102 = ~n2711 ;
  assign y103 = ~n2725 ;
  assign y104 = ~n2737 ;
  assign y105 = ~n2749 ;
  assign y106 = ~n2761 ;
  assign y107 = ~n2773 ;
  assign y108 = ~n2785 ;
  assign y109 = ~n2805 ;
  assign y110 = ~n2827 ;
  assign y111 = ~n2839 ;
  assign y112 = ~n2851 ;
  assign y113 = ~n2863 ;
  assign y114 = ~n2875 ;
  assign y115 = ~n2887 ;
  assign y116 = ~n2927 ;
  assign y117 = ~n2961 ;
  assign y118 = ~n2995 ;
  assign y119 = ~n3029 ;
  assign y120 = ~n3069 ;
  assign y121 = ~n3083 ;
  assign y122 = ~n3123 ;
  assign y123 = ~n3163 ;
  assign y124 = ~n3177 ;
  assign y125 = ~n3191 ;
  assign y126 = ~n3211 ;
  assign y127 = ~n3227 ;
  assign y128 = ~n3243 ;
  assign y129 = ~n3247 ;
  assign y130 = ~n3263 ;
  assign y131 = ~n3279 ;
  assign y132 = ~n3285 ;
  assign y133 = ~n3299 ;
  assign y134 = ~n3305 ;
  assign y135 = ~n3317 ;
  assign y136 = ~n3325 ;
  assign y137 = ~n3331 ;
  assign y138 = ~n3337 ;
  assign y139 = ~n3343 ;
  assign y140 = ~n3353 ;
  assign y141 = ~n3361 ;
endmodule
